magic
tech gf180mcuD
timestamp 1759194789
<< properties >>
string GDS_END 1928558
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1927594
<< end >>
