magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
use M1_NACTIVE4310590878120_256x8m81  M1_NACTIVE4310590878120_256x8m81_0
timestamp 1762296095
transform 1 0 1337 0 1 4210
box 0 0 1 1
use M1_POLY24310590878153_256x8m81  M1_POLY24310590878153_256x8m81_0
timestamp 1762296095
transform 1 0 865 0 1 7450
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1762296095
transform -1 0 824 0 1 4092
box 0 0 1 1
use M2_M1$$43376684_256x8m81  M2_M1$$43376684_256x8m81_0
timestamp 1762296095
transform -1 0 599 0 1 2099
box 0 0 1 1
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_0
timestamp 1762296095
transform 1 0 1113 0 1 10532
box 0 0 1 1
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_1
timestamp 1762296095
transform 1 0 881 0 1 10532
box 0 0 1 1
use M2_M1$$43379756_256x8m81  M2_M1$$43379756_256x8m81_2
timestamp 1762296095
transform 1 0 441 0 1 10532
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_0
timestamp 1762296095
transform 1 0 441 0 1 9494
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_1
timestamp 1762296095
transform 1 0 889 0 1 9494
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_2
timestamp 1762296095
transform 1 0 1337 0 1 9494
box 0 0 1 1
use M2_M1$$47500332_256x8m81  M2_M1$$47500332_256x8m81_0
timestamp 1762296095
transform 1 0 1054 0 1 6153
box 0 0 1 1
use M2_M1$$47500332_256x8m81  M2_M1$$47500332_256x8m81_1
timestamp 1762296095
transform 1 0 602 0 1 6153
box 0 0 1 1
use M2_M1$$47500332_256x8m81  M2_M1$$47500332_256x8m81_2
timestamp 1762296095
transform 1 0 1337 0 1 6153
box 0 0 1 1
use M2_M1$$47640620_256x8m81  M2_M1$$47640620_256x8m81_0
timestamp 1762296095
transform 1 0 1337 0 1 1526
box 0 0 1 1
use M2_M1$$47640620_256x8m81  M2_M1$$47640620_256x8m81_1
timestamp 1762296095
transform 1 0 1054 0 1 1526
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_0
timestamp 1762296095
transform 1 0 1337 0 1 2505
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_1
timestamp 1762296095
transform 1 0 1054 0 1 2505
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_2
timestamp 1762296095
transform 1 0 441 0 1 9494
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_3
timestamp 1762296095
transform 1 0 889 0 1 9494
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_4
timestamp 1762296095
transform 1 0 1337 0 1 9494
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_0
timestamp 1762296095
transform 1 0 1337 0 1 438
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_1
timestamp 1762296095
transform 1 0 1054 0 1 438
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_2
timestamp 1762296095
transform 1 0 881 0 1 10532
box 0 0 1 1
use M3_M2$$47333420_256x8m81  M3_M2$$47333420_256x8m81_3
timestamp 1762296095
transform 1 0 441 0 1 10532
box 0 0 1 1
use M3_M2$$47644716_256x8m81  M3_M2$$47644716_256x8m81_0
timestamp 1762296095
transform 1 0 1054 0 1 6153
box 0 0 1 1
use M3_M2$$47644716_256x8m81  M3_M2$$47644716_256x8m81_1
timestamp 1762296095
transform 1 0 602 0 1 6153
box 0 0 1 1
use M3_M2$$47644716_256x8m81  M3_M2$$47644716_256x8m81_2
timestamp 1762296095
transform 1 0 1337 0 1 6153
box 0 0 1 1
use nmos_1p2$$47641644_256x8m81  nmos_1p2$$47641644_256x8m81_0
timestamp 1762296095
transform -1 0 1254 0 -1 11038
box -31 0 -30 1
use nmos_1p2$$47641644_256x8m81  nmos_1p2$$47641644_256x8m81_1
timestamp 1762296095
transform -1 0 806 0 -1 11038
box -31 0 -30 1
use nmos_1p2$$47641644_256x8m81  nmos_1p2$$47641644_256x8m81_2
timestamp 1762296095
transform -1 0 582 0 -1 11038
box -31 0 -30 1
use nmos_1p2$$47641644_256x8m81  nmos_1p2$$47641644_256x8m81_3
timestamp 1762296095
transform -1 0 1030 0 -1 11038
box -31 0 -30 1
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_0
timestamp 1762296095
transform -1 0 1030 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_1
timestamp 1762296095
transform -1 0 806 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_2
timestamp 1762296095
transform -1 0 582 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47513644_256x8m81  pmos_1p2$$47513644_256x8m81_3
timestamp 1762296095
transform -1 0 1254 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47642668_256x8m81  pmos_1p2$$47642668_256x8m81_0
timestamp 1762296095
transform -1 0 964 0 1 3908
box -31 0 -30 1
use pmos_1p2$$47643692_256x8m81  pmos_1p2$$47643692_256x8m81_0
timestamp 1762296095
transform -1 0 740 0 1 3908
box -31 0 -30 1
<< properties >>
string GDS_END 585702
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 577364
<< end >>
