magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< nwell >>
rect 13512 13500 70089 70434
<< obsm1 >>
rect 13108 13108 71000 71000
<< obsm2 >>
rect 13606 13594 70901 70890
<< metal3 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 40272 70213 40328 70269
rect 41872 70219 41928 70275
rect 54672 70194 54728 70250
rect 56272 70196 56328 70252
rect 59472 70201 59528 70257
rect 61072 70204 61128 70260
rect 62672 70205 62728 70261
rect 65874 70210 65930 70266
rect 67472 70214 67528 70270
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70412 42800 70488 45799
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< obsm3 >>
rect 17060 70740 17140 70890
rect 20260 70740 20340 70890
rect 23460 70740 23540 70890
rect 25060 70740 25140 70890
rect 26660 70740 26740 70890
rect 29860 70740 29940 70890
rect 33060 70740 33140 70890
rect 36260 70740 36340 70890
rect 39460 70740 39540 70890
rect 41060 70740 41140 70890
rect 42660 70740 42740 70890
rect 45860 70740 45940 70890
rect 49060 70740 49140 70890
rect 50660 70740 50740 70890
rect 52260 70740 52340 70890
rect 53860 70740 53940 70890
rect 55460 70740 55540 70890
rect 57060 70740 57140 70890
rect 58660 70740 58740 70890
rect 60260 70740 60340 70890
rect 61860 70740 61940 70890
rect 63460 70740 63540 70890
rect 65060 70740 65140 70890
rect 66660 70740 66740 70890
rect 68260 70740 68340 70890
rect 69738 70740 71000 70890
rect 14000 70275 71000 70740
rect 14000 70269 41872 70275
rect 14000 70213 40272 70269
rect 40328 70219 41872 70269
rect 41928 70270 71000 70275
rect 41928 70266 67472 70270
rect 41928 70261 65874 70266
rect 41928 70260 62672 70261
rect 41928 70257 61072 70260
rect 41928 70252 59472 70257
rect 41928 70250 56272 70252
rect 41928 70219 54672 70250
rect 40328 70213 54672 70219
rect 14000 70194 54672 70213
rect 54728 70196 56272 70250
rect 56328 70201 59472 70252
rect 59528 70204 61072 70257
rect 61128 70205 62672 70260
rect 62728 70210 65874 70261
rect 65930 70214 67472 70266
rect 67528 70214 71000 70270
rect 65930 70210 71000 70214
rect 62728 70205 71000 70210
rect 61128 70204 71000 70205
rect 59528 70201 71000 70204
rect 56328 70196 71000 70201
rect 54728 70194 71000 70196
rect 14000 69738 71000 70194
rect 14000 68340 70740 69738
rect 14000 68260 71000 68340
rect 14000 66740 70740 68260
rect 14000 66660 71000 66740
rect 14000 65140 70740 66660
rect 14000 65060 71000 65140
rect 14000 63540 70740 65060
rect 14000 63460 71000 63540
rect 14000 61940 70740 63460
rect 14000 61860 71000 61940
rect 14000 60340 70740 61860
rect 14000 60260 71000 60340
rect 14000 58740 70740 60260
rect 14000 58660 71000 58740
rect 14000 57140 70740 58660
rect 14000 57060 71000 57140
rect 14000 55540 70740 57060
rect 14000 55460 71000 55540
rect 14000 53940 70740 55460
rect 14000 53860 71000 53940
rect 14000 52340 70740 53860
rect 14000 52260 71000 52340
rect 14000 50740 70740 52260
rect 14000 50660 71000 50740
rect 14000 49140 70740 50660
rect 14000 49060 71000 49140
rect 14000 45940 70740 49060
rect 14000 45859 71000 45940
rect 14000 42740 70352 45859
rect 70548 42740 71000 45859
rect 14000 42660 71000 42740
rect 14000 41140 70740 42660
rect 14000 41060 71000 41140
rect 14000 39540 70740 41060
rect 14000 39460 71000 39540
rect 14000 36340 70740 39460
rect 14000 36260 71000 36340
rect 14000 33140 70740 36260
rect 14000 33060 71000 33140
rect 14000 29940 70740 33060
rect 14000 29860 71000 29940
rect 14000 26740 70740 29860
rect 14000 26660 71000 26740
rect 14000 25140 70740 26660
rect 14000 25060 71000 25140
rect 14000 23540 70740 25060
rect 14000 23460 71000 23540
rect 14000 20340 70740 23460
rect 14000 20260 71000 20340
rect 14000 17140 70740 20260
rect 14000 17060 71000 17140
rect 14000 14000 70740 17060
<< metal4 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 15396 47287 15472 70800
rect 18596 48623 18672 70800
rect 20400 70151 23400 70227
rect 23600 70160 25000 70236
rect 25200 70164 26600 70240
rect 28064 52629 28140 70800
rect 31264 53967 31340 70800
rect 34408 70196 34464 70252
rect 37664 56640 37740 70800
rect 40272 70213 40328 70269
rect 41872 70219 41928 70275
rect 42800 70148 45800 70224
rect 46000 70171 49000 70247
rect 49200 70176 50600 70252
rect 50800 70177 52200 70253
rect 52400 70182 53800 70258
rect 54672 70194 54728 70250
rect 56272 70196 56328 70252
rect 57928 64675 57938 70800
rect 59472 70201 59528 70257
rect 61072 70204 61128 70260
rect 62672 70205 62728 70261
rect 64327 70219 64329 70221
rect 65874 70210 65930 70266
rect 67472 70214 67528 70270
rect 69001 69258 69077 70800
rect 70395 68400 70471 69678
rect 70800 68400 71000 69678
rect 70402 66800 70478 68200
rect 70800 66800 71000 68200
rect 70400 65200 70476 66600
rect 70800 65200 71000 66600
rect 70399 63600 70475 65000
rect 70800 63600 71000 65000
rect 70393 62000 70469 63400
rect 70800 62000 71000 63400
rect 70391 60400 70467 61800
rect 70800 60400 71000 61800
rect 70389 58800 70465 60200
rect 70800 58800 71000 60200
rect 70386 57200 70462 58600
rect 70800 57200 71000 58600
rect 70384 55600 70460 57000
rect 70800 55600 71000 57000
rect 70382 54000 70458 55400
rect 70800 54000 71000 55400
rect 70390 53138 70446 53194
rect 70800 52400 71000 53800
rect 70517 51406 70573 51462
rect 70800 50800 71000 52200
rect 70516 49938 70572 49994
rect 70800 49200 71000 50600
rect 70800 47604 71000 49000
rect 60617 47528 71000 47604
rect 70800 46000 71000 47528
rect 70412 42800 70488 45799
rect 70407 41200 70483 42600
rect 70800 41200 71000 42600
rect 70401 39600 70477 41000
rect 70800 39600 71000 41000
rect 70394 36400 70470 39400
rect 70800 36400 71000 39400
rect 70384 33200 70460 36200
rect 70800 33200 71000 36200
rect 70800 31604 71000 33000
rect 58681 31528 71000 31604
rect 70800 30000 71000 31528
rect 70800 28404 71000 29800
rect 58681 28328 71000 28404
rect 70800 26800 71000 28328
rect 70428 25200 70504 26600
rect 70800 25200 71000 26600
rect 70424 23600 70500 25000
rect 70800 23600 71000 25000
rect 70415 20969 70491 22751
rect 70800 20400 71000 23400
rect 70800 18936 71000 20200
rect 58405 18860 71000 18936
rect 70800 17200 71000 18860
rect 70404 14000 70480 17000
rect 70800 14000 71000 17000
<< obsm4 >>
rect 14000 47227 15336 70740
rect 17060 70740 17140 70800
rect 15532 48563 18536 70740
rect 20260 70740 20340 70800
rect 23460 70740 23540 70800
rect 25060 70740 25140 70800
rect 26660 70740 26740 70800
rect 18732 70300 28004 70740
rect 18732 70296 25140 70300
rect 18732 70287 23540 70296
rect 18732 70091 20340 70287
rect 23460 70100 23540 70287
rect 25060 70104 25140 70296
rect 26660 70104 28004 70300
rect 25060 70100 28004 70104
rect 23460 70091 28004 70100
rect 18732 52569 28004 70091
rect 29860 70740 29940 70800
rect 28200 53907 31204 70740
rect 33060 70740 33140 70800
rect 36260 70740 36340 70800
rect 31400 70252 37604 70740
rect 31400 70196 34408 70252
rect 34464 70196 37604 70252
rect 31400 56580 37604 70196
rect 39460 70740 39540 70800
rect 41060 70740 41140 70800
rect 42660 70740 42740 70800
rect 45860 70740 45940 70800
rect 49060 70740 49140 70800
rect 50660 70740 50740 70800
rect 52260 70740 52340 70800
rect 53860 70740 53940 70800
rect 55460 70740 55540 70800
rect 57060 70740 57140 70800
rect 37800 70335 57868 70740
rect 37800 70329 41812 70335
rect 37800 70153 40212 70329
rect 40388 70159 41812 70329
rect 41988 70318 57868 70335
rect 41988 70313 52340 70318
rect 41988 70312 50740 70313
rect 41988 70307 49140 70312
rect 41988 70284 45940 70307
rect 41988 70159 42740 70284
rect 40388 70153 42740 70159
rect 37800 70088 42740 70153
rect 45860 70111 45940 70284
rect 49060 70116 49140 70307
rect 50660 70117 50740 70312
rect 52260 70122 52340 70313
rect 53860 70312 57868 70318
rect 53860 70310 56212 70312
rect 53860 70134 54612 70310
rect 54788 70136 56212 70310
rect 56388 70136 57868 70312
rect 54788 70134 57868 70136
rect 53860 70122 57868 70134
rect 52260 70117 57868 70122
rect 50660 70116 57868 70117
rect 49060 70111 57868 70116
rect 45860 70088 57868 70111
rect 37800 64615 57868 70088
rect 58660 70740 58740 70800
rect 60260 70740 60340 70800
rect 61860 70740 61940 70800
rect 63460 70740 63540 70800
rect 65060 70740 65140 70800
rect 66660 70740 66740 70800
rect 68260 70740 68340 70800
rect 57998 70330 68941 70740
rect 57998 70326 67412 70330
rect 57998 70321 65814 70326
rect 57998 70320 62612 70321
rect 57998 70317 61012 70320
rect 57998 70141 59412 70317
rect 59588 70144 61012 70317
rect 61188 70145 62612 70320
rect 62788 70281 65814 70321
rect 62788 70159 64267 70281
rect 64389 70159 65814 70281
rect 62788 70150 65814 70159
rect 65990 70154 67412 70326
rect 67588 70154 68941 70330
rect 65990 70150 68941 70154
rect 62788 70145 68941 70150
rect 61188 70144 68941 70145
rect 59588 70141 68941 70144
rect 57998 69198 68941 70141
rect 69738 70740 71000 70800
rect 69137 69738 71000 70740
rect 69137 69198 70335 69738
rect 57998 68340 70335 69198
rect 70531 68340 70740 69738
rect 57998 68260 71000 68340
rect 57998 66740 70342 68260
rect 70538 66740 70740 68260
rect 57998 66660 71000 66740
rect 57998 65140 70340 66660
rect 70536 65140 70740 66660
rect 57998 65060 71000 65140
rect 57998 64615 70339 65060
rect 37800 63540 70339 64615
rect 70535 63540 70740 65060
rect 37800 63460 71000 63540
rect 37800 61940 70333 63460
rect 70529 61940 70740 63460
rect 37800 61860 71000 61940
rect 37800 60340 70331 61860
rect 70527 60340 70740 61860
rect 37800 60260 71000 60340
rect 37800 58740 70329 60260
rect 70525 58740 70740 60260
rect 37800 58660 71000 58740
rect 37800 57140 70326 58660
rect 70522 57140 70740 58660
rect 37800 57060 71000 57140
rect 37800 56580 70324 57060
rect 31400 55540 70324 56580
rect 70520 55540 70740 57060
rect 31400 55460 71000 55540
rect 31400 53940 70322 55460
rect 70518 53940 70740 55460
rect 31400 53907 71000 53940
rect 28200 53860 71000 53907
rect 28200 53254 70740 53860
rect 28200 53078 70330 53254
rect 70506 53078 70740 53254
rect 28200 52569 70740 53078
rect 18732 52340 70740 52569
rect 18732 52260 71000 52340
rect 18732 51462 70740 52260
rect 18732 51406 70517 51462
rect 70573 51406 70740 51462
rect 18732 50740 70740 51406
rect 18732 50660 71000 50740
rect 18732 49994 70740 50660
rect 18732 49938 70516 49994
rect 70572 49938 70740 49994
rect 18732 49140 70740 49938
rect 18732 49060 71000 49140
rect 18732 48563 70740 49060
rect 15532 47664 70740 48563
rect 15532 47468 60557 47664
rect 15532 47227 70740 47468
rect 14000 45940 70740 47227
rect 14000 45859 71000 45940
rect 14000 42740 70352 45859
rect 70548 42740 71000 45859
rect 14000 42660 71000 42740
rect 14000 41140 70347 42660
rect 70543 41140 70740 42660
rect 14000 41060 71000 41140
rect 14000 39540 70341 41060
rect 70537 39540 70740 41060
rect 14000 39460 71000 39540
rect 14000 36340 70334 39460
rect 70530 36340 70740 39460
rect 14000 36260 71000 36340
rect 14000 33140 70324 36260
rect 70520 33140 70740 36260
rect 14000 33060 71000 33140
rect 14000 31664 70740 33060
rect 14000 31468 58621 31664
rect 14000 29940 70740 31468
rect 14000 29860 71000 29940
rect 14000 28464 70740 29860
rect 14000 28268 58621 28464
rect 14000 26740 70740 28268
rect 14000 26660 71000 26740
rect 14000 25140 70368 26660
rect 70564 25140 70740 26660
rect 14000 25060 71000 25140
rect 14000 23540 70364 25060
rect 70560 23540 70740 25060
rect 14000 23460 71000 23540
rect 14000 22811 70740 23460
rect 14000 20909 70355 22811
rect 70551 20909 70740 22811
rect 14000 20340 70740 20909
rect 14000 20260 71000 20340
rect 14000 18996 70740 20260
rect 14000 18800 58345 18996
rect 14000 17140 70740 18800
rect 14000 17060 71000 17140
rect 14000 14000 70344 17060
rect 70540 14000 70740 17060
<< metal5 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 15396 47287 15472 70800
rect 18596 48623 18672 70800
rect 20400 70151 23400 70227
rect 23600 70160 25000 70236
rect 25200 70164 26600 70240
rect 28064 52629 28140 70800
rect 31264 53967 31340 70800
rect 34408 70196 34464 70252
rect 37664 56640 37740 70800
rect 49200 70176 50600 70252
rect 51462 61435 51538 70800
rect 54662 62769 54738 70800
rect 56262 63432 56338 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 62662 66090 62738 70800
rect 64262 66762 64338 70800
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70393 62000 70469 63400
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70390 53138 70446 53194
rect 70800 52400 71000 53800
rect 70517 51406 70573 51462
rect 70800 50800 71000 52200
rect 70516 49938 70572 49994
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70407 41200 70483 42600
rect 70800 41200 71000 42600
rect 70401 39600 70477 41000
rect 70800 39600 71000 41000
rect 70394 36400 70470 39400
rect 70800 36400 71000 39400
rect 70384 33200 70460 36200
rect 70800 33200 71000 36200
rect 70800 31604 71000 33000
rect 58681 31528 71000 31604
rect 70800 30000 71000 31528
rect 70800 28404 71000 29800
rect 58681 28328 71000 28404
rect 70800 26800 71000 28328
rect 70800 26070 71000 26600
rect 51293 25994 71000 26070
rect 70800 25200 71000 25994
rect 70424 23600 70500 25000
rect 70800 23600 71000 25000
rect 70415 20400 70491 23400
rect 70800 20400 71000 23400
rect 70800 18936 71000 20200
rect 58405 18860 71000 18936
rect 70800 17200 71000 18860
rect 70404 14000 70480 17000
rect 70800 14000 71000 17000
<< obsm5 >>
rect 14000 47167 15276 70680
rect 15592 48503 18476 70680
rect 18792 70360 27944 70680
rect 18792 70356 25080 70360
rect 18792 70347 23480 70356
rect 18792 70031 20280 70347
rect 26720 70044 27944 70360
rect 25120 70040 27944 70044
rect 23520 70031 27944 70040
rect 18792 52509 27944 70031
rect 28260 53847 31144 70680
rect 31460 70372 37544 70680
rect 31460 70076 34288 70372
rect 34584 70076 37544 70372
rect 31460 56520 37544 70076
rect 37860 70372 51342 70680
rect 37860 70056 49080 70372
rect 50720 70056 51342 70372
rect 37860 61315 51342 70056
rect 51658 62649 54542 70680
rect 55520 70680 56142 71000
rect 54858 63312 56142 70680
rect 56458 70680 57080 71000
rect 56458 65970 62542 70680
rect 62858 66642 64142 70680
rect 69798 70680 71000 71000
rect 64458 69798 71000 70680
rect 64458 66642 70680 69798
rect 62858 65970 70680 66642
rect 56458 63520 70680 65970
rect 56458 63312 70273 63520
rect 54858 62649 70273 63312
rect 51658 61880 70273 62649
rect 70589 61880 70680 63520
rect 51658 61315 70680 61880
rect 37860 56520 70680 61315
rect 31460 53847 70680 56520
rect 28260 53194 70680 53847
rect 28260 53138 70390 53194
rect 70446 53138 70680 53194
rect 28260 52509 70680 53138
rect 18792 51582 70680 52509
rect 18792 51286 70397 51582
rect 18792 50114 70680 51286
rect 18792 49818 70396 50114
rect 18792 48503 70680 49818
rect 15592 47167 70680 48503
rect 14000 45880 70680 47167
rect 14000 42720 71000 45880
rect 14000 41120 70287 42720
rect 14000 39520 70281 41120
rect 70603 41080 70680 42720
rect 14000 36320 70274 39520
rect 70597 39480 70680 41080
rect 14000 33080 70264 36320
rect 70590 36280 70680 39480
rect 70580 33080 70680 36280
rect 14000 31724 70680 33080
rect 14000 31408 58561 31724
rect 14000 28524 70680 31408
rect 14000 28208 58561 28524
rect 14000 26190 70680 28208
rect 14000 25874 51173 26190
rect 14000 25120 70680 25874
rect 14000 23520 70304 25120
rect 14000 20280 70295 23520
rect 70620 23480 70680 25120
rect 70611 20280 70680 23480
rect 14000 19056 70680 20280
rect 14000 18740 58285 19056
rect 14000 17120 70680 18740
rect 14000 14000 70284 17120
rect 70600 14000 70680 17120
<< labels >>
rlabel metal3 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70412 42800 70488 45799 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 55600 70800 57000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 56262 63432 56338 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 66800 70800 68200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 66800 71000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58800 70800 60200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 58800 71000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 55600 71000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54000 70800 55400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 54000 71000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 52400 70800 53800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 52400 71000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 42800 70800 45800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54662 62769 54738 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 41200 70800 42600 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 41200 71000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 36400 70800 39400 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 36400 71000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 33200 70800 36200 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 33200 71000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 30000 70800 33000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 30000 71000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 26800 70800 29800 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 26800 71000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70800 25000 71000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 23600 71000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 34408 70196 34464 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 34408 70196 34464 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70160 25000 70236 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 28064 52629 28140 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 31264 53967 31340 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 37664 56640 37740 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70394 36400 70470 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70407 41200 70483 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58681 31528 70800 31604 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70384 33200 70460 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70424 23600 70500 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 58681 28328 70800 28404 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 59472 70201 59528 70257 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 59472 70201 59528 70257 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 56272 70196 56328 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 56272 70196 56328 70252 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 52400 70182 53800 70258 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 42800 70148 45800 70224 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 28064 52629 28140 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 23600 70160 25000 70236 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70402 66800 70478 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70389 58800 70465 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70382 54000 70458 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70412 42800 70488 45799 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70394 36400 70470 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 58681 31528 70800 31604 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70424 23600 70500 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 67472 70214 67528 70270 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 67472 70214 67528 70270 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 54672 70194 54728 70250 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 54672 70194 54728 70250 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 41872 70219 41928 70275 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 41872 70219 41928 70275 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 37664 56640 37740 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 31264 53967 31340 70800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70384 55600 70460 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70390 53138 70446 53194 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70390 53138 70446 53194 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70407 41200 70483 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70384 33200 70460 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 58681 28328 70800 28404 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 68400 70800 69678 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 68400 71000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 65200 70800 66600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 65200 71000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 60400 70800 61800 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 60400 71000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 57200 70800 58600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 57200 71000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 46000 70800 49000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 46000 71000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 39600 70800 41000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 39600 71000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70800 26600 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 25200 71000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 20400 70800 23400 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 20400 71000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 17200 70800 20200 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 17200 71000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14000 70800 17000 71000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 14000 71000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70164 26600 70240 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 15396 47287 15472 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 18596 48623 18672 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 20400 70151 23400 70227 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 58405 18860 70800 18936 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70404 14000 70480 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70415 20400 70491 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 51293 25994 70800 26070 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70401 39600 70477 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 69001 69258 69077 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 65874 70210 65930 70266 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 65874 70210 65930 70266 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 40272 70213 40328 70269 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 40272 70213 40328 70269 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 18596 48623 18672 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70395 68400 70471 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70391 60400 70467 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 60617 47528 70800 47604 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70428 25200 70504 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70404 14000 70480 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 61072 70204 61128 70260 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 61072 70204 61128 70260 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 57928 64675 57938 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 46000 70171 49000 70247 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 25200 70164 26600 70240 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 20400 70151 23400 70227 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 15396 47287 15472 70800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70400 65200 70476 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70386 57200 70462 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70401 39600 70477 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70415 20969 70491 22751 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 58405 18860 70800 18936 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 62000 70800 63400 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 62000 71000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 50800 70800 52200 71000 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 50800 71000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70517 51406 70573 51462 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70517 51406 70573 51462 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70393 62000 70469 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 51462 61435 51538 70800 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 62662 66090 62738 70800 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 62672 70205 62728 70261 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 62672 70205 62728 70261 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 50800 70177 52200 70253 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70393 62000 70469 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 63600 70800 65000 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 63600 71000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 49200 70800 50600 71000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 49200 71000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70516 49938 70572 49994 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70516 49938 70572 49994 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 49200 70176 50600 70252 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 64262 66762 64338 70800 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 49200 70176 50600 70252 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 64327 70219 64329 70221 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70399 63600 70475 65000 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string LEFclass ENDCAP BOTTOMLEFT
string LEFsite GF_COR_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 17526940
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17516202
<< end >>
