magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
<< metal1 >>
rect 3 3059 203 3071
rect 3 3007 15 3059
rect 67 3007 139 3059
rect 191 3007 203 3059
rect 3 2935 203 3007
rect 3 2883 15 2935
rect 67 2883 139 2935
rect 191 2883 203 2935
rect 3 2811 203 2883
rect 3 2759 15 2811
rect 67 2759 139 2811
rect 191 2759 203 2811
rect 3 2687 203 2759
rect 3 2635 15 2687
rect 67 2635 139 2687
rect 191 2635 203 2687
rect 3 2563 203 2635
rect 3 2511 15 2563
rect 67 2511 139 2563
rect 191 2511 203 2563
rect 3 2439 203 2511
rect 3 2387 15 2439
rect 67 2387 139 2439
rect 191 2387 203 2439
rect 3 2315 203 2387
rect 3 2263 15 2315
rect 67 2263 139 2315
rect 191 2263 203 2315
rect 3 2191 203 2263
rect 3 2139 15 2191
rect 67 2139 139 2191
rect 191 2139 203 2191
rect 3 2127 203 2139
rect 1020 3059 1220 3071
rect 1020 3007 1032 3059
rect 1084 3007 1156 3059
rect 1208 3007 1220 3059
rect 1020 2935 1220 3007
rect 1020 2883 1032 2935
rect 1084 2883 1156 2935
rect 1208 2883 1220 2935
rect 1020 2811 1220 2883
rect 1020 2759 1032 2811
rect 1084 2759 1156 2811
rect 1208 2759 1220 2811
rect 1020 2687 1220 2759
rect 1020 2635 1032 2687
rect 1084 2635 1156 2687
rect 1208 2635 1220 2687
rect 1020 2563 1220 2635
rect 1020 2511 1032 2563
rect 1084 2511 1156 2563
rect 1208 2511 1220 2563
rect 1020 2439 1220 2511
rect 1020 2387 1032 2439
rect 1084 2387 1156 2439
rect 1208 2387 1220 2439
rect 1020 2315 1220 2387
rect 1020 2263 1032 2315
rect 1084 2263 1156 2315
rect 1208 2263 1220 2315
rect 1020 2191 1220 2263
rect 1020 2139 1032 2191
rect 1084 2139 1156 2191
rect 1208 2139 1220 2191
rect 1020 2127 1220 2139
<< via1 >>
rect 15 3007 67 3059
rect 139 3007 191 3059
rect 15 2883 67 2935
rect 139 2883 191 2935
rect 15 2759 67 2811
rect 139 2759 191 2811
rect 15 2635 67 2687
rect 139 2635 191 2687
rect 15 2511 67 2563
rect 139 2511 191 2563
rect 15 2387 67 2439
rect 139 2387 191 2439
rect 15 2263 67 2315
rect 139 2263 191 2315
rect 15 2139 67 2191
rect 139 2139 191 2191
rect 1032 3007 1084 3059
rect 1156 3007 1208 3059
rect 1032 2883 1084 2935
rect 1156 2883 1208 2935
rect 1032 2759 1084 2811
rect 1156 2759 1208 2811
rect 1032 2635 1084 2687
rect 1156 2635 1208 2687
rect 1032 2511 1084 2563
rect 1156 2511 1208 2563
rect 1032 2387 1084 2439
rect 1156 2387 1208 2439
rect 1032 2263 1084 2315
rect 1156 2263 1208 2315
rect 1032 2139 1084 2191
rect 1156 2139 1208 2191
<< metal2 >>
rect -7 18269 217 18431
rect -7 18213 16 18269
rect 72 18213 140 18269
rect 196 18213 217 18269
rect -7 18145 217 18213
rect -7 18089 16 18145
rect 72 18089 140 18145
rect 196 18089 217 18145
rect -7 18021 217 18089
rect -7 17965 16 18021
rect 72 17965 140 18021
rect 196 17965 217 18021
rect -7 17897 217 17965
rect -7 17841 16 17897
rect 72 17841 140 17897
rect 196 17841 217 17897
rect -7 17773 217 17841
rect -7 17717 16 17773
rect 72 17717 140 17773
rect 196 17717 217 17773
rect -7 17582 217 17717
rect -7 17526 16 17582
rect 72 17526 140 17582
rect 196 17526 217 17582
rect -7 17458 217 17526
rect -7 17402 16 17458
rect 72 17402 140 17458
rect 196 17402 217 17458
rect -7 17334 217 17402
rect -7 17278 16 17334
rect 72 17278 140 17334
rect 196 17278 217 17334
rect -7 17210 217 17278
rect -7 17154 16 17210
rect 72 17154 140 17210
rect 196 17154 217 17210
rect -7 17086 217 17154
rect -7 17030 16 17086
rect 72 17030 140 17086
rect 196 17030 217 17086
rect -7 16898 217 17030
rect -7 16842 16 16898
rect 72 16842 140 16898
rect 196 16842 217 16898
rect -7 16774 217 16842
rect -7 16718 16 16774
rect 72 16718 140 16774
rect 196 16718 217 16774
rect -7 16650 217 16718
rect -7 16594 16 16650
rect 72 16594 140 16650
rect 196 16594 217 16650
rect -7 16526 217 16594
rect -7 16470 16 16526
rect 72 16470 140 16526
rect 196 16470 217 16526
rect -7 16402 217 16470
rect -7 16346 16 16402
rect 72 16346 140 16402
rect 196 16346 217 16402
rect -7 13292 217 16346
rect 1010 18269 1234 18431
rect 1010 18213 1033 18269
rect 1089 18213 1157 18269
rect 1213 18213 1234 18269
rect 1010 18145 1234 18213
rect 1010 18089 1033 18145
rect 1089 18089 1157 18145
rect 1213 18089 1234 18145
rect 1010 18021 1234 18089
rect 1010 17965 1033 18021
rect 1089 17965 1157 18021
rect 1213 17965 1234 18021
rect 1010 17897 1234 17965
rect 1010 17841 1033 17897
rect 1089 17841 1157 17897
rect 1213 17841 1234 17897
rect 1010 17773 1234 17841
rect 1010 17717 1033 17773
rect 1089 17717 1157 17773
rect 1213 17717 1234 17773
rect 1010 17582 1234 17717
rect 1010 17526 1033 17582
rect 1089 17526 1157 17582
rect 1213 17526 1234 17582
rect 1010 17458 1234 17526
rect 1010 17402 1033 17458
rect 1089 17402 1157 17458
rect 1213 17402 1234 17458
rect 1010 17334 1234 17402
rect 1010 17278 1033 17334
rect 1089 17278 1157 17334
rect 1213 17278 1234 17334
rect 1010 17210 1234 17278
rect 1010 17154 1033 17210
rect 1089 17154 1157 17210
rect 1213 17154 1234 17210
rect 1010 17086 1234 17154
rect 1010 17030 1033 17086
rect 1089 17030 1157 17086
rect 1213 17030 1234 17086
rect 1010 16898 1234 17030
rect 1010 16842 1033 16898
rect 1089 16842 1157 16898
rect 1213 16842 1234 16898
rect 1010 16774 1234 16842
rect 1010 16718 1033 16774
rect 1089 16718 1157 16774
rect 1213 16718 1234 16774
rect 1010 16650 1234 16718
rect 1010 16594 1033 16650
rect 1089 16594 1157 16650
rect 1213 16594 1234 16650
rect 1010 16526 1234 16594
rect 1010 16470 1033 16526
rect 1089 16470 1157 16526
rect 1213 16470 1234 16526
rect 1010 16402 1234 16470
rect 1010 16346 1033 16402
rect 1089 16346 1157 16402
rect 1213 16346 1234 16402
rect -7 13236 16 13292
rect 72 13236 140 13292
rect 196 13236 217 13292
rect -7 13168 217 13236
rect -7 13112 16 13168
rect 72 13112 140 13168
rect 196 13112 217 13168
rect -7 13044 217 13112
rect -7 12988 16 13044
rect 72 12988 140 13044
rect 196 12988 217 13044
rect -7 12920 217 12988
rect -7 12864 16 12920
rect 72 12864 140 12920
rect 196 12864 217 12920
rect -7 12796 217 12864
rect -7 12740 16 12796
rect 72 12740 140 12796
rect 196 12740 217 12796
rect -7 12605 217 12740
rect -7 12549 16 12605
rect 72 12549 140 12605
rect 196 12549 217 12605
rect -7 12481 217 12549
rect -7 12425 16 12481
rect 72 12425 140 12481
rect 196 12425 217 12481
rect -7 12357 217 12425
rect -7 12301 16 12357
rect 72 12301 140 12357
rect 196 12301 217 12357
rect -7 12233 217 12301
rect -7 12177 16 12233
rect 72 12177 140 12233
rect 196 12177 217 12233
rect -7 12109 217 12177
rect -7 12053 16 12109
rect 72 12053 140 12109
rect 196 12053 217 12109
rect -7 9403 217 12053
rect -7 9347 16 9403
rect 72 9347 140 9403
rect 196 9347 217 9403
rect -7 9279 217 9347
rect -7 9223 16 9279
rect 72 9223 140 9279
rect 196 9223 217 9279
rect -7 9155 217 9223
rect -7 9099 16 9155
rect 72 9099 140 9155
rect 196 9099 217 9155
rect -7 9031 217 9099
rect -7 8975 16 9031
rect 72 8975 140 9031
rect 196 8975 217 9031
rect -7 8907 217 8975
rect -7 8851 16 8907
rect 72 8851 140 8907
rect 196 8851 217 8907
rect -7 7964 217 8851
rect -7 7908 16 7964
rect 72 7908 140 7964
rect 196 7908 217 7964
rect -7 7840 217 7908
rect -7 7784 16 7840
rect 72 7784 140 7840
rect 196 7784 217 7840
rect -7 7716 217 7784
rect -7 7660 16 7716
rect 72 7660 140 7716
rect 196 7660 217 7716
rect -7 5680 217 7660
rect -7 5624 16 5680
rect 72 5624 140 5680
rect 196 5624 217 5680
rect -7 5556 217 5624
rect -7 5500 16 5556
rect 72 5500 140 5556
rect 196 5500 217 5556
rect -7 5432 217 5500
rect -7 5376 16 5432
rect 72 5376 140 5432
rect 196 5376 217 5432
rect -7 4667 217 5376
rect -7 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 217 4667
rect -7 4543 217 4611
rect -7 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 217 4543
rect -7 4419 217 4487
rect -7 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 217 4419
rect -7 3059 217 4363
rect 495 15840 719 16012
rect 495 15784 516 15840
rect 572 15784 640 15840
rect 696 15784 719 15840
rect 495 15716 719 15784
rect 495 15660 516 15716
rect 572 15660 640 15716
rect 696 15660 719 15716
rect 495 15592 719 15660
rect 495 15536 516 15592
rect 572 15536 640 15592
rect 696 15536 719 15592
rect 495 15468 719 15536
rect 495 15412 516 15468
rect 572 15412 640 15468
rect 696 15412 719 15468
rect 495 15344 719 15412
rect 495 15288 516 15344
rect 572 15288 640 15344
rect 696 15288 719 15344
rect 495 15220 719 15288
rect 495 15164 516 15220
rect 572 15164 640 15220
rect 696 15164 719 15220
rect 495 15096 719 15164
rect 495 15040 516 15096
rect 572 15040 640 15096
rect 696 15040 719 15096
rect 495 14972 719 15040
rect 495 14916 516 14972
rect 572 14916 640 14972
rect 696 14916 719 14972
rect 495 14848 719 14916
rect 495 14792 516 14848
rect 572 14792 640 14848
rect 696 14792 719 14848
rect 495 14724 719 14792
rect 495 14668 516 14724
rect 572 14668 640 14724
rect 696 14668 719 14724
rect 495 14600 719 14668
rect 495 14544 516 14600
rect 572 14544 640 14600
rect 696 14544 719 14600
rect 495 14476 719 14544
rect 495 14420 516 14476
rect 572 14420 640 14476
rect 696 14420 719 14476
rect 495 14352 719 14420
rect 495 14296 516 14352
rect 572 14296 640 14352
rect 696 14296 719 14352
rect 495 14228 719 14296
rect 495 14172 516 14228
rect 572 14172 640 14228
rect 696 14172 719 14228
rect 495 14104 719 14172
rect 495 14048 516 14104
rect 572 14048 640 14104
rect 696 14048 719 14104
rect 495 11233 719 14048
rect 495 11177 516 11233
rect 572 11177 640 11233
rect 696 11177 719 11233
rect 495 11109 719 11177
rect 495 11053 516 11109
rect 572 11053 640 11109
rect 696 11053 719 11109
rect 495 10985 719 11053
rect 495 10929 516 10985
rect 572 10929 640 10985
rect 696 10929 719 10985
rect 495 10861 719 10929
rect 495 10805 516 10861
rect 572 10805 640 10861
rect 696 10805 719 10861
rect 495 10737 719 10805
rect 495 10681 516 10737
rect 572 10681 640 10737
rect 696 10681 719 10737
rect 495 10613 719 10681
rect 495 10557 516 10613
rect 572 10557 640 10613
rect 696 10557 719 10613
rect 495 10489 719 10557
rect 495 10433 516 10489
rect 572 10433 640 10489
rect 696 10433 719 10489
rect 495 10365 719 10433
rect 495 10309 516 10365
rect 572 10309 640 10365
rect 696 10309 719 10365
rect 495 10241 719 10309
rect 495 10185 516 10241
rect 572 10185 640 10241
rect 696 10185 719 10241
rect 495 10117 719 10185
rect 495 10061 516 10117
rect 572 10061 640 10117
rect 696 10061 719 10117
rect 495 7366 719 10061
rect 495 7310 516 7366
rect 572 7310 640 7366
rect 696 7310 719 7366
rect 495 7242 719 7310
rect 495 7186 516 7242
rect 572 7186 640 7242
rect 696 7186 719 7242
rect 495 7118 719 7186
rect 495 7062 516 7118
rect 572 7062 640 7118
rect 696 7062 719 7118
rect 495 6403 719 7062
rect 495 6347 516 6403
rect 572 6347 640 6403
rect 696 6347 719 6403
rect 495 6279 719 6347
rect 495 6223 516 6279
rect 572 6223 640 6279
rect 696 6223 719 6279
rect 495 6155 719 6223
rect 495 6099 516 6155
rect 572 6099 640 6155
rect 696 6099 719 6155
rect 495 4037 719 6099
rect 495 3981 516 4037
rect 572 3981 640 4037
rect 696 3981 719 4037
rect 495 3913 719 3981
rect 495 3857 516 3913
rect 572 3857 640 3913
rect 696 3857 719 3913
rect 495 3789 719 3857
rect 495 3733 516 3789
rect 572 3733 640 3789
rect 696 3733 719 3789
rect 495 3665 719 3733
rect 495 3609 516 3665
rect 572 3609 640 3665
rect 696 3609 719 3665
rect 495 3541 719 3609
rect 495 3485 516 3541
rect 572 3485 640 3541
rect 696 3485 719 3541
rect 495 3417 719 3485
rect 495 3361 516 3417
rect 572 3361 640 3417
rect 696 3361 719 3417
rect 495 3293 719 3361
rect 495 3237 516 3293
rect 572 3237 640 3293
rect 696 3237 719 3293
rect 495 3169 719 3237
rect 495 3113 516 3169
rect 572 3113 640 3169
rect 696 3113 719 3169
rect 495 3065 719 3113
rect 1010 13292 1234 16346
rect 1010 13236 1033 13292
rect 1089 13236 1157 13292
rect 1213 13236 1234 13292
rect 1010 13168 1234 13236
rect 1010 13112 1033 13168
rect 1089 13112 1157 13168
rect 1213 13112 1234 13168
rect 1010 13044 1234 13112
rect 1010 12988 1033 13044
rect 1089 12988 1157 13044
rect 1213 12988 1234 13044
rect 1010 12920 1234 12988
rect 1010 12864 1033 12920
rect 1089 12864 1157 12920
rect 1213 12864 1234 12920
rect 1010 12796 1234 12864
rect 1010 12740 1033 12796
rect 1089 12740 1157 12796
rect 1213 12740 1234 12796
rect 1010 12605 1234 12740
rect 1010 12549 1033 12605
rect 1089 12549 1157 12605
rect 1213 12549 1234 12605
rect 1010 12481 1234 12549
rect 1010 12425 1033 12481
rect 1089 12425 1157 12481
rect 1213 12425 1234 12481
rect 1010 12357 1234 12425
rect 1010 12301 1033 12357
rect 1089 12301 1157 12357
rect 1213 12301 1234 12357
rect 1010 12233 1234 12301
rect 1010 12177 1033 12233
rect 1089 12177 1157 12233
rect 1213 12177 1234 12233
rect 1010 12109 1234 12177
rect 1010 12053 1033 12109
rect 1089 12053 1157 12109
rect 1213 12053 1234 12109
rect 1010 9403 1234 12053
rect 1010 9347 1033 9403
rect 1089 9347 1157 9403
rect 1213 9347 1234 9403
rect 1010 9279 1234 9347
rect 1010 9223 1033 9279
rect 1089 9223 1157 9279
rect 1213 9223 1234 9279
rect 1010 9155 1234 9223
rect 1010 9099 1033 9155
rect 1089 9099 1157 9155
rect 1213 9099 1234 9155
rect 1010 9031 1234 9099
rect 1010 8975 1033 9031
rect 1089 8975 1157 9031
rect 1213 8975 1234 9031
rect 1010 8907 1234 8975
rect 1010 8851 1033 8907
rect 1089 8851 1157 8907
rect 1213 8851 1234 8907
rect 1010 7964 1234 8851
rect 1010 7908 1033 7964
rect 1089 7908 1157 7964
rect 1213 7908 1234 7964
rect 1010 7840 1234 7908
rect 1010 7784 1033 7840
rect 1089 7784 1157 7840
rect 1213 7784 1234 7840
rect 1010 7716 1234 7784
rect 1010 7660 1033 7716
rect 1089 7660 1157 7716
rect 1213 7660 1234 7716
rect 1010 5680 1234 7660
rect 1010 5624 1033 5680
rect 1089 5624 1157 5680
rect 1213 5624 1234 5680
rect 1010 5556 1234 5624
rect 1010 5500 1033 5556
rect 1089 5500 1157 5556
rect 1213 5500 1234 5556
rect 1010 5432 1234 5500
rect 1010 5376 1033 5432
rect 1089 5376 1157 5432
rect 1213 5376 1234 5432
rect 1010 4667 1234 5376
rect 1010 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1234 4667
rect 1010 4543 1234 4611
rect 1010 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1234 4543
rect 1010 4419 1234 4487
rect 1010 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1234 4419
rect -7 3007 15 3059
rect 67 3007 139 3059
rect 191 3007 217 3059
rect -7 2935 217 3007
rect -7 2883 15 2935
rect 67 2883 139 2935
rect 191 2883 217 2935
rect -7 2811 217 2883
rect -7 2759 15 2811
rect 67 2759 139 2811
rect 191 2759 217 2811
rect -7 2687 217 2759
rect -7 2635 15 2687
rect 67 2635 139 2687
rect 191 2635 217 2687
rect -7 2563 217 2635
rect -7 2511 15 2563
rect 67 2511 139 2563
rect 191 2511 217 2563
rect -7 2439 217 2511
rect -7 2387 15 2439
rect 67 2387 139 2439
rect 191 2387 217 2439
rect -7 2315 217 2387
rect -7 2263 15 2315
rect 67 2263 139 2315
rect 191 2263 217 2315
rect -7 2191 217 2263
rect -7 2139 15 2191
rect 67 2139 139 2191
rect 191 2139 217 2191
rect -7 2115 217 2139
rect 1010 3059 1234 4363
rect 1010 3007 1032 3059
rect 1084 3007 1156 3059
rect 1208 3007 1234 3059
rect 1010 2935 1234 3007
rect 1010 2883 1032 2935
rect 1084 2883 1156 2935
rect 1208 2883 1234 2935
rect 1010 2811 1234 2883
rect 1010 2759 1032 2811
rect 1084 2759 1156 2811
rect 1208 2759 1234 2811
rect 1010 2687 1234 2759
rect 1010 2635 1032 2687
rect 1084 2635 1156 2687
rect 1208 2635 1234 2687
rect 1010 2563 1234 2635
rect 1010 2511 1032 2563
rect 1084 2511 1156 2563
rect 1208 2511 1234 2563
rect 1010 2439 1234 2511
rect 1010 2387 1032 2439
rect 1084 2387 1156 2439
rect 1208 2387 1234 2439
rect 1010 2315 1234 2387
rect 1010 2263 1032 2315
rect 1084 2263 1156 2315
rect 1208 2263 1234 2315
rect 1010 2191 1234 2263
rect 1010 2139 1032 2191
rect 1084 2139 1156 2191
rect 1208 2139 1234 2191
rect 1010 2115 1234 2139
<< via2 >>
rect 16 18213 72 18269
rect 140 18213 196 18269
rect 16 18089 72 18145
rect 140 18089 196 18145
rect 16 17965 72 18021
rect 140 17965 196 18021
rect 16 17841 72 17897
rect 140 17841 196 17897
rect 16 17717 72 17773
rect 140 17717 196 17773
rect 16 17526 72 17582
rect 140 17526 196 17582
rect 16 17402 72 17458
rect 140 17402 196 17458
rect 16 17278 72 17334
rect 140 17278 196 17334
rect 16 17154 72 17210
rect 140 17154 196 17210
rect 16 17030 72 17086
rect 140 17030 196 17086
rect 16 16842 72 16898
rect 140 16842 196 16898
rect 16 16718 72 16774
rect 140 16718 196 16774
rect 16 16594 72 16650
rect 140 16594 196 16650
rect 16 16470 72 16526
rect 140 16470 196 16526
rect 16 16346 72 16402
rect 140 16346 196 16402
rect 1033 18213 1089 18269
rect 1157 18213 1213 18269
rect 1033 18089 1089 18145
rect 1157 18089 1213 18145
rect 1033 17965 1089 18021
rect 1157 17965 1213 18021
rect 1033 17841 1089 17897
rect 1157 17841 1213 17897
rect 1033 17717 1089 17773
rect 1157 17717 1213 17773
rect 1033 17526 1089 17582
rect 1157 17526 1213 17582
rect 1033 17402 1089 17458
rect 1157 17402 1213 17458
rect 1033 17278 1089 17334
rect 1157 17278 1213 17334
rect 1033 17154 1089 17210
rect 1157 17154 1213 17210
rect 1033 17030 1089 17086
rect 1157 17030 1213 17086
rect 1033 16842 1089 16898
rect 1157 16842 1213 16898
rect 1033 16718 1089 16774
rect 1157 16718 1213 16774
rect 1033 16594 1089 16650
rect 1157 16594 1213 16650
rect 1033 16470 1089 16526
rect 1157 16470 1213 16526
rect 1033 16346 1089 16402
rect 1157 16346 1213 16402
rect 16 13236 72 13292
rect 140 13236 196 13292
rect 16 13112 72 13168
rect 140 13112 196 13168
rect 16 12988 72 13044
rect 140 12988 196 13044
rect 16 12864 72 12920
rect 140 12864 196 12920
rect 16 12740 72 12796
rect 140 12740 196 12796
rect 16 12549 72 12605
rect 140 12549 196 12605
rect 16 12425 72 12481
rect 140 12425 196 12481
rect 16 12301 72 12357
rect 140 12301 196 12357
rect 16 12177 72 12233
rect 140 12177 196 12233
rect 16 12053 72 12109
rect 140 12053 196 12109
rect 16 9347 72 9403
rect 140 9347 196 9403
rect 16 9223 72 9279
rect 140 9223 196 9279
rect 16 9099 72 9155
rect 140 9099 196 9155
rect 16 8975 72 9031
rect 140 8975 196 9031
rect 16 8851 72 8907
rect 140 8851 196 8907
rect 16 7908 72 7964
rect 140 7908 196 7964
rect 16 7784 72 7840
rect 140 7784 196 7840
rect 16 7660 72 7716
rect 140 7660 196 7716
rect 16 5624 72 5680
rect 140 5624 196 5680
rect 16 5500 72 5556
rect 140 5500 196 5556
rect 16 5376 72 5432
rect 140 5376 196 5432
rect 16 4611 72 4667
rect 140 4611 196 4667
rect 16 4487 72 4543
rect 140 4487 196 4543
rect 16 4363 72 4419
rect 140 4363 196 4419
rect 516 15784 572 15840
rect 640 15784 696 15840
rect 516 15660 572 15716
rect 640 15660 696 15716
rect 516 15536 572 15592
rect 640 15536 696 15592
rect 516 15412 572 15468
rect 640 15412 696 15468
rect 516 15288 572 15344
rect 640 15288 696 15344
rect 516 15164 572 15220
rect 640 15164 696 15220
rect 516 15040 572 15096
rect 640 15040 696 15096
rect 516 14916 572 14972
rect 640 14916 696 14972
rect 516 14792 572 14848
rect 640 14792 696 14848
rect 516 14668 572 14724
rect 640 14668 696 14724
rect 516 14544 572 14600
rect 640 14544 696 14600
rect 516 14420 572 14476
rect 640 14420 696 14476
rect 516 14296 572 14352
rect 640 14296 696 14352
rect 516 14172 572 14228
rect 640 14172 696 14228
rect 516 14048 572 14104
rect 640 14048 696 14104
rect 516 11177 572 11233
rect 640 11177 696 11233
rect 516 11053 572 11109
rect 640 11053 696 11109
rect 516 10929 572 10985
rect 640 10929 696 10985
rect 516 10805 572 10861
rect 640 10805 696 10861
rect 516 10681 572 10737
rect 640 10681 696 10737
rect 516 10557 572 10613
rect 640 10557 696 10613
rect 516 10433 572 10489
rect 640 10433 696 10489
rect 516 10309 572 10365
rect 640 10309 696 10365
rect 516 10185 572 10241
rect 640 10185 696 10241
rect 516 10061 572 10117
rect 640 10061 696 10117
rect 516 7310 572 7366
rect 640 7310 696 7366
rect 516 7186 572 7242
rect 640 7186 696 7242
rect 516 7062 572 7118
rect 640 7062 696 7118
rect 516 6347 572 6403
rect 640 6347 696 6403
rect 516 6223 572 6279
rect 640 6223 696 6279
rect 516 6099 572 6155
rect 640 6099 696 6155
rect 516 3981 572 4037
rect 640 3981 696 4037
rect 516 3857 572 3913
rect 640 3857 696 3913
rect 516 3733 572 3789
rect 640 3733 696 3789
rect 516 3609 572 3665
rect 640 3609 696 3665
rect 516 3485 572 3541
rect 640 3485 696 3541
rect 516 3361 572 3417
rect 640 3361 696 3417
rect 516 3237 572 3293
rect 640 3237 696 3293
rect 516 3113 572 3169
rect 640 3113 696 3169
rect 1033 13236 1089 13292
rect 1157 13236 1213 13292
rect 1033 13112 1089 13168
rect 1157 13112 1213 13168
rect 1033 12988 1089 13044
rect 1157 12988 1213 13044
rect 1033 12864 1089 12920
rect 1157 12864 1213 12920
rect 1033 12740 1089 12796
rect 1157 12740 1213 12796
rect 1033 12549 1089 12605
rect 1157 12549 1213 12605
rect 1033 12425 1089 12481
rect 1157 12425 1213 12481
rect 1033 12301 1089 12357
rect 1157 12301 1213 12357
rect 1033 12177 1089 12233
rect 1157 12177 1213 12233
rect 1033 12053 1089 12109
rect 1157 12053 1213 12109
rect 1033 9347 1089 9403
rect 1157 9347 1213 9403
rect 1033 9223 1089 9279
rect 1157 9223 1213 9279
rect 1033 9099 1089 9155
rect 1157 9099 1213 9155
rect 1033 8975 1089 9031
rect 1157 8975 1213 9031
rect 1033 8851 1089 8907
rect 1157 8851 1213 8907
rect 1033 7908 1089 7964
rect 1157 7908 1213 7964
rect 1033 7784 1089 7840
rect 1157 7784 1213 7840
rect 1033 7660 1089 7716
rect 1157 7660 1213 7716
rect 1033 5624 1089 5680
rect 1157 5624 1213 5680
rect 1033 5500 1089 5556
rect 1157 5500 1213 5556
rect 1033 5376 1089 5432
rect 1157 5376 1213 5432
rect 1033 4611 1089 4667
rect 1157 4611 1213 4667
rect 1033 4487 1089 4543
rect 1157 4487 1213 4543
rect 1033 4363 1089 4419
rect 1157 4363 1213 4419
<< metal3 >>
rect 6 18269 206 18279
rect 6 18213 16 18269
rect 72 18213 140 18269
rect 196 18213 206 18269
rect 6 18145 206 18213
rect 6 18089 16 18145
rect 72 18089 140 18145
rect 196 18089 206 18145
rect 6 18021 206 18089
rect 6 17965 16 18021
rect 72 17965 140 18021
rect 196 17965 206 18021
rect 6 17897 206 17965
rect 6 17841 16 17897
rect 72 17841 140 17897
rect 196 17841 206 17897
rect 6 17773 206 17841
rect 6 17717 16 17773
rect 72 17717 140 17773
rect 196 17717 206 17773
rect 6 17707 206 17717
rect 1023 18269 1223 18279
rect 1023 18213 1033 18269
rect 1089 18213 1157 18269
rect 1213 18213 1223 18269
rect 1023 18145 1223 18213
rect 1023 18089 1033 18145
rect 1089 18089 1157 18145
rect 1213 18089 1223 18145
rect 1023 18021 1223 18089
rect 1023 17965 1033 18021
rect 1089 17965 1157 18021
rect 1213 17965 1223 18021
rect 1023 17897 1223 17965
rect 1023 17841 1033 17897
rect 1089 17841 1157 17897
rect 1213 17841 1223 17897
rect 1023 17773 1223 17841
rect 1023 17717 1033 17773
rect 1089 17717 1157 17773
rect 1213 17717 1223 17773
rect 1023 17707 1223 17717
rect 6 17582 206 17592
rect 6 17526 16 17582
rect 72 17526 140 17582
rect 196 17526 206 17582
rect 6 17458 206 17526
rect 6 17402 16 17458
rect 72 17402 140 17458
rect 196 17402 206 17458
rect 6 17334 206 17402
rect 6 17278 16 17334
rect 72 17278 140 17334
rect 196 17278 206 17334
rect 6 17210 206 17278
rect 6 17154 16 17210
rect 72 17154 140 17210
rect 196 17154 206 17210
rect 6 17086 206 17154
rect 6 17030 16 17086
rect 72 17030 140 17086
rect 196 17030 206 17086
rect 6 17020 206 17030
rect 1023 17582 1223 17592
rect 1023 17526 1033 17582
rect 1089 17526 1157 17582
rect 1213 17526 1223 17582
rect 1023 17458 1223 17526
rect 1023 17402 1033 17458
rect 1089 17402 1157 17458
rect 1213 17402 1223 17458
rect 1023 17334 1223 17402
rect 1023 17278 1033 17334
rect 1089 17278 1157 17334
rect 1213 17278 1223 17334
rect 1023 17210 1223 17278
rect 1023 17154 1033 17210
rect 1089 17154 1157 17210
rect 1213 17154 1223 17210
rect 1023 17086 1223 17154
rect 1023 17030 1033 17086
rect 1089 17030 1157 17086
rect 1213 17030 1223 17086
rect 1023 17020 1223 17030
rect 6 16898 206 16908
rect 6 16842 16 16898
rect 72 16842 140 16898
rect 196 16842 206 16898
rect 6 16774 206 16842
rect 6 16718 16 16774
rect 72 16718 140 16774
rect 196 16718 206 16774
rect 6 16650 206 16718
rect 6 16594 16 16650
rect 72 16594 140 16650
rect 196 16594 206 16650
rect 6 16526 206 16594
rect 6 16470 16 16526
rect 72 16470 140 16526
rect 196 16470 206 16526
rect 6 16402 206 16470
rect 6 16346 16 16402
rect 72 16346 140 16402
rect 196 16346 206 16402
rect 6 16336 206 16346
rect 1023 16898 1223 16908
rect 1023 16842 1033 16898
rect 1089 16842 1157 16898
rect 1213 16842 1223 16898
rect 1023 16774 1223 16842
rect 1023 16718 1033 16774
rect 1089 16718 1157 16774
rect 1213 16718 1223 16774
rect 1023 16650 1223 16718
rect 1023 16594 1033 16650
rect 1089 16594 1157 16650
rect 1213 16594 1223 16650
rect 1023 16526 1223 16594
rect 1023 16470 1033 16526
rect 1089 16470 1157 16526
rect 1213 16470 1223 16526
rect 1023 16402 1223 16470
rect 1023 16346 1033 16402
rect 1089 16346 1157 16402
rect 1213 16346 1223 16402
rect 1023 16336 1223 16346
rect 506 15840 706 15850
rect 506 15784 516 15840
rect 572 15784 640 15840
rect 696 15784 706 15840
rect 506 15716 706 15784
rect 506 15660 516 15716
rect 572 15660 640 15716
rect 696 15660 706 15716
rect 506 15592 706 15660
rect 506 15536 516 15592
rect 572 15536 640 15592
rect 696 15536 706 15592
rect 506 15468 706 15536
rect 506 15412 516 15468
rect 572 15412 640 15468
rect 696 15412 706 15468
rect 506 15344 706 15412
rect 506 15288 516 15344
rect 572 15288 640 15344
rect 696 15288 706 15344
rect 506 15220 706 15288
rect 506 15164 516 15220
rect 572 15164 640 15220
rect 696 15164 706 15220
rect 506 15096 706 15164
rect 506 15040 516 15096
rect 572 15040 640 15096
rect 696 15040 706 15096
rect 506 14972 706 15040
rect 506 14916 516 14972
rect 572 14916 640 14972
rect 696 14916 706 14972
rect 506 14848 706 14916
rect 506 14792 516 14848
rect 572 14792 640 14848
rect 696 14792 706 14848
rect 506 14724 706 14792
rect 506 14668 516 14724
rect 572 14668 640 14724
rect 696 14668 706 14724
rect 506 14600 706 14668
rect 506 14544 516 14600
rect 572 14544 640 14600
rect 696 14544 706 14600
rect 506 14476 706 14544
rect 506 14420 516 14476
rect 572 14420 640 14476
rect 696 14420 706 14476
rect 506 14352 706 14420
rect 506 14296 516 14352
rect 572 14296 640 14352
rect 696 14296 706 14352
rect 506 14228 706 14296
rect 506 14172 516 14228
rect 572 14172 640 14228
rect 696 14172 706 14228
rect 506 14104 706 14172
rect 506 14048 516 14104
rect 572 14048 640 14104
rect 696 14048 706 14104
rect 506 14038 706 14048
rect 6 13292 206 13302
rect 6 13236 16 13292
rect 72 13236 140 13292
rect 196 13236 206 13292
rect 6 13168 206 13236
rect 6 13112 16 13168
rect 72 13112 140 13168
rect 196 13112 206 13168
rect 6 13044 206 13112
rect 6 12988 16 13044
rect 72 12988 140 13044
rect 196 12988 206 13044
rect 6 12920 206 12988
rect 6 12864 16 12920
rect 72 12864 140 12920
rect 196 12864 206 12920
rect 6 12796 206 12864
rect 6 12740 16 12796
rect 72 12740 140 12796
rect 196 12740 206 12796
rect 6 12730 206 12740
rect 1023 13292 1223 13302
rect 1023 13236 1033 13292
rect 1089 13236 1157 13292
rect 1213 13236 1223 13292
rect 1023 13168 1223 13236
rect 1023 13112 1033 13168
rect 1089 13112 1157 13168
rect 1213 13112 1223 13168
rect 1023 13044 1223 13112
rect 1023 12988 1033 13044
rect 1089 12988 1157 13044
rect 1213 12988 1223 13044
rect 1023 12920 1223 12988
rect 1023 12864 1033 12920
rect 1089 12864 1157 12920
rect 1213 12864 1223 12920
rect 1023 12796 1223 12864
rect 1023 12740 1033 12796
rect 1089 12740 1157 12796
rect 1213 12740 1223 12796
rect 1023 12730 1223 12740
rect 6 12605 206 12615
rect 6 12549 16 12605
rect 72 12549 140 12605
rect 196 12549 206 12605
rect 6 12481 206 12549
rect 6 12425 16 12481
rect 72 12425 140 12481
rect 196 12425 206 12481
rect 6 12357 206 12425
rect 6 12301 16 12357
rect 72 12301 140 12357
rect 196 12301 206 12357
rect 6 12233 206 12301
rect 6 12177 16 12233
rect 72 12177 140 12233
rect 196 12177 206 12233
rect 6 12109 206 12177
rect 6 12053 16 12109
rect 72 12053 140 12109
rect 196 12053 206 12109
rect 6 12043 206 12053
rect 1023 12605 1223 12615
rect 1023 12549 1033 12605
rect 1089 12549 1157 12605
rect 1213 12549 1223 12605
rect 1023 12481 1223 12549
rect 1023 12425 1033 12481
rect 1089 12425 1157 12481
rect 1213 12425 1223 12481
rect 1023 12357 1223 12425
rect 1023 12301 1033 12357
rect 1089 12301 1157 12357
rect 1213 12301 1223 12357
rect 1023 12233 1223 12301
rect 1023 12177 1033 12233
rect 1089 12177 1157 12233
rect 1213 12177 1223 12233
rect 1023 12109 1223 12177
rect 1023 12053 1033 12109
rect 1089 12053 1157 12109
rect 1213 12053 1223 12109
rect 1023 12043 1223 12053
rect 506 11233 706 11243
rect 506 11177 516 11233
rect 572 11177 640 11233
rect 696 11177 706 11233
rect 506 11109 706 11177
rect 506 11053 516 11109
rect 572 11053 640 11109
rect 696 11053 706 11109
rect 506 10985 706 11053
rect 506 10929 516 10985
rect 572 10929 640 10985
rect 696 10929 706 10985
rect 506 10861 706 10929
rect 506 10805 516 10861
rect 572 10805 640 10861
rect 696 10805 706 10861
rect 506 10737 706 10805
rect 506 10681 516 10737
rect 572 10681 640 10737
rect 696 10681 706 10737
rect 506 10613 706 10681
rect 506 10557 516 10613
rect 572 10557 640 10613
rect 696 10557 706 10613
rect 506 10489 706 10557
rect 506 10433 516 10489
rect 572 10433 640 10489
rect 696 10433 706 10489
rect 506 10365 706 10433
rect 506 10309 516 10365
rect 572 10309 640 10365
rect 696 10309 706 10365
rect 506 10241 706 10309
rect 506 10185 516 10241
rect 572 10185 640 10241
rect 696 10185 706 10241
rect 506 10117 706 10185
rect 506 10061 516 10117
rect 572 10061 640 10117
rect 696 10061 706 10117
rect 506 10051 706 10061
rect 6 9403 206 9413
rect 6 9347 16 9403
rect 72 9347 140 9403
rect 196 9347 206 9403
rect 6 9279 206 9347
rect 6 9223 16 9279
rect 72 9223 140 9279
rect 196 9223 206 9279
rect 6 9155 206 9223
rect 6 9099 16 9155
rect 72 9099 140 9155
rect 196 9099 206 9155
rect 6 9031 206 9099
rect 6 8975 16 9031
rect 72 8975 140 9031
rect 196 8975 206 9031
rect 6 8907 206 8975
rect 6 8851 16 8907
rect 72 8851 140 8907
rect 196 8851 206 8907
rect 6 8841 206 8851
rect 1023 9403 1223 9413
rect 1023 9347 1033 9403
rect 1089 9347 1157 9403
rect 1213 9347 1223 9403
rect 1023 9279 1223 9347
rect 1023 9223 1033 9279
rect 1089 9223 1157 9279
rect 1213 9223 1223 9279
rect 1023 9155 1223 9223
rect 1023 9099 1033 9155
rect 1089 9099 1157 9155
rect 1213 9099 1223 9155
rect 1023 9031 1223 9099
rect 1023 8975 1033 9031
rect 1089 8975 1157 9031
rect 1213 8975 1223 9031
rect 1023 8907 1223 8975
rect 1023 8851 1033 8907
rect 1089 8851 1157 8907
rect 1213 8851 1223 8907
rect 1023 8841 1223 8851
rect 6 7964 206 7974
rect 6 7908 16 7964
rect 72 7908 140 7964
rect 196 7908 206 7964
rect 6 7840 206 7908
rect 6 7784 16 7840
rect 72 7784 140 7840
rect 196 7784 206 7840
rect 6 7716 206 7784
rect 6 7660 16 7716
rect 72 7660 140 7716
rect 196 7660 206 7716
rect 6 7650 206 7660
rect 1023 7964 1223 7974
rect 1023 7908 1033 7964
rect 1089 7908 1157 7964
rect 1213 7908 1223 7964
rect 1023 7840 1223 7908
rect 1023 7784 1033 7840
rect 1089 7784 1157 7840
rect 1213 7784 1223 7840
rect 1023 7716 1223 7784
rect 1023 7660 1033 7716
rect 1089 7660 1157 7716
rect 1213 7660 1223 7716
rect 1023 7650 1223 7660
rect 506 7366 706 7376
rect 506 7310 516 7366
rect 572 7310 640 7366
rect 696 7310 706 7366
rect 506 7242 706 7310
rect 506 7186 516 7242
rect 572 7186 640 7242
rect 696 7186 706 7242
rect 506 7118 706 7186
rect 506 7062 516 7118
rect 572 7062 640 7118
rect 696 7062 706 7118
rect 506 7052 706 7062
rect 506 6403 706 6413
rect 506 6347 516 6403
rect 572 6347 640 6403
rect 696 6347 706 6403
rect 506 6279 706 6347
rect 506 6223 516 6279
rect 572 6223 640 6279
rect 696 6223 706 6279
rect 506 6155 706 6223
rect 506 6099 516 6155
rect 572 6099 640 6155
rect 696 6099 706 6155
rect 506 6089 706 6099
rect 6 5680 206 5690
rect 6 5624 16 5680
rect 72 5624 140 5680
rect 196 5624 206 5680
rect 6 5556 206 5624
rect 6 5500 16 5556
rect 72 5500 140 5556
rect 196 5500 206 5556
rect 6 5432 206 5500
rect 6 5376 16 5432
rect 72 5376 140 5432
rect 196 5376 206 5432
rect 6 5366 206 5376
rect 1023 5680 1223 5690
rect 1023 5624 1033 5680
rect 1089 5624 1157 5680
rect 1213 5624 1223 5680
rect 1023 5556 1223 5624
rect 1023 5500 1033 5556
rect 1089 5500 1157 5556
rect 1213 5500 1223 5556
rect 1023 5432 1223 5500
rect 1023 5376 1033 5432
rect 1089 5376 1157 5432
rect 1213 5376 1223 5432
rect 1023 5366 1223 5376
rect 6 4667 206 4677
rect 6 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 206 4667
rect 6 4543 206 4611
rect 6 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 206 4543
rect 6 4419 206 4487
rect 6 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 206 4419
rect 6 4353 206 4363
rect 1023 4667 1223 4677
rect 1023 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1223 4667
rect 1023 4543 1223 4611
rect 1023 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1223 4543
rect 1023 4419 1223 4487
rect 1023 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1223 4419
rect 1023 4353 1223 4363
rect 506 4037 706 4047
rect 506 3981 516 4037
rect 572 3981 640 4037
rect 696 3981 706 4037
rect 506 3913 706 3981
rect 506 3857 516 3913
rect 572 3857 640 3913
rect 696 3857 706 3913
rect 506 3789 706 3857
rect 506 3733 516 3789
rect 572 3733 640 3789
rect 696 3733 706 3789
rect 506 3665 706 3733
rect 506 3609 516 3665
rect 572 3609 640 3665
rect 696 3609 706 3665
rect 506 3541 706 3609
rect 506 3485 516 3541
rect 572 3485 640 3541
rect 696 3485 706 3541
rect 506 3417 706 3485
rect 506 3361 516 3417
rect 572 3361 640 3417
rect 696 3361 706 3417
rect 506 3293 706 3361
rect 506 3237 516 3293
rect 572 3237 640 3293
rect 696 3237 706 3293
rect 506 3169 706 3237
rect 506 3113 516 3169
rect 572 3113 640 3169
rect 696 3113 706 3169
rect 506 3103 706 3113
use M2_M14310589983294_64x8m81  M2_M14310589983294_64x8m81_0
timestamp 1762296095
transform 1 0 1120 0 1 2599
box 0 0 1 1
use M2_M14310589983294_64x8m81  M2_M14310589983294_64x8m81_1
timestamp 1762296095
transform 1 0 103 0 1 2599
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_0
timestamp 1762296095
transform 1 0 606 0 1 6251
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_1
timestamp 1762296095
transform 1 0 1123 0 1 4515
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_2
timestamp 1762296095
transform 1 0 106 0 1 5528
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_3
timestamp 1762296095
transform 1 0 1123 0 1 5528
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_4
timestamp 1762296095
transform 1 0 606 0 1 7214
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_5
timestamp 1762296095
transform 1 0 1123 0 1 7812
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_6
timestamp 1762296095
transform 1 0 106 0 1 7812
box 0 0 1 1
use M3_M24310589983292_64x8m81  M3_M24310589983292_64x8m81_7
timestamp 1762296095
transform 1 0 106 0 1 4515
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_0
timestamp 1762296095
transform 1 0 106 0 1 9127
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_1
timestamp 1762296095
transform 1 0 106 0 1 13016
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_2
timestamp 1762296095
transform 1 0 1123 0 1 13016
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_3
timestamp 1762296095
transform 1 0 106 0 1 12329
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_4
timestamp 1762296095
transform 1 0 1123 0 1 12329
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_5
timestamp 1762296095
transform 1 0 106 0 1 17993
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_6
timestamp 1762296095
transform 1 0 1123 0 1 17993
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_7
timestamp 1762296095
transform 1 0 106 0 1 17306
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_8
timestamp 1762296095
transform 1 0 1123 0 1 17306
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_9
timestamp 1762296095
transform 1 0 106 0 1 16622
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_10
timestamp 1762296095
transform 1 0 1123 0 1 16622
box 0 0 1 1
use M3_M24310589983295_64x8m81  M3_M24310589983295_64x8m81_11
timestamp 1762296095
transform 1 0 1123 0 1 9127
box 0 0 1 1
use M3_M24310589983296_64x8m81  M3_M24310589983296_64x8m81_0
timestamp 1762296095
transform 1 0 606 0 1 14944
box 0 0 1 1
use M3_M24310589983297_64x8m81  M3_M24310589983297_64x8m81_0
timestamp 1762296095
transform 1 0 606 0 1 10647
box 0 0 1 1
use M3_M24310589983298_64x8m81  M3_M24310589983298_64x8m81_0
timestamp 1762296095
transform 1 0 606 0 1 3575
box 0 0 1 1
<< properties >>
string GDS_END 1438056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1436610
<< end >>
