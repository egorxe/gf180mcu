magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< nwell >>
rect -83 1281 2361 2575
<< mvnmos >>
rect 462 354 602 654
rect 878 354 1018 654
rect 1294 354 1434 654
rect 1710 354 1850 654
<< mvpmos >>
rect 462 1486 602 2086
rect 878 1486 1018 2086
rect 1294 1486 1434 2086
rect 1710 1486 1850 2086
<< mvndiff >>
rect 374 641 462 654
rect 374 595 387 641
rect 433 595 462 641
rect 374 527 462 595
rect 374 481 387 527
rect 433 481 462 527
rect 374 413 462 481
rect 374 367 387 413
rect 433 367 462 413
rect 374 354 462 367
rect 602 641 690 654
rect 602 595 631 641
rect 677 595 690 641
rect 602 527 690 595
rect 602 481 631 527
rect 677 481 690 527
rect 602 413 690 481
rect 602 367 631 413
rect 677 367 690 413
rect 602 354 690 367
rect 790 641 878 654
rect 790 595 803 641
rect 849 595 878 641
rect 790 527 878 595
rect 790 481 803 527
rect 849 481 878 527
rect 790 413 878 481
rect 790 367 803 413
rect 849 367 878 413
rect 790 354 878 367
rect 1018 641 1106 654
rect 1018 595 1047 641
rect 1093 595 1106 641
rect 1018 527 1106 595
rect 1018 481 1047 527
rect 1093 481 1106 527
rect 1018 413 1106 481
rect 1018 367 1047 413
rect 1093 367 1106 413
rect 1018 354 1106 367
rect 1206 641 1294 654
rect 1206 595 1219 641
rect 1265 595 1294 641
rect 1206 527 1294 595
rect 1206 481 1219 527
rect 1265 481 1294 527
rect 1206 413 1294 481
rect 1206 367 1219 413
rect 1265 367 1294 413
rect 1206 354 1294 367
rect 1434 641 1522 654
rect 1434 595 1463 641
rect 1509 595 1522 641
rect 1434 527 1522 595
rect 1434 481 1463 527
rect 1509 481 1522 527
rect 1434 413 1522 481
rect 1434 367 1463 413
rect 1509 367 1522 413
rect 1434 354 1522 367
rect 1622 641 1710 654
rect 1622 595 1635 641
rect 1681 595 1710 641
rect 1622 527 1710 595
rect 1622 481 1635 527
rect 1681 481 1710 527
rect 1622 413 1710 481
rect 1622 367 1635 413
rect 1681 367 1710 413
rect 1622 354 1710 367
rect 1850 641 1938 654
rect 1850 595 1879 641
rect 1925 595 1938 641
rect 1850 527 1938 595
rect 1850 481 1879 527
rect 1925 481 1938 527
rect 1850 413 1938 481
rect 1850 367 1879 413
rect 1925 367 1938 413
rect 1850 354 1938 367
<< mvpdiff >>
rect 374 2073 462 2086
rect 374 2027 387 2073
rect 433 2027 462 2073
rect 374 1968 462 2027
rect 374 1922 387 1968
rect 433 1922 462 1968
rect 374 1863 462 1922
rect 374 1817 387 1863
rect 433 1817 462 1863
rect 374 1757 462 1817
rect 374 1711 387 1757
rect 433 1711 462 1757
rect 374 1651 462 1711
rect 374 1605 387 1651
rect 433 1605 462 1651
rect 374 1545 462 1605
rect 374 1499 387 1545
rect 433 1499 462 1545
rect 374 1486 462 1499
rect 602 2073 690 2086
rect 602 2027 631 2073
rect 677 2027 690 2073
rect 602 1968 690 2027
rect 602 1922 631 1968
rect 677 1922 690 1968
rect 602 1863 690 1922
rect 602 1817 631 1863
rect 677 1817 690 1863
rect 602 1757 690 1817
rect 602 1711 631 1757
rect 677 1711 690 1757
rect 602 1651 690 1711
rect 602 1605 631 1651
rect 677 1605 690 1651
rect 602 1545 690 1605
rect 602 1499 631 1545
rect 677 1499 690 1545
rect 602 1486 690 1499
rect 790 2073 878 2086
rect 790 2027 803 2073
rect 849 2027 878 2073
rect 790 1968 878 2027
rect 790 1922 803 1968
rect 849 1922 878 1968
rect 790 1863 878 1922
rect 790 1817 803 1863
rect 849 1817 878 1863
rect 790 1757 878 1817
rect 790 1711 803 1757
rect 849 1711 878 1757
rect 790 1651 878 1711
rect 790 1605 803 1651
rect 849 1605 878 1651
rect 790 1545 878 1605
rect 790 1499 803 1545
rect 849 1499 878 1545
rect 790 1486 878 1499
rect 1018 2073 1106 2086
rect 1018 2027 1047 2073
rect 1093 2027 1106 2073
rect 1018 1968 1106 2027
rect 1018 1922 1047 1968
rect 1093 1922 1106 1968
rect 1018 1863 1106 1922
rect 1018 1817 1047 1863
rect 1093 1817 1106 1863
rect 1018 1757 1106 1817
rect 1018 1711 1047 1757
rect 1093 1711 1106 1757
rect 1018 1651 1106 1711
rect 1018 1605 1047 1651
rect 1093 1605 1106 1651
rect 1018 1545 1106 1605
rect 1018 1499 1047 1545
rect 1093 1499 1106 1545
rect 1018 1486 1106 1499
rect 1206 2073 1294 2086
rect 1206 2027 1219 2073
rect 1265 2027 1294 2073
rect 1206 1967 1294 2027
rect 1206 1921 1219 1967
rect 1265 1921 1294 1967
rect 1206 1861 1294 1921
rect 1206 1815 1219 1861
rect 1265 1815 1294 1861
rect 1206 1755 1294 1815
rect 1206 1709 1219 1755
rect 1265 1709 1294 1755
rect 1206 1650 1294 1709
rect 1206 1604 1219 1650
rect 1265 1604 1294 1650
rect 1206 1545 1294 1604
rect 1206 1499 1219 1545
rect 1265 1499 1294 1545
rect 1206 1486 1294 1499
rect 1434 2073 1522 2086
rect 1434 2027 1463 2073
rect 1509 2027 1522 2073
rect 1434 1967 1522 2027
rect 1434 1921 1463 1967
rect 1509 1921 1522 1967
rect 1434 1861 1522 1921
rect 1434 1815 1463 1861
rect 1509 1815 1522 1861
rect 1434 1755 1522 1815
rect 1434 1709 1463 1755
rect 1509 1709 1522 1755
rect 1434 1650 1522 1709
rect 1434 1604 1463 1650
rect 1509 1604 1522 1650
rect 1434 1545 1522 1604
rect 1434 1499 1463 1545
rect 1509 1499 1522 1545
rect 1434 1486 1522 1499
rect 1622 2073 1710 2086
rect 1622 2027 1635 2073
rect 1681 2027 1710 2073
rect 1622 1967 1710 2027
rect 1622 1921 1635 1967
rect 1681 1921 1710 1967
rect 1622 1861 1710 1921
rect 1622 1815 1635 1861
rect 1681 1815 1710 1861
rect 1622 1755 1710 1815
rect 1622 1709 1635 1755
rect 1681 1709 1710 1755
rect 1622 1650 1710 1709
rect 1622 1604 1635 1650
rect 1681 1604 1710 1650
rect 1622 1545 1710 1604
rect 1622 1499 1635 1545
rect 1681 1499 1710 1545
rect 1622 1486 1710 1499
rect 1850 2073 1938 2086
rect 1850 2027 1879 2073
rect 1925 2027 1938 2073
rect 1850 1967 1938 2027
rect 1850 1921 1879 1967
rect 1925 1921 1938 1967
rect 1850 1861 1938 1921
rect 1850 1815 1879 1861
rect 1925 1815 1938 1861
rect 1850 1755 1938 1815
rect 1850 1709 1879 1755
rect 1925 1709 1938 1755
rect 1850 1650 1938 1709
rect 1850 1604 1879 1650
rect 1925 1604 1938 1650
rect 1850 1545 1938 1604
rect 1850 1499 1879 1545
rect 1925 1499 1938 1545
rect 1850 1486 1938 1499
<< mvndiffc >>
rect 387 595 433 641
rect 387 481 433 527
rect 387 367 433 413
rect 631 595 677 641
rect 631 481 677 527
rect 631 367 677 413
rect 803 595 849 641
rect 803 481 849 527
rect 803 367 849 413
rect 1047 595 1093 641
rect 1047 481 1093 527
rect 1047 367 1093 413
rect 1219 595 1265 641
rect 1219 481 1265 527
rect 1219 367 1265 413
rect 1463 595 1509 641
rect 1463 481 1509 527
rect 1463 367 1509 413
rect 1635 595 1681 641
rect 1635 481 1681 527
rect 1635 367 1681 413
rect 1879 595 1925 641
rect 1879 481 1925 527
rect 1879 367 1925 413
<< mvpdiffc >>
rect 387 2027 433 2073
rect 387 1922 433 1968
rect 387 1817 433 1863
rect 387 1711 433 1757
rect 387 1605 433 1651
rect 387 1499 433 1545
rect 631 2027 677 2073
rect 631 1922 677 1968
rect 631 1817 677 1863
rect 631 1711 677 1757
rect 631 1605 677 1651
rect 631 1499 677 1545
rect 803 2027 849 2073
rect 803 1922 849 1968
rect 803 1817 849 1863
rect 803 1711 849 1757
rect 803 1605 849 1651
rect 803 1499 849 1545
rect 1047 2027 1093 2073
rect 1047 1922 1093 1968
rect 1047 1817 1093 1863
rect 1047 1711 1093 1757
rect 1047 1605 1093 1651
rect 1047 1499 1093 1545
rect 1219 2027 1265 2073
rect 1219 1921 1265 1967
rect 1219 1815 1265 1861
rect 1219 1709 1265 1755
rect 1219 1604 1265 1650
rect 1219 1499 1265 1545
rect 1463 2027 1509 2073
rect 1463 1921 1509 1967
rect 1463 1815 1509 1861
rect 1463 1709 1509 1755
rect 1463 1604 1509 1650
rect 1463 1499 1509 1545
rect 1635 2027 1681 2073
rect 1635 1921 1681 1967
rect 1635 1815 1681 1861
rect 1635 1709 1681 1755
rect 1635 1604 1681 1650
rect 1635 1499 1681 1545
rect 1879 2027 1925 2073
rect 1879 1921 1925 1967
rect 1879 1815 1925 1861
rect 1879 1709 1925 1755
rect 1879 1604 1925 1650
rect 1879 1499 1925 1545
<< psubdiff >>
rect 0 1008 90 1030
rect 0 22 22 1008
rect 68 90 90 1008
rect 2188 1008 2278 1030
rect 2188 90 2210 1008
rect 68 68 2210 90
rect 68 22 176 68
rect 2102 22 2210 68
rect 2256 22 2278 1008
rect 0 0 2278 22
<< nsubdiff >>
rect 0 2470 2278 2492
rect 0 1484 22 2470
rect 68 2424 176 2470
rect 2102 2424 2210 2470
rect 68 2402 2210 2424
rect 68 1484 90 2402
rect 0 1462 90 1484
rect 2188 1484 2210 2402
rect 2256 1484 2278 2470
rect 2188 1462 2278 1484
<< psubdiffcont >>
rect 22 22 68 1008
rect 176 22 2102 68
rect 2210 22 2256 1008
<< nsubdiffcont >>
rect 22 1484 68 2470
rect 176 2424 2102 2470
rect 2210 1484 2256 2470
<< polysilicon >>
rect 462 2086 602 2130
rect 878 2086 1018 2130
rect 1294 2086 1434 2130
rect 1710 2086 1850 2130
rect 462 1079 602 1486
rect 878 1301 1018 1486
rect 878 1161 925 1301
rect 971 1161 1018 1301
rect 878 1142 1018 1161
rect 1294 1301 1434 1486
rect 1294 1161 1341 1301
rect 1387 1161 1434 1301
rect 1294 1142 1434 1161
rect 1710 1301 1850 1486
rect 1710 1161 1757 1301
rect 1803 1161 1850 1301
rect 462 939 509 1079
rect 555 939 602 1079
rect 1710 995 1850 1161
rect 462 654 602 939
rect 878 976 1018 995
rect 878 836 925 976
rect 971 836 1018 976
rect 878 654 1018 836
rect 1294 817 1850 995
rect 1294 654 1434 817
rect 1710 654 1850 817
rect 462 310 602 354
rect 878 310 1018 354
rect 1294 310 1434 354
rect 1710 310 1850 354
<< polycontact >>
rect 925 1161 971 1301
rect 1341 1161 1387 1301
rect 1757 1161 1803 1301
rect 509 939 555 1079
rect 925 836 971 976
<< metal1 >>
rect 11 2470 2267 2481
rect 11 1484 22 2470
rect 68 2424 176 2470
rect 2102 2424 2210 2470
rect 68 2413 2210 2424
rect 68 1484 79 2413
rect 372 2073 448 2413
rect 372 2027 387 2073
rect 433 2027 448 2073
rect 372 1968 448 2027
rect 372 1922 387 1968
rect 433 1922 448 1968
rect 372 1863 448 1922
rect 372 1817 387 1863
rect 433 1817 448 1863
rect 372 1757 448 1817
rect 372 1711 387 1757
rect 433 1711 448 1757
rect 372 1651 448 1711
rect 372 1605 387 1651
rect 433 1605 448 1651
rect 372 1545 448 1605
rect 372 1499 387 1545
rect 433 1499 448 1545
rect 372 1486 448 1499
rect 616 2186 1524 2262
rect 616 2073 692 2186
rect 616 2027 631 2073
rect 677 2027 692 2073
rect 616 1968 692 2027
rect 616 1922 631 1968
rect 677 1922 692 1968
rect 616 1863 692 1922
rect 616 1817 631 1863
rect 677 1817 692 1863
rect 616 1757 692 1817
rect 616 1711 631 1757
rect 677 1711 692 1757
rect 616 1654 692 1711
rect 616 1498 628 1654
rect 680 1498 692 1654
rect 616 1486 692 1498
rect 788 2073 864 2086
rect 788 2027 803 2073
rect 849 2027 864 2073
rect 788 1968 864 2027
rect 788 1922 803 1968
rect 849 1922 864 1968
rect 788 1863 864 1922
rect 788 1817 803 1863
rect 849 1817 864 1863
rect 788 1757 864 1817
rect 788 1711 803 1757
rect 849 1711 864 1757
rect 788 1651 864 1711
rect 788 1605 803 1651
rect 849 1605 864 1651
rect 788 1545 864 1605
rect 788 1499 803 1545
rect 849 1499 864 1545
rect 11 1473 79 1484
rect 788 1090 864 1499
rect 1032 2073 1280 2086
rect 1032 2027 1047 2073
rect 1093 2027 1219 2073
rect 1265 2027 1280 2073
rect 1032 1968 1280 2027
rect 1032 1922 1047 1968
rect 1093 1967 1280 1968
rect 1093 1922 1219 1967
rect 1032 1921 1219 1922
rect 1265 1921 1280 1967
rect 1032 1863 1280 1921
rect 1032 1817 1047 1863
rect 1093 1861 1280 1863
rect 1093 1817 1219 1861
rect 1032 1815 1219 1817
rect 1265 1815 1280 1861
rect 1032 1757 1280 1815
rect 1032 1711 1047 1757
rect 1093 1755 1280 1757
rect 1093 1711 1219 1755
rect 1032 1709 1219 1711
rect 1265 1709 1280 1755
rect 1032 1654 1280 1709
rect 1032 1498 1044 1654
rect 1096 1650 1280 1654
rect 1096 1604 1219 1650
rect 1265 1604 1280 1650
rect 1096 1545 1280 1604
rect 1096 1499 1219 1545
rect 1265 1499 1280 1545
rect 1096 1498 1280 1499
rect 1032 1486 1280 1498
rect 1448 2073 1524 2186
rect 1448 2027 1463 2073
rect 1509 2027 1524 2073
rect 1448 1967 1524 2027
rect 1448 1921 1463 1967
rect 1509 1921 1524 1967
rect 1448 1861 1524 1921
rect 1448 1815 1463 1861
rect 1509 1815 1524 1861
rect 1448 1755 1524 1815
rect 1448 1709 1463 1755
rect 1509 1709 1524 1755
rect 1448 1650 1524 1709
rect 1448 1604 1463 1650
rect 1509 1604 1524 1650
rect 1448 1545 1524 1604
rect 1448 1499 1463 1545
rect 1509 1499 1524 1545
rect 1448 1486 1524 1499
rect 1620 2073 1696 2086
rect 1620 2027 1635 2073
rect 1681 2027 1696 2073
rect 1620 1967 1696 2027
rect 1620 1921 1635 1967
rect 1681 1921 1696 1967
rect 1620 1861 1696 1921
rect 1620 1815 1635 1861
rect 1681 1815 1696 1861
rect 1620 1755 1696 1815
rect 1620 1709 1635 1755
rect 1681 1709 1696 1755
rect 1620 1650 1696 1709
rect 1620 1604 1635 1650
rect 1681 1604 1696 1650
rect 1620 1545 1696 1604
rect 1620 1499 1635 1545
rect 1681 1499 1696 1545
rect 914 1309 990 1321
rect 914 1301 926 1309
rect 914 1161 925 1301
rect 914 1153 926 1161
rect 978 1153 990 1309
rect 914 1141 990 1153
rect 1326 1301 1402 1312
rect 1326 1161 1341 1301
rect 1387 1161 1402 1301
rect 498 1079 864 1090
rect 11 1008 79 1019
rect 11 22 22 1008
rect 68 79 79 1008
rect 498 939 509 1079
rect 555 939 864 1079
rect 1326 987 1402 1161
rect 1620 987 1696 1499
rect 1864 2073 1940 2413
rect 1864 2027 1879 2073
rect 1925 2027 1940 2073
rect 1864 1967 1940 2027
rect 1864 1921 1879 1967
rect 1925 1921 1940 1967
rect 1864 1861 1940 1921
rect 1864 1815 1879 1861
rect 1925 1815 1940 1861
rect 1864 1755 1940 1815
rect 1864 1709 1879 1755
rect 1925 1709 1940 1755
rect 1864 1650 1940 1709
rect 1864 1604 1879 1650
rect 1925 1604 1940 1650
rect 1864 1545 1940 1604
rect 1864 1499 1879 1545
rect 1925 1499 1940 1545
rect 1864 1486 1940 1499
rect 2199 1484 2210 2413
rect 2256 1484 2267 2470
rect 2199 1473 2267 1484
rect 1746 1309 1822 1321
rect 1746 1301 1758 1309
rect 1746 1161 1757 1301
rect 1746 1153 1758 1161
rect 1810 1153 1822 1309
rect 1746 1141 1822 1153
rect 498 928 864 939
rect 372 641 448 654
rect 372 595 387 641
rect 433 595 448 641
rect 372 527 448 595
rect 372 481 387 527
rect 433 481 448 527
rect 372 413 448 481
rect 372 367 387 413
rect 433 367 448 413
rect 372 79 448 367
rect 616 642 692 654
rect 616 486 628 642
rect 680 486 692 642
rect 616 481 631 486
rect 677 481 692 486
rect 616 413 692 481
rect 616 367 631 413
rect 677 367 692 413
rect 616 254 692 367
rect 788 641 864 928
rect 914 976 1696 987
rect 914 836 925 976
rect 971 836 1696 976
rect 914 825 1696 836
rect 788 595 803 641
rect 849 595 864 641
rect 788 527 864 595
rect 788 481 803 527
rect 849 481 864 527
rect 788 413 864 481
rect 788 367 803 413
rect 849 367 864 413
rect 788 354 864 367
rect 1032 642 1280 654
rect 1032 486 1044 642
rect 1096 641 1280 642
rect 1096 595 1219 641
rect 1265 595 1280 641
rect 1096 527 1280 595
rect 1096 486 1219 527
rect 1032 481 1047 486
rect 1093 481 1219 486
rect 1265 481 1280 527
rect 1032 413 1280 481
rect 1032 367 1047 413
rect 1093 367 1219 413
rect 1265 367 1280 413
rect 1032 354 1280 367
rect 1448 641 1524 654
rect 1448 595 1463 641
rect 1509 595 1524 641
rect 1448 527 1524 595
rect 1448 481 1463 527
rect 1509 481 1524 527
rect 1448 413 1524 481
rect 1448 367 1463 413
rect 1509 367 1524 413
rect 1448 254 1524 367
rect 1620 641 1696 825
rect 2199 1008 2267 1019
rect 1620 595 1635 641
rect 1681 595 1696 641
rect 1620 527 1696 595
rect 1620 481 1635 527
rect 1681 481 1696 527
rect 1620 413 1696 481
rect 1620 367 1635 413
rect 1681 367 1696 413
rect 1620 354 1696 367
rect 1864 641 1940 654
rect 1864 595 1879 641
rect 1925 595 1940 641
rect 1864 527 1940 595
rect 1864 481 1879 527
rect 1925 481 1940 527
rect 1864 413 1940 481
rect 1864 367 1879 413
rect 1925 367 1940 413
rect 616 178 1524 254
rect 1864 79 1940 367
rect 2199 79 2210 1008
rect 68 68 2210 79
rect 68 22 176 68
rect 2102 22 2210 68
rect 2256 22 2267 1008
rect 11 11 2267 22
<< via1 >>
rect 628 1651 680 1654
rect 628 1605 631 1651
rect 631 1605 677 1651
rect 677 1605 680 1651
rect 628 1545 680 1605
rect 628 1499 631 1545
rect 631 1499 677 1545
rect 677 1499 680 1545
rect 628 1498 680 1499
rect 1044 1651 1096 1654
rect 1044 1605 1047 1651
rect 1047 1605 1093 1651
rect 1093 1605 1096 1651
rect 1044 1545 1096 1605
rect 1044 1499 1047 1545
rect 1047 1499 1093 1545
rect 1093 1499 1096 1545
rect 1044 1498 1096 1499
rect 926 1301 978 1309
rect 926 1161 971 1301
rect 971 1161 978 1301
rect 926 1153 978 1161
rect 1758 1301 1810 1309
rect 1758 1161 1803 1301
rect 1803 1161 1810 1301
rect 1758 1153 1810 1161
rect 628 641 680 642
rect 628 595 631 641
rect 631 595 677 641
rect 677 595 680 641
rect 628 527 680 595
rect 628 486 631 527
rect 631 486 677 527
rect 677 486 680 527
rect 1044 641 1096 642
rect 1044 595 1047 641
rect 1047 595 1093 641
rect 1093 595 1096 641
rect 1044 527 1096 595
rect 1044 486 1047 527
rect 1047 486 1093 527
rect 1093 486 1096 527
<< metal2 >>
rect 616 1654 692 1666
rect 616 1498 628 1654
rect 680 1498 692 1654
rect 616 642 692 1498
rect 616 486 628 642
rect 680 486 692 642
rect 616 474 692 486
rect 752 1654 1108 1666
rect 752 1498 1044 1654
rect 1096 1498 1108 1654
rect 752 1486 1108 1498
rect 752 654 828 1486
rect 914 1309 1822 1321
rect 914 1153 926 1309
rect 978 1153 1758 1309
rect 1810 1153 1822 1309
rect 914 1141 1822 1153
rect 752 642 1108 654
rect 752 486 1044 642
rect 1096 486 1108 642
rect 752 474 1108 486
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_0
timestamp 1759194789
transform 1 0 45 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661953145315  M1_NWELL_CDNS_40661953145315_1
timestamp 1759194789
transform 1 0 2233 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661953145323  M1_NWELL_CDNS_40661953145323_0
timestamp 1759194789
transform 1 0 1139 0 1 2447
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_0
timestamp 1759194789
transform 1 0 948 0 1 906
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_1
timestamp 1759194789
transform 1 0 1364 0 1 1231
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_2
timestamp 1759194789
transform 1 0 948 0 1 1231
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_3
timestamp 1759194789
transform 1 0 1780 0 1 1231
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_4
timestamp 1759194789
transform 1 0 532 0 1 1009
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_0
timestamp 1759194789
transform 1 0 45 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_1
timestamp 1759194789
transform 1 0 2233 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145324  M1_PSUB_CDNS_40661953145324_0
timestamp 1759194789
transform 1 0 1139 0 -1 45
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1759194789
transform 1 0 654 0 1 1576
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1759194789
transform 1 0 654 0 1 564
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1759194789
transform 1 0 1070 0 1 564
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_3
timestamp 1759194789
transform 1 0 1070 0 1 1576
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_4
timestamp 1759194789
transform 1 0 952 0 1 1231
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_5
timestamp 1759194789
transform 1 0 1784 0 1 1231
box 0 0 1 1
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1759194789
transform -1 0 1850 0 -1 654
box 0 0 1 1
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_1
timestamp 1759194789
transform -1 0 1018 0 -1 654
box 0 0 1 1
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_2
timestamp 1759194789
transform 1 0 1294 0 1 354
box 0 0 1 1
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_3
timestamp 1759194789
transform 1 0 462 0 1 354
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1759194789
transform -1 0 1018 0 1 1486
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1759194789
transform 1 0 1294 0 -1 2086
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_2
timestamp 1759194789
transform -1 0 1850 0 -1 2086
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_3
timestamp 1759194789
transform 1 0 462 0 1 1486
box 0 0 1 1
<< labels >>
rlabel metal2 s 1507 1222 1507 1222 4 B
port 1 nsew
rlabel metal2 s 783 1222 783 1222 4 Z
port 2 nsew
rlabel metal1 s 270 2452 270 2452 4 VDD
port 3 nsew
rlabel metal1 s 244 45 244 45 4 VSS
port 4 nsew
rlabel metal1 s 533 1012 533 1012 4 A
port 5 nsew
rlabel metal1 s 1781 1234 1781 1234 4 B
port 1 nsew
<< properties >>
string GDS_END 1531538
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1527460
string path 31.050 37.150 31.050 52.150 
<< end >>
