VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__cor
  CLASS ENDCAP BOTTOMLEFT ;
  FOREIGN gf180mcu_fd_io__cor ;
  ORIGIN 0.000 0.000 ;
  SIZE 355.000 BY 355.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_COR_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 334.000 354.000 341.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 294.000 354.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 278.000 354.000 285.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 270.000 354.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 262.000 354.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 214.000 354.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 352.060 214.000 352.440 228.995 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 206.000 354.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 182.000 354.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 166.000 354.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 150.000 354.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 134.000 354.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 118.000 354.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 334.000 354.000 341.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 294.000 354.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 278.000 354.000 285.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 270.000 354.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.000 354.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.000 354.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 281.310 317.160 281.690 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.000 354.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 182.000 354.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 166.000 354.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.000 354.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 134.000 354.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.000 354.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 334.000 354.000 341.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 334.000 355.000 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 294.000 354.000 301.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 294.000 355.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 278.000 355.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 270.000 354.000 277.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 270.000 355.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 262.000 354.000 269.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 262.000 355.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 214.000 354.000 229.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 273.310 313.845 273.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 206.000 354.000 213.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 206.000 355.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 182.000 354.000 197.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 182.000 355.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 166.000 354.000 181.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 166.000 355.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 150.000 354.000 165.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 150.000 355.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 134.000 354.000 149.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 134.000 355.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 118.000 354.000 125.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 118.000 355.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.040 350.980 172.320 351.260 ;
      LAYER Metal5 ;
        RECT 172.040 350.980 172.320 351.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 118.000 350.800 125.000 351.180 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 140.320 263.145 140.700 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 156.320 269.835 156.700 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 188.320 283.200 188.700 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.970 182.000 352.350 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.035 206.000 352.415 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 293.405 157.640 354.000 158.020 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.920 166.000 352.300 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.120 118.000 352.500 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 293.405 141.640 354.000 142.020 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 297.360 351.005 297.640 351.285 ;
      LAYER Metal4 ;
        RECT 297.360 351.005 297.640 351.285 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 281.360 350.980 281.640 351.260 ;
      LAYER Metal4 ;
        RECT 281.360 350.980 281.640 351.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.000 350.910 269.000 351.290 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 214.000 350.740 229.000 351.120 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 140.320 263.145 140.700 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 118.000 350.800 125.000 351.180 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.010 334.000 352.390 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.945 294.000 352.325 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.910 270.000 352.290 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.060 214.000 352.440 228.995 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.970 182.000 352.350 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 293.405 157.640 354.000 158.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.120 118.000 352.500 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 337.360 351.070 337.640 351.350 ;
      LAYER Metal4 ;
        RECT 337.360 351.070 337.640 351.350 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 273.360 350.970 273.640 351.250 ;
      LAYER Metal4 ;
        RECT 273.360 350.970 273.640 351.250 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 209.360 351.095 209.640 351.375 ;
      LAYER Metal4 ;
        RECT 209.360 351.095 209.640 351.375 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 188.320 283.200 188.700 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.320 269.835 156.700 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.920 278.000 352.300 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.950 265.690 352.230 265.970 ;
      LAYER Metal5 ;
        RECT 351.950 265.690 352.230 265.970 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.035 206.000 352.415 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.920 166.000 352.300 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 293.405 141.640 354.000 142.020 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 342.000 354.000 348.390 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 326.000 354.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 302.000 354.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 286.000 354.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 230.000 354.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 198.000 354.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 126.000 354.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 102.000 354.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 86.000 354.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 354.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 342.000 354.000 348.390 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 326.000 354.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.000 354.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 286.000 354.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 230.000 354.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 198.000 354.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126.000 354.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.000 354.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 86.000 354.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 70.000 354.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 342.000 354.000 348.390 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 342.000 355.000 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 326.000 354.000 333.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 326.000 355.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 302.000 354.000 309.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 302.000 355.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 286.000 354.000 293.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 286.000 355.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 230.000 354.000 245.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 230.000 355.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 198.000 354.000 205.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 198.000 355.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 126.000 354.000 133.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 126.000 355.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 102.000 354.000 117.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 102.000 355.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 86.000 354.000 101.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 86.000 355.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 70.000 354.000 85.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 70.000 355.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 126.000 350.820 133.000 351.200 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 76.980 236.435 77.360 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 92.980 243.115 93.360 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 102.000 350.755 117.000 351.135 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 292.025 94.300 354.000 94.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.020 70.000 352.400 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.075 102.000 352.455 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 256.465 129.970 354.000 130.350 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 352.005 198.000 352.385 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 345.005 346.290 345.385 354.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 329.370 351.050 329.650 351.330 ;
      LAYER Metal4 ;
        RECT 329.370 351.050 329.650 351.330 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 201.360 351.065 201.640 351.345 ;
      LAYER Metal4 ;
        RECT 201.360 351.065 201.640 351.345 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 92.980 243.115 93.360 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.975 342.000 352.355 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.955 302.000 352.335 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 303.085 237.640 354.000 238.020 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.140 126.000 352.520 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.020 70.000 352.400 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 305.360 351.020 305.640 351.300 ;
      LAYER Metal4 ;
        RECT 305.360 351.020 305.640 351.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 289.640 323.375 289.690 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 230.000 350.855 245.000 351.235 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 126.000 350.820 133.000 351.200 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.000 350.755 117.000 351.135 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 76.980 236.435 77.360 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.000 326.000 352.380 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.930 286.000 352.310 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.005 198.000 352.385 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.075 104.845 352.455 113.755 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 292.025 94.300 354.000 94.680 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 310.000 354.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 254.000 354.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 310.000 354.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 254.000 354.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 310.000 354.000 317.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 310.000 355.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 254.000 354.000 261.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 254.000 355.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 254.000 355.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 254.000 355.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.585 257.030 352.865 257.310 ;
      LAYER Metal5 ;
        RECT 352.585 257.030 352.865 257.310 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 351.965 310.000 352.345 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 257.310 307.175 257.690 354.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 313.310 330.450 313.690 354.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 313.360 351.025 313.640 351.305 ;
      LAYER Metal4 ;
        RECT 313.360 351.025 313.640 351.305 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 254.000 350.885 261.000 351.265 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.965 310.000 352.345 317.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 318.000 354.000 325.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 318.000 355.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 246.000 354.000 253.000 355.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 354.000 246.000 355.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.580 249.690 352.860 249.970 ;
      LAYER Metal5 ;
        RECT 352.580 249.690 352.860 249.970 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 246.000 350.880 253.000 351.260 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 321.310 333.810 321.690 354.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.000 350.880 253.000 351.260 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 321.635 351.095 321.645 351.105 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 351.995 318.000 352.375 325.000 ;
    END
  END VSS
  OBS
      LAYER Nwell ;
        RECT 67.560 67.500 350.445 352.170 ;
      LAYER Metal1 ;
        RECT 65.540 65.540 355.000 355.000 ;
      LAYER Metal2 ;
        RECT 68.030 67.970 354.505 354.450 ;
      LAYER Metal3 ;
        RECT 85.300 353.700 85.700 354.450 ;
        RECT 101.300 353.700 101.700 354.450 ;
        RECT 117.300 353.700 117.700 354.450 ;
        RECT 125.300 353.700 125.700 354.450 ;
        RECT 133.300 353.700 133.700 354.450 ;
        RECT 149.300 353.700 149.700 354.450 ;
        RECT 165.300 353.700 165.700 354.450 ;
        RECT 181.300 353.700 181.700 354.450 ;
        RECT 197.300 353.700 197.700 354.450 ;
        RECT 205.300 353.700 205.700 354.450 ;
        RECT 213.300 353.700 213.700 354.450 ;
        RECT 229.300 353.700 229.700 354.450 ;
        RECT 245.300 353.700 245.700 354.450 ;
        RECT 253.300 353.700 253.700 354.450 ;
        RECT 261.300 353.700 261.700 354.450 ;
        RECT 269.300 353.700 269.700 354.450 ;
        RECT 277.300 353.700 277.700 354.450 ;
        RECT 285.300 353.700 285.700 354.450 ;
        RECT 293.300 353.700 293.700 354.450 ;
        RECT 301.300 353.700 301.700 354.450 ;
        RECT 309.300 353.700 309.700 354.450 ;
        RECT 317.300 353.700 317.700 354.450 ;
        RECT 325.300 353.700 325.700 354.450 ;
        RECT 333.300 353.700 333.700 354.450 ;
        RECT 341.300 353.700 341.700 354.450 ;
        RECT 348.690 353.700 355.000 354.450 ;
        RECT 70.000 348.690 355.000 353.700 ;
        RECT 70.000 341.700 353.700 348.690 ;
        RECT 70.000 341.300 355.000 341.700 ;
        RECT 70.000 333.700 353.700 341.300 ;
        RECT 70.000 333.300 355.000 333.700 ;
        RECT 70.000 325.700 353.700 333.300 ;
        RECT 70.000 325.300 355.000 325.700 ;
        RECT 70.000 317.700 353.700 325.300 ;
        RECT 70.000 317.300 355.000 317.700 ;
        RECT 70.000 309.700 353.700 317.300 ;
        RECT 70.000 309.300 355.000 309.700 ;
        RECT 70.000 301.700 353.700 309.300 ;
        RECT 70.000 301.300 355.000 301.700 ;
        RECT 70.000 293.700 353.700 301.300 ;
        RECT 70.000 293.300 355.000 293.700 ;
        RECT 70.000 285.700 353.700 293.300 ;
        RECT 70.000 285.300 355.000 285.700 ;
        RECT 70.000 277.700 353.700 285.300 ;
        RECT 70.000 277.300 355.000 277.700 ;
        RECT 70.000 269.700 353.700 277.300 ;
        RECT 70.000 269.300 355.000 269.700 ;
        RECT 70.000 261.700 353.700 269.300 ;
        RECT 70.000 261.300 355.000 261.700 ;
        RECT 70.000 253.700 353.700 261.300 ;
        RECT 70.000 253.300 355.000 253.700 ;
        RECT 70.000 245.700 353.700 253.300 ;
        RECT 70.000 245.300 355.000 245.700 ;
        RECT 70.000 229.700 353.700 245.300 ;
        RECT 70.000 229.295 355.000 229.700 ;
        RECT 70.000 213.700 351.760 229.295 ;
        RECT 352.740 213.700 355.000 229.295 ;
        RECT 70.000 213.300 355.000 213.700 ;
        RECT 70.000 205.700 353.700 213.300 ;
        RECT 70.000 205.300 355.000 205.700 ;
        RECT 70.000 197.700 353.700 205.300 ;
        RECT 70.000 197.300 355.000 197.700 ;
        RECT 70.000 181.700 353.700 197.300 ;
        RECT 70.000 181.300 355.000 181.700 ;
        RECT 70.000 165.700 353.700 181.300 ;
        RECT 70.000 165.300 355.000 165.700 ;
        RECT 70.000 149.700 353.700 165.300 ;
        RECT 70.000 149.300 355.000 149.700 ;
        RECT 70.000 133.700 353.700 149.300 ;
        RECT 70.000 133.300 355.000 133.700 ;
        RECT 70.000 125.700 353.700 133.300 ;
        RECT 70.000 125.300 355.000 125.700 ;
        RECT 70.000 117.700 353.700 125.300 ;
        RECT 70.000 117.300 355.000 117.700 ;
        RECT 70.000 101.700 353.700 117.300 ;
        RECT 70.000 101.300 355.000 101.700 ;
        RECT 70.000 85.700 353.700 101.300 ;
        RECT 70.000 85.300 355.000 85.700 ;
        RECT 70.000 70.000 353.700 85.300 ;
      LAYER Metal4 ;
        RECT 85.300 353.700 85.700 354.000 ;
        RECT 101.300 353.700 101.700 354.000 ;
        RECT 117.300 353.700 117.700 354.000 ;
        RECT 125.300 353.700 125.700 354.000 ;
        RECT 133.300 353.700 133.700 354.000 ;
        RECT 149.300 353.700 149.700 354.000 ;
        RECT 165.300 353.700 165.700 354.000 ;
        RECT 181.300 353.700 181.700 354.000 ;
        RECT 197.300 353.700 197.700 354.000 ;
        RECT 205.300 353.700 205.700 354.000 ;
        RECT 213.300 353.700 213.700 354.000 ;
        RECT 229.300 353.700 229.700 354.000 ;
        RECT 245.300 353.700 245.700 354.000 ;
        RECT 253.300 353.700 253.700 354.000 ;
        RECT 261.300 353.700 261.700 354.000 ;
        RECT 269.300 353.700 269.700 354.000 ;
        RECT 277.300 353.700 277.700 354.000 ;
        RECT 285.300 353.700 285.700 354.000 ;
        RECT 293.300 353.700 293.700 354.000 ;
        RECT 301.300 353.700 301.700 354.000 ;
        RECT 309.300 353.700 309.700 354.000 ;
        RECT 317.300 353.700 317.700 354.000 ;
        RECT 325.300 353.700 325.700 354.000 ;
        RECT 333.300 353.700 333.700 354.000 ;
        RECT 341.300 353.700 341.700 354.000 ;
        RECT 348.690 353.700 355.000 354.000 ;
        RECT 70.000 236.135 76.680 353.700 ;
        RECT 77.660 242.815 92.680 353.700 ;
        RECT 93.660 351.500 140.020 353.700 ;
        RECT 93.660 351.480 125.700 351.500 ;
        RECT 93.660 351.435 117.700 351.480 ;
        RECT 93.660 350.455 101.700 351.435 ;
        RECT 117.300 350.500 117.700 351.435 ;
        RECT 125.300 350.520 125.700 351.480 ;
        RECT 133.300 350.520 140.020 351.500 ;
        RECT 125.300 350.500 140.020 350.520 ;
        RECT 117.300 350.455 140.020 350.500 ;
        RECT 93.660 262.845 140.020 350.455 ;
        RECT 141.000 269.535 156.020 353.700 ;
        RECT 157.000 282.900 188.020 353.700 ;
        RECT 189.000 351.675 289.340 353.700 ;
        RECT 189.000 351.645 209.060 351.675 ;
        RECT 189.000 350.765 201.060 351.645 ;
        RECT 201.940 350.795 209.060 351.645 ;
        RECT 209.940 351.590 289.340 351.675 ;
        RECT 209.940 351.565 261.700 351.590 ;
        RECT 209.940 351.560 253.700 351.565 ;
        RECT 209.940 351.535 245.700 351.560 ;
        RECT 209.940 351.420 229.700 351.535 ;
        RECT 209.940 350.795 213.700 351.420 ;
        RECT 201.940 350.765 213.700 350.795 ;
        RECT 189.000 350.440 213.700 350.765 ;
        RECT 229.300 350.555 229.700 351.420 ;
        RECT 245.300 350.580 245.700 351.535 ;
        RECT 253.300 350.585 253.700 351.560 ;
        RECT 261.300 350.610 261.700 351.565 ;
        RECT 269.300 351.560 289.340 351.590 ;
        RECT 269.300 351.550 281.060 351.560 ;
        RECT 269.300 350.670 273.060 351.550 ;
        RECT 273.940 350.680 281.060 351.550 ;
        RECT 281.940 350.680 289.340 351.560 ;
        RECT 273.940 350.670 289.340 350.680 ;
        RECT 269.300 350.610 289.340 350.670 ;
        RECT 261.300 350.585 289.340 350.610 ;
        RECT 253.300 350.580 289.340 350.585 ;
        RECT 245.300 350.555 289.340 350.580 ;
        RECT 229.300 350.440 289.340 350.555 ;
        RECT 189.000 323.075 289.340 350.440 ;
        RECT 289.990 351.650 344.705 353.700 ;
        RECT 289.990 351.630 337.060 351.650 ;
        RECT 289.990 351.605 329.070 351.630 ;
        RECT 289.990 351.600 313.060 351.605 ;
        RECT 289.990 351.585 305.060 351.600 ;
        RECT 289.990 350.705 297.060 351.585 ;
        RECT 297.940 350.720 305.060 351.585 ;
        RECT 305.940 350.725 313.060 351.600 ;
        RECT 313.940 351.405 329.070 351.605 ;
        RECT 313.940 350.795 321.335 351.405 ;
        RECT 321.945 350.795 329.070 351.405 ;
        RECT 313.940 350.750 329.070 350.795 ;
        RECT 329.950 350.770 337.060 351.630 ;
        RECT 337.940 350.770 344.705 351.650 ;
        RECT 329.950 350.750 344.705 350.770 ;
        RECT 313.940 350.725 344.705 350.750 ;
        RECT 305.940 350.720 344.705 350.725 ;
        RECT 297.940 350.705 344.705 350.720 ;
        RECT 289.990 345.990 344.705 350.705 ;
        RECT 345.685 348.690 355.000 353.700 ;
        RECT 345.685 345.990 351.675 348.690 ;
        RECT 289.990 341.700 351.675 345.990 ;
        RECT 352.655 341.700 353.700 348.690 ;
        RECT 289.990 341.300 355.000 341.700 ;
        RECT 289.990 333.700 351.710 341.300 ;
        RECT 352.690 333.700 353.700 341.300 ;
        RECT 289.990 333.300 355.000 333.700 ;
        RECT 289.990 325.700 351.700 333.300 ;
        RECT 352.680 325.700 353.700 333.300 ;
        RECT 289.990 325.300 355.000 325.700 ;
        RECT 289.990 323.075 351.695 325.300 ;
        RECT 189.000 317.700 351.695 323.075 ;
        RECT 352.675 317.700 353.700 325.300 ;
        RECT 189.000 317.300 355.000 317.700 ;
        RECT 189.000 309.700 351.665 317.300 ;
        RECT 352.645 309.700 353.700 317.300 ;
        RECT 189.000 309.300 355.000 309.700 ;
        RECT 189.000 301.700 351.655 309.300 ;
        RECT 352.635 301.700 353.700 309.300 ;
        RECT 189.000 301.300 355.000 301.700 ;
        RECT 189.000 293.700 351.645 301.300 ;
        RECT 352.625 293.700 353.700 301.300 ;
        RECT 189.000 293.300 355.000 293.700 ;
        RECT 189.000 285.700 351.630 293.300 ;
        RECT 352.610 285.700 353.700 293.300 ;
        RECT 189.000 285.300 355.000 285.700 ;
        RECT 189.000 282.900 351.620 285.300 ;
        RECT 157.000 277.700 351.620 282.900 ;
        RECT 352.600 277.700 353.700 285.300 ;
        RECT 157.000 277.300 355.000 277.700 ;
        RECT 157.000 269.700 351.610 277.300 ;
        RECT 352.590 269.700 353.700 277.300 ;
        RECT 157.000 269.535 355.000 269.700 ;
        RECT 141.000 269.300 355.000 269.535 ;
        RECT 141.000 266.270 353.700 269.300 ;
        RECT 141.000 265.390 351.650 266.270 ;
        RECT 352.530 265.390 353.700 266.270 ;
        RECT 141.000 262.845 353.700 265.390 ;
        RECT 93.660 261.700 353.700 262.845 ;
        RECT 93.660 261.300 355.000 261.700 ;
        RECT 93.660 253.700 353.700 261.300 ;
        RECT 93.660 253.300 355.000 253.700 ;
        RECT 93.660 245.700 353.700 253.300 ;
        RECT 93.660 245.300 355.000 245.700 ;
        RECT 93.660 242.815 353.700 245.300 ;
        RECT 77.660 238.320 353.700 242.815 ;
        RECT 77.660 237.340 302.785 238.320 ;
        RECT 77.660 236.135 353.700 237.340 ;
        RECT 70.000 229.700 353.700 236.135 ;
        RECT 70.000 229.295 355.000 229.700 ;
        RECT 70.000 213.700 351.760 229.295 ;
        RECT 352.740 213.700 355.000 229.295 ;
        RECT 70.000 213.300 355.000 213.700 ;
        RECT 70.000 205.700 351.735 213.300 ;
        RECT 352.715 205.700 353.700 213.300 ;
        RECT 70.000 205.300 355.000 205.700 ;
        RECT 70.000 197.700 351.705 205.300 ;
        RECT 352.685 197.700 353.700 205.300 ;
        RECT 70.000 197.300 355.000 197.700 ;
        RECT 70.000 181.700 351.670 197.300 ;
        RECT 352.650 181.700 353.700 197.300 ;
        RECT 70.000 181.300 355.000 181.700 ;
        RECT 70.000 165.700 351.620 181.300 ;
        RECT 352.600 165.700 353.700 181.300 ;
        RECT 70.000 165.300 355.000 165.700 ;
        RECT 70.000 158.320 353.700 165.300 ;
        RECT 70.000 157.340 293.105 158.320 ;
        RECT 70.000 149.700 353.700 157.340 ;
        RECT 70.000 149.300 355.000 149.700 ;
        RECT 70.000 142.320 353.700 149.300 ;
        RECT 70.000 141.340 293.105 142.320 ;
        RECT 70.000 133.700 353.700 141.340 ;
        RECT 70.000 133.300 355.000 133.700 ;
        RECT 70.000 125.700 351.840 133.300 ;
        RECT 352.820 125.700 353.700 133.300 ;
        RECT 70.000 125.300 355.000 125.700 ;
        RECT 70.000 117.700 351.820 125.300 ;
        RECT 352.800 117.700 353.700 125.300 ;
        RECT 70.000 117.300 355.000 117.700 ;
        RECT 70.000 114.055 353.700 117.300 ;
        RECT 70.000 104.545 351.775 114.055 ;
        RECT 352.755 104.545 353.700 114.055 ;
        RECT 70.000 101.700 353.700 104.545 ;
        RECT 70.000 101.300 355.000 101.700 ;
        RECT 70.000 94.980 353.700 101.300 ;
        RECT 70.000 94.000 291.725 94.980 ;
        RECT 70.000 85.700 353.700 94.000 ;
        RECT 70.000 85.300 355.000 85.700 ;
        RECT 70.000 70.000 351.720 85.300 ;
        RECT 352.700 70.000 353.700 85.300 ;
      LAYER Metal5 ;
        RECT 277.600 353.400 280.710 355.000 ;
        RECT 70.000 235.835 76.380 353.400 ;
        RECT 77.960 242.515 92.380 353.400 ;
        RECT 93.960 351.800 139.720 353.400 ;
        RECT 93.960 351.780 125.400 351.800 ;
        RECT 93.960 351.735 117.400 351.780 ;
        RECT 93.960 350.155 101.400 351.735 ;
        RECT 133.600 350.220 139.720 351.800 ;
        RECT 125.600 350.200 139.720 350.220 ;
        RECT 117.600 350.155 139.720 350.200 ;
        RECT 93.960 262.545 139.720 350.155 ;
        RECT 141.300 269.235 155.720 353.400 ;
        RECT 157.300 351.860 187.720 353.400 ;
        RECT 157.300 350.380 171.440 351.860 ;
        RECT 172.920 350.380 187.720 351.860 ;
        RECT 157.300 282.600 187.720 350.380 ;
        RECT 189.300 351.860 256.710 353.400 ;
        RECT 189.300 350.280 245.400 351.860 ;
        RECT 253.600 350.280 256.710 351.860 ;
        RECT 189.300 306.575 256.710 350.280 ;
        RECT 258.290 313.245 272.710 353.400 ;
        RECT 274.290 316.560 280.710 353.400 ;
        RECT 282.290 353.400 285.400 355.000 ;
        RECT 348.990 353.400 355.000 355.000 ;
        RECT 282.290 329.850 312.710 353.400 ;
        RECT 314.290 333.210 320.710 353.400 ;
        RECT 322.290 348.990 355.000 353.400 ;
        RECT 322.290 333.210 353.400 348.990 ;
        RECT 314.290 329.850 353.400 333.210 ;
        RECT 282.290 317.600 353.400 329.850 ;
        RECT 282.290 316.560 351.365 317.600 ;
        RECT 274.290 313.245 351.365 316.560 ;
        RECT 258.290 309.400 351.365 313.245 ;
        RECT 352.945 309.400 353.400 317.600 ;
        RECT 258.290 306.575 353.400 309.400 ;
        RECT 189.300 282.600 353.400 306.575 ;
        RECT 157.300 269.235 353.400 282.600 ;
        RECT 141.300 262.545 353.400 269.235 ;
        RECT 93.960 257.910 353.400 262.545 ;
        RECT 93.960 256.430 351.985 257.910 ;
        RECT 93.960 250.570 353.400 256.430 ;
        RECT 93.960 249.090 351.980 250.570 ;
        RECT 93.960 242.515 353.400 249.090 ;
        RECT 77.960 235.835 353.400 242.515 ;
        RECT 70.000 229.400 353.400 235.835 ;
        RECT 70.000 213.600 355.000 229.400 ;
        RECT 70.000 205.600 351.435 213.600 ;
        RECT 70.000 197.600 351.405 205.600 ;
        RECT 353.015 205.400 353.400 213.600 ;
        RECT 70.000 181.600 351.370 197.600 ;
        RECT 352.985 197.400 353.400 205.400 ;
        RECT 70.000 165.400 351.320 181.600 ;
        RECT 352.950 181.400 353.400 197.400 ;
        RECT 352.900 165.400 353.400 181.400 ;
        RECT 70.000 158.620 353.400 165.400 ;
        RECT 70.000 157.040 292.805 158.620 ;
        RECT 70.000 142.620 353.400 157.040 ;
        RECT 70.000 141.040 292.805 142.620 ;
        RECT 70.000 130.950 353.400 141.040 ;
        RECT 70.000 129.370 255.865 130.950 ;
        RECT 70.000 125.600 353.400 129.370 ;
        RECT 70.000 117.600 351.520 125.600 ;
        RECT 70.000 101.400 351.475 117.600 ;
        RECT 353.100 117.400 353.400 125.600 ;
        RECT 353.055 101.400 353.400 117.400 ;
        RECT 70.000 95.280 353.400 101.400 ;
        RECT 70.000 93.700 291.425 95.280 ;
        RECT 70.000 85.600 353.400 93.700 ;
        RECT 70.000 70.000 351.420 85.600 ;
        RECT 353.000 70.000 353.400 85.600 ;
  END
END gf180mcu_fd_io__cor
END LIBRARY

