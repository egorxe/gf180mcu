magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< isosubstrate >>
rect 1197 -83 2889 2911
<< nwell >>
rect -83 1213 857 2911
rect 1197 1213 2889 2911
<< mvnmos >>
rect 317 354 457 654
rect 1605 354 1745 654
rect 1849 354 1989 654
rect 2093 354 2233 654
rect 2337 354 2477 654
<< mvpmos >>
rect 317 1622 457 2222
rect 1605 1622 1745 2222
rect 1849 1622 1989 2222
rect 2093 1622 2233 2222
rect 2337 1622 2477 2222
<< mvndiff >>
rect 229 641 317 654
rect 229 595 242 641
rect 288 595 317 641
rect 229 527 317 595
rect 229 481 242 527
rect 288 481 317 527
rect 229 413 317 481
rect 229 367 242 413
rect 288 367 317 413
rect 229 354 317 367
rect 457 641 545 654
rect 457 595 486 641
rect 532 595 545 641
rect 457 527 545 595
rect 457 481 486 527
rect 532 481 545 527
rect 457 413 545 481
rect 457 367 486 413
rect 532 367 545 413
rect 457 354 545 367
rect 1517 641 1605 654
rect 1517 595 1530 641
rect 1576 595 1605 641
rect 1517 527 1605 595
rect 1517 481 1530 527
rect 1576 481 1605 527
rect 1517 413 1605 481
rect 1517 367 1530 413
rect 1576 367 1605 413
rect 1517 354 1605 367
rect 1745 641 1849 654
rect 1745 595 1774 641
rect 1820 595 1849 641
rect 1745 527 1849 595
rect 1745 481 1774 527
rect 1820 481 1849 527
rect 1745 413 1849 481
rect 1745 367 1774 413
rect 1820 367 1849 413
rect 1745 354 1849 367
rect 1989 641 2093 654
rect 1989 595 2018 641
rect 2064 595 2093 641
rect 1989 527 2093 595
rect 1989 481 2018 527
rect 2064 481 2093 527
rect 1989 413 2093 481
rect 1989 367 2018 413
rect 2064 367 2093 413
rect 1989 354 2093 367
rect 2233 641 2337 654
rect 2233 595 2262 641
rect 2308 595 2337 641
rect 2233 527 2337 595
rect 2233 481 2262 527
rect 2308 481 2337 527
rect 2233 413 2337 481
rect 2233 367 2262 413
rect 2308 367 2337 413
rect 2233 354 2337 367
rect 2477 641 2565 654
rect 2477 595 2506 641
rect 2552 595 2565 641
rect 2477 527 2565 595
rect 2477 481 2506 527
rect 2552 481 2565 527
rect 2477 413 2565 481
rect 2477 367 2506 413
rect 2552 367 2565 413
rect 2477 354 2565 367
<< mvpdiff >>
rect 229 2209 317 2222
rect 229 2163 242 2209
rect 288 2163 317 2209
rect 229 2104 317 2163
rect 229 2058 242 2104
rect 288 2058 317 2104
rect 229 1999 317 2058
rect 229 1953 242 1999
rect 288 1953 317 1999
rect 229 1893 317 1953
rect 229 1847 242 1893
rect 288 1847 317 1893
rect 229 1787 317 1847
rect 229 1741 242 1787
rect 288 1741 317 1787
rect 229 1681 317 1741
rect 229 1635 242 1681
rect 288 1635 317 1681
rect 229 1622 317 1635
rect 457 2209 545 2222
rect 457 2163 486 2209
rect 532 2163 545 2209
rect 457 2104 545 2163
rect 457 2058 486 2104
rect 532 2058 545 2104
rect 457 1999 545 2058
rect 457 1953 486 1999
rect 532 1953 545 1999
rect 457 1893 545 1953
rect 457 1847 486 1893
rect 532 1847 545 1893
rect 457 1787 545 1847
rect 457 1741 486 1787
rect 532 1741 545 1787
rect 457 1681 545 1741
rect 457 1635 486 1681
rect 532 1635 545 1681
rect 457 1622 545 1635
rect 1517 2209 1605 2222
rect 1517 2163 1530 2209
rect 1576 2163 1605 2209
rect 1517 2104 1605 2163
rect 1517 2058 1530 2104
rect 1576 2058 1605 2104
rect 1517 1999 1605 2058
rect 1517 1953 1530 1999
rect 1576 1953 1605 1999
rect 1517 1893 1605 1953
rect 1517 1847 1530 1893
rect 1576 1847 1605 1893
rect 1517 1787 1605 1847
rect 1517 1741 1530 1787
rect 1576 1741 1605 1787
rect 1517 1681 1605 1741
rect 1517 1635 1530 1681
rect 1576 1635 1605 1681
rect 1517 1622 1605 1635
rect 1745 2209 1849 2222
rect 1745 2163 1774 2209
rect 1820 2163 1849 2209
rect 1745 2104 1849 2163
rect 1745 2058 1774 2104
rect 1820 2058 1849 2104
rect 1745 1999 1849 2058
rect 1745 1953 1774 1999
rect 1820 1953 1849 1999
rect 1745 1893 1849 1953
rect 1745 1847 1774 1893
rect 1820 1847 1849 1893
rect 1745 1787 1849 1847
rect 1745 1741 1774 1787
rect 1820 1741 1849 1787
rect 1745 1681 1849 1741
rect 1745 1635 1774 1681
rect 1820 1635 1849 1681
rect 1745 1622 1849 1635
rect 1989 2209 2093 2222
rect 1989 2163 2018 2209
rect 2064 2163 2093 2209
rect 1989 2104 2093 2163
rect 1989 2058 2018 2104
rect 2064 2058 2093 2104
rect 1989 1999 2093 2058
rect 1989 1953 2018 1999
rect 2064 1953 2093 1999
rect 1989 1893 2093 1953
rect 1989 1847 2018 1893
rect 2064 1847 2093 1893
rect 1989 1787 2093 1847
rect 1989 1741 2018 1787
rect 2064 1741 2093 1787
rect 1989 1681 2093 1741
rect 1989 1635 2018 1681
rect 2064 1635 2093 1681
rect 1989 1622 2093 1635
rect 2233 2209 2337 2222
rect 2233 2163 2262 2209
rect 2308 2163 2337 2209
rect 2233 2104 2337 2163
rect 2233 2058 2262 2104
rect 2308 2058 2337 2104
rect 2233 1999 2337 2058
rect 2233 1953 2262 1999
rect 2308 1953 2337 1999
rect 2233 1893 2337 1953
rect 2233 1847 2262 1893
rect 2308 1847 2337 1893
rect 2233 1787 2337 1847
rect 2233 1741 2262 1787
rect 2308 1741 2337 1787
rect 2233 1681 2337 1741
rect 2233 1635 2262 1681
rect 2308 1635 2337 1681
rect 2233 1622 2337 1635
rect 2477 2209 2565 2222
rect 2477 2163 2506 2209
rect 2552 2163 2565 2209
rect 2477 2104 2565 2163
rect 2477 2058 2506 2104
rect 2552 2058 2565 2104
rect 2477 1999 2565 2058
rect 2477 1953 2506 1999
rect 2552 1953 2565 1999
rect 2477 1893 2565 1953
rect 2477 1847 2506 1893
rect 2552 1847 2565 1893
rect 2477 1787 2565 1847
rect 2477 1741 2506 1787
rect 2552 1741 2565 1787
rect 2477 1681 2565 1741
rect 2477 1635 2506 1681
rect 2552 1635 2565 1681
rect 2477 1622 2565 1635
<< mvndiffc >>
rect 242 595 288 641
rect 242 481 288 527
rect 242 367 288 413
rect 486 595 532 641
rect 486 481 532 527
rect 486 367 532 413
rect 1530 595 1576 641
rect 1530 481 1576 527
rect 1530 367 1576 413
rect 1774 595 1820 641
rect 1774 481 1820 527
rect 1774 367 1820 413
rect 2018 595 2064 641
rect 2018 481 2064 527
rect 2018 367 2064 413
rect 2262 595 2308 641
rect 2262 481 2308 527
rect 2262 367 2308 413
rect 2506 595 2552 641
rect 2506 481 2552 527
rect 2506 367 2552 413
<< mvpdiffc >>
rect 242 2163 288 2209
rect 242 2058 288 2104
rect 242 1953 288 1999
rect 242 1847 288 1893
rect 242 1741 288 1787
rect 242 1635 288 1681
rect 486 2163 532 2209
rect 486 2058 532 2104
rect 486 1953 532 1999
rect 486 1847 532 1893
rect 486 1741 532 1787
rect 486 1635 532 1681
rect 1530 2163 1576 2209
rect 1530 2058 1576 2104
rect 1530 1953 1576 1999
rect 1530 1847 1576 1893
rect 1530 1741 1576 1787
rect 1530 1635 1576 1681
rect 1774 2163 1820 2209
rect 1774 2058 1820 2104
rect 1774 1953 1820 1999
rect 1774 1847 1820 1893
rect 1774 1741 1820 1787
rect 1774 1635 1820 1681
rect 2018 2163 2064 2209
rect 2018 2058 2064 2104
rect 2018 1953 2064 1999
rect 2018 1847 2064 1893
rect 2018 1741 2064 1787
rect 2018 1635 2064 1681
rect 2262 2163 2308 2209
rect 2262 2058 2308 2104
rect 2262 1953 2308 1999
rect 2262 1847 2308 1893
rect 2262 1741 2308 1787
rect 2262 1635 2308 1681
rect 2506 2163 2552 2209
rect 2506 2058 2552 2104
rect 2506 1953 2552 1999
rect 2506 1847 2552 1893
rect 2506 1741 2552 1787
rect 2506 1635 2552 1681
<< psubdiff >>
rect 0 1008 90 1030
rect 0 22 22 1008
rect 68 90 90 1008
rect 684 914 774 936
rect 684 90 706 914
rect 68 68 706 90
rect 68 22 176 68
rect 598 22 706 68
rect 752 22 774 914
rect 0 0 774 22
rect 1280 914 1370 936
rect 1280 22 1302 914
rect 1348 90 1370 914
rect 2716 1008 2806 1030
rect 2716 90 2738 1008
rect 1348 68 2738 90
rect 1348 22 1456 68
rect 2630 22 2738 68
rect 2784 22 2806 1008
rect 1280 0 2806 22
<< nsubdiff >>
rect 0 2806 774 2828
rect 0 1350 22 2806
rect 68 2760 176 2806
rect 598 2760 706 2806
rect 68 2738 706 2760
rect 68 1350 90 2738
rect 0 1328 90 1350
rect 684 1350 706 2738
rect 752 1350 774 2806
rect 684 1328 774 1350
rect 1280 2806 2806 2828
rect 1280 1350 1302 2806
rect 1348 2760 1456 2806
rect 2630 2760 2738 2806
rect 1348 2738 2738 2760
rect 1348 1350 1370 2738
rect 1280 1328 1370 1350
rect 2716 1350 2738 2738
rect 2784 1350 2806 2806
rect 2716 1328 2806 1350
<< psubdiffcont >>
rect 22 22 68 1008
rect 176 22 598 68
rect 706 22 752 914
rect 1302 22 1348 914
rect 1456 22 2630 68
rect 2738 22 2784 1008
<< nsubdiffcont >>
rect 22 1350 68 2806
rect 176 2760 598 2806
rect 706 1350 752 2806
rect 1302 1350 1348 2806
rect 1456 2760 2630 2806
rect 2738 1350 2784 2806
<< polysilicon >>
rect 317 2222 457 2266
rect 317 1167 457 1622
rect 1605 2222 1745 2266
rect 1849 2222 1989 2266
rect 2093 2222 2233 2266
rect 2337 2222 2477 2266
rect 317 1027 354 1167
rect 400 1027 457 1167
rect 317 654 457 1027
rect 1605 1202 1745 1622
rect 1849 1202 1989 1622
rect 1605 1167 1989 1202
rect 1605 1027 1642 1167
rect 1688 1027 1989 1167
rect 1605 991 1989 1027
rect 317 310 457 354
rect 1605 654 1745 991
rect 1849 654 1989 991
rect 2093 1202 2233 1622
rect 2337 1202 2477 1622
rect 2093 1167 2477 1202
rect 2093 1027 2130 1167
rect 2176 1027 2477 1167
rect 2093 991 2477 1027
rect 2093 654 2233 991
rect 2337 654 2477 991
rect 1605 310 1745 354
rect 1849 310 1989 354
rect 2093 310 2233 354
rect 2337 310 2477 354
<< polycontact >>
rect 354 1027 400 1167
rect 1642 1027 1688 1167
rect 2130 1027 2176 1167
<< metal1 >>
rect 11 2806 763 2817
rect 11 1350 22 2806
rect 68 2760 176 2806
rect 598 2760 706 2806
rect 68 2749 706 2760
rect 68 1350 79 2749
rect 227 2209 303 2749
rect 227 2163 242 2209
rect 288 2163 303 2209
rect 227 2104 303 2163
rect 227 2058 242 2104
rect 288 2058 303 2104
rect 227 1999 303 2058
rect 227 1953 242 1999
rect 288 1953 303 1999
rect 227 1893 303 1953
rect 227 1847 242 1893
rect 288 1847 303 1893
rect 227 1787 303 1847
rect 227 1741 242 1787
rect 288 1741 303 1787
rect 227 1681 303 1741
rect 227 1635 242 1681
rect 288 1635 303 1681
rect 227 1622 303 1635
rect 471 2209 547 2222
rect 471 2163 486 2209
rect 532 2163 547 2209
rect 471 2104 547 2163
rect 471 2058 486 2104
rect 532 2058 547 2104
rect 471 1999 547 2058
rect 471 1953 486 1999
rect 532 1953 547 1999
rect 471 1893 547 1953
rect 471 1847 486 1893
rect 532 1847 547 1893
rect 471 1787 547 1847
rect 471 1741 486 1787
rect 532 1741 547 1787
rect 471 1681 547 1741
rect 471 1635 486 1681
rect 532 1635 547 1681
rect 11 1339 79 1350
rect 471 1186 547 1635
rect 695 1350 706 2749
rect 752 1350 763 2806
rect 695 1339 763 1350
rect 1291 2806 2795 2817
rect 1291 1350 1302 2806
rect 1348 2760 1456 2806
rect 2630 2760 2738 2806
rect 1348 2749 2738 2760
rect 1348 1350 1359 2749
rect 1515 2209 1591 2749
rect 1515 2163 1530 2209
rect 1576 2163 1591 2209
rect 1515 2104 1591 2163
rect 1515 2058 1530 2104
rect 1576 2058 1591 2104
rect 1515 1999 1591 2058
rect 1515 1953 1530 1999
rect 1576 1953 1591 1999
rect 1515 1893 1591 1953
rect 1515 1847 1530 1893
rect 1576 1847 1591 1893
rect 1515 1787 1591 1847
rect 1515 1741 1530 1787
rect 1576 1741 1591 1787
rect 1515 1681 1591 1741
rect 1515 1635 1530 1681
rect 1576 1635 1591 1681
rect 1515 1622 1591 1635
rect 1759 2209 1835 2222
rect 1759 2163 1774 2209
rect 1820 2163 1835 2209
rect 1759 2104 1835 2163
rect 1759 2058 1774 2104
rect 1820 2058 1835 2104
rect 1759 1999 1835 2058
rect 1759 1953 1774 1999
rect 1820 1953 1835 1999
rect 1759 1893 1835 1953
rect 1759 1847 1774 1893
rect 1820 1847 1835 1893
rect 1759 1787 1835 1847
rect 1759 1741 1774 1787
rect 1820 1741 1835 1787
rect 1759 1681 1835 1741
rect 1759 1635 1774 1681
rect 1820 1635 1835 1681
rect 1291 1339 1359 1350
rect 1759 1186 1835 1635
rect 2003 2209 2079 2749
rect 2003 2163 2018 2209
rect 2064 2163 2079 2209
rect 2003 2104 2079 2163
rect 2003 2058 2018 2104
rect 2064 2058 2079 2104
rect 2003 1999 2079 2058
rect 2003 1953 2018 1999
rect 2064 1953 2079 1999
rect 2003 1893 2079 1953
rect 2003 1847 2018 1893
rect 2064 1847 2079 1893
rect 2003 1787 2079 1847
rect 2003 1741 2018 1787
rect 2064 1741 2079 1787
rect 2003 1681 2079 1741
rect 2003 1635 2018 1681
rect 2064 1635 2079 1681
rect 2003 1622 2079 1635
rect 2247 2209 2323 2222
rect 2247 2163 2262 2209
rect 2308 2163 2323 2209
rect 2247 2104 2323 2163
rect 2247 2058 2262 2104
rect 2308 2058 2323 2104
rect 2247 1999 2323 2058
rect 2247 1953 2262 1999
rect 2308 1953 2323 1999
rect 2247 1893 2323 1953
rect 2247 1847 2262 1893
rect 2308 1847 2323 1893
rect 2247 1787 2323 1847
rect 2247 1741 2262 1787
rect 2308 1741 2323 1787
rect 2247 1681 2323 1741
rect 2247 1635 2262 1681
rect 2308 1635 2323 1681
rect 343 1167 411 1178
rect 343 1027 354 1167
rect 400 1027 411 1167
rect 11 1008 79 1019
rect 343 1016 411 1027
rect 471 1167 1699 1186
rect 471 1027 1642 1167
rect 1688 1027 1699 1167
rect 11 22 22 1008
rect 68 79 79 1008
rect 471 1008 1699 1027
rect 1759 1167 2187 1186
rect 1759 1027 2130 1167
rect 2176 1027 2187 1167
rect 1759 1008 2187 1027
rect 227 641 303 654
rect 227 595 242 641
rect 288 595 303 641
rect 227 527 303 595
rect 227 481 242 527
rect 288 481 303 527
rect 227 413 303 481
rect 227 367 242 413
rect 288 367 303 413
rect 227 79 303 367
rect 471 641 547 1008
rect 471 595 486 641
rect 532 595 547 641
rect 471 527 547 595
rect 471 481 486 527
rect 532 481 547 527
rect 471 413 547 481
rect 471 367 486 413
rect 532 367 547 413
rect 471 354 547 367
rect 695 914 763 925
rect 695 79 706 914
rect 68 68 706 79
rect 68 22 176 68
rect 598 22 706 68
rect 752 22 763 914
rect 11 11 763 22
rect 1291 914 1359 925
rect 1291 22 1302 914
rect 1348 79 1359 914
rect 1515 641 1591 654
rect 1515 595 1530 641
rect 1576 595 1591 641
rect 1515 527 1591 595
rect 1515 481 1530 527
rect 1576 481 1591 527
rect 1515 413 1591 481
rect 1515 367 1530 413
rect 1576 367 1591 413
rect 1515 79 1591 367
rect 1759 641 1835 1008
rect 1759 595 1774 641
rect 1820 595 1835 641
rect 1759 527 1835 595
rect 1759 481 1774 527
rect 1820 481 1835 527
rect 1759 413 1835 481
rect 1759 367 1774 413
rect 1820 367 1835 413
rect 1759 354 1835 367
rect 2003 641 2079 654
rect 2003 595 2018 641
rect 2064 595 2079 641
rect 2003 527 2079 595
rect 2003 481 2018 527
rect 2064 481 2079 527
rect 2003 413 2079 481
rect 2003 367 2018 413
rect 2064 367 2079 413
rect 2003 79 2079 367
rect 2247 641 2323 1635
rect 2491 2209 2567 2749
rect 2491 2163 2506 2209
rect 2552 2163 2567 2209
rect 2491 2104 2567 2163
rect 2491 2058 2506 2104
rect 2552 2058 2567 2104
rect 2491 1999 2567 2058
rect 2491 1953 2506 1999
rect 2552 1953 2567 1999
rect 2491 1893 2567 1953
rect 2491 1847 2506 1893
rect 2552 1847 2567 1893
rect 2491 1787 2567 1847
rect 2491 1741 2506 1787
rect 2552 1741 2567 1787
rect 2491 1681 2567 1741
rect 2491 1635 2506 1681
rect 2552 1635 2567 1681
rect 2491 1622 2567 1635
rect 2727 1350 2738 2749
rect 2784 1350 2795 2806
rect 2727 1339 2795 1350
rect 2727 1008 2795 1019
rect 2247 595 2262 641
rect 2308 595 2323 641
rect 2247 527 2323 595
rect 2247 481 2262 527
rect 2308 481 2323 527
rect 2247 413 2323 481
rect 2247 367 2262 413
rect 2308 367 2323 413
rect 2247 354 2323 367
rect 2491 641 2567 654
rect 2491 595 2506 641
rect 2552 595 2567 641
rect 2491 527 2567 595
rect 2491 481 2506 527
rect 2552 481 2567 527
rect 2491 413 2567 481
rect 2491 367 2506 413
rect 2552 367 2567 413
rect 2491 79 2567 367
rect 2727 79 2738 1008
rect 1348 68 2738 79
rect 1348 22 1456 68
rect 2630 22 2738 68
rect 2784 22 2795 1008
rect 1291 11 2795 22
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_0
timestamp 1759194789
transform 1 0 2761 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_1
timestamp 1759194789
transform 1 0 45 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_2
timestamp 1759194789
transform 1 0 729 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_3
timestamp 1759194789
transform 1 0 1325 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145273  M1_NWELL_CDNS_40661953145273_0
timestamp 1759194789
transform 1 0 387 0 1 2783
box 0 0 1 1
use M1_NWELL_CDNS_40661953145274  M1_NWELL_CDNS_40661953145274_0
timestamp 1759194789
transform 1 0 2043 0 1 2783
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_0
timestamp 1759194789
transform 1 0 2153 0 1 1097
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_1
timestamp 1759194789
transform 1 0 1665 0 1 1097
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_2
timestamp 1759194789
transform 1 0 377 0 1 1097
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_0
timestamp 1759194789
transform 1 0 45 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_1
timestamp 1759194789
transform 1 0 2761 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145228  M1_PSUB_CDNS_40661953145228_0
timestamp 1759194789
transform 1 0 729 0 -1 468
box 0 0 1 1
use M1_PSUB_CDNS_40661953145228  M1_PSUB_CDNS_40661953145228_1
timestamp 1759194789
transform 1 0 1325 0 -1 468
box 0 0 1 1
use M1_PSUB_CDNS_40661953145237  M1_PSUB_CDNS_40661953145237_0
timestamp 1759194789
transform 1 0 387 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661953145275  M1_PSUB_CDNS_40661953145275_0
timestamp 1759194789
transform 1 0 2043 0 -1 45
box 0 0 1 1
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1759194789
transform 1 0 317 0 1 354
box 0 0 1 1
use nmos_6p0_CDNS_4066195314531  nmos_6p0_CDNS_4066195314531_0
timestamp 1759194789
transform 1 0 2093 0 1 354
box 0 0 1 1
use nmos_6p0_CDNS_4066195314531  nmos_6p0_CDNS_4066195314531_1
timestamp 1759194789
transform 1 0 1605 0 1 354
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1759194789
transform 1 0 317 0 1 1622
box 0 0 1 1
use pmos_6p0_CDNS_4066195314529  pmos_6p0_CDNS_4066195314529_0
timestamp 1759194789
transform 1 0 2093 0 1 1622
box 0 0 1 1
use pmos_6p0_CDNS_4066195314529  pmos_6p0_CDNS_4066195314529_1
timestamp 1759194789
transform 1 0 1605 0 1 1622
box 0 0 1 1
<< labels >>
rlabel metal1 s 2031 1098 2031 1098 4 Z
port 1 nsew
rlabel metal1 s 263 45 263 45 4 VSS
port 2 nsew
rlabel metal1 s 2433 45 2433 45 4 DVSS
port 3 nsew
rlabel metal1 s 2442 2788 2442 2788 4 DVDD
port 4 nsew
rlabel metal1 s 377 1098 377 1098 4 A
port 5 nsew
rlabel metal1 s 350 2788 350 2788 4 VDD
port 6 nsew
rlabel metal1 s 2286 1098 2286 1098 4 ZB
port 7 nsew
<< properties >>
string GDS_END 1794310
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1790390
string path 44.925 8.850 44.925 55.550 
<< end >>
