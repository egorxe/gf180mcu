magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< isosubstrate >>
rect 294 20724 14770 56850
rect 1350 15369 13714 20724
<< nwell >>
rect 2400 20168 12664 20724
rect 2400 16224 2956 20168
rect 12108 16224 12664 20168
rect 2400 15668 12664 16224
<< pwell >>
rect 790 53248 3966 56248
rect 4226 53248 7402 56248
rect 7662 53248 10838 56248
rect 11098 53248 14274 56248
rect 790 49300 3966 52300
rect 4226 49300 7402 52300
rect 7662 49300 10838 52300
rect 11098 49300 14274 52300
rect 790 45352 3966 48352
rect 4226 45352 7402 48352
rect 7662 45352 10838 48352
rect 11098 45352 14274 48352
rect 790 41404 3966 44404
rect 4226 41404 7402 44404
rect 7662 41404 10838 44404
rect 11098 41404 14274 44404
rect 790 37456 3966 40456
rect 4226 37456 7402 40456
rect 7662 37456 10838 40456
rect 11098 37456 14274 40456
rect 790 33508 3966 36508
rect 4226 33508 7402 36508
rect 7662 33508 10838 36508
rect 11098 33508 14274 36508
rect 790 29560 3966 32560
rect 4226 29560 7402 32560
rect 7662 29560 10838 32560
rect 11098 29560 14274 32560
rect 790 25612 3966 28612
rect 4226 25612 7402 28612
rect 7662 25612 10838 28612
rect 11098 25612 14274 28612
rect 790 21664 3966 24664
rect 4226 21664 7402 24664
rect 7662 21664 10838 24664
rect 11098 21664 14274 24664
<< mvndiff >>
rect 790 56211 878 56248
rect 790 53285 803 56211
rect 849 53285 878 56211
rect 790 53248 878 53285
rect 3878 56211 3966 56248
rect 3878 53285 3907 56211
rect 3953 53285 3966 56211
rect 3878 53248 3966 53285
rect 4226 56211 4314 56248
rect 4226 53285 4239 56211
rect 4285 53285 4314 56211
rect 4226 53248 4314 53285
rect 7314 56211 7402 56248
rect 7314 53285 7343 56211
rect 7389 53285 7402 56211
rect 7314 53248 7402 53285
rect 7662 56211 7750 56248
rect 7662 53285 7675 56211
rect 7721 53285 7750 56211
rect 7662 53248 7750 53285
rect 10750 56211 10838 56248
rect 10750 53285 10779 56211
rect 10825 53285 10838 56211
rect 10750 53248 10838 53285
rect 11098 56211 11186 56248
rect 11098 53285 11111 56211
rect 11157 53285 11186 56211
rect 11098 53248 11186 53285
rect 14186 56211 14274 56248
rect 14186 53285 14215 56211
rect 14261 53285 14274 56211
rect 14186 53248 14274 53285
rect 790 52263 878 52300
rect 790 49337 803 52263
rect 849 49337 878 52263
rect 790 49300 878 49337
rect 3878 52263 3966 52300
rect 3878 49337 3907 52263
rect 3953 49337 3966 52263
rect 3878 49300 3966 49337
rect 4226 52263 4314 52300
rect 4226 49337 4239 52263
rect 4285 49337 4314 52263
rect 4226 49300 4314 49337
rect 7314 52263 7402 52300
rect 7314 49337 7343 52263
rect 7389 49337 7402 52263
rect 7314 49300 7402 49337
rect 7662 52263 7750 52300
rect 7662 49337 7675 52263
rect 7721 49337 7750 52263
rect 7662 49300 7750 49337
rect 10750 52263 10838 52300
rect 10750 49337 10779 52263
rect 10825 49337 10838 52263
rect 10750 49300 10838 49337
rect 11098 52263 11186 52300
rect 11098 49337 11111 52263
rect 11157 49337 11186 52263
rect 11098 49300 11186 49337
rect 14186 52263 14274 52300
rect 14186 49337 14215 52263
rect 14261 49337 14274 52263
rect 14186 49300 14274 49337
rect 790 48315 878 48352
rect 790 45389 803 48315
rect 849 45389 878 48315
rect 790 45352 878 45389
rect 3878 48315 3966 48352
rect 3878 45389 3907 48315
rect 3953 45389 3966 48315
rect 3878 45352 3966 45389
rect 4226 48315 4314 48352
rect 4226 45389 4239 48315
rect 4285 45389 4314 48315
rect 4226 45352 4314 45389
rect 7314 48315 7402 48352
rect 7314 45389 7343 48315
rect 7389 45389 7402 48315
rect 7314 45352 7402 45389
rect 7662 48315 7750 48352
rect 7662 45389 7675 48315
rect 7721 45389 7750 48315
rect 7662 45352 7750 45389
rect 10750 48315 10838 48352
rect 10750 45389 10779 48315
rect 10825 45389 10838 48315
rect 10750 45352 10838 45389
rect 11098 48315 11186 48352
rect 11098 45389 11111 48315
rect 11157 45389 11186 48315
rect 11098 45352 11186 45389
rect 14186 48315 14274 48352
rect 14186 45389 14215 48315
rect 14261 45389 14274 48315
rect 14186 45352 14274 45389
rect 790 44367 878 44404
rect 790 41441 803 44367
rect 849 41441 878 44367
rect 790 41404 878 41441
rect 3878 44367 3966 44404
rect 3878 41441 3907 44367
rect 3953 41441 3966 44367
rect 3878 41404 3966 41441
rect 4226 44367 4314 44404
rect 4226 41441 4239 44367
rect 4285 41441 4314 44367
rect 4226 41404 4314 41441
rect 7314 44367 7402 44404
rect 7314 41441 7343 44367
rect 7389 41441 7402 44367
rect 7314 41404 7402 41441
rect 7662 44367 7750 44404
rect 7662 41441 7675 44367
rect 7721 41441 7750 44367
rect 7662 41404 7750 41441
rect 10750 44367 10838 44404
rect 10750 41441 10779 44367
rect 10825 41441 10838 44367
rect 10750 41404 10838 41441
rect 11098 44367 11186 44404
rect 11098 41441 11111 44367
rect 11157 41441 11186 44367
rect 11098 41404 11186 41441
rect 14186 44367 14274 44404
rect 14186 41441 14215 44367
rect 14261 41441 14274 44367
rect 14186 41404 14274 41441
rect 790 40419 878 40456
rect 790 37493 803 40419
rect 849 37493 878 40419
rect 790 37456 878 37493
rect 3878 40419 3966 40456
rect 3878 37493 3907 40419
rect 3953 37493 3966 40419
rect 3878 37456 3966 37493
rect 4226 40419 4314 40456
rect 4226 37493 4239 40419
rect 4285 37493 4314 40419
rect 4226 37456 4314 37493
rect 7314 40419 7402 40456
rect 7314 37493 7343 40419
rect 7389 37493 7402 40419
rect 7314 37456 7402 37493
rect 7662 40419 7750 40456
rect 7662 37493 7675 40419
rect 7721 37493 7750 40419
rect 7662 37456 7750 37493
rect 10750 40419 10838 40456
rect 10750 37493 10779 40419
rect 10825 37493 10838 40419
rect 10750 37456 10838 37493
rect 11098 40419 11186 40456
rect 11098 37493 11111 40419
rect 11157 37493 11186 40419
rect 11098 37456 11186 37493
rect 14186 40419 14274 40456
rect 14186 37493 14215 40419
rect 14261 37493 14274 40419
rect 14186 37456 14274 37493
rect 790 36471 878 36508
rect 790 33545 803 36471
rect 849 33545 878 36471
rect 790 33508 878 33545
rect 3878 36471 3966 36508
rect 3878 33545 3907 36471
rect 3953 33545 3966 36471
rect 3878 33508 3966 33545
rect 4226 36471 4314 36508
rect 4226 33545 4239 36471
rect 4285 33545 4314 36471
rect 4226 33508 4314 33545
rect 7314 36471 7402 36508
rect 7314 33545 7343 36471
rect 7389 33545 7402 36471
rect 7314 33508 7402 33545
rect 7662 36471 7750 36508
rect 7662 33545 7675 36471
rect 7721 33545 7750 36471
rect 7662 33508 7750 33545
rect 10750 36471 10838 36508
rect 10750 33545 10779 36471
rect 10825 33545 10838 36471
rect 10750 33508 10838 33545
rect 11098 36471 11186 36508
rect 11098 33545 11111 36471
rect 11157 33545 11186 36471
rect 11098 33508 11186 33545
rect 14186 36471 14274 36508
rect 14186 33545 14215 36471
rect 14261 33545 14274 36471
rect 14186 33508 14274 33545
rect 790 32523 878 32560
rect 790 29597 803 32523
rect 849 29597 878 32523
rect 790 29560 878 29597
rect 3878 32523 3966 32560
rect 3878 29597 3907 32523
rect 3953 29597 3966 32523
rect 3878 29560 3966 29597
rect 4226 32523 4314 32560
rect 4226 29597 4239 32523
rect 4285 29597 4314 32523
rect 4226 29560 4314 29597
rect 7314 32523 7402 32560
rect 7314 29597 7343 32523
rect 7389 29597 7402 32523
rect 7314 29560 7402 29597
rect 7662 32523 7750 32560
rect 7662 29597 7675 32523
rect 7721 29597 7750 32523
rect 7662 29560 7750 29597
rect 10750 32523 10838 32560
rect 10750 29597 10779 32523
rect 10825 29597 10838 32523
rect 10750 29560 10838 29597
rect 11098 32523 11186 32560
rect 11098 29597 11111 32523
rect 11157 29597 11186 32523
rect 11098 29560 11186 29597
rect 14186 32523 14274 32560
rect 14186 29597 14215 32523
rect 14261 29597 14274 32523
rect 14186 29560 14274 29597
rect 790 28575 878 28612
rect 790 25649 803 28575
rect 849 25649 878 28575
rect 790 25612 878 25649
rect 3878 28575 3966 28612
rect 3878 25649 3907 28575
rect 3953 25649 3966 28575
rect 3878 25612 3966 25649
rect 4226 28575 4314 28612
rect 4226 25649 4239 28575
rect 4285 25649 4314 28575
rect 4226 25612 4314 25649
rect 7314 28575 7402 28612
rect 7314 25649 7343 28575
rect 7389 25649 7402 28575
rect 7314 25612 7402 25649
rect 7662 28575 7750 28612
rect 7662 25649 7675 28575
rect 7721 25649 7750 28575
rect 7662 25612 7750 25649
rect 10750 28575 10838 28612
rect 10750 25649 10779 28575
rect 10825 25649 10838 28575
rect 10750 25612 10838 25649
rect 11098 28575 11186 28612
rect 11098 25649 11111 28575
rect 11157 25649 11186 28575
rect 11098 25612 11186 25649
rect 14186 28575 14274 28612
rect 14186 25649 14215 28575
rect 14261 25649 14274 28575
rect 14186 25612 14274 25649
rect 790 24627 878 24664
rect 790 21701 803 24627
rect 849 21701 878 24627
rect 790 21664 878 21701
rect 3878 24627 3966 24664
rect 3878 21701 3907 24627
rect 3953 21701 3966 24627
rect 3878 21664 3966 21701
rect 4226 24627 4314 24664
rect 4226 21701 4239 24627
rect 4285 21701 4314 24627
rect 4226 21664 4314 21701
rect 7314 24627 7402 24664
rect 7314 21701 7343 24627
rect 7389 21701 7402 24627
rect 7314 21664 7402 21701
rect 7662 24627 7750 24664
rect 7662 21701 7675 24627
rect 7721 21701 7750 24627
rect 7662 21664 7750 21701
rect 10750 24627 10838 24664
rect 10750 21701 10779 24627
rect 10825 21701 10838 24627
rect 10750 21664 10838 21701
rect 11098 24627 11186 24664
rect 11098 21701 11111 24627
rect 11157 21701 11186 24627
rect 11098 21664 11186 21701
rect 14186 24627 14274 24664
rect 14186 21701 14215 24627
rect 14261 21701 14274 24627
rect 14186 21664 14274 21701
<< mvndiffc >>
rect 803 53285 849 56211
rect 3907 53285 3953 56211
rect 4239 53285 4285 56211
rect 7343 53285 7389 56211
rect 7675 53285 7721 56211
rect 10779 53285 10825 56211
rect 11111 53285 11157 56211
rect 14215 53285 14261 56211
rect 803 49337 849 52263
rect 3907 49337 3953 52263
rect 4239 49337 4285 52263
rect 7343 49337 7389 52263
rect 7675 49337 7721 52263
rect 10779 49337 10825 52263
rect 11111 49337 11157 52263
rect 14215 49337 14261 52263
rect 803 45389 849 48315
rect 3907 45389 3953 48315
rect 4239 45389 4285 48315
rect 7343 45389 7389 48315
rect 7675 45389 7721 48315
rect 10779 45389 10825 48315
rect 11111 45389 11157 48315
rect 14215 45389 14261 48315
rect 803 41441 849 44367
rect 3907 41441 3953 44367
rect 4239 41441 4285 44367
rect 7343 41441 7389 44367
rect 7675 41441 7721 44367
rect 10779 41441 10825 44367
rect 11111 41441 11157 44367
rect 14215 41441 14261 44367
rect 803 37493 849 40419
rect 3907 37493 3953 40419
rect 4239 37493 4285 40419
rect 7343 37493 7389 40419
rect 7675 37493 7721 40419
rect 10779 37493 10825 40419
rect 11111 37493 11157 40419
rect 14215 37493 14261 40419
rect 803 33545 849 36471
rect 3907 33545 3953 36471
rect 4239 33545 4285 36471
rect 7343 33545 7389 36471
rect 7675 33545 7721 36471
rect 10779 33545 10825 36471
rect 11111 33545 11157 36471
rect 14215 33545 14261 36471
rect 803 29597 849 32523
rect 3907 29597 3953 32523
rect 4239 29597 4285 32523
rect 7343 29597 7389 32523
rect 7675 29597 7721 32523
rect 10779 29597 10825 32523
rect 11111 29597 11157 32523
rect 14215 29597 14261 32523
rect 803 25649 849 28575
rect 3907 25649 3953 28575
rect 4239 25649 4285 28575
rect 7343 25649 7389 28575
rect 7675 25649 7721 28575
rect 10779 25649 10825 28575
rect 11111 25649 11157 28575
rect 14215 25649 14261 28575
rect 803 21701 849 24627
rect 3907 21701 3953 24627
rect 4239 21701 4285 24627
rect 7343 21701 7389 24627
rect 7675 21701 7721 24627
rect 10779 21701 10825 24627
rect 11111 21701 11157 24627
rect 14215 21701 14261 24627
<< psubdiff >>
rect 377 56745 14687 56767
rect 377 21167 399 56745
rect 445 56699 553 56745
rect 14511 56699 14619 56745
rect 445 56677 14619 56699
rect 445 21235 467 56677
rect 531 52797 14533 52819
rect 531 52751 553 52797
rect 14511 52751 14533 52797
rect 531 52729 14533 52751
rect 531 48849 14533 48871
rect 531 48803 553 48849
rect 14511 48803 14533 48849
rect 531 48781 14533 48803
rect 531 44901 14533 44923
rect 531 44855 553 44901
rect 14511 44855 14533 44901
rect 531 44833 14533 44855
rect 531 40953 14533 40975
rect 531 40907 553 40953
rect 14511 40907 14533 40953
rect 531 40885 14533 40907
rect 531 37005 14533 37027
rect 531 36959 553 37005
rect 14511 36959 14533 37005
rect 531 36937 14533 36959
rect 531 33057 14533 33079
rect 531 33011 553 33057
rect 14511 33011 14533 33057
rect 531 32989 14533 33011
rect 531 29109 14533 29131
rect 531 29063 553 29109
rect 14511 29063 14533 29109
rect 531 29041 14533 29063
rect 531 25161 14533 25183
rect 531 25115 553 25161
rect 14511 25115 14533 25161
rect 531 25093 14533 25115
rect 14597 21235 14619 56677
rect 445 21213 14619 21235
rect 445 21167 553 21213
rect 14511 21167 14619 21213
rect 14665 21167 14687 56745
rect 377 21145 14687 21167
rect 289 20357 1079 20379
rect 289 911 311 20357
rect 1057 911 1079 20357
rect 3116 19971 11948 19993
rect 3116 19925 3138 19971
rect 11926 19925 11948 19971
rect 3116 19817 11948 19925
rect 3116 16575 3138 19817
rect 3184 19809 3467 19817
rect 3184 19199 3292 19809
rect 3338 19771 3467 19809
rect 11597 19809 11880 19817
rect 11597 19771 11726 19809
rect 3338 19749 11726 19771
rect 3338 19267 3360 19749
rect 11704 19267 11726 19749
rect 3338 19245 11726 19267
rect 3338 19199 3467 19245
rect 11597 19199 11726 19245
rect 11772 19199 11880 19809
rect 3184 19091 11880 19199
rect 3184 19045 3326 19091
rect 11738 19045 11880 19091
rect 3184 18937 11880 19045
rect 3184 18327 3292 18937
rect 3338 18891 3467 18937
rect 11597 18891 11726 18937
rect 3338 18869 11726 18891
rect 3338 18395 3360 18869
rect 11704 18395 11726 18869
rect 3338 18373 11726 18395
rect 3338 18327 3467 18373
rect 11597 18327 11726 18373
rect 11772 18327 11880 18937
rect 3184 18219 11880 18327
rect 3184 18173 3326 18219
rect 11738 18173 11880 18219
rect 3184 18065 11880 18173
rect 3184 17455 3292 18065
rect 3338 18019 3467 18065
rect 11597 18019 11726 18065
rect 3338 17997 11726 18019
rect 3338 17523 3360 17997
rect 11704 17523 11726 17997
rect 3338 17501 11726 17523
rect 3338 17455 3467 17501
rect 11597 17455 11726 17501
rect 11772 17455 11880 18065
rect 3184 17347 11880 17455
rect 3184 17301 3326 17347
rect 11738 17301 11880 17347
rect 3184 17193 11880 17301
rect 3184 16583 3292 17193
rect 3338 17147 3467 17193
rect 11597 17147 11726 17193
rect 3338 17125 11726 17147
rect 3338 16643 3360 17125
rect 11704 16643 11726 17125
rect 3338 16621 11726 16643
rect 3338 16583 3467 16621
rect 3184 16575 3467 16583
rect 11597 16583 11726 16621
rect 11772 16583 11880 17193
rect 11597 16575 11880 16583
rect 11926 16575 11948 19817
rect 3116 16467 11948 16575
rect 3116 16421 3138 16467
rect 11926 16421 11948 16467
rect 3116 16399 11948 16421
rect 13985 20357 14775 20379
rect 289 889 1079 911
rect 13985 911 14007 20357
rect 14753 911 14775 20357
rect 13985 889 14775 911
<< nsubdiff >>
rect 2483 20619 12581 20641
rect 2483 15773 2505 20619
rect 2851 20273 2959 20619
rect 12105 20273 12213 20619
rect 2851 20251 12213 20273
rect 2851 16141 2873 20251
rect 12191 16141 12213 20251
rect 2851 16119 12213 16141
rect 2851 15773 2959 16119
rect 12105 15773 12213 16119
rect 12559 15773 12581 20619
rect 2483 15751 12581 15773
<< psubdiffcont >>
rect 399 21167 445 56745
rect 553 56699 14511 56745
rect 553 52751 14511 52797
rect 553 48803 14511 48849
rect 553 44855 14511 44901
rect 553 40907 14511 40953
rect 553 36959 14511 37005
rect 553 33011 14511 33057
rect 553 29063 14511 29109
rect 553 25115 14511 25161
rect 553 21167 14511 21213
rect 14619 21167 14665 56745
rect 311 911 1057 20357
rect 3138 19925 11926 19971
rect 3138 16575 3184 19817
rect 3292 19199 3338 19809
rect 3467 19771 11597 19817
rect 3467 19199 11597 19245
rect 11726 19199 11772 19809
rect 3326 19045 11738 19091
rect 3292 18327 3338 18937
rect 3467 18891 11597 18937
rect 3467 18327 11597 18373
rect 11726 18327 11772 18937
rect 3326 18173 11738 18219
rect 3292 17455 3338 18065
rect 3467 18019 11597 18065
rect 3467 17455 11597 17501
rect 11726 17455 11772 18065
rect 3326 17301 11738 17347
rect 3292 16583 3338 17193
rect 3467 17147 11597 17193
rect 3467 16575 11597 16621
rect 11726 16583 11772 17193
rect 11880 16575 11926 19817
rect 3138 16421 11926 16467
rect 14007 911 14753 20357
<< nsubdiffcont >>
rect 2505 15773 2851 20619
rect 2959 20273 12105 20619
rect 2959 15773 12105 16119
rect 12213 15773 12559 20619
<< mvnmoscap >>
rect 878 53248 3878 56248
rect 4314 53248 7314 56248
rect 7750 53248 10750 56248
rect 11186 53248 14186 56248
rect 878 49300 3878 52300
rect 4314 49300 7314 52300
rect 7750 49300 10750 52300
rect 11186 49300 14186 52300
rect 878 45352 3878 48352
rect 4314 45352 7314 48352
rect 7750 45352 10750 48352
rect 11186 45352 14186 48352
rect 878 41404 3878 44404
rect 4314 41404 7314 44404
rect 7750 41404 10750 44404
rect 11186 41404 14186 44404
rect 878 37456 3878 40456
rect 4314 37456 7314 40456
rect 7750 37456 10750 40456
rect 11186 37456 14186 40456
rect 878 33508 3878 36508
rect 4314 33508 7314 36508
rect 7750 33508 10750 36508
rect 11186 33508 14186 36508
rect 878 29560 3878 32560
rect 4314 29560 7314 32560
rect 7750 29560 10750 32560
rect 11186 29560 14186 32560
rect 878 25612 3878 28612
rect 4314 25612 7314 28612
rect 7750 25612 10750 28612
rect 11186 25612 14186 28612
rect 878 21664 3878 24664
rect 4314 21664 7314 24664
rect 7750 21664 10750 24664
rect 11186 21664 14186 24664
<< polysilicon >>
rect 878 56327 3878 56340
rect 878 56281 931 56327
rect 3825 56281 3878 56327
rect 878 56248 3878 56281
rect 4314 56327 7314 56340
rect 4314 56281 4367 56327
rect 7261 56281 7314 56327
rect 4314 56248 7314 56281
rect 7750 56327 10750 56340
rect 7750 56281 7803 56327
rect 10697 56281 10750 56327
rect 7750 56248 10750 56281
rect 11186 56327 14186 56340
rect 11186 56281 11239 56327
rect 14133 56281 14186 56327
rect 11186 56248 14186 56281
rect 878 53215 3878 53248
rect 878 53169 931 53215
rect 3825 53169 3878 53215
rect 878 53156 3878 53169
rect 4314 53215 7314 53248
rect 4314 53169 4367 53215
rect 7261 53169 7314 53215
rect 4314 53156 7314 53169
rect 7750 53215 10750 53248
rect 7750 53169 7803 53215
rect 10697 53169 10750 53215
rect 7750 53156 10750 53169
rect 11186 53215 14186 53248
rect 11186 53169 11239 53215
rect 14133 53169 14186 53215
rect 11186 53156 14186 53169
rect 878 52379 3878 52392
rect 878 52333 931 52379
rect 3825 52333 3878 52379
rect 878 52300 3878 52333
rect 4314 52379 7314 52392
rect 4314 52333 4367 52379
rect 7261 52333 7314 52379
rect 4314 52300 7314 52333
rect 7750 52379 10750 52392
rect 7750 52333 7803 52379
rect 10697 52333 10750 52379
rect 7750 52300 10750 52333
rect 11186 52379 14186 52392
rect 11186 52333 11239 52379
rect 14133 52333 14186 52379
rect 11186 52300 14186 52333
rect 878 49267 3878 49300
rect 878 49221 931 49267
rect 3825 49221 3878 49267
rect 878 49208 3878 49221
rect 4314 49267 7314 49300
rect 4314 49221 4367 49267
rect 7261 49221 7314 49267
rect 4314 49208 7314 49221
rect 7750 49267 10750 49300
rect 7750 49221 7803 49267
rect 10697 49221 10750 49267
rect 7750 49208 10750 49221
rect 11186 49267 14186 49300
rect 11186 49221 11239 49267
rect 14133 49221 14186 49267
rect 11186 49208 14186 49221
rect 878 48431 3878 48444
rect 878 48385 931 48431
rect 3825 48385 3878 48431
rect 878 48352 3878 48385
rect 4314 48431 7314 48444
rect 4314 48385 4367 48431
rect 7261 48385 7314 48431
rect 4314 48352 7314 48385
rect 7750 48431 10750 48444
rect 7750 48385 7803 48431
rect 10697 48385 10750 48431
rect 7750 48352 10750 48385
rect 11186 48431 14186 48444
rect 11186 48385 11239 48431
rect 14133 48385 14186 48431
rect 11186 48352 14186 48385
rect 878 45319 3878 45352
rect 878 45273 931 45319
rect 3825 45273 3878 45319
rect 878 45260 3878 45273
rect 4314 45319 7314 45352
rect 4314 45273 4367 45319
rect 7261 45273 7314 45319
rect 4314 45260 7314 45273
rect 7750 45319 10750 45352
rect 7750 45273 7803 45319
rect 10697 45273 10750 45319
rect 7750 45260 10750 45273
rect 11186 45319 14186 45352
rect 11186 45273 11239 45319
rect 14133 45273 14186 45319
rect 11186 45260 14186 45273
rect 878 44483 3878 44496
rect 878 44437 931 44483
rect 3825 44437 3878 44483
rect 878 44404 3878 44437
rect 4314 44483 7314 44496
rect 4314 44437 4367 44483
rect 7261 44437 7314 44483
rect 4314 44404 7314 44437
rect 7750 44483 10750 44496
rect 7750 44437 7803 44483
rect 10697 44437 10750 44483
rect 7750 44404 10750 44437
rect 11186 44483 14186 44496
rect 11186 44437 11239 44483
rect 14133 44437 14186 44483
rect 11186 44404 14186 44437
rect 878 41371 3878 41404
rect 878 41325 931 41371
rect 3825 41325 3878 41371
rect 878 41312 3878 41325
rect 4314 41371 7314 41404
rect 4314 41325 4367 41371
rect 7261 41325 7314 41371
rect 4314 41312 7314 41325
rect 7750 41371 10750 41404
rect 7750 41325 7803 41371
rect 10697 41325 10750 41371
rect 7750 41312 10750 41325
rect 11186 41371 14186 41404
rect 11186 41325 11239 41371
rect 14133 41325 14186 41371
rect 11186 41312 14186 41325
rect 878 40535 3878 40548
rect 878 40489 931 40535
rect 3825 40489 3878 40535
rect 878 40456 3878 40489
rect 4314 40535 7314 40548
rect 4314 40489 4367 40535
rect 7261 40489 7314 40535
rect 4314 40456 7314 40489
rect 7750 40535 10750 40548
rect 7750 40489 7803 40535
rect 10697 40489 10750 40535
rect 7750 40456 10750 40489
rect 11186 40535 14186 40548
rect 11186 40489 11239 40535
rect 14133 40489 14186 40535
rect 11186 40456 14186 40489
rect 878 37423 3878 37456
rect 878 37377 931 37423
rect 3825 37377 3878 37423
rect 878 37364 3878 37377
rect 4314 37423 7314 37456
rect 4314 37377 4367 37423
rect 7261 37377 7314 37423
rect 4314 37364 7314 37377
rect 7750 37423 10750 37456
rect 7750 37377 7803 37423
rect 10697 37377 10750 37423
rect 7750 37364 10750 37377
rect 11186 37423 14186 37456
rect 11186 37377 11239 37423
rect 14133 37377 14186 37423
rect 11186 37364 14186 37377
rect 878 36587 3878 36600
rect 878 36541 931 36587
rect 3825 36541 3878 36587
rect 878 36508 3878 36541
rect 4314 36587 7314 36600
rect 4314 36541 4367 36587
rect 7261 36541 7314 36587
rect 4314 36508 7314 36541
rect 7750 36587 10750 36600
rect 7750 36541 7803 36587
rect 10697 36541 10750 36587
rect 7750 36508 10750 36541
rect 11186 36587 14186 36600
rect 11186 36541 11239 36587
rect 14133 36541 14186 36587
rect 11186 36508 14186 36541
rect 878 33475 3878 33508
rect 878 33429 931 33475
rect 3825 33429 3878 33475
rect 878 33416 3878 33429
rect 4314 33475 7314 33508
rect 4314 33429 4367 33475
rect 7261 33429 7314 33475
rect 4314 33416 7314 33429
rect 7750 33475 10750 33508
rect 7750 33429 7803 33475
rect 10697 33429 10750 33475
rect 7750 33416 10750 33429
rect 11186 33475 14186 33508
rect 11186 33429 11239 33475
rect 14133 33429 14186 33475
rect 11186 33416 14186 33429
rect 878 32639 3878 32652
rect 878 32593 931 32639
rect 3825 32593 3878 32639
rect 878 32560 3878 32593
rect 4314 32639 7314 32652
rect 4314 32593 4367 32639
rect 7261 32593 7314 32639
rect 4314 32560 7314 32593
rect 7750 32639 10750 32652
rect 7750 32593 7803 32639
rect 10697 32593 10750 32639
rect 7750 32560 10750 32593
rect 11186 32639 14186 32652
rect 11186 32593 11239 32639
rect 14133 32593 14186 32639
rect 11186 32560 14186 32593
rect 878 29527 3878 29560
rect 878 29481 931 29527
rect 3825 29481 3878 29527
rect 878 29468 3878 29481
rect 4314 29527 7314 29560
rect 4314 29481 4367 29527
rect 7261 29481 7314 29527
rect 4314 29468 7314 29481
rect 7750 29527 10750 29560
rect 7750 29481 7803 29527
rect 10697 29481 10750 29527
rect 7750 29468 10750 29481
rect 11186 29527 14186 29560
rect 11186 29481 11239 29527
rect 14133 29481 14186 29527
rect 11186 29468 14186 29481
rect 878 28691 3878 28704
rect 878 28645 931 28691
rect 3825 28645 3878 28691
rect 878 28612 3878 28645
rect 4314 28691 7314 28704
rect 4314 28645 4367 28691
rect 7261 28645 7314 28691
rect 4314 28612 7314 28645
rect 7750 28691 10750 28704
rect 7750 28645 7803 28691
rect 10697 28645 10750 28691
rect 7750 28612 10750 28645
rect 11186 28691 14186 28704
rect 11186 28645 11239 28691
rect 14133 28645 14186 28691
rect 11186 28612 14186 28645
rect 878 25579 3878 25612
rect 878 25533 931 25579
rect 3825 25533 3878 25579
rect 878 25520 3878 25533
rect 4314 25579 7314 25612
rect 4314 25533 4367 25579
rect 7261 25533 7314 25579
rect 4314 25520 7314 25533
rect 7750 25579 10750 25612
rect 7750 25533 7803 25579
rect 10697 25533 10750 25579
rect 7750 25520 10750 25533
rect 11186 25579 14186 25612
rect 11186 25533 11239 25579
rect 14133 25533 14186 25579
rect 11186 25520 14186 25533
rect 878 24743 3878 24756
rect 878 24697 931 24743
rect 3825 24697 3878 24743
rect 878 24664 3878 24697
rect 4314 24743 7314 24756
rect 4314 24697 4367 24743
rect 7261 24697 7314 24743
rect 4314 24664 7314 24697
rect 7750 24743 10750 24756
rect 7750 24697 7803 24743
rect 10697 24697 10750 24743
rect 7750 24664 10750 24697
rect 11186 24743 14186 24756
rect 11186 24697 11239 24743
rect 14133 24697 14186 24743
rect 11186 24664 14186 24697
rect 878 21631 3878 21664
rect 878 21585 931 21631
rect 3825 21585 3878 21631
rect 878 21572 3878 21585
rect 4314 21631 7314 21664
rect 4314 21585 4367 21631
rect 7261 21585 7314 21631
rect 4314 21572 7314 21585
rect 7750 21631 10750 21664
rect 7750 21585 7803 21631
rect 10697 21585 10750 21631
rect 7750 21572 10750 21585
rect 11186 21631 14186 21664
rect 11186 21585 11239 21631
rect 14133 21585 14186 21631
rect 11186 21572 14186 21585
<< polycontact >>
rect 931 56281 3825 56327
rect 4367 56281 7261 56327
rect 7803 56281 10697 56327
rect 11239 56281 14133 56327
rect 931 53169 3825 53215
rect 4367 53169 7261 53215
rect 7803 53169 10697 53215
rect 11239 53169 14133 53215
rect 931 52333 3825 52379
rect 4367 52333 7261 52379
rect 7803 52333 10697 52379
rect 11239 52333 14133 52379
rect 931 49221 3825 49267
rect 4367 49221 7261 49267
rect 7803 49221 10697 49267
rect 11239 49221 14133 49267
rect 931 48385 3825 48431
rect 4367 48385 7261 48431
rect 7803 48385 10697 48431
rect 11239 48385 14133 48431
rect 931 45273 3825 45319
rect 4367 45273 7261 45319
rect 7803 45273 10697 45319
rect 11239 45273 14133 45319
rect 931 44437 3825 44483
rect 4367 44437 7261 44483
rect 7803 44437 10697 44483
rect 11239 44437 14133 44483
rect 931 41325 3825 41371
rect 4367 41325 7261 41371
rect 7803 41325 10697 41371
rect 11239 41325 14133 41371
rect 931 40489 3825 40535
rect 4367 40489 7261 40535
rect 7803 40489 10697 40535
rect 11239 40489 14133 40535
rect 931 37377 3825 37423
rect 4367 37377 7261 37423
rect 7803 37377 10697 37423
rect 11239 37377 14133 37423
rect 931 36541 3825 36587
rect 4367 36541 7261 36587
rect 7803 36541 10697 36587
rect 11239 36541 14133 36587
rect 931 33429 3825 33475
rect 4367 33429 7261 33475
rect 7803 33429 10697 33475
rect 11239 33429 14133 33475
rect 931 32593 3825 32639
rect 4367 32593 7261 32639
rect 7803 32593 10697 32639
rect 11239 32593 14133 32639
rect 931 29481 3825 29527
rect 4367 29481 7261 29527
rect 7803 29481 10697 29527
rect 11239 29481 14133 29527
rect 931 28645 3825 28691
rect 4367 28645 7261 28691
rect 7803 28645 10697 28691
rect 11239 28645 14133 28691
rect 931 25533 3825 25579
rect 4367 25533 7261 25579
rect 7803 25533 10697 25579
rect 11239 25533 14133 25579
rect 931 24697 3825 24743
rect 4367 24697 7261 24743
rect 7803 24697 10697 24743
rect 11239 24697 14133 24743
rect 931 21585 3825 21631
rect 4367 21585 7261 21631
rect 7803 21585 10697 21631
rect 11239 21585 14133 21631
<< mvndiode >>
rect 3532 19591 11532 19604
rect 3532 19545 3545 19591
rect 11519 19545 11532 19591
rect 3532 19463 11532 19545
rect 3532 19417 3545 19463
rect 11519 19417 11532 19463
rect 3532 19404 11532 19417
rect 3532 18719 11532 18732
rect 3532 18673 3545 18719
rect 11519 18673 11532 18719
rect 3532 18591 11532 18673
rect 3532 18545 3545 18591
rect 11519 18545 11532 18591
rect 3532 18532 11532 18545
rect 3532 17847 11532 17860
rect 3532 17801 3545 17847
rect 11519 17801 11532 17847
rect 3532 17719 11532 17801
rect 3532 17673 3545 17719
rect 11519 17673 11532 17719
rect 3532 17660 11532 17673
rect 3532 16975 11532 16988
rect 3532 16929 3545 16975
rect 11519 16929 11532 16975
rect 3532 16847 11532 16929
rect 3532 16801 3545 16847
rect 11519 16801 11532 16847
rect 3532 16788 11532 16801
<< mvndiodec >>
rect 3545 19545 11519 19591
rect 3545 19417 11519 19463
rect 3545 18673 11519 18719
rect 3545 18545 11519 18591
rect 3545 17801 11519 17847
rect 3545 17673 11519 17719
rect 3545 16929 11519 16975
rect 3545 16801 11519 16847
<< metal1 >>
rect 0 52271 122 57254
rect 0 52219 58 52271
rect 110 52219 122 52271
rect 0 52163 122 52219
rect 0 52111 58 52163
rect 110 52111 122 52163
rect 0 52055 122 52111
rect 0 52003 58 52055
rect 110 52003 122 52055
rect 0 51947 122 52003
rect 0 51895 58 51947
rect 110 51895 122 51947
rect 0 51839 122 51895
rect 0 51787 58 51839
rect 110 51787 122 51839
rect 0 51731 122 51787
rect 0 51679 58 51731
rect 110 51679 122 51731
rect 0 51623 122 51679
rect 0 51571 58 51623
rect 110 51571 122 51623
rect 0 51515 122 51571
rect 0 51463 58 51515
rect 110 51463 122 51515
rect 0 51407 122 51463
rect 0 51355 58 51407
rect 110 51355 122 51407
rect 0 51299 122 51355
rect 0 51247 58 51299
rect 110 51247 122 51299
rect 0 51191 122 51247
rect 0 51139 58 51191
rect 110 51139 122 51191
rect 0 51083 122 51139
rect 0 51031 58 51083
rect 110 51031 122 51083
rect 0 50975 122 51031
rect 0 50923 58 50975
rect 110 50923 122 50975
rect 0 37871 122 50923
rect 0 37819 58 37871
rect 110 37819 122 37871
rect 0 37763 122 37819
rect 0 37711 58 37763
rect 110 37711 122 37763
rect 0 37655 122 37711
rect 0 37603 58 37655
rect 110 37603 122 37655
rect 0 37547 122 37603
rect 0 37495 58 37547
rect 110 37495 122 37547
rect 0 37439 122 37495
rect 0 37387 58 37439
rect 110 37387 122 37439
rect 0 37331 122 37387
rect 0 37279 58 37331
rect 110 37279 122 37331
rect 0 37223 122 37279
rect 0 37171 58 37223
rect 110 37171 122 37223
rect 0 37115 122 37171
rect 0 37063 58 37115
rect 110 37063 122 37115
rect 0 37007 122 37063
rect 0 36955 58 37007
rect 110 36955 122 37007
rect 0 36899 122 36955
rect 0 36847 58 36899
rect 110 36847 122 36899
rect 0 36791 122 36847
rect 0 36739 58 36791
rect 110 36739 122 36791
rect 0 36683 122 36739
rect 0 36631 58 36683
rect 110 36631 122 36683
rect 0 36575 122 36631
rect 0 36523 58 36575
rect 110 36523 122 36575
rect 0 20368 122 36523
rect 388 56745 14676 56756
rect 388 21167 399 56745
rect 445 56711 553 56745
rect 14511 56711 14619 56745
rect 496 56659 552 56711
rect 604 56659 660 56699
rect 712 56659 1408 56699
rect 1460 56659 1516 56699
rect 1568 56659 1624 56699
rect 1676 56659 1732 56699
rect 1784 56659 1840 56699
rect 1892 56659 2544 56699
rect 2596 56659 2652 56699
rect 2704 56659 2760 56699
rect 2812 56659 2868 56699
rect 2920 56659 2976 56699
rect 3028 56659 4816 56699
rect 4868 56659 4924 56699
rect 4976 56659 5032 56699
rect 5084 56659 5140 56699
rect 5192 56659 5248 56699
rect 5300 56659 7101 56699
rect 7153 56659 7209 56699
rect 7261 56659 7317 56699
rect 7369 56659 7425 56699
rect 7477 56659 7587 56699
rect 7639 56659 7695 56699
rect 7747 56659 7803 56699
rect 7855 56659 7911 56699
rect 7963 56659 9764 56699
rect 9816 56659 9872 56699
rect 9924 56659 9980 56699
rect 10032 56659 10088 56699
rect 10140 56659 10196 56699
rect 10248 56659 12036 56699
rect 12088 56659 12144 56699
rect 12196 56659 12252 56699
rect 12304 56659 12360 56699
rect 12412 56659 12468 56699
rect 12520 56659 13172 56699
rect 13224 56659 13280 56699
rect 13332 56659 13388 56699
rect 13440 56659 13496 56699
rect 13548 56659 13604 56699
rect 13656 56659 14352 56699
rect 14404 56659 14460 56699
rect 14512 56659 14568 56711
rect 445 56603 14619 56659
rect 496 56551 552 56603
rect 604 56551 660 56603
rect 712 56551 1408 56603
rect 1460 56551 1516 56603
rect 1568 56551 1624 56603
rect 1676 56551 1732 56603
rect 1784 56551 1840 56603
rect 1892 56551 2544 56603
rect 2596 56551 2652 56603
rect 2704 56551 2760 56603
rect 2812 56551 2868 56603
rect 2920 56551 2976 56603
rect 3028 56551 4816 56603
rect 4868 56551 4924 56603
rect 4976 56551 5032 56603
rect 5084 56551 5140 56603
rect 5192 56551 5248 56603
rect 5300 56551 7101 56603
rect 7153 56551 7209 56603
rect 7261 56551 7317 56603
rect 7369 56551 7425 56603
rect 7477 56551 7587 56603
rect 7639 56551 7695 56603
rect 7747 56551 7803 56603
rect 7855 56551 7911 56603
rect 7963 56551 9764 56603
rect 9816 56551 9872 56603
rect 9924 56551 9980 56603
rect 10032 56551 10088 56603
rect 10140 56551 10196 56603
rect 10248 56551 12036 56603
rect 12088 56551 12144 56603
rect 12196 56551 12252 56603
rect 12304 56551 12360 56603
rect 12412 56551 12468 56603
rect 12520 56551 13172 56603
rect 13224 56551 13280 56603
rect 13332 56551 13388 56603
rect 13440 56551 13496 56603
rect 13548 56551 13604 56603
rect 13656 56551 14352 56603
rect 14404 56551 14460 56603
rect 14512 56551 14568 56603
rect 445 56495 14619 56551
rect 496 56443 552 56495
rect 604 56443 660 56495
rect 712 56443 1408 56495
rect 1460 56443 1516 56495
rect 1568 56443 1624 56495
rect 1676 56443 1732 56495
rect 1784 56443 1840 56495
rect 1892 56443 2544 56495
rect 2596 56443 2652 56495
rect 2704 56443 2760 56495
rect 2812 56443 2868 56495
rect 2920 56443 2976 56495
rect 3028 56443 4816 56495
rect 4868 56443 4924 56495
rect 4976 56443 5032 56495
rect 5084 56443 5140 56495
rect 5192 56443 5248 56495
rect 5300 56443 7101 56495
rect 7153 56443 7209 56495
rect 7261 56443 7317 56495
rect 7369 56443 7425 56495
rect 7477 56443 7587 56495
rect 7639 56443 7695 56495
rect 7747 56443 7803 56495
rect 7855 56443 7911 56495
rect 7963 56443 9764 56495
rect 9816 56443 9872 56495
rect 9924 56443 9980 56495
rect 10032 56443 10088 56495
rect 10140 56443 10196 56495
rect 10248 56443 12036 56495
rect 12088 56443 12144 56495
rect 12196 56443 12252 56495
rect 12304 56443 12360 56495
rect 12412 56443 12468 56495
rect 12520 56443 13172 56495
rect 13224 56443 13280 56495
rect 13332 56443 13388 56495
rect 13440 56443 13496 56495
rect 13548 56443 13604 56495
rect 13656 56443 14352 56495
rect 14404 56443 14460 56495
rect 14512 56443 14568 56495
rect 445 56398 14619 56443
rect 445 53098 456 56398
rect 920 56327 3836 56338
rect 920 56281 931 56327
rect 3825 56281 3836 56327
rect 920 56272 978 56281
rect 1030 56272 1102 56281
rect 1154 56272 1226 56281
rect 1278 56272 3729 56281
rect 920 56270 3729 56272
rect 660 56211 860 56248
rect 660 53285 803 56211
rect 849 53285 860 56211
rect 660 53098 860 53285
rect 920 56200 1920 56270
rect 920 56148 978 56200
rect 1030 56148 1102 56200
rect 1154 56148 1226 56200
rect 1278 56148 1920 56200
rect 920 56076 1920 56148
rect 920 56024 978 56076
rect 1030 56024 1102 56076
rect 1154 56024 1226 56076
rect 1278 56024 1920 56076
rect 920 55952 1920 56024
rect 920 55900 978 55952
rect 1030 55900 1102 55952
rect 1154 55900 1226 55952
rect 1278 55900 1920 55952
rect 920 55828 1920 55900
rect 920 55776 978 55828
rect 1030 55776 1102 55828
rect 1154 55776 1226 55828
rect 1278 55776 1920 55828
rect 920 55704 1920 55776
rect 920 55652 978 55704
rect 1030 55652 1102 55704
rect 1154 55652 1226 55704
rect 1278 55652 1920 55704
rect 920 55580 1920 55652
rect 920 55528 978 55580
rect 1030 55528 1102 55580
rect 1154 55528 1226 55580
rect 1278 55528 1920 55580
rect 920 55456 1920 55528
rect 920 55404 978 55456
rect 1030 55404 1102 55456
rect 1154 55404 1226 55456
rect 1278 55404 1920 55456
rect 920 55332 1920 55404
rect 920 55280 978 55332
rect 1030 55280 1102 55332
rect 1154 55280 1226 55332
rect 1278 55280 1920 55332
rect 920 55208 1920 55280
rect 920 55156 978 55208
rect 1030 55156 1102 55208
rect 1154 55156 1226 55208
rect 1278 55156 1920 55208
rect 920 55084 1920 55156
rect 920 55032 978 55084
rect 1030 55032 1102 55084
rect 1154 55032 1226 55084
rect 1278 55032 1920 55084
rect 920 54960 1920 55032
rect 920 54908 978 54960
rect 1030 54908 1102 54960
rect 1154 54908 1226 54960
rect 1278 54908 1920 54960
rect 920 54836 1920 54908
rect 920 54784 978 54836
rect 1030 54784 1102 54836
rect 1154 54784 1226 54836
rect 1278 54784 1920 54836
rect 920 54712 1920 54784
rect 920 54660 978 54712
rect 1030 54660 1102 54712
rect 1154 54660 1226 54712
rect 1278 54660 1920 54712
rect 920 54588 1920 54660
rect 920 54536 978 54588
rect 1030 54536 1102 54588
rect 1154 54536 1226 54588
rect 1278 54536 1920 54588
rect 920 54464 1920 54536
rect 920 54412 978 54464
rect 1030 54412 1102 54464
rect 1154 54412 1226 54464
rect 1278 54412 1920 54464
rect 920 54340 1920 54412
rect 920 54288 978 54340
rect 1030 54288 1102 54340
rect 1154 54288 1226 54340
rect 1278 54288 1920 54340
rect 920 54216 1920 54288
rect 920 54164 978 54216
rect 1030 54164 1102 54216
rect 1154 54164 1226 54216
rect 1278 54164 1920 54216
rect 920 54092 1920 54164
rect 920 54040 978 54092
rect 1030 54040 1102 54092
rect 1154 54040 1226 54092
rect 1278 54040 1920 54092
rect 920 53968 1920 54040
rect 920 53916 978 53968
rect 1030 53916 1102 53968
rect 1154 53916 1226 53968
rect 1278 53916 1920 53968
rect 920 53844 1920 53916
rect 920 53792 978 53844
rect 1030 53792 1102 53844
rect 1154 53792 1226 53844
rect 1278 53792 1920 53844
rect 920 53720 1920 53792
rect 920 53668 978 53720
rect 1030 53668 1102 53720
rect 1154 53668 1226 53720
rect 1278 53668 1920 53720
rect 920 53596 1920 53668
rect 920 53544 978 53596
rect 1030 53544 1102 53596
rect 1154 53544 1226 53596
rect 1278 53544 1920 53596
rect 920 53472 1920 53544
rect 920 53420 978 53472
rect 1030 53420 1102 53472
rect 1154 53420 1226 53472
rect 1278 53420 1920 53472
rect 920 53348 1920 53420
rect 920 53296 978 53348
rect 1030 53296 1102 53348
rect 1154 53296 1226 53348
rect 1278 53296 1920 53348
rect 920 53226 1920 53296
rect 2836 56234 3729 56270
rect 3781 56234 3836 56281
rect 4356 56327 7272 56338
rect 4356 56281 4367 56327
rect 7261 56281 7272 56327
rect 4356 56270 6335 56281
rect 2836 56178 3836 56234
rect 2836 56126 3729 56178
rect 3781 56126 3836 56178
rect 2836 56070 3836 56126
rect 2836 56018 3729 56070
rect 3781 56018 3836 56070
rect 2836 55962 3836 56018
rect 2836 55910 3729 55962
rect 3781 55910 3836 55962
rect 2836 55854 3836 55910
rect 2836 55802 3729 55854
rect 3781 55802 3836 55854
rect 2836 55746 3836 55802
rect 2836 55694 3729 55746
rect 3781 55694 3836 55746
rect 2836 55638 3836 55694
rect 2836 55586 3729 55638
rect 3781 55586 3836 55638
rect 2836 55530 3836 55586
rect 2836 55478 3729 55530
rect 3781 55478 3836 55530
rect 2836 55422 3836 55478
rect 2836 55370 3729 55422
rect 3781 55370 3836 55422
rect 2836 55314 3836 55370
rect 2836 55262 3729 55314
rect 3781 55262 3836 55314
rect 2836 55206 3836 55262
rect 2836 55154 3729 55206
rect 3781 55154 3836 55206
rect 2836 55098 3836 55154
rect 2836 55046 3729 55098
rect 3781 55046 3836 55098
rect 2836 54990 3836 55046
rect 2836 54938 3729 54990
rect 3781 54938 3836 54990
rect 2836 54882 3836 54938
rect 2836 54830 3729 54882
rect 3781 54830 3836 54882
rect 2836 54774 3836 54830
rect 2836 54722 3729 54774
rect 3781 54722 3836 54774
rect 2836 54666 3836 54722
rect 2836 54614 3729 54666
rect 3781 54614 3836 54666
rect 2836 54558 3836 54614
rect 2836 54506 3729 54558
rect 3781 54506 3836 54558
rect 2836 54450 3836 54506
rect 2836 54398 3729 54450
rect 3781 54398 3836 54450
rect 2836 54342 3836 54398
rect 2836 54290 3729 54342
rect 3781 54290 3836 54342
rect 2836 54234 3836 54290
rect 2836 54182 3729 54234
rect 3781 54182 3836 54234
rect 2836 54126 3836 54182
rect 2836 54074 3729 54126
rect 3781 54074 3836 54126
rect 2836 54018 3836 54074
rect 2836 53966 3729 54018
rect 3781 53966 3836 54018
rect 2836 53910 3836 53966
rect 2836 53858 3729 53910
rect 3781 53858 3836 53910
rect 2836 53802 3836 53858
rect 2836 53750 3729 53802
rect 3781 53750 3836 53802
rect 2836 53694 3836 53750
rect 2836 53642 3729 53694
rect 3781 53642 3836 53694
rect 2836 53586 3836 53642
rect 2836 53534 3729 53586
rect 3781 53534 3836 53586
rect 2836 53478 3836 53534
rect 2836 53426 3729 53478
rect 3781 53426 3836 53478
rect 2836 53370 3836 53426
rect 2836 53318 3729 53370
rect 3781 53318 3836 53370
rect 2836 53262 3836 53318
rect 2836 53226 3729 53262
rect 920 53224 3729 53226
rect 920 53215 978 53224
rect 1030 53215 1102 53224
rect 1154 53215 1226 53224
rect 1278 53215 3729 53224
rect 3781 53215 3836 53262
rect 920 53169 931 53215
rect 3825 53169 3836 53215
rect 920 53158 3836 53169
rect 3896 56211 4296 56248
rect 3896 53285 3907 56211
rect 3953 53285 4239 56211
rect 4285 53285 4296 56211
rect 3896 53098 4296 53285
rect 4356 53226 5356 56270
rect 6272 56234 6335 56270
rect 6387 56234 7272 56281
rect 7792 56327 10708 56338
rect 7792 56281 7803 56327
rect 10697 56281 10708 56327
rect 6272 56178 7272 56234
rect 6272 56126 6335 56178
rect 6387 56126 7272 56178
rect 6272 56070 7272 56126
rect 6272 56018 6335 56070
rect 6387 56018 7272 56070
rect 6272 55962 7272 56018
rect 6272 55910 6335 55962
rect 6387 55910 7272 55962
rect 6272 55854 7272 55910
rect 6272 55802 6335 55854
rect 6387 55802 7272 55854
rect 6272 55746 7272 55802
rect 6272 55694 6335 55746
rect 6387 55694 7272 55746
rect 6272 55638 7272 55694
rect 6272 55586 6335 55638
rect 6387 55586 7272 55638
rect 6272 55530 7272 55586
rect 6272 55478 6335 55530
rect 6387 55478 7272 55530
rect 6272 55422 7272 55478
rect 6272 55370 6335 55422
rect 6387 55370 7272 55422
rect 6272 55314 7272 55370
rect 6272 55262 6335 55314
rect 6387 55262 7272 55314
rect 6272 55206 7272 55262
rect 6272 55154 6335 55206
rect 6387 55154 7272 55206
rect 6272 55098 7272 55154
rect 6272 55046 6335 55098
rect 6387 55046 7272 55098
rect 6272 54990 7272 55046
rect 6272 54938 6335 54990
rect 6387 54938 7272 54990
rect 6272 54882 7272 54938
rect 6272 54830 6335 54882
rect 6387 54830 7272 54882
rect 6272 54774 7272 54830
rect 6272 54722 6335 54774
rect 6387 54722 7272 54774
rect 6272 54666 7272 54722
rect 6272 54614 6335 54666
rect 6387 54614 7272 54666
rect 6272 54558 7272 54614
rect 6272 54506 6335 54558
rect 6387 54506 7272 54558
rect 6272 54450 7272 54506
rect 6272 54398 6335 54450
rect 6387 54398 7272 54450
rect 6272 54342 7272 54398
rect 6272 54290 6335 54342
rect 6387 54290 7272 54342
rect 6272 54234 7272 54290
rect 6272 54182 6335 54234
rect 6387 54182 7272 54234
rect 6272 54126 7272 54182
rect 6272 54074 6335 54126
rect 6387 54074 7272 54126
rect 6272 54018 7272 54074
rect 6272 53966 6335 54018
rect 6387 53966 7272 54018
rect 6272 53910 7272 53966
rect 6272 53858 6335 53910
rect 6387 53858 7272 53910
rect 6272 53802 7272 53858
rect 6272 53750 6335 53802
rect 6387 53750 7272 53802
rect 6272 53694 7272 53750
rect 6272 53642 6335 53694
rect 6387 53642 7272 53694
rect 6272 53586 7272 53642
rect 6272 53534 6335 53586
rect 6387 53534 7272 53586
rect 6272 53478 7272 53534
rect 6272 53426 6335 53478
rect 6387 53426 7272 53478
rect 6272 53370 7272 53426
rect 6272 53318 6335 53370
rect 6387 53318 7272 53370
rect 6272 53262 7272 53318
rect 6272 53226 6335 53262
rect 4356 53215 6335 53226
rect 6387 53215 7272 53262
rect 4356 53169 4367 53215
rect 7261 53169 7272 53215
rect 4356 53158 7272 53169
rect 7332 56232 7732 56248
rect 7332 56211 7388 56232
rect 7332 53285 7343 56211
rect 7440 56180 7624 56232
rect 7676 56211 7732 56232
rect 7389 56124 7675 56180
rect 7440 56072 7624 56124
rect 7389 56016 7675 56072
rect 7440 55964 7624 56016
rect 7389 55908 7675 55964
rect 7440 55856 7624 55908
rect 7389 55800 7675 55856
rect 7440 55748 7624 55800
rect 7389 55692 7675 55748
rect 7440 55640 7624 55692
rect 7389 55584 7675 55640
rect 7440 55532 7624 55584
rect 7389 55476 7675 55532
rect 7440 55424 7624 55476
rect 7389 55368 7675 55424
rect 7440 55316 7624 55368
rect 7389 55260 7675 55316
rect 7440 55208 7624 55260
rect 7389 55152 7675 55208
rect 7440 55100 7624 55152
rect 7389 55044 7675 55100
rect 7440 54992 7624 55044
rect 7389 54936 7675 54992
rect 7440 54884 7624 54936
rect 7389 54828 7675 54884
rect 7440 54776 7624 54828
rect 7389 54720 7675 54776
rect 7440 54668 7624 54720
rect 7389 54612 7675 54668
rect 7440 54560 7624 54612
rect 7389 54504 7675 54560
rect 7440 54452 7624 54504
rect 7389 54396 7675 54452
rect 7440 54344 7624 54396
rect 7389 54288 7675 54344
rect 7440 54236 7624 54288
rect 7389 54180 7675 54236
rect 7440 54128 7624 54180
rect 7389 54072 7675 54128
rect 7440 54020 7624 54072
rect 7389 53964 7675 54020
rect 7440 53912 7624 53964
rect 7389 53856 7675 53912
rect 7440 53804 7624 53856
rect 7389 53748 7675 53804
rect 7440 53696 7624 53748
rect 7389 53640 7675 53696
rect 7440 53588 7624 53640
rect 7389 53532 7675 53588
rect 7440 53480 7624 53532
rect 7389 53424 7675 53480
rect 7440 53372 7624 53424
rect 7389 53316 7675 53372
rect 7332 53264 7388 53285
rect 7440 53264 7624 53316
rect 7721 53285 7732 56211
rect 7676 53264 7732 53285
rect 7332 53098 7732 53264
rect 7792 56234 8677 56281
rect 8729 56270 10708 56281
rect 8729 56234 8792 56270
rect 7792 56178 8792 56234
rect 7792 56126 8677 56178
rect 8729 56126 8792 56178
rect 7792 56070 8792 56126
rect 7792 56018 8677 56070
rect 8729 56018 8792 56070
rect 7792 55962 8792 56018
rect 7792 55910 8677 55962
rect 8729 55910 8792 55962
rect 7792 55854 8792 55910
rect 7792 55802 8677 55854
rect 8729 55802 8792 55854
rect 7792 55746 8792 55802
rect 7792 55694 8677 55746
rect 8729 55694 8792 55746
rect 7792 55638 8792 55694
rect 7792 55586 8677 55638
rect 8729 55586 8792 55638
rect 7792 55530 8792 55586
rect 7792 55478 8677 55530
rect 8729 55478 8792 55530
rect 7792 55422 8792 55478
rect 7792 55370 8677 55422
rect 8729 55370 8792 55422
rect 7792 55314 8792 55370
rect 7792 55262 8677 55314
rect 8729 55262 8792 55314
rect 7792 55206 8792 55262
rect 7792 55154 8677 55206
rect 8729 55154 8792 55206
rect 7792 55098 8792 55154
rect 7792 55046 8677 55098
rect 8729 55046 8792 55098
rect 7792 54990 8792 55046
rect 7792 54938 8677 54990
rect 8729 54938 8792 54990
rect 7792 54882 8792 54938
rect 7792 54830 8677 54882
rect 8729 54830 8792 54882
rect 7792 54774 8792 54830
rect 7792 54722 8677 54774
rect 8729 54722 8792 54774
rect 7792 54666 8792 54722
rect 7792 54614 8677 54666
rect 8729 54614 8792 54666
rect 7792 54558 8792 54614
rect 7792 54506 8677 54558
rect 8729 54506 8792 54558
rect 7792 54450 8792 54506
rect 7792 54398 8677 54450
rect 8729 54398 8792 54450
rect 7792 54342 8792 54398
rect 7792 54290 8677 54342
rect 8729 54290 8792 54342
rect 7792 54234 8792 54290
rect 7792 54182 8677 54234
rect 8729 54182 8792 54234
rect 7792 54126 8792 54182
rect 7792 54074 8677 54126
rect 8729 54074 8792 54126
rect 7792 54018 8792 54074
rect 7792 53966 8677 54018
rect 8729 53966 8792 54018
rect 7792 53910 8792 53966
rect 7792 53858 8677 53910
rect 8729 53858 8792 53910
rect 7792 53802 8792 53858
rect 7792 53750 8677 53802
rect 8729 53750 8792 53802
rect 7792 53694 8792 53750
rect 7792 53642 8677 53694
rect 8729 53642 8792 53694
rect 7792 53586 8792 53642
rect 7792 53534 8677 53586
rect 8729 53534 8792 53586
rect 7792 53478 8792 53534
rect 7792 53426 8677 53478
rect 8729 53426 8792 53478
rect 7792 53370 8792 53426
rect 7792 53318 8677 53370
rect 8729 53318 8792 53370
rect 7792 53262 8792 53318
rect 7792 53215 8677 53262
rect 8729 53226 8792 53262
rect 9708 53226 10708 56270
rect 11228 56327 14144 56338
rect 11228 56281 11239 56327
rect 14133 56281 14144 56327
rect 8729 53215 10708 53226
rect 7792 53169 7803 53215
rect 10697 53169 10708 53215
rect 7792 53158 10708 53169
rect 10768 56211 11168 56248
rect 10768 53285 10779 56211
rect 10825 53285 11111 56211
rect 11157 53285 11168 56211
rect 10768 53098 11168 53285
rect 11228 56234 11283 56281
rect 11335 56272 13786 56281
rect 13838 56272 13910 56281
rect 13962 56272 14034 56281
rect 14086 56272 14144 56281
rect 11335 56270 14144 56272
rect 11335 56234 12228 56270
rect 11228 56178 12228 56234
rect 11228 56126 11283 56178
rect 11335 56126 12228 56178
rect 11228 56070 12228 56126
rect 11228 56018 11283 56070
rect 11335 56018 12228 56070
rect 11228 55962 12228 56018
rect 11228 55910 11283 55962
rect 11335 55910 12228 55962
rect 11228 55854 12228 55910
rect 11228 55802 11283 55854
rect 11335 55802 12228 55854
rect 11228 55746 12228 55802
rect 11228 55694 11283 55746
rect 11335 55694 12228 55746
rect 11228 55638 12228 55694
rect 11228 55586 11283 55638
rect 11335 55586 12228 55638
rect 11228 55530 12228 55586
rect 11228 55478 11283 55530
rect 11335 55478 12228 55530
rect 11228 55422 12228 55478
rect 11228 55370 11283 55422
rect 11335 55370 12228 55422
rect 11228 55314 12228 55370
rect 11228 55262 11283 55314
rect 11335 55262 12228 55314
rect 11228 55206 12228 55262
rect 11228 55154 11283 55206
rect 11335 55154 12228 55206
rect 11228 55098 12228 55154
rect 11228 55046 11283 55098
rect 11335 55046 12228 55098
rect 11228 54990 12228 55046
rect 11228 54938 11283 54990
rect 11335 54938 12228 54990
rect 11228 54882 12228 54938
rect 11228 54830 11283 54882
rect 11335 54830 12228 54882
rect 11228 54774 12228 54830
rect 11228 54722 11283 54774
rect 11335 54722 12228 54774
rect 11228 54666 12228 54722
rect 11228 54614 11283 54666
rect 11335 54614 12228 54666
rect 11228 54558 12228 54614
rect 11228 54506 11283 54558
rect 11335 54506 12228 54558
rect 11228 54450 12228 54506
rect 11228 54398 11283 54450
rect 11335 54398 12228 54450
rect 11228 54342 12228 54398
rect 11228 54290 11283 54342
rect 11335 54290 12228 54342
rect 11228 54234 12228 54290
rect 11228 54182 11283 54234
rect 11335 54182 12228 54234
rect 11228 54126 12228 54182
rect 11228 54074 11283 54126
rect 11335 54074 12228 54126
rect 11228 54018 12228 54074
rect 11228 53966 11283 54018
rect 11335 53966 12228 54018
rect 11228 53910 12228 53966
rect 11228 53858 11283 53910
rect 11335 53858 12228 53910
rect 11228 53802 12228 53858
rect 11228 53750 11283 53802
rect 11335 53750 12228 53802
rect 11228 53694 12228 53750
rect 11228 53642 11283 53694
rect 11335 53642 12228 53694
rect 11228 53586 12228 53642
rect 11228 53534 11283 53586
rect 11335 53534 12228 53586
rect 11228 53478 12228 53534
rect 11228 53426 11283 53478
rect 11335 53426 12228 53478
rect 11228 53370 12228 53426
rect 11228 53318 11283 53370
rect 11335 53318 12228 53370
rect 11228 53262 12228 53318
rect 11228 53215 11283 53262
rect 11335 53226 12228 53262
rect 13144 56200 14144 56270
rect 13144 56148 13786 56200
rect 13838 56148 13910 56200
rect 13962 56148 14034 56200
rect 14086 56148 14144 56200
rect 13144 56076 14144 56148
rect 13144 56024 13786 56076
rect 13838 56024 13910 56076
rect 13962 56024 14034 56076
rect 14086 56024 14144 56076
rect 13144 55952 14144 56024
rect 13144 55900 13786 55952
rect 13838 55900 13910 55952
rect 13962 55900 14034 55952
rect 14086 55900 14144 55952
rect 13144 55828 14144 55900
rect 13144 55776 13786 55828
rect 13838 55776 13910 55828
rect 13962 55776 14034 55828
rect 14086 55776 14144 55828
rect 13144 55704 14144 55776
rect 13144 55652 13786 55704
rect 13838 55652 13910 55704
rect 13962 55652 14034 55704
rect 14086 55652 14144 55704
rect 13144 55580 14144 55652
rect 13144 55528 13786 55580
rect 13838 55528 13910 55580
rect 13962 55528 14034 55580
rect 14086 55528 14144 55580
rect 13144 55456 14144 55528
rect 13144 55404 13786 55456
rect 13838 55404 13910 55456
rect 13962 55404 14034 55456
rect 14086 55404 14144 55456
rect 13144 55332 14144 55404
rect 13144 55280 13786 55332
rect 13838 55280 13910 55332
rect 13962 55280 14034 55332
rect 14086 55280 14144 55332
rect 13144 55208 14144 55280
rect 13144 55156 13786 55208
rect 13838 55156 13910 55208
rect 13962 55156 14034 55208
rect 14086 55156 14144 55208
rect 13144 55084 14144 55156
rect 13144 55032 13786 55084
rect 13838 55032 13910 55084
rect 13962 55032 14034 55084
rect 14086 55032 14144 55084
rect 13144 54960 14144 55032
rect 13144 54908 13786 54960
rect 13838 54908 13910 54960
rect 13962 54908 14034 54960
rect 14086 54908 14144 54960
rect 13144 54836 14144 54908
rect 13144 54784 13786 54836
rect 13838 54784 13910 54836
rect 13962 54784 14034 54836
rect 14086 54784 14144 54836
rect 13144 54712 14144 54784
rect 13144 54660 13786 54712
rect 13838 54660 13910 54712
rect 13962 54660 14034 54712
rect 14086 54660 14144 54712
rect 13144 54588 14144 54660
rect 13144 54536 13786 54588
rect 13838 54536 13910 54588
rect 13962 54536 14034 54588
rect 14086 54536 14144 54588
rect 13144 54464 14144 54536
rect 13144 54412 13786 54464
rect 13838 54412 13910 54464
rect 13962 54412 14034 54464
rect 14086 54412 14144 54464
rect 13144 54340 14144 54412
rect 13144 54288 13786 54340
rect 13838 54288 13910 54340
rect 13962 54288 14034 54340
rect 14086 54288 14144 54340
rect 13144 54216 14144 54288
rect 13144 54164 13786 54216
rect 13838 54164 13910 54216
rect 13962 54164 14034 54216
rect 14086 54164 14144 54216
rect 13144 54092 14144 54164
rect 13144 54040 13786 54092
rect 13838 54040 13910 54092
rect 13962 54040 14034 54092
rect 14086 54040 14144 54092
rect 13144 53968 14144 54040
rect 13144 53916 13786 53968
rect 13838 53916 13910 53968
rect 13962 53916 14034 53968
rect 14086 53916 14144 53968
rect 13144 53844 14144 53916
rect 13144 53792 13786 53844
rect 13838 53792 13910 53844
rect 13962 53792 14034 53844
rect 14086 53792 14144 53844
rect 13144 53720 14144 53792
rect 13144 53668 13786 53720
rect 13838 53668 13910 53720
rect 13962 53668 14034 53720
rect 14086 53668 14144 53720
rect 13144 53596 14144 53668
rect 13144 53544 13786 53596
rect 13838 53544 13910 53596
rect 13962 53544 14034 53596
rect 14086 53544 14144 53596
rect 13144 53472 14144 53544
rect 13144 53420 13786 53472
rect 13838 53420 13910 53472
rect 13962 53420 14034 53472
rect 14086 53420 14144 53472
rect 13144 53348 14144 53420
rect 13144 53296 13786 53348
rect 13838 53296 13910 53348
rect 13962 53296 14034 53348
rect 14086 53296 14144 53348
rect 13144 53226 14144 53296
rect 11335 53224 14144 53226
rect 11335 53215 13786 53224
rect 13838 53215 13910 53224
rect 13962 53215 14034 53224
rect 14086 53215 14144 53224
rect 11228 53169 11239 53215
rect 14133 53169 14144 53215
rect 11228 53158 14144 53169
rect 14204 56211 14404 56248
rect 14204 53285 14215 56211
rect 14261 53285 14404 56211
rect 14204 53098 14404 53285
rect 14608 53098 14619 56398
rect 445 53048 14619 53098
rect 445 53016 1438 53048
rect 496 52964 552 53016
rect 604 52964 660 53016
rect 712 52996 1438 53016
rect 1490 52996 1562 53048
rect 1614 52996 1686 53048
rect 1738 52996 1810 53048
rect 1862 52996 2574 53048
rect 2626 52996 2698 53048
rect 2750 52996 2822 53048
rect 2874 52996 2946 53048
rect 2998 52996 4846 53048
rect 4898 52996 4970 53048
rect 5022 52996 5094 53048
rect 5146 52996 5218 53048
rect 5270 52996 7139 53048
rect 7191 52996 7263 53048
rect 7315 52996 7387 53048
rect 7439 52996 7625 53048
rect 7677 52996 7749 53048
rect 7801 52996 7873 53048
rect 7925 52996 9794 53048
rect 9846 52996 9918 53048
rect 9970 52996 10042 53048
rect 10094 52996 10166 53048
rect 10218 52996 12066 53048
rect 12118 52996 12190 53048
rect 12242 52996 12314 53048
rect 12366 52996 12438 53048
rect 12490 52996 13202 53048
rect 13254 52996 13326 53048
rect 13378 52996 13450 53048
rect 13502 52996 13574 53048
rect 13626 53016 14619 53048
rect 13626 52996 14352 53016
rect 712 52964 14352 52996
rect 14404 52964 14460 53016
rect 14512 52964 14568 53016
rect 445 52924 14619 52964
rect 445 52908 1438 52924
rect 496 52856 552 52908
rect 604 52856 660 52908
rect 712 52872 1438 52908
rect 1490 52872 1562 52924
rect 1614 52872 1686 52924
rect 1738 52872 1810 52924
rect 1862 52872 2574 52924
rect 2626 52872 2698 52924
rect 2750 52872 2822 52924
rect 2874 52872 2946 52924
rect 2998 52872 4846 52924
rect 4898 52872 4970 52924
rect 5022 52872 5094 52924
rect 5146 52872 5218 52924
rect 5270 52872 7139 52924
rect 7191 52872 7263 52924
rect 7315 52872 7387 52924
rect 7439 52872 7625 52924
rect 7677 52872 7749 52924
rect 7801 52872 7873 52924
rect 7925 52872 9794 52924
rect 9846 52872 9918 52924
rect 9970 52872 10042 52924
rect 10094 52872 10166 52924
rect 10218 52872 12066 52924
rect 12118 52872 12190 52924
rect 12242 52872 12314 52924
rect 12366 52872 12438 52924
rect 12490 52872 13202 52924
rect 13254 52872 13326 52924
rect 13378 52872 13450 52924
rect 13502 52872 13574 52924
rect 13626 52908 14619 52924
rect 13626 52872 14352 52908
rect 712 52856 14352 52872
rect 14404 52856 14460 52908
rect 14512 52856 14568 52908
rect 445 52800 14619 52856
rect 496 52748 552 52800
rect 604 52797 660 52800
rect 712 52797 1438 52800
rect 1490 52797 1562 52800
rect 1614 52797 1686 52800
rect 1738 52797 1810 52800
rect 1862 52797 2574 52800
rect 2626 52797 2698 52800
rect 2750 52797 2822 52800
rect 2874 52797 2946 52800
rect 2998 52797 4846 52800
rect 4898 52797 4970 52800
rect 5022 52797 5094 52800
rect 5146 52797 5218 52800
rect 5270 52797 7139 52800
rect 7191 52797 7263 52800
rect 7315 52797 7387 52800
rect 7439 52797 7625 52800
rect 7677 52797 7749 52800
rect 7801 52797 7873 52800
rect 7925 52797 9794 52800
rect 9846 52797 9918 52800
rect 9970 52797 10042 52800
rect 10094 52797 10166 52800
rect 10218 52797 12066 52800
rect 12118 52797 12190 52800
rect 12242 52797 12314 52800
rect 12366 52797 12438 52800
rect 12490 52797 13202 52800
rect 13254 52797 13326 52800
rect 13378 52797 13450 52800
rect 13502 52797 13574 52800
rect 13626 52797 14352 52800
rect 14404 52797 14460 52800
rect 604 52748 660 52751
rect 712 52748 1438 52751
rect 1490 52748 1562 52751
rect 1614 52748 1686 52751
rect 1738 52748 1810 52751
rect 1862 52748 2574 52751
rect 2626 52748 2698 52751
rect 2750 52748 2822 52751
rect 2874 52748 2946 52751
rect 2998 52748 4846 52751
rect 4898 52748 4970 52751
rect 5022 52748 5094 52751
rect 5146 52748 5218 52751
rect 5270 52748 7139 52751
rect 7191 52748 7263 52751
rect 7315 52748 7387 52751
rect 7439 52748 7625 52751
rect 7677 52748 7749 52751
rect 7801 52748 7873 52751
rect 7925 52748 9794 52751
rect 9846 52748 9918 52751
rect 9970 52748 10042 52751
rect 10094 52748 10166 52751
rect 10218 52748 12066 52751
rect 12118 52748 12190 52751
rect 12242 52748 12314 52751
rect 12366 52748 12438 52751
rect 12490 52748 13202 52751
rect 13254 52748 13326 52751
rect 13378 52748 13450 52751
rect 13502 52748 13574 52751
rect 13626 52748 14352 52751
rect 14404 52748 14460 52751
rect 14512 52748 14568 52800
rect 445 52692 14619 52748
rect 496 52640 552 52692
rect 604 52640 660 52692
rect 712 52676 14352 52692
rect 712 52640 1438 52676
rect 445 52624 1438 52640
rect 1490 52624 1562 52676
rect 1614 52624 1686 52676
rect 1738 52624 1810 52676
rect 1862 52624 2574 52676
rect 2626 52624 2698 52676
rect 2750 52624 2822 52676
rect 2874 52624 2946 52676
rect 2998 52624 4846 52676
rect 4898 52624 4970 52676
rect 5022 52624 5094 52676
rect 5146 52624 5218 52676
rect 5270 52624 7139 52676
rect 7191 52624 7263 52676
rect 7315 52624 7387 52676
rect 7439 52624 7625 52676
rect 7677 52624 7749 52676
rect 7801 52624 7873 52676
rect 7925 52624 9794 52676
rect 9846 52624 9918 52676
rect 9970 52624 10042 52676
rect 10094 52624 10166 52676
rect 10218 52624 12066 52676
rect 12118 52624 12190 52676
rect 12242 52624 12314 52676
rect 12366 52624 12438 52676
rect 12490 52624 13202 52676
rect 13254 52624 13326 52676
rect 13378 52624 13450 52676
rect 13502 52624 13574 52676
rect 13626 52640 14352 52676
rect 14404 52640 14460 52692
rect 14512 52640 14568 52692
rect 13626 52624 14619 52640
rect 445 52584 14619 52624
rect 496 52532 552 52584
rect 604 52532 660 52584
rect 712 52552 14352 52584
rect 712 52532 1438 52552
rect 445 52500 1438 52532
rect 1490 52500 1562 52552
rect 1614 52500 1686 52552
rect 1738 52500 1810 52552
rect 1862 52500 2574 52552
rect 2626 52500 2698 52552
rect 2750 52500 2822 52552
rect 2874 52500 2946 52552
rect 2998 52500 4846 52552
rect 4898 52500 4970 52552
rect 5022 52500 5094 52552
rect 5146 52500 5218 52552
rect 5270 52500 7139 52552
rect 7191 52500 7263 52552
rect 7315 52500 7387 52552
rect 7439 52500 7625 52552
rect 7677 52500 7749 52552
rect 7801 52500 7873 52552
rect 7925 52500 9794 52552
rect 9846 52500 9918 52552
rect 9970 52500 10042 52552
rect 10094 52500 10166 52552
rect 10218 52500 12066 52552
rect 12118 52500 12190 52552
rect 12242 52500 12314 52552
rect 12366 52500 12438 52552
rect 12490 52500 13202 52552
rect 13254 52500 13326 52552
rect 13378 52500 13450 52552
rect 13502 52500 13574 52552
rect 13626 52532 14352 52552
rect 14404 52532 14460 52584
rect 14512 52532 14568 52584
rect 13626 52500 14619 52532
rect 445 52450 14619 52500
rect 445 49150 456 52450
rect 920 52379 3836 52390
rect 920 52333 931 52379
rect 3825 52333 3836 52379
rect 920 52324 1148 52333
rect 1200 52324 1272 52333
rect 1324 52324 3729 52333
rect 920 52322 3729 52324
rect 660 52263 860 52300
rect 660 49337 803 52263
rect 849 49337 860 52263
rect 660 49150 860 49337
rect 920 52252 1920 52322
rect 920 52200 1148 52252
rect 1200 52200 1272 52252
rect 1324 52200 1920 52252
rect 920 52128 1920 52200
rect 920 52076 1148 52128
rect 1200 52076 1272 52128
rect 1324 52076 1920 52128
rect 920 52004 1920 52076
rect 920 51952 1148 52004
rect 1200 51952 1272 52004
rect 1324 51952 1920 52004
rect 920 51880 1920 51952
rect 920 51828 1148 51880
rect 1200 51828 1272 51880
rect 1324 51828 1920 51880
rect 920 51756 1920 51828
rect 920 51704 1148 51756
rect 1200 51704 1272 51756
rect 1324 51704 1920 51756
rect 920 51632 1920 51704
rect 920 51580 1148 51632
rect 1200 51580 1272 51632
rect 1324 51580 1920 51632
rect 920 51508 1920 51580
rect 920 51456 1148 51508
rect 1200 51456 1272 51508
rect 1324 51456 1920 51508
rect 920 51384 1920 51456
rect 920 51332 1148 51384
rect 1200 51332 1272 51384
rect 1324 51332 1920 51384
rect 920 51260 1920 51332
rect 920 51208 1148 51260
rect 1200 51208 1272 51260
rect 1324 51208 1920 51260
rect 920 51136 1920 51208
rect 920 51084 1148 51136
rect 1200 51084 1272 51136
rect 1324 51084 1920 51136
rect 920 51012 1920 51084
rect 920 50960 1148 51012
rect 1200 50960 1272 51012
rect 1324 50960 1920 51012
rect 920 50888 1920 50960
rect 920 50836 1148 50888
rect 1200 50836 1272 50888
rect 1324 50836 1920 50888
rect 920 50764 1920 50836
rect 920 50712 1148 50764
rect 1200 50712 1272 50764
rect 1324 50712 1920 50764
rect 920 50640 1920 50712
rect 920 50588 1148 50640
rect 1200 50588 1272 50640
rect 1324 50588 1920 50640
rect 920 50516 1920 50588
rect 920 50464 1148 50516
rect 1200 50464 1272 50516
rect 1324 50464 1920 50516
rect 920 50392 1920 50464
rect 920 50340 1148 50392
rect 1200 50340 1272 50392
rect 1324 50340 1920 50392
rect 920 50268 1920 50340
rect 920 50216 1148 50268
rect 1200 50216 1272 50268
rect 1324 50216 1920 50268
rect 920 50144 1920 50216
rect 920 50092 1148 50144
rect 1200 50092 1272 50144
rect 1324 50092 1920 50144
rect 920 50020 1920 50092
rect 920 49968 1148 50020
rect 1200 49968 1272 50020
rect 1324 49968 1920 50020
rect 920 49896 1920 49968
rect 920 49844 1148 49896
rect 1200 49844 1272 49896
rect 1324 49844 1920 49896
rect 920 49772 1920 49844
rect 920 49720 1148 49772
rect 1200 49720 1272 49772
rect 1324 49720 1920 49772
rect 920 49648 1920 49720
rect 920 49596 1148 49648
rect 1200 49596 1272 49648
rect 1324 49596 1920 49648
rect 920 49524 1920 49596
rect 920 49472 1148 49524
rect 1200 49472 1272 49524
rect 1324 49472 1920 49524
rect 920 49400 1920 49472
rect 920 49348 1148 49400
rect 1200 49348 1272 49400
rect 1324 49348 1920 49400
rect 920 49278 1920 49348
rect 2836 52286 3729 52322
rect 3781 52286 3836 52333
rect 4356 52379 7272 52390
rect 4356 52333 4367 52379
rect 7261 52333 7272 52379
rect 4356 52322 6335 52333
rect 2836 52230 3836 52286
rect 2836 52178 3729 52230
rect 3781 52178 3836 52230
rect 2836 52122 3836 52178
rect 2836 52070 3729 52122
rect 3781 52070 3836 52122
rect 2836 52014 3836 52070
rect 2836 51962 3729 52014
rect 3781 51962 3836 52014
rect 2836 51906 3836 51962
rect 2836 51854 3729 51906
rect 3781 51854 3836 51906
rect 2836 51798 3836 51854
rect 2836 51746 3729 51798
rect 3781 51746 3836 51798
rect 2836 51690 3836 51746
rect 2836 51638 3729 51690
rect 3781 51638 3836 51690
rect 2836 51582 3836 51638
rect 2836 51530 3729 51582
rect 3781 51530 3836 51582
rect 2836 51474 3836 51530
rect 2836 51422 3729 51474
rect 3781 51422 3836 51474
rect 2836 51366 3836 51422
rect 2836 51314 3729 51366
rect 3781 51314 3836 51366
rect 2836 51258 3836 51314
rect 2836 51206 3729 51258
rect 3781 51206 3836 51258
rect 2836 51150 3836 51206
rect 2836 51098 3729 51150
rect 3781 51098 3836 51150
rect 2836 51042 3836 51098
rect 2836 50990 3729 51042
rect 3781 50990 3836 51042
rect 2836 50934 3836 50990
rect 2836 50882 3729 50934
rect 3781 50882 3836 50934
rect 2836 50826 3836 50882
rect 2836 50774 3729 50826
rect 3781 50774 3836 50826
rect 2836 50718 3836 50774
rect 2836 50666 3729 50718
rect 3781 50666 3836 50718
rect 2836 50610 3836 50666
rect 2836 50558 3729 50610
rect 3781 50558 3836 50610
rect 2836 50502 3836 50558
rect 2836 50450 3729 50502
rect 3781 50450 3836 50502
rect 2836 50394 3836 50450
rect 2836 50342 3729 50394
rect 3781 50342 3836 50394
rect 2836 50286 3836 50342
rect 2836 50234 3729 50286
rect 3781 50234 3836 50286
rect 2836 50178 3836 50234
rect 2836 50126 3729 50178
rect 3781 50126 3836 50178
rect 2836 50070 3836 50126
rect 2836 50018 3729 50070
rect 3781 50018 3836 50070
rect 2836 49962 3836 50018
rect 2836 49910 3729 49962
rect 3781 49910 3836 49962
rect 2836 49854 3836 49910
rect 2836 49802 3729 49854
rect 3781 49802 3836 49854
rect 2836 49746 3836 49802
rect 2836 49694 3729 49746
rect 3781 49694 3836 49746
rect 2836 49638 3836 49694
rect 2836 49586 3729 49638
rect 3781 49586 3836 49638
rect 2836 49530 3836 49586
rect 2836 49478 3729 49530
rect 3781 49478 3836 49530
rect 2836 49422 3836 49478
rect 2836 49370 3729 49422
rect 3781 49370 3836 49422
rect 2836 49314 3836 49370
rect 2836 49278 3729 49314
rect 920 49276 3729 49278
rect 920 49267 1148 49276
rect 1200 49267 1272 49276
rect 1324 49267 3729 49276
rect 3781 49267 3836 49314
rect 920 49221 931 49267
rect 3825 49221 3836 49267
rect 920 49210 3836 49221
rect 3896 52263 4296 52300
rect 3896 49337 3907 52263
rect 3953 49337 4239 52263
rect 4285 49337 4296 52263
rect 3896 49150 4296 49337
rect 4356 49278 5356 52322
rect 6272 52286 6335 52322
rect 6387 52286 7272 52333
rect 7792 52379 10708 52390
rect 7792 52333 7803 52379
rect 10697 52333 10708 52379
rect 6272 52230 7272 52286
rect 6272 52178 6335 52230
rect 6387 52178 7272 52230
rect 6272 52122 7272 52178
rect 6272 52070 6335 52122
rect 6387 52070 7272 52122
rect 6272 52014 7272 52070
rect 6272 51962 6335 52014
rect 6387 51962 7272 52014
rect 6272 51906 7272 51962
rect 6272 51854 6335 51906
rect 6387 51854 7272 51906
rect 6272 51798 7272 51854
rect 6272 51746 6335 51798
rect 6387 51746 7272 51798
rect 6272 51690 7272 51746
rect 6272 51638 6335 51690
rect 6387 51638 7272 51690
rect 6272 51582 7272 51638
rect 6272 51530 6335 51582
rect 6387 51530 7272 51582
rect 6272 51474 7272 51530
rect 6272 51422 6335 51474
rect 6387 51422 7272 51474
rect 6272 51366 7272 51422
rect 6272 51314 6335 51366
rect 6387 51314 7272 51366
rect 6272 51258 7272 51314
rect 6272 51206 6335 51258
rect 6387 51206 7272 51258
rect 6272 51150 7272 51206
rect 6272 51098 6335 51150
rect 6387 51098 7272 51150
rect 6272 51042 7272 51098
rect 6272 50990 6335 51042
rect 6387 50990 7272 51042
rect 6272 50934 7272 50990
rect 6272 50882 6335 50934
rect 6387 50882 7272 50934
rect 6272 50826 7272 50882
rect 6272 50774 6335 50826
rect 6387 50774 7272 50826
rect 6272 50718 7272 50774
rect 6272 50666 6335 50718
rect 6387 50666 7272 50718
rect 6272 50610 7272 50666
rect 6272 50558 6335 50610
rect 6387 50558 7272 50610
rect 6272 50502 7272 50558
rect 6272 50450 6335 50502
rect 6387 50450 7272 50502
rect 6272 50394 7272 50450
rect 6272 50342 6335 50394
rect 6387 50342 7272 50394
rect 6272 50286 7272 50342
rect 6272 50234 6335 50286
rect 6387 50234 7272 50286
rect 6272 50178 7272 50234
rect 6272 50126 6335 50178
rect 6387 50126 7272 50178
rect 6272 50070 7272 50126
rect 6272 50018 6335 50070
rect 6387 50018 7272 50070
rect 6272 49962 7272 50018
rect 6272 49910 6335 49962
rect 6387 49910 7272 49962
rect 6272 49854 7272 49910
rect 6272 49802 6335 49854
rect 6387 49802 7272 49854
rect 6272 49746 7272 49802
rect 6272 49694 6335 49746
rect 6387 49694 7272 49746
rect 6272 49638 7272 49694
rect 6272 49586 6335 49638
rect 6387 49586 7272 49638
rect 6272 49530 7272 49586
rect 6272 49478 6335 49530
rect 6387 49478 7272 49530
rect 6272 49422 7272 49478
rect 6272 49370 6335 49422
rect 6387 49370 7272 49422
rect 6272 49314 7272 49370
rect 6272 49278 6335 49314
rect 4356 49267 6335 49278
rect 6387 49267 7272 49314
rect 4356 49221 4367 49267
rect 7261 49221 7272 49267
rect 4356 49210 7272 49221
rect 7332 52284 7732 52300
rect 7332 52263 7388 52284
rect 7332 49337 7343 52263
rect 7440 52232 7624 52284
rect 7676 52263 7732 52284
rect 7389 52176 7675 52232
rect 7440 52124 7624 52176
rect 7389 52068 7675 52124
rect 7440 52016 7624 52068
rect 7389 51960 7675 52016
rect 7440 51908 7624 51960
rect 7389 51852 7675 51908
rect 7440 51800 7624 51852
rect 7389 51744 7675 51800
rect 7440 51692 7624 51744
rect 7389 51636 7675 51692
rect 7440 51584 7624 51636
rect 7389 51528 7675 51584
rect 7440 51476 7624 51528
rect 7389 51420 7675 51476
rect 7440 51368 7624 51420
rect 7389 51312 7675 51368
rect 7440 51260 7624 51312
rect 7389 51204 7675 51260
rect 7440 51152 7624 51204
rect 7389 51096 7675 51152
rect 7440 51044 7624 51096
rect 7389 50988 7675 51044
rect 7440 50936 7624 50988
rect 7389 50880 7675 50936
rect 7440 50828 7624 50880
rect 7389 50772 7675 50828
rect 7440 50720 7624 50772
rect 7389 50664 7675 50720
rect 7440 50612 7624 50664
rect 7389 50556 7675 50612
rect 7440 50504 7624 50556
rect 7389 50448 7675 50504
rect 7440 50396 7624 50448
rect 7389 50340 7675 50396
rect 7440 50288 7624 50340
rect 7389 50232 7675 50288
rect 7440 50180 7624 50232
rect 7389 50124 7675 50180
rect 7440 50072 7624 50124
rect 7389 50016 7675 50072
rect 7440 49964 7624 50016
rect 7389 49908 7675 49964
rect 7440 49856 7624 49908
rect 7389 49800 7675 49856
rect 7440 49748 7624 49800
rect 7389 49692 7675 49748
rect 7440 49640 7624 49692
rect 7389 49584 7675 49640
rect 7440 49532 7624 49584
rect 7389 49476 7675 49532
rect 7440 49424 7624 49476
rect 7389 49368 7675 49424
rect 7332 49316 7388 49337
rect 7440 49316 7624 49368
rect 7721 49337 7732 52263
rect 7676 49316 7732 49337
rect 7332 49150 7732 49316
rect 7792 52286 8677 52333
rect 8729 52322 10708 52333
rect 8729 52286 8792 52322
rect 7792 52230 8792 52286
rect 7792 52178 8677 52230
rect 8729 52178 8792 52230
rect 7792 52122 8792 52178
rect 7792 52070 8677 52122
rect 8729 52070 8792 52122
rect 7792 52014 8792 52070
rect 7792 51962 8677 52014
rect 8729 51962 8792 52014
rect 7792 51906 8792 51962
rect 7792 51854 8677 51906
rect 8729 51854 8792 51906
rect 7792 51798 8792 51854
rect 7792 51746 8677 51798
rect 8729 51746 8792 51798
rect 7792 51690 8792 51746
rect 7792 51638 8677 51690
rect 8729 51638 8792 51690
rect 7792 51582 8792 51638
rect 7792 51530 8677 51582
rect 8729 51530 8792 51582
rect 7792 51474 8792 51530
rect 7792 51422 8677 51474
rect 8729 51422 8792 51474
rect 7792 51366 8792 51422
rect 7792 51314 8677 51366
rect 8729 51314 8792 51366
rect 7792 51258 8792 51314
rect 7792 51206 8677 51258
rect 8729 51206 8792 51258
rect 7792 51150 8792 51206
rect 7792 51098 8677 51150
rect 8729 51098 8792 51150
rect 7792 51042 8792 51098
rect 7792 50990 8677 51042
rect 8729 50990 8792 51042
rect 7792 50934 8792 50990
rect 7792 50882 8677 50934
rect 8729 50882 8792 50934
rect 7792 50826 8792 50882
rect 7792 50774 8677 50826
rect 8729 50774 8792 50826
rect 7792 50718 8792 50774
rect 7792 50666 8677 50718
rect 8729 50666 8792 50718
rect 7792 50610 8792 50666
rect 7792 50558 8677 50610
rect 8729 50558 8792 50610
rect 7792 50502 8792 50558
rect 7792 50450 8677 50502
rect 8729 50450 8792 50502
rect 7792 50394 8792 50450
rect 7792 50342 8677 50394
rect 8729 50342 8792 50394
rect 7792 50286 8792 50342
rect 7792 50234 8677 50286
rect 8729 50234 8792 50286
rect 7792 50178 8792 50234
rect 7792 50126 8677 50178
rect 8729 50126 8792 50178
rect 7792 50070 8792 50126
rect 7792 50018 8677 50070
rect 8729 50018 8792 50070
rect 7792 49962 8792 50018
rect 7792 49910 8677 49962
rect 8729 49910 8792 49962
rect 7792 49854 8792 49910
rect 7792 49802 8677 49854
rect 8729 49802 8792 49854
rect 7792 49746 8792 49802
rect 7792 49694 8677 49746
rect 8729 49694 8792 49746
rect 7792 49638 8792 49694
rect 7792 49586 8677 49638
rect 8729 49586 8792 49638
rect 7792 49530 8792 49586
rect 7792 49478 8677 49530
rect 8729 49478 8792 49530
rect 7792 49422 8792 49478
rect 7792 49370 8677 49422
rect 8729 49370 8792 49422
rect 7792 49314 8792 49370
rect 7792 49267 8677 49314
rect 8729 49278 8792 49314
rect 9708 49278 10708 52322
rect 11228 52379 14144 52390
rect 11228 52333 11239 52379
rect 14133 52333 14144 52379
rect 8729 49267 10708 49278
rect 7792 49221 7803 49267
rect 10697 49221 10708 49267
rect 7792 49210 10708 49221
rect 10768 52263 11168 52300
rect 10768 49337 10779 52263
rect 10825 49337 11111 52263
rect 11157 49337 11168 52263
rect 10768 49150 11168 49337
rect 11228 52286 11283 52333
rect 11335 52324 13786 52333
rect 13838 52324 13910 52333
rect 13962 52324 14034 52333
rect 14086 52324 14144 52333
rect 11335 52322 14144 52324
rect 11335 52286 12228 52322
rect 11228 52230 12228 52286
rect 11228 52178 11283 52230
rect 11335 52178 12228 52230
rect 11228 52122 12228 52178
rect 11228 52070 11283 52122
rect 11335 52070 12228 52122
rect 11228 52014 12228 52070
rect 11228 51962 11283 52014
rect 11335 51962 12228 52014
rect 11228 51906 12228 51962
rect 11228 51854 11283 51906
rect 11335 51854 12228 51906
rect 11228 51798 12228 51854
rect 11228 51746 11283 51798
rect 11335 51746 12228 51798
rect 11228 51690 12228 51746
rect 11228 51638 11283 51690
rect 11335 51638 12228 51690
rect 11228 51582 12228 51638
rect 11228 51530 11283 51582
rect 11335 51530 12228 51582
rect 11228 51474 12228 51530
rect 11228 51422 11283 51474
rect 11335 51422 12228 51474
rect 11228 51366 12228 51422
rect 11228 51314 11283 51366
rect 11335 51314 12228 51366
rect 11228 51258 12228 51314
rect 11228 51206 11283 51258
rect 11335 51206 12228 51258
rect 11228 51150 12228 51206
rect 11228 51098 11283 51150
rect 11335 51098 12228 51150
rect 11228 51042 12228 51098
rect 11228 50990 11283 51042
rect 11335 50990 12228 51042
rect 11228 50934 12228 50990
rect 11228 50882 11283 50934
rect 11335 50882 12228 50934
rect 11228 50826 12228 50882
rect 11228 50774 11283 50826
rect 11335 50774 12228 50826
rect 11228 50718 12228 50774
rect 11228 50666 11283 50718
rect 11335 50666 12228 50718
rect 11228 50610 12228 50666
rect 11228 50558 11283 50610
rect 11335 50558 12228 50610
rect 11228 50502 12228 50558
rect 11228 50450 11283 50502
rect 11335 50450 12228 50502
rect 11228 50394 12228 50450
rect 11228 50342 11283 50394
rect 11335 50342 12228 50394
rect 11228 50286 12228 50342
rect 11228 50234 11283 50286
rect 11335 50234 12228 50286
rect 11228 50178 12228 50234
rect 11228 50126 11283 50178
rect 11335 50126 12228 50178
rect 11228 50070 12228 50126
rect 11228 50018 11283 50070
rect 11335 50018 12228 50070
rect 11228 49962 12228 50018
rect 11228 49910 11283 49962
rect 11335 49910 12228 49962
rect 11228 49854 12228 49910
rect 11228 49802 11283 49854
rect 11335 49802 12228 49854
rect 11228 49746 12228 49802
rect 11228 49694 11283 49746
rect 11335 49694 12228 49746
rect 11228 49638 12228 49694
rect 11228 49586 11283 49638
rect 11335 49586 12228 49638
rect 11228 49530 12228 49586
rect 11228 49478 11283 49530
rect 11335 49478 12228 49530
rect 11228 49422 12228 49478
rect 11228 49370 11283 49422
rect 11335 49370 12228 49422
rect 11228 49314 12228 49370
rect 11228 49267 11283 49314
rect 11335 49278 12228 49314
rect 13144 52252 14144 52322
rect 13144 52200 13786 52252
rect 13838 52200 13910 52252
rect 13962 52200 14034 52252
rect 14086 52200 14144 52252
rect 13144 52128 14144 52200
rect 13144 52076 13786 52128
rect 13838 52076 13910 52128
rect 13962 52076 14034 52128
rect 14086 52076 14144 52128
rect 13144 52004 14144 52076
rect 13144 51952 13786 52004
rect 13838 51952 13910 52004
rect 13962 51952 14034 52004
rect 14086 51952 14144 52004
rect 13144 51880 14144 51952
rect 13144 51828 13786 51880
rect 13838 51828 13910 51880
rect 13962 51828 14034 51880
rect 14086 51828 14144 51880
rect 13144 51756 14144 51828
rect 13144 51704 13786 51756
rect 13838 51704 13910 51756
rect 13962 51704 14034 51756
rect 14086 51704 14144 51756
rect 13144 51632 14144 51704
rect 13144 51580 13786 51632
rect 13838 51580 13910 51632
rect 13962 51580 14034 51632
rect 14086 51580 14144 51632
rect 13144 51508 14144 51580
rect 13144 51456 13786 51508
rect 13838 51456 13910 51508
rect 13962 51456 14034 51508
rect 14086 51456 14144 51508
rect 13144 51384 14144 51456
rect 13144 51332 13786 51384
rect 13838 51332 13910 51384
rect 13962 51332 14034 51384
rect 14086 51332 14144 51384
rect 13144 51260 14144 51332
rect 13144 51208 13786 51260
rect 13838 51208 13910 51260
rect 13962 51208 14034 51260
rect 14086 51208 14144 51260
rect 13144 51136 14144 51208
rect 13144 51084 13786 51136
rect 13838 51084 13910 51136
rect 13962 51084 14034 51136
rect 14086 51084 14144 51136
rect 13144 51012 14144 51084
rect 13144 50960 13786 51012
rect 13838 50960 13910 51012
rect 13962 50960 14034 51012
rect 14086 50960 14144 51012
rect 13144 50888 14144 50960
rect 13144 50836 13786 50888
rect 13838 50836 13910 50888
rect 13962 50836 14034 50888
rect 14086 50836 14144 50888
rect 13144 50764 14144 50836
rect 13144 50712 13786 50764
rect 13838 50712 13910 50764
rect 13962 50712 14034 50764
rect 14086 50712 14144 50764
rect 13144 50640 14144 50712
rect 13144 50588 13786 50640
rect 13838 50588 13910 50640
rect 13962 50588 14034 50640
rect 14086 50588 14144 50640
rect 13144 50516 14144 50588
rect 13144 50464 13786 50516
rect 13838 50464 13910 50516
rect 13962 50464 14034 50516
rect 14086 50464 14144 50516
rect 13144 50392 14144 50464
rect 13144 50340 13786 50392
rect 13838 50340 13910 50392
rect 13962 50340 14034 50392
rect 14086 50340 14144 50392
rect 13144 50268 14144 50340
rect 13144 50216 13786 50268
rect 13838 50216 13910 50268
rect 13962 50216 14034 50268
rect 14086 50216 14144 50268
rect 13144 50144 14144 50216
rect 13144 50092 13786 50144
rect 13838 50092 13910 50144
rect 13962 50092 14034 50144
rect 14086 50092 14144 50144
rect 13144 50020 14144 50092
rect 13144 49968 13786 50020
rect 13838 49968 13910 50020
rect 13962 49968 14034 50020
rect 14086 49968 14144 50020
rect 13144 49896 14144 49968
rect 13144 49844 13786 49896
rect 13838 49844 13910 49896
rect 13962 49844 14034 49896
rect 14086 49844 14144 49896
rect 13144 49772 14144 49844
rect 13144 49720 13786 49772
rect 13838 49720 13910 49772
rect 13962 49720 14034 49772
rect 14086 49720 14144 49772
rect 13144 49648 14144 49720
rect 13144 49596 13786 49648
rect 13838 49596 13910 49648
rect 13962 49596 14034 49648
rect 14086 49596 14144 49648
rect 13144 49524 14144 49596
rect 13144 49472 13786 49524
rect 13838 49472 13910 49524
rect 13962 49472 14034 49524
rect 14086 49472 14144 49524
rect 13144 49400 14144 49472
rect 13144 49348 13786 49400
rect 13838 49348 13910 49400
rect 13962 49348 14034 49400
rect 14086 49348 14144 49400
rect 13144 49278 14144 49348
rect 11335 49276 14144 49278
rect 11335 49267 13786 49276
rect 13838 49267 13910 49276
rect 13962 49267 14034 49276
rect 14086 49267 14144 49276
rect 11228 49221 11239 49267
rect 14133 49221 14144 49267
rect 11228 49210 14144 49221
rect 14204 52263 14404 52300
rect 14204 49337 14215 52263
rect 14261 49337 14404 52263
rect 14204 49150 14404 49337
rect 14608 49150 14619 52450
rect 445 49100 14619 49150
rect 445 49068 1438 49100
rect 496 49016 552 49068
rect 604 49016 660 49068
rect 712 49048 1438 49068
rect 1490 49048 1562 49100
rect 1614 49048 1686 49100
rect 1738 49048 1810 49100
rect 1862 49048 2574 49100
rect 2626 49048 2698 49100
rect 2750 49048 2822 49100
rect 2874 49048 2946 49100
rect 2998 49048 4846 49100
rect 4898 49048 4970 49100
rect 5022 49048 5094 49100
rect 5146 49048 5218 49100
rect 5270 49048 7139 49100
rect 7191 49048 7263 49100
rect 7315 49048 7387 49100
rect 7439 49048 7625 49100
rect 7677 49048 7749 49100
rect 7801 49048 7873 49100
rect 7925 49048 9794 49100
rect 9846 49048 9918 49100
rect 9970 49048 10042 49100
rect 10094 49048 10166 49100
rect 10218 49048 12066 49100
rect 12118 49048 12190 49100
rect 12242 49048 12314 49100
rect 12366 49048 12438 49100
rect 12490 49048 13480 49100
rect 13532 49048 13604 49100
rect 13656 49068 14619 49100
rect 13656 49048 14352 49068
rect 712 49016 14352 49048
rect 14404 49016 14460 49068
rect 14512 49016 14568 49068
rect 445 48976 14619 49016
rect 445 48960 1438 48976
rect 496 48908 552 48960
rect 604 48908 660 48960
rect 712 48924 1438 48960
rect 1490 48924 1562 48976
rect 1614 48924 1686 48976
rect 1738 48924 1810 48976
rect 1862 48924 2574 48976
rect 2626 48924 2698 48976
rect 2750 48924 2822 48976
rect 2874 48924 2946 48976
rect 2998 48924 4846 48976
rect 4898 48924 4970 48976
rect 5022 48924 5094 48976
rect 5146 48924 5218 48976
rect 5270 48924 7139 48976
rect 7191 48924 7263 48976
rect 7315 48924 7387 48976
rect 7439 48924 7625 48976
rect 7677 48924 7749 48976
rect 7801 48924 7873 48976
rect 7925 48924 9794 48976
rect 9846 48924 9918 48976
rect 9970 48924 10042 48976
rect 10094 48924 10166 48976
rect 10218 48924 12066 48976
rect 12118 48924 12190 48976
rect 12242 48924 12314 48976
rect 12366 48924 12438 48976
rect 12490 48924 13480 48976
rect 13532 48924 13604 48976
rect 13656 48960 14619 48976
rect 13656 48924 14352 48960
rect 712 48908 14352 48924
rect 14404 48908 14460 48960
rect 14512 48908 14568 48960
rect 445 48852 14619 48908
rect 496 48800 552 48852
rect 604 48849 660 48852
rect 712 48849 1438 48852
rect 1490 48849 1562 48852
rect 1614 48849 1686 48852
rect 1738 48849 1810 48852
rect 1862 48849 2574 48852
rect 2626 48849 2698 48852
rect 2750 48849 2822 48852
rect 2874 48849 2946 48852
rect 2998 48849 4846 48852
rect 4898 48849 4970 48852
rect 5022 48849 5094 48852
rect 5146 48849 5218 48852
rect 5270 48849 7139 48852
rect 7191 48849 7263 48852
rect 7315 48849 7387 48852
rect 7439 48849 7625 48852
rect 7677 48849 7749 48852
rect 7801 48849 7873 48852
rect 7925 48849 9794 48852
rect 9846 48849 9918 48852
rect 9970 48849 10042 48852
rect 10094 48849 10166 48852
rect 10218 48849 12066 48852
rect 12118 48849 12190 48852
rect 12242 48849 12314 48852
rect 12366 48849 12438 48852
rect 12490 48849 13480 48852
rect 13532 48849 13604 48852
rect 13656 48849 14352 48852
rect 14404 48849 14460 48852
rect 604 48800 660 48803
rect 712 48800 1438 48803
rect 1490 48800 1562 48803
rect 1614 48800 1686 48803
rect 1738 48800 1810 48803
rect 1862 48800 2574 48803
rect 2626 48800 2698 48803
rect 2750 48800 2822 48803
rect 2874 48800 2946 48803
rect 2998 48800 4846 48803
rect 4898 48800 4970 48803
rect 5022 48800 5094 48803
rect 5146 48800 5218 48803
rect 5270 48800 7139 48803
rect 7191 48800 7263 48803
rect 7315 48800 7387 48803
rect 7439 48800 7625 48803
rect 7677 48800 7749 48803
rect 7801 48800 7873 48803
rect 7925 48800 9794 48803
rect 9846 48800 9918 48803
rect 9970 48800 10042 48803
rect 10094 48800 10166 48803
rect 10218 48800 12066 48803
rect 12118 48800 12190 48803
rect 12242 48800 12314 48803
rect 12366 48800 12438 48803
rect 12490 48800 13480 48803
rect 13532 48800 13604 48803
rect 13656 48800 14352 48803
rect 14404 48800 14460 48803
rect 14512 48800 14568 48852
rect 445 48744 14619 48800
rect 496 48692 552 48744
rect 604 48692 660 48744
rect 712 48728 14352 48744
rect 712 48692 1438 48728
rect 445 48676 1438 48692
rect 1490 48676 1562 48728
rect 1614 48676 1686 48728
rect 1738 48676 1810 48728
rect 1862 48676 2574 48728
rect 2626 48676 2698 48728
rect 2750 48676 2822 48728
rect 2874 48676 2946 48728
rect 2998 48676 4846 48728
rect 4898 48676 4970 48728
rect 5022 48676 5094 48728
rect 5146 48676 5218 48728
rect 5270 48676 7139 48728
rect 7191 48676 7263 48728
rect 7315 48676 7387 48728
rect 7439 48676 7625 48728
rect 7677 48676 7749 48728
rect 7801 48676 7873 48728
rect 7925 48676 9794 48728
rect 9846 48676 9918 48728
rect 9970 48676 10042 48728
rect 10094 48676 10166 48728
rect 10218 48676 12066 48728
rect 12118 48676 12190 48728
rect 12242 48676 12314 48728
rect 12366 48676 12438 48728
rect 12490 48676 13480 48728
rect 13532 48676 13604 48728
rect 13656 48692 14352 48728
rect 14404 48692 14460 48744
rect 14512 48692 14568 48744
rect 13656 48676 14619 48692
rect 445 48636 14619 48676
rect 496 48584 552 48636
rect 604 48584 660 48636
rect 712 48604 14352 48636
rect 712 48584 1438 48604
rect 445 48552 1438 48584
rect 1490 48552 1562 48604
rect 1614 48552 1686 48604
rect 1738 48552 1810 48604
rect 1862 48552 2574 48604
rect 2626 48552 2698 48604
rect 2750 48552 2822 48604
rect 2874 48552 2946 48604
rect 2998 48552 4846 48604
rect 4898 48552 4970 48604
rect 5022 48552 5094 48604
rect 5146 48552 5218 48604
rect 5270 48552 7139 48604
rect 7191 48552 7263 48604
rect 7315 48552 7387 48604
rect 7439 48552 7625 48604
rect 7677 48552 7749 48604
rect 7801 48552 7873 48604
rect 7925 48552 9794 48604
rect 9846 48552 9918 48604
rect 9970 48552 10042 48604
rect 10094 48552 10166 48604
rect 10218 48552 12066 48604
rect 12118 48552 12190 48604
rect 12242 48552 12314 48604
rect 12366 48552 12438 48604
rect 12490 48552 13480 48604
rect 13532 48552 13604 48604
rect 13656 48584 14352 48604
rect 14404 48584 14460 48636
rect 14512 48584 14568 48636
rect 13656 48552 14619 48584
rect 445 48502 14619 48552
rect 445 45202 456 48502
rect 920 48431 3836 48442
rect 920 48385 931 48431
rect 3825 48385 3836 48431
rect 920 48376 1148 48385
rect 1200 48376 1272 48385
rect 1324 48376 3729 48385
rect 920 48374 3729 48376
rect 660 48315 860 48352
rect 660 45389 803 48315
rect 849 45389 860 48315
rect 660 45202 860 45389
rect 920 48304 1920 48374
rect 920 48252 1148 48304
rect 1200 48252 1272 48304
rect 1324 48252 1920 48304
rect 920 48180 1920 48252
rect 920 48128 1148 48180
rect 1200 48128 1272 48180
rect 1324 48128 1920 48180
rect 920 48056 1920 48128
rect 920 48004 1148 48056
rect 1200 48004 1272 48056
rect 1324 48004 1920 48056
rect 920 47932 1920 48004
rect 920 47880 1148 47932
rect 1200 47880 1272 47932
rect 1324 47880 1920 47932
rect 920 47808 1920 47880
rect 920 47756 1148 47808
rect 1200 47756 1272 47808
rect 1324 47756 1920 47808
rect 920 47684 1920 47756
rect 920 47632 1148 47684
rect 1200 47632 1272 47684
rect 1324 47632 1920 47684
rect 920 47560 1920 47632
rect 920 47508 1148 47560
rect 1200 47508 1272 47560
rect 1324 47508 1920 47560
rect 920 47436 1920 47508
rect 920 47384 1148 47436
rect 1200 47384 1272 47436
rect 1324 47384 1920 47436
rect 920 47312 1920 47384
rect 920 47260 1148 47312
rect 1200 47260 1272 47312
rect 1324 47260 1920 47312
rect 920 47188 1920 47260
rect 920 47136 1148 47188
rect 1200 47136 1272 47188
rect 1324 47136 1920 47188
rect 920 47064 1920 47136
rect 920 47012 1148 47064
rect 1200 47012 1272 47064
rect 1324 47012 1920 47064
rect 920 46940 1920 47012
rect 920 46888 1148 46940
rect 1200 46888 1272 46940
rect 1324 46888 1920 46940
rect 920 46816 1920 46888
rect 920 46764 1148 46816
rect 1200 46764 1272 46816
rect 1324 46764 1920 46816
rect 920 46692 1920 46764
rect 920 46640 1148 46692
rect 1200 46640 1272 46692
rect 1324 46640 1920 46692
rect 920 46568 1920 46640
rect 920 46516 1148 46568
rect 1200 46516 1272 46568
rect 1324 46516 1920 46568
rect 920 46444 1920 46516
rect 920 46392 1148 46444
rect 1200 46392 1272 46444
rect 1324 46392 1920 46444
rect 920 46320 1920 46392
rect 920 46268 1148 46320
rect 1200 46268 1272 46320
rect 1324 46268 1920 46320
rect 920 46196 1920 46268
rect 920 46144 1148 46196
rect 1200 46144 1272 46196
rect 1324 46144 1920 46196
rect 920 46072 1920 46144
rect 920 46020 1148 46072
rect 1200 46020 1272 46072
rect 1324 46020 1920 46072
rect 920 45948 1920 46020
rect 920 45896 1148 45948
rect 1200 45896 1272 45948
rect 1324 45896 1920 45948
rect 920 45824 1920 45896
rect 920 45772 1148 45824
rect 1200 45772 1272 45824
rect 1324 45772 1920 45824
rect 920 45700 1920 45772
rect 920 45648 1148 45700
rect 1200 45648 1272 45700
rect 1324 45648 1920 45700
rect 920 45576 1920 45648
rect 920 45524 1148 45576
rect 1200 45524 1272 45576
rect 1324 45524 1920 45576
rect 920 45452 1920 45524
rect 920 45400 1148 45452
rect 1200 45400 1272 45452
rect 1324 45400 1920 45452
rect 920 45330 1920 45400
rect 2836 48338 3729 48374
rect 3781 48338 3836 48385
rect 4356 48431 7272 48442
rect 4356 48385 4367 48431
rect 7261 48385 7272 48431
rect 4356 48374 6335 48385
rect 2836 48282 3836 48338
rect 2836 48230 3729 48282
rect 3781 48230 3836 48282
rect 2836 48174 3836 48230
rect 2836 48122 3729 48174
rect 3781 48122 3836 48174
rect 2836 48066 3836 48122
rect 2836 48014 3729 48066
rect 3781 48014 3836 48066
rect 2836 47958 3836 48014
rect 2836 47906 3729 47958
rect 3781 47906 3836 47958
rect 2836 47850 3836 47906
rect 2836 47798 3729 47850
rect 3781 47798 3836 47850
rect 2836 47742 3836 47798
rect 2836 47690 3729 47742
rect 3781 47690 3836 47742
rect 2836 47634 3836 47690
rect 2836 47582 3729 47634
rect 3781 47582 3836 47634
rect 2836 47526 3836 47582
rect 2836 47474 3729 47526
rect 3781 47474 3836 47526
rect 2836 47418 3836 47474
rect 2836 47366 3729 47418
rect 3781 47366 3836 47418
rect 2836 47310 3836 47366
rect 2836 47258 3729 47310
rect 3781 47258 3836 47310
rect 2836 47202 3836 47258
rect 2836 47150 3729 47202
rect 3781 47150 3836 47202
rect 2836 47094 3836 47150
rect 2836 47042 3729 47094
rect 3781 47042 3836 47094
rect 2836 46986 3836 47042
rect 2836 46934 3729 46986
rect 3781 46934 3836 46986
rect 2836 46878 3836 46934
rect 2836 46826 3729 46878
rect 3781 46826 3836 46878
rect 2836 46770 3836 46826
rect 2836 46718 3729 46770
rect 3781 46718 3836 46770
rect 2836 46662 3836 46718
rect 2836 46610 3729 46662
rect 3781 46610 3836 46662
rect 2836 46554 3836 46610
rect 2836 46502 3729 46554
rect 3781 46502 3836 46554
rect 2836 46446 3836 46502
rect 2836 46394 3729 46446
rect 3781 46394 3836 46446
rect 2836 46338 3836 46394
rect 2836 46286 3729 46338
rect 3781 46286 3836 46338
rect 2836 46230 3836 46286
rect 2836 46178 3729 46230
rect 3781 46178 3836 46230
rect 2836 46122 3836 46178
rect 2836 46070 3729 46122
rect 3781 46070 3836 46122
rect 2836 46014 3836 46070
rect 2836 45962 3729 46014
rect 3781 45962 3836 46014
rect 2836 45906 3836 45962
rect 2836 45854 3729 45906
rect 3781 45854 3836 45906
rect 2836 45798 3836 45854
rect 2836 45746 3729 45798
rect 3781 45746 3836 45798
rect 2836 45690 3836 45746
rect 2836 45638 3729 45690
rect 3781 45638 3836 45690
rect 2836 45582 3836 45638
rect 2836 45530 3729 45582
rect 3781 45530 3836 45582
rect 2836 45474 3836 45530
rect 2836 45422 3729 45474
rect 3781 45422 3836 45474
rect 2836 45366 3836 45422
rect 2836 45330 3729 45366
rect 920 45328 3729 45330
rect 920 45319 1148 45328
rect 1200 45319 1272 45328
rect 1324 45319 3729 45328
rect 3781 45319 3836 45366
rect 920 45273 931 45319
rect 3825 45273 3836 45319
rect 920 45262 3836 45273
rect 3896 48315 4296 48352
rect 3896 45389 3907 48315
rect 3953 45389 4239 48315
rect 4285 45389 4296 48315
rect 3896 45202 4296 45389
rect 4356 45330 5356 48374
rect 6272 48338 6335 48374
rect 6387 48338 7272 48385
rect 7792 48431 10708 48442
rect 7792 48385 7803 48431
rect 10697 48385 10708 48431
rect 6272 48282 7272 48338
rect 6272 48230 6335 48282
rect 6387 48230 7272 48282
rect 6272 48174 7272 48230
rect 6272 48122 6335 48174
rect 6387 48122 7272 48174
rect 6272 48066 7272 48122
rect 6272 48014 6335 48066
rect 6387 48014 7272 48066
rect 6272 47958 7272 48014
rect 6272 47906 6335 47958
rect 6387 47906 7272 47958
rect 6272 47850 7272 47906
rect 6272 47798 6335 47850
rect 6387 47798 7272 47850
rect 6272 47742 7272 47798
rect 6272 47690 6335 47742
rect 6387 47690 7272 47742
rect 6272 47634 7272 47690
rect 6272 47582 6335 47634
rect 6387 47582 7272 47634
rect 6272 47526 7272 47582
rect 6272 47474 6335 47526
rect 6387 47474 7272 47526
rect 6272 47418 7272 47474
rect 6272 47366 6335 47418
rect 6387 47366 7272 47418
rect 6272 47310 7272 47366
rect 6272 47258 6335 47310
rect 6387 47258 7272 47310
rect 6272 47202 7272 47258
rect 6272 47150 6335 47202
rect 6387 47150 7272 47202
rect 6272 47094 7272 47150
rect 6272 47042 6335 47094
rect 6387 47042 7272 47094
rect 6272 46986 7272 47042
rect 6272 46934 6335 46986
rect 6387 46934 7272 46986
rect 6272 46878 7272 46934
rect 6272 46826 6335 46878
rect 6387 46826 7272 46878
rect 6272 46770 7272 46826
rect 6272 46718 6335 46770
rect 6387 46718 7272 46770
rect 6272 46662 7272 46718
rect 6272 46610 6335 46662
rect 6387 46610 7272 46662
rect 6272 46554 7272 46610
rect 6272 46502 6335 46554
rect 6387 46502 7272 46554
rect 6272 46446 7272 46502
rect 6272 46394 6335 46446
rect 6387 46394 7272 46446
rect 6272 46338 7272 46394
rect 6272 46286 6335 46338
rect 6387 46286 7272 46338
rect 6272 46230 7272 46286
rect 6272 46178 6335 46230
rect 6387 46178 7272 46230
rect 6272 46122 7272 46178
rect 6272 46070 6335 46122
rect 6387 46070 7272 46122
rect 6272 46014 7272 46070
rect 6272 45962 6335 46014
rect 6387 45962 7272 46014
rect 6272 45906 7272 45962
rect 6272 45854 6335 45906
rect 6387 45854 7272 45906
rect 6272 45798 7272 45854
rect 6272 45746 6335 45798
rect 6387 45746 7272 45798
rect 6272 45690 7272 45746
rect 6272 45638 6335 45690
rect 6387 45638 7272 45690
rect 6272 45582 7272 45638
rect 6272 45530 6335 45582
rect 6387 45530 7272 45582
rect 6272 45474 7272 45530
rect 6272 45422 6335 45474
rect 6387 45422 7272 45474
rect 6272 45366 7272 45422
rect 6272 45330 6335 45366
rect 4356 45319 6335 45330
rect 6387 45319 7272 45366
rect 4356 45273 4367 45319
rect 7261 45273 7272 45319
rect 4356 45262 7272 45273
rect 7332 48336 7732 48352
rect 7332 48315 7388 48336
rect 7332 45389 7343 48315
rect 7440 48284 7624 48336
rect 7676 48315 7732 48336
rect 7389 48228 7675 48284
rect 7440 48176 7624 48228
rect 7389 48120 7675 48176
rect 7440 48068 7624 48120
rect 7389 48012 7675 48068
rect 7440 47960 7624 48012
rect 7389 47904 7675 47960
rect 7440 47852 7624 47904
rect 7389 47796 7675 47852
rect 7440 47744 7624 47796
rect 7389 47688 7675 47744
rect 7440 47636 7624 47688
rect 7389 47580 7675 47636
rect 7440 47528 7624 47580
rect 7389 47472 7675 47528
rect 7440 47420 7624 47472
rect 7389 47364 7675 47420
rect 7440 47312 7624 47364
rect 7389 47256 7675 47312
rect 7440 47204 7624 47256
rect 7389 47148 7675 47204
rect 7440 47096 7624 47148
rect 7389 47040 7675 47096
rect 7440 46988 7624 47040
rect 7389 46932 7675 46988
rect 7440 46880 7624 46932
rect 7389 46824 7675 46880
rect 7440 46772 7624 46824
rect 7389 46716 7675 46772
rect 7440 46664 7624 46716
rect 7389 46608 7675 46664
rect 7440 46556 7624 46608
rect 7389 46500 7675 46556
rect 7440 46448 7624 46500
rect 7389 46392 7675 46448
rect 7440 46340 7624 46392
rect 7389 46284 7675 46340
rect 7440 46232 7624 46284
rect 7389 46176 7675 46232
rect 7440 46124 7624 46176
rect 7389 46068 7675 46124
rect 7440 46016 7624 46068
rect 7389 45960 7675 46016
rect 7440 45908 7624 45960
rect 7389 45852 7675 45908
rect 7440 45800 7624 45852
rect 7389 45744 7675 45800
rect 7440 45692 7624 45744
rect 7389 45636 7675 45692
rect 7440 45584 7624 45636
rect 7389 45528 7675 45584
rect 7440 45476 7624 45528
rect 7389 45420 7675 45476
rect 7332 45368 7388 45389
rect 7440 45368 7624 45420
rect 7721 45389 7732 48315
rect 7676 45368 7732 45389
rect 7332 45202 7732 45368
rect 7792 48338 8677 48385
rect 8729 48374 10708 48385
rect 8729 48338 8792 48374
rect 7792 48282 8792 48338
rect 7792 48230 8677 48282
rect 8729 48230 8792 48282
rect 7792 48174 8792 48230
rect 7792 48122 8677 48174
rect 8729 48122 8792 48174
rect 7792 48066 8792 48122
rect 7792 48014 8677 48066
rect 8729 48014 8792 48066
rect 7792 47958 8792 48014
rect 7792 47906 8677 47958
rect 8729 47906 8792 47958
rect 7792 47850 8792 47906
rect 7792 47798 8677 47850
rect 8729 47798 8792 47850
rect 7792 47742 8792 47798
rect 7792 47690 8677 47742
rect 8729 47690 8792 47742
rect 7792 47634 8792 47690
rect 7792 47582 8677 47634
rect 8729 47582 8792 47634
rect 7792 47526 8792 47582
rect 7792 47474 8677 47526
rect 8729 47474 8792 47526
rect 7792 47418 8792 47474
rect 7792 47366 8677 47418
rect 8729 47366 8792 47418
rect 7792 47310 8792 47366
rect 7792 47258 8677 47310
rect 8729 47258 8792 47310
rect 7792 47202 8792 47258
rect 7792 47150 8677 47202
rect 8729 47150 8792 47202
rect 7792 47094 8792 47150
rect 7792 47042 8677 47094
rect 8729 47042 8792 47094
rect 7792 46986 8792 47042
rect 7792 46934 8677 46986
rect 8729 46934 8792 46986
rect 7792 46878 8792 46934
rect 7792 46826 8677 46878
rect 8729 46826 8792 46878
rect 7792 46770 8792 46826
rect 7792 46718 8677 46770
rect 8729 46718 8792 46770
rect 7792 46662 8792 46718
rect 7792 46610 8677 46662
rect 8729 46610 8792 46662
rect 7792 46554 8792 46610
rect 7792 46502 8677 46554
rect 8729 46502 8792 46554
rect 7792 46446 8792 46502
rect 7792 46394 8677 46446
rect 8729 46394 8792 46446
rect 7792 46338 8792 46394
rect 7792 46286 8677 46338
rect 8729 46286 8792 46338
rect 7792 46230 8792 46286
rect 7792 46178 8677 46230
rect 8729 46178 8792 46230
rect 7792 46122 8792 46178
rect 7792 46070 8677 46122
rect 8729 46070 8792 46122
rect 7792 46014 8792 46070
rect 7792 45962 8677 46014
rect 8729 45962 8792 46014
rect 7792 45906 8792 45962
rect 7792 45854 8677 45906
rect 8729 45854 8792 45906
rect 7792 45798 8792 45854
rect 7792 45746 8677 45798
rect 8729 45746 8792 45798
rect 7792 45690 8792 45746
rect 7792 45638 8677 45690
rect 8729 45638 8792 45690
rect 7792 45582 8792 45638
rect 7792 45530 8677 45582
rect 8729 45530 8792 45582
rect 7792 45474 8792 45530
rect 7792 45422 8677 45474
rect 8729 45422 8792 45474
rect 7792 45366 8792 45422
rect 7792 45319 8677 45366
rect 8729 45330 8792 45366
rect 9708 45330 10708 48374
rect 11228 48431 14144 48442
rect 11228 48385 11239 48431
rect 14133 48385 14144 48431
rect 8729 45319 10708 45330
rect 7792 45273 7803 45319
rect 10697 45273 10708 45319
rect 7792 45262 10708 45273
rect 10768 48315 11168 48352
rect 10768 45389 10779 48315
rect 10825 45389 11111 48315
rect 11157 45389 11168 48315
rect 10768 45202 11168 45389
rect 11228 48338 11283 48385
rect 11335 48376 13786 48385
rect 13838 48376 13910 48385
rect 13962 48376 14034 48385
rect 14086 48376 14144 48385
rect 11335 48374 14144 48376
rect 11335 48338 12228 48374
rect 11228 48282 12228 48338
rect 11228 48230 11283 48282
rect 11335 48230 12228 48282
rect 11228 48174 12228 48230
rect 11228 48122 11283 48174
rect 11335 48122 12228 48174
rect 11228 48066 12228 48122
rect 11228 48014 11283 48066
rect 11335 48014 12228 48066
rect 11228 47958 12228 48014
rect 11228 47906 11283 47958
rect 11335 47906 12228 47958
rect 11228 47850 12228 47906
rect 11228 47798 11283 47850
rect 11335 47798 12228 47850
rect 11228 47742 12228 47798
rect 11228 47690 11283 47742
rect 11335 47690 12228 47742
rect 11228 47634 12228 47690
rect 11228 47582 11283 47634
rect 11335 47582 12228 47634
rect 11228 47526 12228 47582
rect 11228 47474 11283 47526
rect 11335 47474 12228 47526
rect 11228 47418 12228 47474
rect 11228 47366 11283 47418
rect 11335 47366 12228 47418
rect 11228 47310 12228 47366
rect 11228 47258 11283 47310
rect 11335 47258 12228 47310
rect 11228 47202 12228 47258
rect 11228 47150 11283 47202
rect 11335 47150 12228 47202
rect 11228 47094 12228 47150
rect 11228 47042 11283 47094
rect 11335 47042 12228 47094
rect 11228 46986 12228 47042
rect 11228 46934 11283 46986
rect 11335 46934 12228 46986
rect 11228 46878 12228 46934
rect 11228 46826 11283 46878
rect 11335 46826 12228 46878
rect 11228 46770 12228 46826
rect 11228 46718 11283 46770
rect 11335 46718 12228 46770
rect 11228 46662 12228 46718
rect 11228 46610 11283 46662
rect 11335 46610 12228 46662
rect 11228 46554 12228 46610
rect 11228 46502 11283 46554
rect 11335 46502 12228 46554
rect 11228 46446 12228 46502
rect 11228 46394 11283 46446
rect 11335 46394 12228 46446
rect 11228 46338 12228 46394
rect 11228 46286 11283 46338
rect 11335 46286 12228 46338
rect 11228 46230 12228 46286
rect 11228 46178 11283 46230
rect 11335 46178 12228 46230
rect 11228 46122 12228 46178
rect 11228 46070 11283 46122
rect 11335 46070 12228 46122
rect 11228 46014 12228 46070
rect 11228 45962 11283 46014
rect 11335 45962 12228 46014
rect 11228 45906 12228 45962
rect 11228 45854 11283 45906
rect 11335 45854 12228 45906
rect 11228 45798 12228 45854
rect 11228 45746 11283 45798
rect 11335 45746 12228 45798
rect 11228 45690 12228 45746
rect 11228 45638 11283 45690
rect 11335 45638 12228 45690
rect 11228 45582 12228 45638
rect 11228 45530 11283 45582
rect 11335 45530 12228 45582
rect 11228 45474 12228 45530
rect 11228 45422 11283 45474
rect 11335 45422 12228 45474
rect 11228 45366 12228 45422
rect 11228 45319 11283 45366
rect 11335 45330 12228 45366
rect 13144 48304 14144 48374
rect 13144 48252 13786 48304
rect 13838 48252 13910 48304
rect 13962 48252 14034 48304
rect 14086 48252 14144 48304
rect 13144 48180 14144 48252
rect 13144 48128 13786 48180
rect 13838 48128 13910 48180
rect 13962 48128 14034 48180
rect 14086 48128 14144 48180
rect 13144 48056 14144 48128
rect 13144 48004 13786 48056
rect 13838 48004 13910 48056
rect 13962 48004 14034 48056
rect 14086 48004 14144 48056
rect 13144 47932 14144 48004
rect 13144 47880 13786 47932
rect 13838 47880 13910 47932
rect 13962 47880 14034 47932
rect 14086 47880 14144 47932
rect 13144 47808 14144 47880
rect 13144 47756 13786 47808
rect 13838 47756 13910 47808
rect 13962 47756 14034 47808
rect 14086 47756 14144 47808
rect 13144 47684 14144 47756
rect 13144 47632 13786 47684
rect 13838 47632 13910 47684
rect 13962 47632 14034 47684
rect 14086 47632 14144 47684
rect 13144 47560 14144 47632
rect 13144 47508 13786 47560
rect 13838 47508 13910 47560
rect 13962 47508 14034 47560
rect 14086 47508 14144 47560
rect 13144 47436 14144 47508
rect 13144 47384 13786 47436
rect 13838 47384 13910 47436
rect 13962 47384 14034 47436
rect 14086 47384 14144 47436
rect 13144 47312 14144 47384
rect 13144 47260 13786 47312
rect 13838 47260 13910 47312
rect 13962 47260 14034 47312
rect 14086 47260 14144 47312
rect 13144 47188 14144 47260
rect 13144 47136 13786 47188
rect 13838 47136 13910 47188
rect 13962 47136 14034 47188
rect 14086 47136 14144 47188
rect 13144 47064 14144 47136
rect 13144 47012 13786 47064
rect 13838 47012 13910 47064
rect 13962 47012 14034 47064
rect 14086 47012 14144 47064
rect 13144 46940 14144 47012
rect 13144 46888 13786 46940
rect 13838 46888 13910 46940
rect 13962 46888 14034 46940
rect 14086 46888 14144 46940
rect 13144 46816 14144 46888
rect 13144 46764 13786 46816
rect 13838 46764 13910 46816
rect 13962 46764 14034 46816
rect 14086 46764 14144 46816
rect 13144 46692 14144 46764
rect 13144 46640 13786 46692
rect 13838 46640 13910 46692
rect 13962 46640 14034 46692
rect 14086 46640 14144 46692
rect 13144 46568 14144 46640
rect 13144 46516 13786 46568
rect 13838 46516 13910 46568
rect 13962 46516 14034 46568
rect 14086 46516 14144 46568
rect 13144 46444 14144 46516
rect 13144 46392 13786 46444
rect 13838 46392 13910 46444
rect 13962 46392 14034 46444
rect 14086 46392 14144 46444
rect 13144 46320 14144 46392
rect 13144 46268 13786 46320
rect 13838 46268 13910 46320
rect 13962 46268 14034 46320
rect 14086 46268 14144 46320
rect 13144 46196 14144 46268
rect 13144 46144 13786 46196
rect 13838 46144 13910 46196
rect 13962 46144 14034 46196
rect 14086 46144 14144 46196
rect 13144 46072 14144 46144
rect 13144 46020 13786 46072
rect 13838 46020 13910 46072
rect 13962 46020 14034 46072
rect 14086 46020 14144 46072
rect 13144 45948 14144 46020
rect 13144 45896 13786 45948
rect 13838 45896 13910 45948
rect 13962 45896 14034 45948
rect 14086 45896 14144 45948
rect 13144 45824 14144 45896
rect 13144 45772 13786 45824
rect 13838 45772 13910 45824
rect 13962 45772 14034 45824
rect 14086 45772 14144 45824
rect 13144 45700 14144 45772
rect 13144 45648 13786 45700
rect 13838 45648 13910 45700
rect 13962 45648 14034 45700
rect 14086 45648 14144 45700
rect 13144 45576 14144 45648
rect 13144 45524 13786 45576
rect 13838 45524 13910 45576
rect 13962 45524 14034 45576
rect 14086 45524 14144 45576
rect 13144 45452 14144 45524
rect 13144 45400 13786 45452
rect 13838 45400 13910 45452
rect 13962 45400 14034 45452
rect 14086 45400 14144 45452
rect 13144 45330 14144 45400
rect 11335 45328 14144 45330
rect 11335 45319 13786 45328
rect 13838 45319 13910 45328
rect 13962 45319 14034 45328
rect 14086 45319 14144 45328
rect 11228 45273 11239 45319
rect 14133 45273 14144 45319
rect 11228 45262 14144 45273
rect 14204 48315 14404 48352
rect 14204 45389 14215 48315
rect 14261 45389 14404 48315
rect 14204 45202 14404 45389
rect 14608 45202 14619 48502
rect 445 45152 14619 45202
rect 445 45120 1438 45152
rect 496 45068 552 45120
rect 604 45068 660 45120
rect 712 45100 1438 45120
rect 1490 45100 1562 45152
rect 1614 45100 1686 45152
rect 1738 45100 1810 45152
rect 1862 45100 2574 45152
rect 2626 45100 2698 45152
rect 2750 45100 2822 45152
rect 2874 45100 2946 45152
rect 2998 45100 4846 45152
rect 4898 45100 4970 45152
rect 5022 45100 5094 45152
rect 5146 45100 5218 45152
rect 5270 45100 7139 45152
rect 7191 45100 7263 45152
rect 7315 45100 7387 45152
rect 7439 45100 7625 45152
rect 7677 45100 7749 45152
rect 7801 45100 7873 45152
rect 7925 45100 9794 45152
rect 9846 45100 9918 45152
rect 9970 45100 10042 45152
rect 10094 45100 10166 45152
rect 10218 45100 12066 45152
rect 12118 45100 12190 45152
rect 12242 45100 12314 45152
rect 12366 45100 12438 45152
rect 12490 45100 13480 45152
rect 13532 45100 13604 45152
rect 13656 45120 14619 45152
rect 13656 45100 14352 45120
rect 712 45068 14352 45100
rect 14404 45068 14460 45120
rect 14512 45068 14568 45120
rect 445 45028 14619 45068
rect 445 45012 1438 45028
rect 496 44960 552 45012
rect 604 44960 660 45012
rect 712 44976 1438 45012
rect 1490 44976 1562 45028
rect 1614 44976 1686 45028
rect 1738 44976 1810 45028
rect 1862 44976 2574 45028
rect 2626 44976 2698 45028
rect 2750 44976 2822 45028
rect 2874 44976 2946 45028
rect 2998 44976 4846 45028
rect 4898 44976 4970 45028
rect 5022 44976 5094 45028
rect 5146 44976 5218 45028
rect 5270 44976 7139 45028
rect 7191 44976 7263 45028
rect 7315 44976 7387 45028
rect 7439 44976 7625 45028
rect 7677 44976 7749 45028
rect 7801 44976 7873 45028
rect 7925 44976 9794 45028
rect 9846 44976 9918 45028
rect 9970 44976 10042 45028
rect 10094 44976 10166 45028
rect 10218 44976 12066 45028
rect 12118 44976 12190 45028
rect 12242 44976 12314 45028
rect 12366 44976 12438 45028
rect 12490 44976 13480 45028
rect 13532 44976 13604 45028
rect 13656 45012 14619 45028
rect 13656 44976 14352 45012
rect 712 44960 14352 44976
rect 14404 44960 14460 45012
rect 14512 44960 14568 45012
rect 445 44904 14619 44960
rect 496 44852 552 44904
rect 604 44901 660 44904
rect 712 44901 1438 44904
rect 1490 44901 1562 44904
rect 1614 44901 1686 44904
rect 1738 44901 1810 44904
rect 1862 44901 2574 44904
rect 2626 44901 2698 44904
rect 2750 44901 2822 44904
rect 2874 44901 2946 44904
rect 2998 44901 4846 44904
rect 4898 44901 4970 44904
rect 5022 44901 5094 44904
rect 5146 44901 5218 44904
rect 5270 44901 7139 44904
rect 7191 44901 7263 44904
rect 7315 44901 7387 44904
rect 7439 44901 7625 44904
rect 7677 44901 7749 44904
rect 7801 44901 7873 44904
rect 7925 44901 9794 44904
rect 9846 44901 9918 44904
rect 9970 44901 10042 44904
rect 10094 44901 10166 44904
rect 10218 44901 12066 44904
rect 12118 44901 12190 44904
rect 12242 44901 12314 44904
rect 12366 44901 12438 44904
rect 12490 44901 13480 44904
rect 13532 44901 13604 44904
rect 13656 44901 14352 44904
rect 14404 44901 14460 44904
rect 604 44852 660 44855
rect 712 44852 1438 44855
rect 1490 44852 1562 44855
rect 1614 44852 1686 44855
rect 1738 44852 1810 44855
rect 1862 44852 2574 44855
rect 2626 44852 2698 44855
rect 2750 44852 2822 44855
rect 2874 44852 2946 44855
rect 2998 44852 4846 44855
rect 4898 44852 4970 44855
rect 5022 44852 5094 44855
rect 5146 44852 5218 44855
rect 5270 44852 7139 44855
rect 7191 44852 7263 44855
rect 7315 44852 7387 44855
rect 7439 44852 7625 44855
rect 7677 44852 7749 44855
rect 7801 44852 7873 44855
rect 7925 44852 9794 44855
rect 9846 44852 9918 44855
rect 9970 44852 10042 44855
rect 10094 44852 10166 44855
rect 10218 44852 12066 44855
rect 12118 44852 12190 44855
rect 12242 44852 12314 44855
rect 12366 44852 12438 44855
rect 12490 44852 13480 44855
rect 13532 44852 13604 44855
rect 13656 44852 14352 44855
rect 14404 44852 14460 44855
rect 14512 44852 14568 44904
rect 445 44796 14619 44852
rect 496 44744 552 44796
rect 604 44744 660 44796
rect 712 44780 14352 44796
rect 712 44744 1438 44780
rect 445 44728 1438 44744
rect 1490 44728 1562 44780
rect 1614 44728 1686 44780
rect 1738 44728 1810 44780
rect 1862 44728 2574 44780
rect 2626 44728 2698 44780
rect 2750 44728 2822 44780
rect 2874 44728 2946 44780
rect 2998 44728 4846 44780
rect 4898 44728 4970 44780
rect 5022 44728 5094 44780
rect 5146 44728 5218 44780
rect 5270 44728 7139 44780
rect 7191 44728 7263 44780
rect 7315 44728 7387 44780
rect 7439 44728 7625 44780
rect 7677 44728 7749 44780
rect 7801 44728 7873 44780
rect 7925 44728 9794 44780
rect 9846 44728 9918 44780
rect 9970 44728 10042 44780
rect 10094 44728 10166 44780
rect 10218 44728 12066 44780
rect 12118 44728 12190 44780
rect 12242 44728 12314 44780
rect 12366 44728 12438 44780
rect 12490 44728 13480 44780
rect 13532 44728 13604 44780
rect 13656 44744 14352 44780
rect 14404 44744 14460 44796
rect 14512 44744 14568 44796
rect 13656 44728 14619 44744
rect 445 44688 14619 44728
rect 496 44636 552 44688
rect 604 44636 660 44688
rect 712 44656 14352 44688
rect 712 44636 1438 44656
rect 445 44604 1438 44636
rect 1490 44604 1562 44656
rect 1614 44604 1686 44656
rect 1738 44604 1810 44656
rect 1862 44604 2574 44656
rect 2626 44604 2698 44656
rect 2750 44604 2822 44656
rect 2874 44604 2946 44656
rect 2998 44604 4846 44656
rect 4898 44604 4970 44656
rect 5022 44604 5094 44656
rect 5146 44604 5218 44656
rect 5270 44604 7139 44656
rect 7191 44604 7263 44656
rect 7315 44604 7387 44656
rect 7439 44604 7625 44656
rect 7677 44604 7749 44656
rect 7801 44604 7873 44656
rect 7925 44604 9794 44656
rect 9846 44604 9918 44656
rect 9970 44604 10042 44656
rect 10094 44604 10166 44656
rect 10218 44604 12066 44656
rect 12118 44604 12190 44656
rect 12242 44604 12314 44656
rect 12366 44604 12438 44656
rect 12490 44604 13480 44656
rect 13532 44604 13604 44656
rect 13656 44636 14352 44656
rect 14404 44636 14460 44688
rect 14512 44636 14568 44688
rect 13656 44604 14619 44636
rect 445 44554 14619 44604
rect 445 41254 456 44554
rect 920 44483 3836 44494
rect 920 44437 931 44483
rect 3825 44437 3836 44483
rect 920 44428 1148 44437
rect 1200 44428 1272 44437
rect 1324 44428 3729 44437
rect 920 44426 3729 44428
rect 660 44367 860 44404
rect 660 41441 803 44367
rect 849 41441 860 44367
rect 660 41254 860 41441
rect 920 44356 1920 44426
rect 920 44304 1148 44356
rect 1200 44304 1272 44356
rect 1324 44304 1920 44356
rect 920 44232 1920 44304
rect 920 44180 1148 44232
rect 1200 44180 1272 44232
rect 1324 44180 1920 44232
rect 920 44108 1920 44180
rect 920 44056 1148 44108
rect 1200 44056 1272 44108
rect 1324 44056 1920 44108
rect 920 43984 1920 44056
rect 920 43932 1148 43984
rect 1200 43932 1272 43984
rect 1324 43932 1920 43984
rect 920 43860 1920 43932
rect 920 43808 1148 43860
rect 1200 43808 1272 43860
rect 1324 43808 1920 43860
rect 920 43736 1920 43808
rect 920 43684 1148 43736
rect 1200 43684 1272 43736
rect 1324 43684 1920 43736
rect 920 43612 1920 43684
rect 920 43560 1148 43612
rect 1200 43560 1272 43612
rect 1324 43560 1920 43612
rect 920 43488 1920 43560
rect 920 43436 1148 43488
rect 1200 43436 1272 43488
rect 1324 43436 1920 43488
rect 920 43364 1920 43436
rect 920 43312 1148 43364
rect 1200 43312 1272 43364
rect 1324 43312 1920 43364
rect 920 43240 1920 43312
rect 920 43188 1148 43240
rect 1200 43188 1272 43240
rect 1324 43188 1920 43240
rect 920 43116 1920 43188
rect 920 43064 1148 43116
rect 1200 43064 1272 43116
rect 1324 43064 1920 43116
rect 920 42992 1920 43064
rect 920 42940 1148 42992
rect 1200 42940 1272 42992
rect 1324 42940 1920 42992
rect 920 42868 1920 42940
rect 920 42816 1148 42868
rect 1200 42816 1272 42868
rect 1324 42816 1920 42868
rect 920 42744 1920 42816
rect 920 42692 1148 42744
rect 1200 42692 1272 42744
rect 1324 42692 1920 42744
rect 920 42620 1920 42692
rect 920 42568 1148 42620
rect 1200 42568 1272 42620
rect 1324 42568 1920 42620
rect 920 42496 1920 42568
rect 920 42444 1148 42496
rect 1200 42444 1272 42496
rect 1324 42444 1920 42496
rect 920 42372 1920 42444
rect 920 42320 1148 42372
rect 1200 42320 1272 42372
rect 1324 42320 1920 42372
rect 920 42248 1920 42320
rect 920 42196 1148 42248
rect 1200 42196 1272 42248
rect 1324 42196 1920 42248
rect 920 42124 1920 42196
rect 920 42072 1148 42124
rect 1200 42072 1272 42124
rect 1324 42072 1920 42124
rect 920 42000 1920 42072
rect 920 41948 1148 42000
rect 1200 41948 1272 42000
rect 1324 41948 1920 42000
rect 920 41876 1920 41948
rect 920 41824 1148 41876
rect 1200 41824 1272 41876
rect 1324 41824 1920 41876
rect 920 41752 1920 41824
rect 920 41700 1148 41752
rect 1200 41700 1272 41752
rect 1324 41700 1920 41752
rect 920 41628 1920 41700
rect 920 41576 1148 41628
rect 1200 41576 1272 41628
rect 1324 41576 1920 41628
rect 920 41504 1920 41576
rect 920 41452 1148 41504
rect 1200 41452 1272 41504
rect 1324 41452 1920 41504
rect 920 41382 1920 41452
rect 2836 44390 3729 44426
rect 3781 44390 3836 44437
rect 4356 44483 7272 44494
rect 4356 44437 4367 44483
rect 7261 44437 7272 44483
rect 4356 44426 6335 44437
rect 2836 44334 3836 44390
rect 2836 44282 3729 44334
rect 3781 44282 3836 44334
rect 2836 44226 3836 44282
rect 2836 44174 3729 44226
rect 3781 44174 3836 44226
rect 2836 44118 3836 44174
rect 2836 44066 3729 44118
rect 3781 44066 3836 44118
rect 2836 44010 3836 44066
rect 2836 43958 3729 44010
rect 3781 43958 3836 44010
rect 2836 43902 3836 43958
rect 2836 43850 3729 43902
rect 3781 43850 3836 43902
rect 2836 43794 3836 43850
rect 2836 43742 3729 43794
rect 3781 43742 3836 43794
rect 2836 43686 3836 43742
rect 2836 43634 3729 43686
rect 3781 43634 3836 43686
rect 2836 43578 3836 43634
rect 2836 43526 3729 43578
rect 3781 43526 3836 43578
rect 2836 43470 3836 43526
rect 2836 43418 3729 43470
rect 3781 43418 3836 43470
rect 2836 43362 3836 43418
rect 2836 43310 3729 43362
rect 3781 43310 3836 43362
rect 2836 43254 3836 43310
rect 2836 43202 3729 43254
rect 3781 43202 3836 43254
rect 2836 43146 3836 43202
rect 2836 43094 3729 43146
rect 3781 43094 3836 43146
rect 2836 43038 3836 43094
rect 2836 42986 3729 43038
rect 3781 42986 3836 43038
rect 2836 42930 3836 42986
rect 2836 42878 3729 42930
rect 3781 42878 3836 42930
rect 2836 42822 3836 42878
rect 2836 42770 3729 42822
rect 3781 42770 3836 42822
rect 2836 42714 3836 42770
rect 2836 42662 3729 42714
rect 3781 42662 3836 42714
rect 2836 42606 3836 42662
rect 2836 42554 3729 42606
rect 3781 42554 3836 42606
rect 2836 42498 3836 42554
rect 2836 42446 3729 42498
rect 3781 42446 3836 42498
rect 2836 42390 3836 42446
rect 2836 42338 3729 42390
rect 3781 42338 3836 42390
rect 2836 42282 3836 42338
rect 2836 42230 3729 42282
rect 3781 42230 3836 42282
rect 2836 42174 3836 42230
rect 2836 42122 3729 42174
rect 3781 42122 3836 42174
rect 2836 42066 3836 42122
rect 2836 42014 3729 42066
rect 3781 42014 3836 42066
rect 2836 41958 3836 42014
rect 2836 41906 3729 41958
rect 3781 41906 3836 41958
rect 2836 41850 3836 41906
rect 2836 41798 3729 41850
rect 3781 41798 3836 41850
rect 2836 41742 3836 41798
rect 2836 41690 3729 41742
rect 3781 41690 3836 41742
rect 2836 41634 3836 41690
rect 2836 41582 3729 41634
rect 3781 41582 3836 41634
rect 2836 41526 3836 41582
rect 2836 41474 3729 41526
rect 3781 41474 3836 41526
rect 2836 41418 3836 41474
rect 2836 41382 3729 41418
rect 920 41380 3729 41382
rect 920 41371 1148 41380
rect 1200 41371 1272 41380
rect 1324 41371 3729 41380
rect 3781 41371 3836 41418
rect 920 41325 931 41371
rect 3825 41325 3836 41371
rect 920 41314 3836 41325
rect 3896 44367 4296 44404
rect 3896 41441 3907 44367
rect 3953 41441 4239 44367
rect 4285 41441 4296 44367
rect 3896 41254 4296 41441
rect 4356 41382 5356 44426
rect 6272 44390 6335 44426
rect 6387 44390 7272 44437
rect 7792 44483 10708 44494
rect 7792 44437 7803 44483
rect 10697 44437 10708 44483
rect 6272 44334 7272 44390
rect 6272 44282 6335 44334
rect 6387 44282 7272 44334
rect 6272 44226 7272 44282
rect 6272 44174 6335 44226
rect 6387 44174 7272 44226
rect 6272 44118 7272 44174
rect 6272 44066 6335 44118
rect 6387 44066 7272 44118
rect 6272 44010 7272 44066
rect 6272 43958 6335 44010
rect 6387 43958 7272 44010
rect 6272 43902 7272 43958
rect 6272 43850 6335 43902
rect 6387 43850 7272 43902
rect 6272 43794 7272 43850
rect 6272 43742 6335 43794
rect 6387 43742 7272 43794
rect 6272 43686 7272 43742
rect 6272 43634 6335 43686
rect 6387 43634 7272 43686
rect 6272 43578 7272 43634
rect 6272 43526 6335 43578
rect 6387 43526 7272 43578
rect 6272 43470 7272 43526
rect 6272 43418 6335 43470
rect 6387 43418 7272 43470
rect 6272 43362 7272 43418
rect 6272 43310 6335 43362
rect 6387 43310 7272 43362
rect 6272 43254 7272 43310
rect 6272 43202 6335 43254
rect 6387 43202 7272 43254
rect 6272 43146 7272 43202
rect 6272 43094 6335 43146
rect 6387 43094 7272 43146
rect 6272 43038 7272 43094
rect 6272 42986 6335 43038
rect 6387 42986 7272 43038
rect 6272 42930 7272 42986
rect 6272 42878 6335 42930
rect 6387 42878 7272 42930
rect 6272 42822 7272 42878
rect 6272 42770 6335 42822
rect 6387 42770 7272 42822
rect 6272 42714 7272 42770
rect 6272 42662 6335 42714
rect 6387 42662 7272 42714
rect 6272 42606 7272 42662
rect 6272 42554 6335 42606
rect 6387 42554 7272 42606
rect 6272 42498 7272 42554
rect 6272 42446 6335 42498
rect 6387 42446 7272 42498
rect 6272 42390 7272 42446
rect 6272 42338 6335 42390
rect 6387 42338 7272 42390
rect 6272 42282 7272 42338
rect 6272 42230 6335 42282
rect 6387 42230 7272 42282
rect 6272 42174 7272 42230
rect 6272 42122 6335 42174
rect 6387 42122 7272 42174
rect 6272 42066 7272 42122
rect 6272 42014 6335 42066
rect 6387 42014 7272 42066
rect 6272 41958 7272 42014
rect 6272 41906 6335 41958
rect 6387 41906 7272 41958
rect 6272 41850 7272 41906
rect 6272 41798 6335 41850
rect 6387 41798 7272 41850
rect 6272 41742 7272 41798
rect 6272 41690 6335 41742
rect 6387 41690 7272 41742
rect 6272 41634 7272 41690
rect 6272 41582 6335 41634
rect 6387 41582 7272 41634
rect 6272 41526 7272 41582
rect 6272 41474 6335 41526
rect 6387 41474 7272 41526
rect 6272 41418 7272 41474
rect 6272 41382 6335 41418
rect 4356 41371 6335 41382
rect 6387 41371 7272 41418
rect 4356 41325 4367 41371
rect 7261 41325 7272 41371
rect 4356 41314 7272 41325
rect 7332 44388 7732 44404
rect 7332 44367 7388 44388
rect 7332 41441 7343 44367
rect 7440 44336 7624 44388
rect 7676 44367 7732 44388
rect 7389 44280 7675 44336
rect 7440 44228 7624 44280
rect 7389 44172 7675 44228
rect 7440 44120 7624 44172
rect 7389 44064 7675 44120
rect 7440 44012 7624 44064
rect 7389 43956 7675 44012
rect 7440 43904 7624 43956
rect 7389 43848 7675 43904
rect 7440 43796 7624 43848
rect 7389 43740 7675 43796
rect 7440 43688 7624 43740
rect 7389 43632 7675 43688
rect 7440 43580 7624 43632
rect 7389 43524 7675 43580
rect 7440 43472 7624 43524
rect 7389 43416 7675 43472
rect 7440 43364 7624 43416
rect 7389 43308 7675 43364
rect 7440 43256 7624 43308
rect 7389 43200 7675 43256
rect 7440 43148 7624 43200
rect 7389 43092 7675 43148
rect 7440 43040 7624 43092
rect 7389 42984 7675 43040
rect 7440 42932 7624 42984
rect 7389 42876 7675 42932
rect 7440 42824 7624 42876
rect 7389 42768 7675 42824
rect 7440 42716 7624 42768
rect 7389 42660 7675 42716
rect 7440 42608 7624 42660
rect 7389 42552 7675 42608
rect 7440 42500 7624 42552
rect 7389 42444 7675 42500
rect 7440 42392 7624 42444
rect 7389 42336 7675 42392
rect 7440 42284 7624 42336
rect 7389 42228 7675 42284
rect 7440 42176 7624 42228
rect 7389 42120 7675 42176
rect 7440 42068 7624 42120
rect 7389 42012 7675 42068
rect 7440 41960 7624 42012
rect 7389 41904 7675 41960
rect 7440 41852 7624 41904
rect 7389 41796 7675 41852
rect 7440 41744 7624 41796
rect 7389 41688 7675 41744
rect 7440 41636 7624 41688
rect 7389 41580 7675 41636
rect 7440 41528 7624 41580
rect 7389 41472 7675 41528
rect 7332 41420 7388 41441
rect 7440 41420 7624 41472
rect 7721 41441 7732 44367
rect 7676 41420 7732 41441
rect 7332 41254 7732 41420
rect 7792 44390 8677 44437
rect 8729 44426 10708 44437
rect 8729 44390 8792 44426
rect 7792 44334 8792 44390
rect 7792 44282 8677 44334
rect 8729 44282 8792 44334
rect 7792 44226 8792 44282
rect 7792 44174 8677 44226
rect 8729 44174 8792 44226
rect 7792 44118 8792 44174
rect 7792 44066 8677 44118
rect 8729 44066 8792 44118
rect 7792 44010 8792 44066
rect 7792 43958 8677 44010
rect 8729 43958 8792 44010
rect 7792 43902 8792 43958
rect 7792 43850 8677 43902
rect 8729 43850 8792 43902
rect 7792 43794 8792 43850
rect 7792 43742 8677 43794
rect 8729 43742 8792 43794
rect 7792 43686 8792 43742
rect 7792 43634 8677 43686
rect 8729 43634 8792 43686
rect 7792 43578 8792 43634
rect 7792 43526 8677 43578
rect 8729 43526 8792 43578
rect 7792 43470 8792 43526
rect 7792 43418 8677 43470
rect 8729 43418 8792 43470
rect 7792 43362 8792 43418
rect 7792 43310 8677 43362
rect 8729 43310 8792 43362
rect 7792 43254 8792 43310
rect 7792 43202 8677 43254
rect 8729 43202 8792 43254
rect 7792 43146 8792 43202
rect 7792 43094 8677 43146
rect 8729 43094 8792 43146
rect 7792 43038 8792 43094
rect 7792 42986 8677 43038
rect 8729 42986 8792 43038
rect 7792 42930 8792 42986
rect 7792 42878 8677 42930
rect 8729 42878 8792 42930
rect 7792 42822 8792 42878
rect 7792 42770 8677 42822
rect 8729 42770 8792 42822
rect 7792 42714 8792 42770
rect 7792 42662 8677 42714
rect 8729 42662 8792 42714
rect 7792 42606 8792 42662
rect 7792 42554 8677 42606
rect 8729 42554 8792 42606
rect 7792 42498 8792 42554
rect 7792 42446 8677 42498
rect 8729 42446 8792 42498
rect 7792 42390 8792 42446
rect 7792 42338 8677 42390
rect 8729 42338 8792 42390
rect 7792 42282 8792 42338
rect 7792 42230 8677 42282
rect 8729 42230 8792 42282
rect 7792 42174 8792 42230
rect 7792 42122 8677 42174
rect 8729 42122 8792 42174
rect 7792 42066 8792 42122
rect 7792 42014 8677 42066
rect 8729 42014 8792 42066
rect 7792 41958 8792 42014
rect 7792 41906 8677 41958
rect 8729 41906 8792 41958
rect 7792 41850 8792 41906
rect 7792 41798 8677 41850
rect 8729 41798 8792 41850
rect 7792 41742 8792 41798
rect 7792 41690 8677 41742
rect 8729 41690 8792 41742
rect 7792 41634 8792 41690
rect 7792 41582 8677 41634
rect 8729 41582 8792 41634
rect 7792 41526 8792 41582
rect 7792 41474 8677 41526
rect 8729 41474 8792 41526
rect 7792 41418 8792 41474
rect 7792 41371 8677 41418
rect 8729 41382 8792 41418
rect 9708 41382 10708 44426
rect 11228 44483 14144 44494
rect 11228 44437 11239 44483
rect 14133 44437 14144 44483
rect 8729 41371 10708 41382
rect 7792 41325 7803 41371
rect 10697 41325 10708 41371
rect 7792 41314 10708 41325
rect 10768 44367 11168 44404
rect 10768 41441 10779 44367
rect 10825 41441 11111 44367
rect 11157 41441 11168 44367
rect 10768 41254 11168 41441
rect 11228 44390 11283 44437
rect 11335 44428 13786 44437
rect 13838 44428 13910 44437
rect 13962 44428 14034 44437
rect 14086 44428 14144 44437
rect 11335 44426 14144 44428
rect 11335 44390 12228 44426
rect 11228 44334 12228 44390
rect 11228 44282 11283 44334
rect 11335 44282 12228 44334
rect 11228 44226 12228 44282
rect 11228 44174 11283 44226
rect 11335 44174 12228 44226
rect 11228 44118 12228 44174
rect 11228 44066 11283 44118
rect 11335 44066 12228 44118
rect 11228 44010 12228 44066
rect 11228 43958 11283 44010
rect 11335 43958 12228 44010
rect 11228 43902 12228 43958
rect 11228 43850 11283 43902
rect 11335 43850 12228 43902
rect 11228 43794 12228 43850
rect 11228 43742 11283 43794
rect 11335 43742 12228 43794
rect 11228 43686 12228 43742
rect 11228 43634 11283 43686
rect 11335 43634 12228 43686
rect 11228 43578 12228 43634
rect 11228 43526 11283 43578
rect 11335 43526 12228 43578
rect 11228 43470 12228 43526
rect 11228 43418 11283 43470
rect 11335 43418 12228 43470
rect 11228 43362 12228 43418
rect 11228 43310 11283 43362
rect 11335 43310 12228 43362
rect 11228 43254 12228 43310
rect 11228 43202 11283 43254
rect 11335 43202 12228 43254
rect 11228 43146 12228 43202
rect 11228 43094 11283 43146
rect 11335 43094 12228 43146
rect 11228 43038 12228 43094
rect 11228 42986 11283 43038
rect 11335 42986 12228 43038
rect 11228 42930 12228 42986
rect 11228 42878 11283 42930
rect 11335 42878 12228 42930
rect 11228 42822 12228 42878
rect 11228 42770 11283 42822
rect 11335 42770 12228 42822
rect 11228 42714 12228 42770
rect 11228 42662 11283 42714
rect 11335 42662 12228 42714
rect 11228 42606 12228 42662
rect 11228 42554 11283 42606
rect 11335 42554 12228 42606
rect 11228 42498 12228 42554
rect 11228 42446 11283 42498
rect 11335 42446 12228 42498
rect 11228 42390 12228 42446
rect 11228 42338 11283 42390
rect 11335 42338 12228 42390
rect 11228 42282 12228 42338
rect 11228 42230 11283 42282
rect 11335 42230 12228 42282
rect 11228 42174 12228 42230
rect 11228 42122 11283 42174
rect 11335 42122 12228 42174
rect 11228 42066 12228 42122
rect 11228 42014 11283 42066
rect 11335 42014 12228 42066
rect 11228 41958 12228 42014
rect 11228 41906 11283 41958
rect 11335 41906 12228 41958
rect 11228 41850 12228 41906
rect 11228 41798 11283 41850
rect 11335 41798 12228 41850
rect 11228 41742 12228 41798
rect 11228 41690 11283 41742
rect 11335 41690 12228 41742
rect 11228 41634 12228 41690
rect 11228 41582 11283 41634
rect 11335 41582 12228 41634
rect 11228 41526 12228 41582
rect 11228 41474 11283 41526
rect 11335 41474 12228 41526
rect 11228 41418 12228 41474
rect 11228 41371 11283 41418
rect 11335 41382 12228 41418
rect 13144 44356 14144 44426
rect 13144 44304 13786 44356
rect 13838 44304 13910 44356
rect 13962 44304 14034 44356
rect 14086 44304 14144 44356
rect 13144 44232 14144 44304
rect 13144 44180 13786 44232
rect 13838 44180 13910 44232
rect 13962 44180 14034 44232
rect 14086 44180 14144 44232
rect 13144 44108 14144 44180
rect 13144 44056 13786 44108
rect 13838 44056 13910 44108
rect 13962 44056 14034 44108
rect 14086 44056 14144 44108
rect 13144 43984 14144 44056
rect 13144 43932 13786 43984
rect 13838 43932 13910 43984
rect 13962 43932 14034 43984
rect 14086 43932 14144 43984
rect 13144 43860 14144 43932
rect 13144 43808 13786 43860
rect 13838 43808 13910 43860
rect 13962 43808 14034 43860
rect 14086 43808 14144 43860
rect 13144 43736 14144 43808
rect 13144 43684 13786 43736
rect 13838 43684 13910 43736
rect 13962 43684 14034 43736
rect 14086 43684 14144 43736
rect 13144 43612 14144 43684
rect 13144 43560 13786 43612
rect 13838 43560 13910 43612
rect 13962 43560 14034 43612
rect 14086 43560 14144 43612
rect 13144 43488 14144 43560
rect 13144 43436 13786 43488
rect 13838 43436 13910 43488
rect 13962 43436 14034 43488
rect 14086 43436 14144 43488
rect 13144 43364 14144 43436
rect 13144 43312 13786 43364
rect 13838 43312 13910 43364
rect 13962 43312 14034 43364
rect 14086 43312 14144 43364
rect 13144 43240 14144 43312
rect 13144 43188 13786 43240
rect 13838 43188 13910 43240
rect 13962 43188 14034 43240
rect 14086 43188 14144 43240
rect 13144 43116 14144 43188
rect 13144 43064 13786 43116
rect 13838 43064 13910 43116
rect 13962 43064 14034 43116
rect 14086 43064 14144 43116
rect 13144 42992 14144 43064
rect 13144 42940 13786 42992
rect 13838 42940 13910 42992
rect 13962 42940 14034 42992
rect 14086 42940 14144 42992
rect 13144 42868 14144 42940
rect 13144 42816 13786 42868
rect 13838 42816 13910 42868
rect 13962 42816 14034 42868
rect 14086 42816 14144 42868
rect 13144 42744 14144 42816
rect 13144 42692 13786 42744
rect 13838 42692 13910 42744
rect 13962 42692 14034 42744
rect 14086 42692 14144 42744
rect 13144 42620 14144 42692
rect 13144 42568 13786 42620
rect 13838 42568 13910 42620
rect 13962 42568 14034 42620
rect 14086 42568 14144 42620
rect 13144 42496 14144 42568
rect 13144 42444 13786 42496
rect 13838 42444 13910 42496
rect 13962 42444 14034 42496
rect 14086 42444 14144 42496
rect 13144 42372 14144 42444
rect 13144 42320 13786 42372
rect 13838 42320 13910 42372
rect 13962 42320 14034 42372
rect 14086 42320 14144 42372
rect 13144 42248 14144 42320
rect 13144 42196 13786 42248
rect 13838 42196 13910 42248
rect 13962 42196 14034 42248
rect 14086 42196 14144 42248
rect 13144 42124 14144 42196
rect 13144 42072 13786 42124
rect 13838 42072 13910 42124
rect 13962 42072 14034 42124
rect 14086 42072 14144 42124
rect 13144 42000 14144 42072
rect 13144 41948 13786 42000
rect 13838 41948 13910 42000
rect 13962 41948 14034 42000
rect 14086 41948 14144 42000
rect 13144 41876 14144 41948
rect 13144 41824 13786 41876
rect 13838 41824 13910 41876
rect 13962 41824 14034 41876
rect 14086 41824 14144 41876
rect 13144 41752 14144 41824
rect 13144 41700 13786 41752
rect 13838 41700 13910 41752
rect 13962 41700 14034 41752
rect 14086 41700 14144 41752
rect 13144 41628 14144 41700
rect 13144 41576 13786 41628
rect 13838 41576 13910 41628
rect 13962 41576 14034 41628
rect 14086 41576 14144 41628
rect 13144 41504 14144 41576
rect 13144 41452 13786 41504
rect 13838 41452 13910 41504
rect 13962 41452 14034 41504
rect 14086 41452 14144 41504
rect 13144 41382 14144 41452
rect 11335 41380 14144 41382
rect 11335 41371 13786 41380
rect 13838 41371 13910 41380
rect 13962 41371 14034 41380
rect 14086 41371 14144 41380
rect 11228 41325 11239 41371
rect 14133 41325 14144 41371
rect 11228 41314 14144 41325
rect 14204 44367 14404 44404
rect 14204 41441 14215 44367
rect 14261 41441 14404 44367
rect 14204 41254 14404 41441
rect 14608 41254 14619 44554
rect 445 41204 14619 41254
rect 445 41172 1438 41204
rect 496 41120 552 41172
rect 604 41120 660 41172
rect 712 41152 1438 41172
rect 1490 41152 1562 41204
rect 1614 41152 1686 41204
rect 1738 41152 1810 41204
rect 1862 41152 2574 41204
rect 2626 41152 2698 41204
rect 2750 41152 2822 41204
rect 2874 41152 2946 41204
rect 2998 41152 4846 41204
rect 4898 41152 4970 41204
rect 5022 41152 5094 41204
rect 5146 41152 5218 41204
rect 5270 41152 7139 41204
rect 7191 41152 7263 41204
rect 7315 41152 7387 41204
rect 7439 41152 7625 41204
rect 7677 41152 7749 41204
rect 7801 41152 7873 41204
rect 7925 41152 9794 41204
rect 9846 41152 9918 41204
rect 9970 41152 10042 41204
rect 10094 41152 10166 41204
rect 10218 41152 12066 41204
rect 12118 41152 12190 41204
rect 12242 41152 12314 41204
rect 12366 41152 12438 41204
rect 12490 41152 13480 41204
rect 13532 41152 13604 41204
rect 13656 41172 14619 41204
rect 13656 41152 14352 41172
rect 712 41120 14352 41152
rect 14404 41120 14460 41172
rect 14512 41120 14568 41172
rect 445 41080 14619 41120
rect 445 41064 1438 41080
rect 496 41012 552 41064
rect 604 41012 660 41064
rect 712 41028 1438 41064
rect 1490 41028 1562 41080
rect 1614 41028 1686 41080
rect 1738 41028 1810 41080
rect 1862 41028 2574 41080
rect 2626 41028 2698 41080
rect 2750 41028 2822 41080
rect 2874 41028 2946 41080
rect 2998 41028 4846 41080
rect 4898 41028 4970 41080
rect 5022 41028 5094 41080
rect 5146 41028 5218 41080
rect 5270 41028 7139 41080
rect 7191 41028 7263 41080
rect 7315 41028 7387 41080
rect 7439 41028 7625 41080
rect 7677 41028 7749 41080
rect 7801 41028 7873 41080
rect 7925 41028 9794 41080
rect 9846 41028 9918 41080
rect 9970 41028 10042 41080
rect 10094 41028 10166 41080
rect 10218 41028 12066 41080
rect 12118 41028 12190 41080
rect 12242 41028 12314 41080
rect 12366 41028 12438 41080
rect 12490 41028 13480 41080
rect 13532 41028 13604 41080
rect 13656 41064 14619 41080
rect 13656 41028 14352 41064
rect 712 41012 14352 41028
rect 14404 41012 14460 41064
rect 14512 41012 14568 41064
rect 445 40956 14619 41012
rect 496 40904 552 40956
rect 604 40953 660 40956
rect 712 40953 1438 40956
rect 1490 40953 1562 40956
rect 1614 40953 1686 40956
rect 1738 40953 1810 40956
rect 1862 40953 2574 40956
rect 2626 40953 2698 40956
rect 2750 40953 2822 40956
rect 2874 40953 2946 40956
rect 2998 40953 4846 40956
rect 4898 40953 4970 40956
rect 5022 40953 5094 40956
rect 5146 40953 5218 40956
rect 5270 40953 7139 40956
rect 7191 40953 7263 40956
rect 7315 40953 7387 40956
rect 7439 40953 7625 40956
rect 7677 40953 7749 40956
rect 7801 40953 7873 40956
rect 7925 40953 9794 40956
rect 9846 40953 9918 40956
rect 9970 40953 10042 40956
rect 10094 40953 10166 40956
rect 10218 40953 12066 40956
rect 12118 40953 12190 40956
rect 12242 40953 12314 40956
rect 12366 40953 12438 40956
rect 12490 40953 13480 40956
rect 13532 40953 13604 40956
rect 13656 40953 14352 40956
rect 14404 40953 14460 40956
rect 604 40904 660 40907
rect 712 40904 1438 40907
rect 1490 40904 1562 40907
rect 1614 40904 1686 40907
rect 1738 40904 1810 40907
rect 1862 40904 2574 40907
rect 2626 40904 2698 40907
rect 2750 40904 2822 40907
rect 2874 40904 2946 40907
rect 2998 40904 4846 40907
rect 4898 40904 4970 40907
rect 5022 40904 5094 40907
rect 5146 40904 5218 40907
rect 5270 40904 7139 40907
rect 7191 40904 7263 40907
rect 7315 40904 7387 40907
rect 7439 40904 7625 40907
rect 7677 40904 7749 40907
rect 7801 40904 7873 40907
rect 7925 40904 9794 40907
rect 9846 40904 9918 40907
rect 9970 40904 10042 40907
rect 10094 40904 10166 40907
rect 10218 40904 12066 40907
rect 12118 40904 12190 40907
rect 12242 40904 12314 40907
rect 12366 40904 12438 40907
rect 12490 40904 13480 40907
rect 13532 40904 13604 40907
rect 13656 40904 14352 40907
rect 14404 40904 14460 40907
rect 14512 40904 14568 40956
rect 445 40848 14619 40904
rect 496 40796 552 40848
rect 604 40796 660 40848
rect 712 40832 14352 40848
rect 712 40796 1438 40832
rect 445 40780 1438 40796
rect 1490 40780 1562 40832
rect 1614 40780 1686 40832
rect 1738 40780 1810 40832
rect 1862 40780 2574 40832
rect 2626 40780 2698 40832
rect 2750 40780 2822 40832
rect 2874 40780 2946 40832
rect 2998 40780 4846 40832
rect 4898 40780 4970 40832
rect 5022 40780 5094 40832
rect 5146 40780 5218 40832
rect 5270 40780 7139 40832
rect 7191 40780 7263 40832
rect 7315 40780 7387 40832
rect 7439 40780 7625 40832
rect 7677 40780 7749 40832
rect 7801 40780 7873 40832
rect 7925 40780 9794 40832
rect 9846 40780 9918 40832
rect 9970 40780 10042 40832
rect 10094 40780 10166 40832
rect 10218 40780 12066 40832
rect 12118 40780 12190 40832
rect 12242 40780 12314 40832
rect 12366 40780 12438 40832
rect 12490 40780 13480 40832
rect 13532 40780 13604 40832
rect 13656 40796 14352 40832
rect 14404 40796 14460 40848
rect 14512 40796 14568 40848
rect 13656 40780 14619 40796
rect 445 40740 14619 40780
rect 496 40688 552 40740
rect 604 40688 660 40740
rect 712 40708 14352 40740
rect 712 40688 1438 40708
rect 445 40656 1438 40688
rect 1490 40656 1562 40708
rect 1614 40656 1686 40708
rect 1738 40656 1810 40708
rect 1862 40656 2574 40708
rect 2626 40656 2698 40708
rect 2750 40656 2822 40708
rect 2874 40656 2946 40708
rect 2998 40656 4846 40708
rect 4898 40656 4970 40708
rect 5022 40656 5094 40708
rect 5146 40656 5218 40708
rect 5270 40656 7139 40708
rect 7191 40656 7263 40708
rect 7315 40656 7387 40708
rect 7439 40656 7625 40708
rect 7677 40656 7749 40708
rect 7801 40656 7873 40708
rect 7925 40656 9794 40708
rect 9846 40656 9918 40708
rect 9970 40656 10042 40708
rect 10094 40656 10166 40708
rect 10218 40656 12066 40708
rect 12118 40656 12190 40708
rect 12242 40656 12314 40708
rect 12366 40656 12438 40708
rect 12490 40656 13480 40708
rect 13532 40656 13604 40708
rect 13656 40688 14352 40708
rect 14404 40688 14460 40740
rect 14512 40688 14568 40740
rect 13656 40656 14619 40688
rect 445 40606 14619 40656
rect 445 37306 456 40606
rect 920 40535 3836 40546
rect 920 40489 931 40535
rect 3825 40489 3836 40535
rect 920 40480 1148 40489
rect 1200 40480 1272 40489
rect 1324 40480 3729 40489
rect 920 40478 3729 40480
rect 660 40419 860 40456
rect 660 37493 803 40419
rect 849 37493 860 40419
rect 660 37306 860 37493
rect 920 40408 1920 40478
rect 920 40356 1148 40408
rect 1200 40356 1272 40408
rect 1324 40356 1920 40408
rect 920 40284 1920 40356
rect 920 40232 1148 40284
rect 1200 40232 1272 40284
rect 1324 40232 1920 40284
rect 920 40160 1920 40232
rect 920 40108 1148 40160
rect 1200 40108 1272 40160
rect 1324 40108 1920 40160
rect 920 40036 1920 40108
rect 920 39984 1148 40036
rect 1200 39984 1272 40036
rect 1324 39984 1920 40036
rect 920 39912 1920 39984
rect 920 39860 1148 39912
rect 1200 39860 1272 39912
rect 1324 39860 1920 39912
rect 920 39788 1920 39860
rect 920 39736 1148 39788
rect 1200 39736 1272 39788
rect 1324 39736 1920 39788
rect 920 39664 1920 39736
rect 920 39612 1148 39664
rect 1200 39612 1272 39664
rect 1324 39612 1920 39664
rect 920 39540 1920 39612
rect 920 39488 1148 39540
rect 1200 39488 1272 39540
rect 1324 39488 1920 39540
rect 920 39416 1920 39488
rect 920 39364 1148 39416
rect 1200 39364 1272 39416
rect 1324 39364 1920 39416
rect 920 39292 1920 39364
rect 920 39240 1148 39292
rect 1200 39240 1272 39292
rect 1324 39240 1920 39292
rect 920 39168 1920 39240
rect 920 39116 1148 39168
rect 1200 39116 1272 39168
rect 1324 39116 1920 39168
rect 920 39044 1920 39116
rect 920 38992 1148 39044
rect 1200 38992 1272 39044
rect 1324 38992 1920 39044
rect 920 38920 1920 38992
rect 920 38868 1148 38920
rect 1200 38868 1272 38920
rect 1324 38868 1920 38920
rect 920 38796 1920 38868
rect 920 38744 1148 38796
rect 1200 38744 1272 38796
rect 1324 38744 1920 38796
rect 920 38672 1920 38744
rect 920 38620 1148 38672
rect 1200 38620 1272 38672
rect 1324 38620 1920 38672
rect 920 38548 1920 38620
rect 920 38496 1148 38548
rect 1200 38496 1272 38548
rect 1324 38496 1920 38548
rect 920 38424 1920 38496
rect 920 38372 1148 38424
rect 1200 38372 1272 38424
rect 1324 38372 1920 38424
rect 920 38300 1920 38372
rect 920 38248 1148 38300
rect 1200 38248 1272 38300
rect 1324 38248 1920 38300
rect 920 38176 1920 38248
rect 920 38124 1148 38176
rect 1200 38124 1272 38176
rect 1324 38124 1920 38176
rect 920 38052 1920 38124
rect 920 38000 1148 38052
rect 1200 38000 1272 38052
rect 1324 38000 1920 38052
rect 920 37928 1920 38000
rect 920 37876 1148 37928
rect 1200 37876 1272 37928
rect 1324 37876 1920 37928
rect 920 37804 1920 37876
rect 920 37752 1148 37804
rect 1200 37752 1272 37804
rect 1324 37752 1920 37804
rect 920 37680 1920 37752
rect 920 37628 1148 37680
rect 1200 37628 1272 37680
rect 1324 37628 1920 37680
rect 920 37556 1920 37628
rect 920 37504 1148 37556
rect 1200 37504 1272 37556
rect 1324 37504 1920 37556
rect 920 37434 1920 37504
rect 2836 40442 3729 40478
rect 3781 40442 3836 40489
rect 4356 40535 7272 40546
rect 4356 40489 4367 40535
rect 7261 40489 7272 40535
rect 4356 40478 6335 40489
rect 2836 40386 3836 40442
rect 2836 40334 3729 40386
rect 3781 40334 3836 40386
rect 2836 40278 3836 40334
rect 2836 40226 3729 40278
rect 3781 40226 3836 40278
rect 2836 40170 3836 40226
rect 2836 40118 3729 40170
rect 3781 40118 3836 40170
rect 2836 40062 3836 40118
rect 2836 40010 3729 40062
rect 3781 40010 3836 40062
rect 2836 39954 3836 40010
rect 2836 39902 3729 39954
rect 3781 39902 3836 39954
rect 2836 39846 3836 39902
rect 2836 39794 3729 39846
rect 3781 39794 3836 39846
rect 2836 39738 3836 39794
rect 2836 39686 3729 39738
rect 3781 39686 3836 39738
rect 2836 39630 3836 39686
rect 2836 39578 3729 39630
rect 3781 39578 3836 39630
rect 2836 39522 3836 39578
rect 2836 39470 3729 39522
rect 3781 39470 3836 39522
rect 2836 39414 3836 39470
rect 2836 39362 3729 39414
rect 3781 39362 3836 39414
rect 2836 39306 3836 39362
rect 2836 39254 3729 39306
rect 3781 39254 3836 39306
rect 2836 39198 3836 39254
rect 2836 39146 3729 39198
rect 3781 39146 3836 39198
rect 2836 39090 3836 39146
rect 2836 39038 3729 39090
rect 3781 39038 3836 39090
rect 2836 38982 3836 39038
rect 2836 38930 3729 38982
rect 3781 38930 3836 38982
rect 2836 38874 3836 38930
rect 2836 38822 3729 38874
rect 3781 38822 3836 38874
rect 2836 38766 3836 38822
rect 2836 38714 3729 38766
rect 3781 38714 3836 38766
rect 2836 38658 3836 38714
rect 2836 38606 3729 38658
rect 3781 38606 3836 38658
rect 2836 38550 3836 38606
rect 2836 38498 3729 38550
rect 3781 38498 3836 38550
rect 2836 38442 3836 38498
rect 2836 38390 3729 38442
rect 3781 38390 3836 38442
rect 2836 38334 3836 38390
rect 2836 38282 3729 38334
rect 3781 38282 3836 38334
rect 2836 38226 3836 38282
rect 2836 38174 3729 38226
rect 3781 38174 3836 38226
rect 2836 38118 3836 38174
rect 2836 38066 3729 38118
rect 3781 38066 3836 38118
rect 2836 38010 3836 38066
rect 2836 37958 3729 38010
rect 3781 37958 3836 38010
rect 2836 37902 3836 37958
rect 2836 37850 3729 37902
rect 3781 37850 3836 37902
rect 2836 37794 3836 37850
rect 2836 37742 3729 37794
rect 3781 37742 3836 37794
rect 2836 37686 3836 37742
rect 2836 37634 3729 37686
rect 3781 37634 3836 37686
rect 2836 37578 3836 37634
rect 2836 37526 3729 37578
rect 3781 37526 3836 37578
rect 2836 37470 3836 37526
rect 2836 37434 3729 37470
rect 920 37432 3729 37434
rect 920 37423 1148 37432
rect 1200 37423 1272 37432
rect 1324 37423 3729 37432
rect 3781 37423 3836 37470
rect 920 37377 931 37423
rect 3825 37377 3836 37423
rect 920 37366 3836 37377
rect 3896 40419 4296 40456
rect 3896 37493 3907 40419
rect 3953 37493 4239 40419
rect 4285 37493 4296 40419
rect 3896 37306 4296 37493
rect 4356 37434 5356 40478
rect 6272 40442 6335 40478
rect 6387 40442 7272 40489
rect 7792 40535 10708 40546
rect 7792 40489 7803 40535
rect 10697 40489 10708 40535
rect 6272 40386 7272 40442
rect 6272 40334 6335 40386
rect 6387 40334 7272 40386
rect 6272 40278 7272 40334
rect 6272 40226 6335 40278
rect 6387 40226 7272 40278
rect 6272 40170 7272 40226
rect 6272 40118 6335 40170
rect 6387 40118 7272 40170
rect 6272 40062 7272 40118
rect 6272 40010 6335 40062
rect 6387 40010 7272 40062
rect 6272 39954 7272 40010
rect 6272 39902 6335 39954
rect 6387 39902 7272 39954
rect 6272 39846 7272 39902
rect 6272 39794 6335 39846
rect 6387 39794 7272 39846
rect 6272 39738 7272 39794
rect 6272 39686 6335 39738
rect 6387 39686 7272 39738
rect 6272 39630 7272 39686
rect 6272 39578 6335 39630
rect 6387 39578 7272 39630
rect 6272 39522 7272 39578
rect 6272 39470 6335 39522
rect 6387 39470 7272 39522
rect 6272 39414 7272 39470
rect 6272 39362 6335 39414
rect 6387 39362 7272 39414
rect 6272 39306 7272 39362
rect 6272 39254 6335 39306
rect 6387 39254 7272 39306
rect 6272 39198 7272 39254
rect 6272 39146 6335 39198
rect 6387 39146 7272 39198
rect 6272 39090 7272 39146
rect 6272 39038 6335 39090
rect 6387 39038 7272 39090
rect 6272 38982 7272 39038
rect 6272 38930 6335 38982
rect 6387 38930 7272 38982
rect 6272 38874 7272 38930
rect 6272 38822 6335 38874
rect 6387 38822 7272 38874
rect 6272 38766 7272 38822
rect 6272 38714 6335 38766
rect 6387 38714 7272 38766
rect 6272 38658 7272 38714
rect 6272 38606 6335 38658
rect 6387 38606 7272 38658
rect 6272 38550 7272 38606
rect 6272 38498 6335 38550
rect 6387 38498 7272 38550
rect 6272 38442 7272 38498
rect 6272 38390 6335 38442
rect 6387 38390 7272 38442
rect 6272 38334 7272 38390
rect 6272 38282 6335 38334
rect 6387 38282 7272 38334
rect 6272 38226 7272 38282
rect 6272 38174 6335 38226
rect 6387 38174 7272 38226
rect 6272 38118 7272 38174
rect 6272 38066 6335 38118
rect 6387 38066 7272 38118
rect 6272 38010 7272 38066
rect 6272 37958 6335 38010
rect 6387 37958 7272 38010
rect 6272 37902 7272 37958
rect 6272 37850 6335 37902
rect 6387 37850 7272 37902
rect 6272 37794 7272 37850
rect 6272 37742 6335 37794
rect 6387 37742 7272 37794
rect 6272 37686 7272 37742
rect 6272 37634 6335 37686
rect 6387 37634 7272 37686
rect 6272 37578 7272 37634
rect 6272 37526 6335 37578
rect 6387 37526 7272 37578
rect 6272 37470 7272 37526
rect 6272 37434 6335 37470
rect 4356 37423 6335 37434
rect 6387 37423 7272 37470
rect 4356 37377 4367 37423
rect 7261 37377 7272 37423
rect 4356 37366 7272 37377
rect 7332 40440 7732 40456
rect 7332 40419 7388 40440
rect 7332 37493 7343 40419
rect 7440 40388 7624 40440
rect 7676 40419 7732 40440
rect 7389 40332 7675 40388
rect 7440 40280 7624 40332
rect 7389 40224 7675 40280
rect 7440 40172 7624 40224
rect 7389 40116 7675 40172
rect 7440 40064 7624 40116
rect 7389 40008 7675 40064
rect 7440 39956 7624 40008
rect 7389 39900 7675 39956
rect 7440 39848 7624 39900
rect 7389 39792 7675 39848
rect 7440 39740 7624 39792
rect 7389 39684 7675 39740
rect 7440 39632 7624 39684
rect 7389 39576 7675 39632
rect 7440 39524 7624 39576
rect 7389 39468 7675 39524
rect 7440 39416 7624 39468
rect 7389 39360 7675 39416
rect 7440 39308 7624 39360
rect 7389 39252 7675 39308
rect 7440 39200 7624 39252
rect 7389 39144 7675 39200
rect 7440 39092 7624 39144
rect 7389 39036 7675 39092
rect 7440 38984 7624 39036
rect 7389 38928 7675 38984
rect 7440 38876 7624 38928
rect 7389 38820 7675 38876
rect 7440 38768 7624 38820
rect 7389 38712 7675 38768
rect 7440 38660 7624 38712
rect 7389 38604 7675 38660
rect 7440 38552 7624 38604
rect 7389 38496 7675 38552
rect 7440 38444 7624 38496
rect 7389 38388 7675 38444
rect 7440 38336 7624 38388
rect 7389 38280 7675 38336
rect 7440 38228 7624 38280
rect 7389 38172 7675 38228
rect 7440 38120 7624 38172
rect 7389 38064 7675 38120
rect 7440 38012 7624 38064
rect 7389 37956 7675 38012
rect 7440 37904 7624 37956
rect 7389 37848 7675 37904
rect 7440 37796 7624 37848
rect 7389 37740 7675 37796
rect 7440 37688 7624 37740
rect 7389 37632 7675 37688
rect 7440 37580 7624 37632
rect 7389 37524 7675 37580
rect 7332 37472 7388 37493
rect 7440 37472 7624 37524
rect 7721 37493 7732 40419
rect 7676 37472 7732 37493
rect 7332 37306 7732 37472
rect 7792 40442 8677 40489
rect 8729 40478 10708 40489
rect 8729 40442 8792 40478
rect 7792 40386 8792 40442
rect 7792 40334 8677 40386
rect 8729 40334 8792 40386
rect 7792 40278 8792 40334
rect 7792 40226 8677 40278
rect 8729 40226 8792 40278
rect 7792 40170 8792 40226
rect 7792 40118 8677 40170
rect 8729 40118 8792 40170
rect 7792 40062 8792 40118
rect 7792 40010 8677 40062
rect 8729 40010 8792 40062
rect 7792 39954 8792 40010
rect 7792 39902 8677 39954
rect 8729 39902 8792 39954
rect 7792 39846 8792 39902
rect 7792 39794 8677 39846
rect 8729 39794 8792 39846
rect 7792 39738 8792 39794
rect 7792 39686 8677 39738
rect 8729 39686 8792 39738
rect 7792 39630 8792 39686
rect 7792 39578 8677 39630
rect 8729 39578 8792 39630
rect 7792 39522 8792 39578
rect 7792 39470 8677 39522
rect 8729 39470 8792 39522
rect 7792 39414 8792 39470
rect 7792 39362 8677 39414
rect 8729 39362 8792 39414
rect 7792 39306 8792 39362
rect 7792 39254 8677 39306
rect 8729 39254 8792 39306
rect 7792 39198 8792 39254
rect 7792 39146 8677 39198
rect 8729 39146 8792 39198
rect 7792 39090 8792 39146
rect 7792 39038 8677 39090
rect 8729 39038 8792 39090
rect 7792 38982 8792 39038
rect 7792 38930 8677 38982
rect 8729 38930 8792 38982
rect 7792 38874 8792 38930
rect 7792 38822 8677 38874
rect 8729 38822 8792 38874
rect 7792 38766 8792 38822
rect 7792 38714 8677 38766
rect 8729 38714 8792 38766
rect 7792 38658 8792 38714
rect 7792 38606 8677 38658
rect 8729 38606 8792 38658
rect 7792 38550 8792 38606
rect 7792 38498 8677 38550
rect 8729 38498 8792 38550
rect 7792 38442 8792 38498
rect 7792 38390 8677 38442
rect 8729 38390 8792 38442
rect 7792 38334 8792 38390
rect 7792 38282 8677 38334
rect 8729 38282 8792 38334
rect 7792 38226 8792 38282
rect 7792 38174 8677 38226
rect 8729 38174 8792 38226
rect 7792 38118 8792 38174
rect 7792 38066 8677 38118
rect 8729 38066 8792 38118
rect 7792 38010 8792 38066
rect 7792 37958 8677 38010
rect 8729 37958 8792 38010
rect 7792 37902 8792 37958
rect 7792 37850 8677 37902
rect 8729 37850 8792 37902
rect 7792 37794 8792 37850
rect 7792 37742 8677 37794
rect 8729 37742 8792 37794
rect 7792 37686 8792 37742
rect 7792 37634 8677 37686
rect 8729 37634 8792 37686
rect 7792 37578 8792 37634
rect 7792 37526 8677 37578
rect 8729 37526 8792 37578
rect 7792 37470 8792 37526
rect 7792 37423 8677 37470
rect 8729 37434 8792 37470
rect 9708 37434 10708 40478
rect 11228 40535 14144 40546
rect 11228 40489 11239 40535
rect 14133 40489 14144 40535
rect 8729 37423 10708 37434
rect 7792 37377 7803 37423
rect 10697 37377 10708 37423
rect 7792 37366 10708 37377
rect 10768 40419 11168 40456
rect 10768 37493 10779 40419
rect 10825 37493 11111 40419
rect 11157 37493 11168 40419
rect 10768 37306 11168 37493
rect 11228 40442 11283 40489
rect 11335 40480 13786 40489
rect 13838 40480 13910 40489
rect 13962 40480 14034 40489
rect 14086 40480 14144 40489
rect 11335 40478 14144 40480
rect 11335 40442 12228 40478
rect 11228 40386 12228 40442
rect 11228 40334 11283 40386
rect 11335 40334 12228 40386
rect 11228 40278 12228 40334
rect 11228 40226 11283 40278
rect 11335 40226 12228 40278
rect 11228 40170 12228 40226
rect 11228 40118 11283 40170
rect 11335 40118 12228 40170
rect 11228 40062 12228 40118
rect 11228 40010 11283 40062
rect 11335 40010 12228 40062
rect 11228 39954 12228 40010
rect 11228 39902 11283 39954
rect 11335 39902 12228 39954
rect 11228 39846 12228 39902
rect 11228 39794 11283 39846
rect 11335 39794 12228 39846
rect 11228 39738 12228 39794
rect 11228 39686 11283 39738
rect 11335 39686 12228 39738
rect 11228 39630 12228 39686
rect 11228 39578 11283 39630
rect 11335 39578 12228 39630
rect 11228 39522 12228 39578
rect 11228 39470 11283 39522
rect 11335 39470 12228 39522
rect 11228 39414 12228 39470
rect 11228 39362 11283 39414
rect 11335 39362 12228 39414
rect 11228 39306 12228 39362
rect 11228 39254 11283 39306
rect 11335 39254 12228 39306
rect 11228 39198 12228 39254
rect 11228 39146 11283 39198
rect 11335 39146 12228 39198
rect 11228 39090 12228 39146
rect 11228 39038 11283 39090
rect 11335 39038 12228 39090
rect 11228 38982 12228 39038
rect 11228 38930 11283 38982
rect 11335 38930 12228 38982
rect 11228 38874 12228 38930
rect 11228 38822 11283 38874
rect 11335 38822 12228 38874
rect 11228 38766 12228 38822
rect 11228 38714 11283 38766
rect 11335 38714 12228 38766
rect 11228 38658 12228 38714
rect 11228 38606 11283 38658
rect 11335 38606 12228 38658
rect 11228 38550 12228 38606
rect 11228 38498 11283 38550
rect 11335 38498 12228 38550
rect 11228 38442 12228 38498
rect 11228 38390 11283 38442
rect 11335 38390 12228 38442
rect 11228 38334 12228 38390
rect 11228 38282 11283 38334
rect 11335 38282 12228 38334
rect 11228 38226 12228 38282
rect 11228 38174 11283 38226
rect 11335 38174 12228 38226
rect 11228 38118 12228 38174
rect 11228 38066 11283 38118
rect 11335 38066 12228 38118
rect 11228 38010 12228 38066
rect 11228 37958 11283 38010
rect 11335 37958 12228 38010
rect 11228 37902 12228 37958
rect 11228 37850 11283 37902
rect 11335 37850 12228 37902
rect 11228 37794 12228 37850
rect 11228 37742 11283 37794
rect 11335 37742 12228 37794
rect 11228 37686 12228 37742
rect 11228 37634 11283 37686
rect 11335 37634 12228 37686
rect 11228 37578 12228 37634
rect 11228 37526 11283 37578
rect 11335 37526 12228 37578
rect 11228 37470 12228 37526
rect 11228 37423 11283 37470
rect 11335 37434 12228 37470
rect 13144 40408 14144 40478
rect 13144 40356 13786 40408
rect 13838 40356 13910 40408
rect 13962 40356 14034 40408
rect 14086 40356 14144 40408
rect 13144 40284 14144 40356
rect 13144 40232 13786 40284
rect 13838 40232 13910 40284
rect 13962 40232 14034 40284
rect 14086 40232 14144 40284
rect 13144 40160 14144 40232
rect 13144 40108 13786 40160
rect 13838 40108 13910 40160
rect 13962 40108 14034 40160
rect 14086 40108 14144 40160
rect 13144 40036 14144 40108
rect 13144 39984 13786 40036
rect 13838 39984 13910 40036
rect 13962 39984 14034 40036
rect 14086 39984 14144 40036
rect 13144 39912 14144 39984
rect 13144 39860 13786 39912
rect 13838 39860 13910 39912
rect 13962 39860 14034 39912
rect 14086 39860 14144 39912
rect 13144 39788 14144 39860
rect 13144 39736 13786 39788
rect 13838 39736 13910 39788
rect 13962 39736 14034 39788
rect 14086 39736 14144 39788
rect 13144 39664 14144 39736
rect 13144 39612 13786 39664
rect 13838 39612 13910 39664
rect 13962 39612 14034 39664
rect 14086 39612 14144 39664
rect 13144 39540 14144 39612
rect 13144 39488 13786 39540
rect 13838 39488 13910 39540
rect 13962 39488 14034 39540
rect 14086 39488 14144 39540
rect 13144 39416 14144 39488
rect 13144 39364 13786 39416
rect 13838 39364 13910 39416
rect 13962 39364 14034 39416
rect 14086 39364 14144 39416
rect 13144 39292 14144 39364
rect 13144 39240 13786 39292
rect 13838 39240 13910 39292
rect 13962 39240 14034 39292
rect 14086 39240 14144 39292
rect 13144 39168 14144 39240
rect 13144 39116 13786 39168
rect 13838 39116 13910 39168
rect 13962 39116 14034 39168
rect 14086 39116 14144 39168
rect 13144 39044 14144 39116
rect 13144 38992 13786 39044
rect 13838 38992 13910 39044
rect 13962 38992 14034 39044
rect 14086 38992 14144 39044
rect 13144 38920 14144 38992
rect 13144 38868 13786 38920
rect 13838 38868 13910 38920
rect 13962 38868 14034 38920
rect 14086 38868 14144 38920
rect 13144 38796 14144 38868
rect 13144 38744 13786 38796
rect 13838 38744 13910 38796
rect 13962 38744 14034 38796
rect 14086 38744 14144 38796
rect 13144 38672 14144 38744
rect 13144 38620 13786 38672
rect 13838 38620 13910 38672
rect 13962 38620 14034 38672
rect 14086 38620 14144 38672
rect 13144 38548 14144 38620
rect 13144 38496 13786 38548
rect 13838 38496 13910 38548
rect 13962 38496 14034 38548
rect 14086 38496 14144 38548
rect 13144 38424 14144 38496
rect 13144 38372 13786 38424
rect 13838 38372 13910 38424
rect 13962 38372 14034 38424
rect 14086 38372 14144 38424
rect 13144 38300 14144 38372
rect 13144 38248 13786 38300
rect 13838 38248 13910 38300
rect 13962 38248 14034 38300
rect 14086 38248 14144 38300
rect 13144 38176 14144 38248
rect 13144 38124 13786 38176
rect 13838 38124 13910 38176
rect 13962 38124 14034 38176
rect 14086 38124 14144 38176
rect 13144 38052 14144 38124
rect 13144 38000 13786 38052
rect 13838 38000 13910 38052
rect 13962 38000 14034 38052
rect 14086 38000 14144 38052
rect 13144 37928 14144 38000
rect 13144 37876 13786 37928
rect 13838 37876 13910 37928
rect 13962 37876 14034 37928
rect 14086 37876 14144 37928
rect 13144 37804 14144 37876
rect 13144 37752 13786 37804
rect 13838 37752 13910 37804
rect 13962 37752 14034 37804
rect 14086 37752 14144 37804
rect 13144 37680 14144 37752
rect 13144 37628 13786 37680
rect 13838 37628 13910 37680
rect 13962 37628 14034 37680
rect 14086 37628 14144 37680
rect 13144 37556 14144 37628
rect 13144 37504 13786 37556
rect 13838 37504 13910 37556
rect 13962 37504 14034 37556
rect 14086 37504 14144 37556
rect 13144 37434 14144 37504
rect 11335 37432 14144 37434
rect 11335 37423 13786 37432
rect 13838 37423 13910 37432
rect 13962 37423 14034 37432
rect 14086 37423 14144 37432
rect 11228 37377 11239 37423
rect 14133 37377 14144 37423
rect 11228 37366 14144 37377
rect 14204 40419 14404 40456
rect 14204 37493 14215 40419
rect 14261 37493 14404 40419
rect 14204 37306 14404 37493
rect 14608 37306 14619 40606
rect 445 37256 14619 37306
rect 445 37224 1438 37256
rect 496 37172 552 37224
rect 604 37172 660 37224
rect 712 37204 1438 37224
rect 1490 37204 1562 37256
rect 1614 37204 1686 37256
rect 1738 37204 1810 37256
rect 1862 37204 2574 37256
rect 2626 37204 2698 37256
rect 2750 37204 2822 37256
rect 2874 37204 2946 37256
rect 2998 37204 4846 37256
rect 4898 37204 4970 37256
rect 5022 37204 5094 37256
rect 5146 37204 5218 37256
rect 5270 37204 7139 37256
rect 7191 37204 7263 37256
rect 7315 37204 7387 37256
rect 7439 37204 7625 37256
rect 7677 37204 7749 37256
rect 7801 37204 7873 37256
rect 7925 37204 9794 37256
rect 9846 37204 9918 37256
rect 9970 37204 10042 37256
rect 10094 37204 10166 37256
rect 10218 37204 12066 37256
rect 12118 37204 12190 37256
rect 12242 37204 12314 37256
rect 12366 37204 12438 37256
rect 12490 37204 13480 37256
rect 13532 37204 13604 37256
rect 13656 37224 14619 37256
rect 13656 37204 14352 37224
rect 712 37172 14352 37204
rect 14404 37172 14460 37224
rect 14512 37172 14568 37224
rect 445 37132 14619 37172
rect 445 37116 1438 37132
rect 496 37064 552 37116
rect 604 37064 660 37116
rect 712 37080 1438 37116
rect 1490 37080 1562 37132
rect 1614 37080 1686 37132
rect 1738 37080 1810 37132
rect 1862 37080 2574 37132
rect 2626 37080 2698 37132
rect 2750 37080 2822 37132
rect 2874 37080 2946 37132
rect 2998 37080 4846 37132
rect 4898 37080 4970 37132
rect 5022 37080 5094 37132
rect 5146 37080 5218 37132
rect 5270 37080 7139 37132
rect 7191 37080 7263 37132
rect 7315 37080 7387 37132
rect 7439 37080 7625 37132
rect 7677 37080 7749 37132
rect 7801 37080 7873 37132
rect 7925 37080 9794 37132
rect 9846 37080 9918 37132
rect 9970 37080 10042 37132
rect 10094 37080 10166 37132
rect 10218 37080 12066 37132
rect 12118 37080 12190 37132
rect 12242 37080 12314 37132
rect 12366 37080 12438 37132
rect 12490 37080 13480 37132
rect 13532 37080 13604 37132
rect 13656 37116 14619 37132
rect 13656 37080 14352 37116
rect 712 37064 14352 37080
rect 14404 37064 14460 37116
rect 14512 37064 14568 37116
rect 445 37008 14619 37064
rect 496 36956 552 37008
rect 604 37005 660 37008
rect 712 37005 1438 37008
rect 1490 37005 1562 37008
rect 1614 37005 1686 37008
rect 1738 37005 1810 37008
rect 1862 37005 2574 37008
rect 2626 37005 2698 37008
rect 2750 37005 2822 37008
rect 2874 37005 2946 37008
rect 2998 37005 4846 37008
rect 4898 37005 4970 37008
rect 5022 37005 5094 37008
rect 5146 37005 5218 37008
rect 5270 37005 7139 37008
rect 7191 37005 7263 37008
rect 7315 37005 7387 37008
rect 7439 37005 7625 37008
rect 7677 37005 7749 37008
rect 7801 37005 7873 37008
rect 7925 37005 9794 37008
rect 9846 37005 9918 37008
rect 9970 37005 10042 37008
rect 10094 37005 10166 37008
rect 10218 37005 12066 37008
rect 12118 37005 12190 37008
rect 12242 37005 12314 37008
rect 12366 37005 12438 37008
rect 12490 37005 13480 37008
rect 13532 37005 13604 37008
rect 13656 37005 14352 37008
rect 14404 37005 14460 37008
rect 604 36956 660 36959
rect 712 36956 1438 36959
rect 1490 36956 1562 36959
rect 1614 36956 1686 36959
rect 1738 36956 1810 36959
rect 1862 36956 2574 36959
rect 2626 36956 2698 36959
rect 2750 36956 2822 36959
rect 2874 36956 2946 36959
rect 2998 36956 4846 36959
rect 4898 36956 4970 36959
rect 5022 36956 5094 36959
rect 5146 36956 5218 36959
rect 5270 36956 7139 36959
rect 7191 36956 7263 36959
rect 7315 36956 7387 36959
rect 7439 36956 7625 36959
rect 7677 36956 7749 36959
rect 7801 36956 7873 36959
rect 7925 36956 9794 36959
rect 9846 36956 9918 36959
rect 9970 36956 10042 36959
rect 10094 36956 10166 36959
rect 10218 36956 12066 36959
rect 12118 36956 12190 36959
rect 12242 36956 12314 36959
rect 12366 36956 12438 36959
rect 12490 36956 13480 36959
rect 13532 36956 13604 36959
rect 13656 36956 14352 36959
rect 14404 36956 14460 36959
rect 14512 36956 14568 37008
rect 445 36900 14619 36956
rect 496 36848 552 36900
rect 604 36848 660 36900
rect 712 36884 14352 36900
rect 712 36848 1438 36884
rect 445 36832 1438 36848
rect 1490 36832 1562 36884
rect 1614 36832 1686 36884
rect 1738 36832 1810 36884
rect 1862 36832 2574 36884
rect 2626 36832 2698 36884
rect 2750 36832 2822 36884
rect 2874 36832 2946 36884
rect 2998 36832 4846 36884
rect 4898 36832 4970 36884
rect 5022 36832 5094 36884
rect 5146 36832 5218 36884
rect 5270 36832 7139 36884
rect 7191 36832 7263 36884
rect 7315 36832 7387 36884
rect 7439 36832 7625 36884
rect 7677 36832 7749 36884
rect 7801 36832 7873 36884
rect 7925 36832 9794 36884
rect 9846 36832 9918 36884
rect 9970 36832 10042 36884
rect 10094 36832 10166 36884
rect 10218 36832 12066 36884
rect 12118 36832 12190 36884
rect 12242 36832 12314 36884
rect 12366 36832 12438 36884
rect 12490 36832 13480 36884
rect 13532 36832 13604 36884
rect 13656 36848 14352 36884
rect 14404 36848 14460 36900
rect 14512 36848 14568 36900
rect 13656 36832 14619 36848
rect 445 36792 14619 36832
rect 496 36740 552 36792
rect 604 36740 660 36792
rect 712 36760 14352 36792
rect 712 36740 1438 36760
rect 445 36708 1438 36740
rect 1490 36708 1562 36760
rect 1614 36708 1686 36760
rect 1738 36708 1810 36760
rect 1862 36708 2574 36760
rect 2626 36708 2698 36760
rect 2750 36708 2822 36760
rect 2874 36708 2946 36760
rect 2998 36708 4846 36760
rect 4898 36708 4970 36760
rect 5022 36708 5094 36760
rect 5146 36708 5218 36760
rect 5270 36708 7139 36760
rect 7191 36708 7263 36760
rect 7315 36708 7387 36760
rect 7439 36708 7625 36760
rect 7677 36708 7749 36760
rect 7801 36708 7873 36760
rect 7925 36708 9794 36760
rect 9846 36708 9918 36760
rect 9970 36708 10042 36760
rect 10094 36708 10166 36760
rect 10218 36708 12066 36760
rect 12118 36708 12190 36760
rect 12242 36708 12314 36760
rect 12366 36708 12438 36760
rect 12490 36708 13480 36760
rect 13532 36708 13604 36760
rect 13656 36740 14352 36760
rect 14404 36740 14460 36792
rect 14512 36740 14568 36792
rect 13656 36708 14619 36740
rect 445 36658 14619 36708
rect 445 33358 456 36658
rect 920 36587 3836 36598
rect 920 36541 931 36587
rect 3825 36541 3836 36587
rect 920 36532 978 36541
rect 1030 36532 1102 36541
rect 1154 36532 1226 36541
rect 1278 36532 3729 36541
rect 920 36530 3729 36532
rect 660 36471 860 36508
rect 660 33545 803 36471
rect 849 33545 860 36471
rect 660 33358 860 33545
rect 920 36460 1920 36530
rect 920 36408 978 36460
rect 1030 36408 1102 36460
rect 1154 36408 1226 36460
rect 1278 36408 1920 36460
rect 920 36336 1920 36408
rect 920 36284 978 36336
rect 1030 36284 1102 36336
rect 1154 36284 1226 36336
rect 1278 36284 1920 36336
rect 920 36212 1920 36284
rect 920 36160 978 36212
rect 1030 36160 1102 36212
rect 1154 36160 1226 36212
rect 1278 36160 1920 36212
rect 920 36088 1920 36160
rect 920 36036 978 36088
rect 1030 36036 1102 36088
rect 1154 36036 1226 36088
rect 1278 36036 1920 36088
rect 920 35964 1920 36036
rect 920 35912 978 35964
rect 1030 35912 1102 35964
rect 1154 35912 1226 35964
rect 1278 35912 1920 35964
rect 920 35840 1920 35912
rect 920 35788 978 35840
rect 1030 35788 1102 35840
rect 1154 35788 1226 35840
rect 1278 35788 1920 35840
rect 920 35716 1920 35788
rect 920 35664 978 35716
rect 1030 35664 1102 35716
rect 1154 35664 1226 35716
rect 1278 35664 1920 35716
rect 920 35592 1920 35664
rect 920 35540 978 35592
rect 1030 35540 1102 35592
rect 1154 35540 1226 35592
rect 1278 35540 1920 35592
rect 920 35468 1920 35540
rect 920 35416 978 35468
rect 1030 35416 1102 35468
rect 1154 35416 1226 35468
rect 1278 35416 1920 35468
rect 920 35344 1920 35416
rect 920 35292 978 35344
rect 1030 35292 1102 35344
rect 1154 35292 1226 35344
rect 1278 35292 1920 35344
rect 920 35220 1920 35292
rect 920 35168 978 35220
rect 1030 35168 1102 35220
rect 1154 35168 1226 35220
rect 1278 35168 1920 35220
rect 920 35096 1920 35168
rect 920 35044 978 35096
rect 1030 35044 1102 35096
rect 1154 35044 1226 35096
rect 1278 35044 1920 35096
rect 920 34972 1920 35044
rect 920 34920 978 34972
rect 1030 34920 1102 34972
rect 1154 34920 1226 34972
rect 1278 34920 1920 34972
rect 920 34848 1920 34920
rect 920 34796 978 34848
rect 1030 34796 1102 34848
rect 1154 34796 1226 34848
rect 1278 34796 1920 34848
rect 920 34724 1920 34796
rect 920 34672 978 34724
rect 1030 34672 1102 34724
rect 1154 34672 1226 34724
rect 1278 34672 1920 34724
rect 920 34600 1920 34672
rect 920 34548 978 34600
rect 1030 34548 1102 34600
rect 1154 34548 1226 34600
rect 1278 34548 1920 34600
rect 920 34476 1920 34548
rect 920 34424 978 34476
rect 1030 34424 1102 34476
rect 1154 34424 1226 34476
rect 1278 34424 1920 34476
rect 920 34352 1920 34424
rect 920 34300 978 34352
rect 1030 34300 1102 34352
rect 1154 34300 1226 34352
rect 1278 34300 1920 34352
rect 920 34228 1920 34300
rect 920 34176 978 34228
rect 1030 34176 1102 34228
rect 1154 34176 1226 34228
rect 1278 34176 1920 34228
rect 920 34104 1920 34176
rect 920 34052 978 34104
rect 1030 34052 1102 34104
rect 1154 34052 1226 34104
rect 1278 34052 1920 34104
rect 920 33980 1920 34052
rect 920 33928 978 33980
rect 1030 33928 1102 33980
rect 1154 33928 1226 33980
rect 1278 33928 1920 33980
rect 920 33856 1920 33928
rect 920 33804 978 33856
rect 1030 33804 1102 33856
rect 1154 33804 1226 33856
rect 1278 33804 1920 33856
rect 920 33732 1920 33804
rect 920 33680 978 33732
rect 1030 33680 1102 33732
rect 1154 33680 1226 33732
rect 1278 33680 1920 33732
rect 920 33608 1920 33680
rect 920 33556 978 33608
rect 1030 33556 1102 33608
rect 1154 33556 1226 33608
rect 1278 33556 1920 33608
rect 920 33486 1920 33556
rect 2836 36494 3729 36530
rect 3781 36494 3836 36541
rect 4356 36587 7272 36598
rect 4356 36541 4367 36587
rect 7261 36541 7272 36587
rect 4356 36530 6335 36541
rect 2836 36438 3836 36494
rect 2836 36386 3729 36438
rect 3781 36386 3836 36438
rect 2836 36330 3836 36386
rect 2836 36278 3729 36330
rect 3781 36278 3836 36330
rect 2836 36222 3836 36278
rect 2836 36170 3729 36222
rect 3781 36170 3836 36222
rect 2836 36114 3836 36170
rect 2836 36062 3729 36114
rect 3781 36062 3836 36114
rect 2836 36006 3836 36062
rect 2836 35954 3729 36006
rect 3781 35954 3836 36006
rect 2836 35898 3836 35954
rect 2836 35846 3729 35898
rect 3781 35846 3836 35898
rect 2836 35790 3836 35846
rect 2836 35738 3729 35790
rect 3781 35738 3836 35790
rect 2836 35682 3836 35738
rect 2836 35630 3729 35682
rect 3781 35630 3836 35682
rect 2836 35574 3836 35630
rect 2836 35522 3729 35574
rect 3781 35522 3836 35574
rect 2836 35466 3836 35522
rect 2836 35414 3729 35466
rect 3781 35414 3836 35466
rect 2836 35358 3836 35414
rect 2836 35306 3729 35358
rect 3781 35306 3836 35358
rect 2836 35250 3836 35306
rect 2836 35198 3729 35250
rect 3781 35198 3836 35250
rect 2836 35142 3836 35198
rect 2836 35090 3729 35142
rect 3781 35090 3836 35142
rect 2836 35034 3836 35090
rect 2836 34982 3729 35034
rect 3781 34982 3836 35034
rect 2836 34926 3836 34982
rect 2836 34874 3729 34926
rect 3781 34874 3836 34926
rect 2836 34818 3836 34874
rect 2836 34766 3729 34818
rect 3781 34766 3836 34818
rect 2836 34710 3836 34766
rect 2836 34658 3729 34710
rect 3781 34658 3836 34710
rect 2836 34602 3836 34658
rect 2836 34550 3729 34602
rect 3781 34550 3836 34602
rect 2836 34494 3836 34550
rect 2836 34442 3729 34494
rect 3781 34442 3836 34494
rect 2836 34386 3836 34442
rect 2836 34334 3729 34386
rect 3781 34334 3836 34386
rect 2836 34278 3836 34334
rect 2836 34226 3729 34278
rect 3781 34226 3836 34278
rect 2836 34170 3836 34226
rect 2836 34118 3729 34170
rect 3781 34118 3836 34170
rect 2836 34062 3836 34118
rect 2836 34010 3729 34062
rect 3781 34010 3836 34062
rect 2836 33954 3836 34010
rect 2836 33902 3729 33954
rect 3781 33902 3836 33954
rect 2836 33846 3836 33902
rect 2836 33794 3729 33846
rect 3781 33794 3836 33846
rect 2836 33738 3836 33794
rect 2836 33686 3729 33738
rect 3781 33686 3836 33738
rect 2836 33630 3836 33686
rect 2836 33578 3729 33630
rect 3781 33578 3836 33630
rect 2836 33522 3836 33578
rect 2836 33486 3729 33522
rect 920 33484 3729 33486
rect 920 33475 978 33484
rect 1030 33475 1102 33484
rect 1154 33475 1226 33484
rect 1278 33475 3729 33484
rect 3781 33475 3836 33522
rect 920 33429 931 33475
rect 3825 33429 3836 33475
rect 920 33418 3836 33429
rect 3896 36471 4296 36508
rect 3896 33545 3907 36471
rect 3953 33545 4239 36471
rect 4285 33545 4296 36471
rect 3896 33358 4296 33545
rect 4356 33486 5356 36530
rect 6272 36494 6335 36530
rect 6387 36494 7272 36541
rect 7792 36587 10708 36598
rect 7792 36541 7803 36587
rect 10697 36541 10708 36587
rect 6272 36438 7272 36494
rect 6272 36386 6335 36438
rect 6387 36386 7272 36438
rect 6272 36330 7272 36386
rect 6272 36278 6335 36330
rect 6387 36278 7272 36330
rect 6272 36222 7272 36278
rect 6272 36170 6335 36222
rect 6387 36170 7272 36222
rect 6272 36114 7272 36170
rect 6272 36062 6335 36114
rect 6387 36062 7272 36114
rect 6272 36006 7272 36062
rect 6272 35954 6335 36006
rect 6387 35954 7272 36006
rect 6272 35898 7272 35954
rect 6272 35846 6335 35898
rect 6387 35846 7272 35898
rect 6272 35790 7272 35846
rect 6272 35738 6335 35790
rect 6387 35738 7272 35790
rect 6272 35682 7272 35738
rect 6272 35630 6335 35682
rect 6387 35630 7272 35682
rect 6272 35574 7272 35630
rect 6272 35522 6335 35574
rect 6387 35522 7272 35574
rect 6272 35466 7272 35522
rect 6272 35414 6335 35466
rect 6387 35414 7272 35466
rect 6272 35358 7272 35414
rect 6272 35306 6335 35358
rect 6387 35306 7272 35358
rect 6272 35250 7272 35306
rect 6272 35198 6335 35250
rect 6387 35198 7272 35250
rect 6272 35142 7272 35198
rect 6272 35090 6335 35142
rect 6387 35090 7272 35142
rect 6272 35034 7272 35090
rect 6272 34982 6335 35034
rect 6387 34982 7272 35034
rect 6272 34926 7272 34982
rect 6272 34874 6335 34926
rect 6387 34874 7272 34926
rect 6272 34818 7272 34874
rect 6272 34766 6335 34818
rect 6387 34766 7272 34818
rect 6272 34710 7272 34766
rect 6272 34658 6335 34710
rect 6387 34658 7272 34710
rect 6272 34602 7272 34658
rect 6272 34550 6335 34602
rect 6387 34550 7272 34602
rect 6272 34494 7272 34550
rect 6272 34442 6335 34494
rect 6387 34442 7272 34494
rect 6272 34386 7272 34442
rect 6272 34334 6335 34386
rect 6387 34334 7272 34386
rect 6272 34278 7272 34334
rect 6272 34226 6335 34278
rect 6387 34226 7272 34278
rect 6272 34170 7272 34226
rect 6272 34118 6335 34170
rect 6387 34118 7272 34170
rect 6272 34062 7272 34118
rect 6272 34010 6335 34062
rect 6387 34010 7272 34062
rect 6272 33954 7272 34010
rect 6272 33902 6335 33954
rect 6387 33902 7272 33954
rect 6272 33846 7272 33902
rect 6272 33794 6335 33846
rect 6387 33794 7272 33846
rect 6272 33738 7272 33794
rect 6272 33686 6335 33738
rect 6387 33686 7272 33738
rect 6272 33630 7272 33686
rect 6272 33578 6335 33630
rect 6387 33578 7272 33630
rect 6272 33522 7272 33578
rect 6272 33486 6335 33522
rect 4356 33475 6335 33486
rect 6387 33475 7272 33522
rect 4356 33429 4367 33475
rect 7261 33429 7272 33475
rect 4356 33418 7272 33429
rect 7332 36492 7732 36508
rect 7332 36471 7388 36492
rect 7332 33545 7343 36471
rect 7440 36440 7624 36492
rect 7676 36471 7732 36492
rect 7389 36384 7675 36440
rect 7440 36332 7624 36384
rect 7389 36276 7675 36332
rect 7440 36224 7624 36276
rect 7389 36168 7675 36224
rect 7440 36116 7624 36168
rect 7389 36060 7675 36116
rect 7440 36008 7624 36060
rect 7389 35952 7675 36008
rect 7440 35900 7624 35952
rect 7389 35844 7675 35900
rect 7440 35792 7624 35844
rect 7389 35736 7675 35792
rect 7440 35684 7624 35736
rect 7389 35628 7675 35684
rect 7440 35576 7624 35628
rect 7389 35520 7675 35576
rect 7440 35468 7624 35520
rect 7389 35412 7675 35468
rect 7440 35360 7624 35412
rect 7389 35304 7675 35360
rect 7440 35252 7624 35304
rect 7389 35196 7675 35252
rect 7440 35144 7624 35196
rect 7389 35088 7675 35144
rect 7440 35036 7624 35088
rect 7389 34980 7675 35036
rect 7440 34928 7624 34980
rect 7389 34872 7675 34928
rect 7440 34820 7624 34872
rect 7389 34764 7675 34820
rect 7440 34712 7624 34764
rect 7389 34656 7675 34712
rect 7440 34604 7624 34656
rect 7389 34548 7675 34604
rect 7440 34496 7624 34548
rect 7389 34440 7675 34496
rect 7440 34388 7624 34440
rect 7389 34332 7675 34388
rect 7440 34280 7624 34332
rect 7389 34224 7675 34280
rect 7440 34172 7624 34224
rect 7389 34116 7675 34172
rect 7440 34064 7624 34116
rect 7389 34008 7675 34064
rect 7440 33956 7624 34008
rect 7389 33900 7675 33956
rect 7440 33848 7624 33900
rect 7389 33792 7675 33848
rect 7440 33740 7624 33792
rect 7389 33684 7675 33740
rect 7440 33632 7624 33684
rect 7389 33576 7675 33632
rect 7332 33524 7388 33545
rect 7440 33524 7624 33576
rect 7721 33545 7732 36471
rect 7676 33524 7732 33545
rect 7332 33358 7732 33524
rect 7792 36494 8677 36541
rect 8729 36530 10708 36541
rect 8729 36494 8792 36530
rect 7792 36438 8792 36494
rect 7792 36386 8677 36438
rect 8729 36386 8792 36438
rect 7792 36330 8792 36386
rect 7792 36278 8677 36330
rect 8729 36278 8792 36330
rect 7792 36222 8792 36278
rect 7792 36170 8677 36222
rect 8729 36170 8792 36222
rect 7792 36114 8792 36170
rect 7792 36062 8677 36114
rect 8729 36062 8792 36114
rect 7792 36006 8792 36062
rect 7792 35954 8677 36006
rect 8729 35954 8792 36006
rect 7792 35898 8792 35954
rect 7792 35846 8677 35898
rect 8729 35846 8792 35898
rect 7792 35790 8792 35846
rect 7792 35738 8677 35790
rect 8729 35738 8792 35790
rect 7792 35682 8792 35738
rect 7792 35630 8677 35682
rect 8729 35630 8792 35682
rect 7792 35574 8792 35630
rect 7792 35522 8677 35574
rect 8729 35522 8792 35574
rect 7792 35466 8792 35522
rect 7792 35414 8677 35466
rect 8729 35414 8792 35466
rect 7792 35358 8792 35414
rect 7792 35306 8677 35358
rect 8729 35306 8792 35358
rect 7792 35250 8792 35306
rect 7792 35198 8677 35250
rect 8729 35198 8792 35250
rect 7792 35142 8792 35198
rect 7792 35090 8677 35142
rect 8729 35090 8792 35142
rect 7792 35034 8792 35090
rect 7792 34982 8677 35034
rect 8729 34982 8792 35034
rect 7792 34926 8792 34982
rect 7792 34874 8677 34926
rect 8729 34874 8792 34926
rect 7792 34818 8792 34874
rect 7792 34766 8677 34818
rect 8729 34766 8792 34818
rect 7792 34710 8792 34766
rect 7792 34658 8677 34710
rect 8729 34658 8792 34710
rect 7792 34602 8792 34658
rect 7792 34550 8677 34602
rect 8729 34550 8792 34602
rect 7792 34494 8792 34550
rect 7792 34442 8677 34494
rect 8729 34442 8792 34494
rect 7792 34386 8792 34442
rect 7792 34334 8677 34386
rect 8729 34334 8792 34386
rect 7792 34278 8792 34334
rect 7792 34226 8677 34278
rect 8729 34226 8792 34278
rect 7792 34170 8792 34226
rect 7792 34118 8677 34170
rect 8729 34118 8792 34170
rect 7792 34062 8792 34118
rect 7792 34010 8677 34062
rect 8729 34010 8792 34062
rect 7792 33954 8792 34010
rect 7792 33902 8677 33954
rect 8729 33902 8792 33954
rect 7792 33846 8792 33902
rect 7792 33794 8677 33846
rect 8729 33794 8792 33846
rect 7792 33738 8792 33794
rect 7792 33686 8677 33738
rect 8729 33686 8792 33738
rect 7792 33630 8792 33686
rect 7792 33578 8677 33630
rect 8729 33578 8792 33630
rect 7792 33522 8792 33578
rect 7792 33475 8677 33522
rect 8729 33486 8792 33522
rect 9708 33486 10708 36530
rect 11228 36587 14144 36598
rect 11228 36541 11239 36587
rect 14133 36541 14144 36587
rect 8729 33475 10708 33486
rect 7792 33429 7803 33475
rect 10697 33429 10708 33475
rect 7792 33418 10708 33429
rect 10768 36471 11168 36508
rect 10768 33545 10779 36471
rect 10825 33545 11111 36471
rect 11157 33545 11168 36471
rect 10768 33358 11168 33545
rect 11228 36494 11283 36541
rect 11335 36532 13786 36541
rect 13838 36532 13910 36541
rect 13962 36532 14034 36541
rect 14086 36532 14144 36541
rect 11335 36530 14144 36532
rect 11335 36494 12228 36530
rect 11228 36438 12228 36494
rect 11228 36386 11283 36438
rect 11335 36386 12228 36438
rect 11228 36330 12228 36386
rect 11228 36278 11283 36330
rect 11335 36278 12228 36330
rect 11228 36222 12228 36278
rect 11228 36170 11283 36222
rect 11335 36170 12228 36222
rect 11228 36114 12228 36170
rect 11228 36062 11283 36114
rect 11335 36062 12228 36114
rect 11228 36006 12228 36062
rect 11228 35954 11283 36006
rect 11335 35954 12228 36006
rect 11228 35898 12228 35954
rect 11228 35846 11283 35898
rect 11335 35846 12228 35898
rect 11228 35790 12228 35846
rect 11228 35738 11283 35790
rect 11335 35738 12228 35790
rect 11228 35682 12228 35738
rect 11228 35630 11283 35682
rect 11335 35630 12228 35682
rect 11228 35574 12228 35630
rect 11228 35522 11283 35574
rect 11335 35522 12228 35574
rect 11228 35466 12228 35522
rect 11228 35414 11283 35466
rect 11335 35414 12228 35466
rect 11228 35358 12228 35414
rect 11228 35306 11283 35358
rect 11335 35306 12228 35358
rect 11228 35250 12228 35306
rect 11228 35198 11283 35250
rect 11335 35198 12228 35250
rect 11228 35142 12228 35198
rect 11228 35090 11283 35142
rect 11335 35090 12228 35142
rect 11228 35034 12228 35090
rect 11228 34982 11283 35034
rect 11335 34982 12228 35034
rect 11228 34926 12228 34982
rect 11228 34874 11283 34926
rect 11335 34874 12228 34926
rect 11228 34818 12228 34874
rect 11228 34766 11283 34818
rect 11335 34766 12228 34818
rect 11228 34710 12228 34766
rect 11228 34658 11283 34710
rect 11335 34658 12228 34710
rect 11228 34602 12228 34658
rect 11228 34550 11283 34602
rect 11335 34550 12228 34602
rect 11228 34494 12228 34550
rect 11228 34442 11283 34494
rect 11335 34442 12228 34494
rect 11228 34386 12228 34442
rect 11228 34334 11283 34386
rect 11335 34334 12228 34386
rect 11228 34278 12228 34334
rect 11228 34226 11283 34278
rect 11335 34226 12228 34278
rect 11228 34170 12228 34226
rect 11228 34118 11283 34170
rect 11335 34118 12228 34170
rect 11228 34062 12228 34118
rect 11228 34010 11283 34062
rect 11335 34010 12228 34062
rect 11228 33954 12228 34010
rect 11228 33902 11283 33954
rect 11335 33902 12228 33954
rect 11228 33846 12228 33902
rect 11228 33794 11283 33846
rect 11335 33794 12228 33846
rect 11228 33738 12228 33794
rect 11228 33686 11283 33738
rect 11335 33686 12228 33738
rect 11228 33630 12228 33686
rect 11228 33578 11283 33630
rect 11335 33578 12228 33630
rect 11228 33522 12228 33578
rect 11228 33475 11283 33522
rect 11335 33486 12228 33522
rect 13144 36460 14144 36530
rect 13144 36408 13786 36460
rect 13838 36408 13910 36460
rect 13962 36408 14034 36460
rect 14086 36408 14144 36460
rect 13144 36336 14144 36408
rect 13144 36284 13786 36336
rect 13838 36284 13910 36336
rect 13962 36284 14034 36336
rect 14086 36284 14144 36336
rect 13144 36212 14144 36284
rect 13144 36160 13786 36212
rect 13838 36160 13910 36212
rect 13962 36160 14034 36212
rect 14086 36160 14144 36212
rect 13144 36088 14144 36160
rect 13144 36036 13786 36088
rect 13838 36036 13910 36088
rect 13962 36036 14034 36088
rect 14086 36036 14144 36088
rect 13144 35964 14144 36036
rect 13144 35912 13786 35964
rect 13838 35912 13910 35964
rect 13962 35912 14034 35964
rect 14086 35912 14144 35964
rect 13144 35840 14144 35912
rect 13144 35788 13786 35840
rect 13838 35788 13910 35840
rect 13962 35788 14034 35840
rect 14086 35788 14144 35840
rect 13144 35716 14144 35788
rect 13144 35664 13786 35716
rect 13838 35664 13910 35716
rect 13962 35664 14034 35716
rect 14086 35664 14144 35716
rect 13144 35592 14144 35664
rect 13144 35540 13786 35592
rect 13838 35540 13910 35592
rect 13962 35540 14034 35592
rect 14086 35540 14144 35592
rect 13144 35468 14144 35540
rect 13144 35416 13786 35468
rect 13838 35416 13910 35468
rect 13962 35416 14034 35468
rect 14086 35416 14144 35468
rect 13144 35344 14144 35416
rect 13144 35292 13786 35344
rect 13838 35292 13910 35344
rect 13962 35292 14034 35344
rect 14086 35292 14144 35344
rect 13144 35220 14144 35292
rect 13144 35168 13786 35220
rect 13838 35168 13910 35220
rect 13962 35168 14034 35220
rect 14086 35168 14144 35220
rect 13144 35096 14144 35168
rect 13144 35044 13786 35096
rect 13838 35044 13910 35096
rect 13962 35044 14034 35096
rect 14086 35044 14144 35096
rect 13144 34972 14144 35044
rect 13144 34920 13786 34972
rect 13838 34920 13910 34972
rect 13962 34920 14034 34972
rect 14086 34920 14144 34972
rect 13144 34848 14144 34920
rect 13144 34796 13786 34848
rect 13838 34796 13910 34848
rect 13962 34796 14034 34848
rect 14086 34796 14144 34848
rect 13144 34724 14144 34796
rect 13144 34672 13786 34724
rect 13838 34672 13910 34724
rect 13962 34672 14034 34724
rect 14086 34672 14144 34724
rect 13144 34600 14144 34672
rect 13144 34548 13786 34600
rect 13838 34548 13910 34600
rect 13962 34548 14034 34600
rect 14086 34548 14144 34600
rect 13144 34476 14144 34548
rect 13144 34424 13786 34476
rect 13838 34424 13910 34476
rect 13962 34424 14034 34476
rect 14086 34424 14144 34476
rect 13144 34352 14144 34424
rect 13144 34300 13786 34352
rect 13838 34300 13910 34352
rect 13962 34300 14034 34352
rect 14086 34300 14144 34352
rect 13144 34228 14144 34300
rect 13144 34176 13786 34228
rect 13838 34176 13910 34228
rect 13962 34176 14034 34228
rect 14086 34176 14144 34228
rect 13144 34104 14144 34176
rect 13144 34052 13786 34104
rect 13838 34052 13910 34104
rect 13962 34052 14034 34104
rect 14086 34052 14144 34104
rect 13144 33980 14144 34052
rect 13144 33928 13786 33980
rect 13838 33928 13910 33980
rect 13962 33928 14034 33980
rect 14086 33928 14144 33980
rect 13144 33856 14144 33928
rect 13144 33804 13786 33856
rect 13838 33804 13910 33856
rect 13962 33804 14034 33856
rect 14086 33804 14144 33856
rect 13144 33732 14144 33804
rect 13144 33680 13786 33732
rect 13838 33680 13910 33732
rect 13962 33680 14034 33732
rect 14086 33680 14144 33732
rect 13144 33608 14144 33680
rect 13144 33556 13786 33608
rect 13838 33556 13910 33608
rect 13962 33556 14034 33608
rect 14086 33556 14144 33608
rect 13144 33486 14144 33556
rect 11335 33484 14144 33486
rect 11335 33475 13786 33484
rect 13838 33475 13910 33484
rect 13962 33475 14034 33484
rect 14086 33475 14144 33484
rect 11228 33429 11239 33475
rect 14133 33429 14144 33475
rect 11228 33418 14144 33429
rect 14204 36471 14404 36508
rect 14204 33545 14215 36471
rect 14261 33545 14404 36471
rect 14204 33358 14404 33545
rect 14608 33358 14619 36658
rect 445 33308 14619 33358
rect 445 33276 1438 33308
rect 496 33224 552 33276
rect 604 33224 660 33276
rect 712 33256 1438 33276
rect 1490 33256 1562 33308
rect 1614 33256 1686 33308
rect 1738 33256 1810 33308
rect 1862 33256 2574 33308
rect 2626 33256 2698 33308
rect 2750 33256 2822 33308
rect 2874 33256 2946 33308
rect 2998 33256 4846 33308
rect 4898 33256 4970 33308
rect 5022 33256 5094 33308
rect 5146 33256 5218 33308
rect 5270 33256 7139 33308
rect 7191 33256 7263 33308
rect 7315 33256 7387 33308
rect 7439 33256 7625 33308
rect 7677 33256 7749 33308
rect 7801 33256 7873 33308
rect 7925 33256 9794 33308
rect 9846 33256 9918 33308
rect 9970 33256 10042 33308
rect 10094 33256 10166 33308
rect 10218 33256 12066 33308
rect 12118 33256 12190 33308
rect 12242 33256 12314 33308
rect 12366 33256 12438 33308
rect 12490 33256 13202 33308
rect 13254 33256 13326 33308
rect 13378 33256 13450 33308
rect 13502 33256 13574 33308
rect 13626 33276 14619 33308
rect 13626 33256 14352 33276
rect 712 33224 14352 33256
rect 14404 33224 14460 33276
rect 14512 33224 14568 33276
rect 445 33184 14619 33224
rect 445 33168 1438 33184
rect 496 33116 552 33168
rect 604 33116 660 33168
rect 712 33132 1438 33168
rect 1490 33132 1562 33184
rect 1614 33132 1686 33184
rect 1738 33132 1810 33184
rect 1862 33132 2574 33184
rect 2626 33132 2698 33184
rect 2750 33132 2822 33184
rect 2874 33132 2946 33184
rect 2998 33132 4846 33184
rect 4898 33132 4970 33184
rect 5022 33132 5094 33184
rect 5146 33132 5218 33184
rect 5270 33132 7139 33184
rect 7191 33132 7263 33184
rect 7315 33132 7387 33184
rect 7439 33132 7625 33184
rect 7677 33132 7749 33184
rect 7801 33132 7873 33184
rect 7925 33132 9794 33184
rect 9846 33132 9918 33184
rect 9970 33132 10042 33184
rect 10094 33132 10166 33184
rect 10218 33132 12066 33184
rect 12118 33132 12190 33184
rect 12242 33132 12314 33184
rect 12366 33132 12438 33184
rect 12490 33132 13202 33184
rect 13254 33132 13326 33184
rect 13378 33132 13450 33184
rect 13502 33132 13574 33184
rect 13626 33168 14619 33184
rect 13626 33132 14352 33168
rect 712 33116 14352 33132
rect 14404 33116 14460 33168
rect 14512 33116 14568 33168
rect 445 33060 14619 33116
rect 496 33008 552 33060
rect 604 33057 660 33060
rect 712 33057 1438 33060
rect 1490 33057 1562 33060
rect 1614 33057 1686 33060
rect 1738 33057 1810 33060
rect 1862 33057 2574 33060
rect 2626 33057 2698 33060
rect 2750 33057 2822 33060
rect 2874 33057 2946 33060
rect 2998 33057 4846 33060
rect 4898 33057 4970 33060
rect 5022 33057 5094 33060
rect 5146 33057 5218 33060
rect 5270 33057 7139 33060
rect 7191 33057 7263 33060
rect 7315 33057 7387 33060
rect 7439 33057 7625 33060
rect 7677 33057 7749 33060
rect 7801 33057 7873 33060
rect 7925 33057 9794 33060
rect 9846 33057 9918 33060
rect 9970 33057 10042 33060
rect 10094 33057 10166 33060
rect 10218 33057 12066 33060
rect 12118 33057 12190 33060
rect 12242 33057 12314 33060
rect 12366 33057 12438 33060
rect 12490 33057 13202 33060
rect 13254 33057 13326 33060
rect 13378 33057 13450 33060
rect 13502 33057 13574 33060
rect 13626 33057 14352 33060
rect 14404 33057 14460 33060
rect 604 33008 660 33011
rect 712 33008 1438 33011
rect 1490 33008 1562 33011
rect 1614 33008 1686 33011
rect 1738 33008 1810 33011
rect 1862 33008 2574 33011
rect 2626 33008 2698 33011
rect 2750 33008 2822 33011
rect 2874 33008 2946 33011
rect 2998 33008 4846 33011
rect 4898 33008 4970 33011
rect 5022 33008 5094 33011
rect 5146 33008 5218 33011
rect 5270 33008 7139 33011
rect 7191 33008 7263 33011
rect 7315 33008 7387 33011
rect 7439 33008 7625 33011
rect 7677 33008 7749 33011
rect 7801 33008 7873 33011
rect 7925 33008 9794 33011
rect 9846 33008 9918 33011
rect 9970 33008 10042 33011
rect 10094 33008 10166 33011
rect 10218 33008 12066 33011
rect 12118 33008 12190 33011
rect 12242 33008 12314 33011
rect 12366 33008 12438 33011
rect 12490 33008 13202 33011
rect 13254 33008 13326 33011
rect 13378 33008 13450 33011
rect 13502 33008 13574 33011
rect 13626 33008 14352 33011
rect 14404 33008 14460 33011
rect 14512 33008 14568 33060
rect 445 32952 14619 33008
rect 496 32900 552 32952
rect 604 32900 660 32952
rect 712 32936 14352 32952
rect 712 32900 1438 32936
rect 445 32884 1438 32900
rect 1490 32884 1562 32936
rect 1614 32884 1686 32936
rect 1738 32884 1810 32936
rect 1862 32884 2574 32936
rect 2626 32884 2698 32936
rect 2750 32884 2822 32936
rect 2874 32884 2946 32936
rect 2998 32884 4846 32936
rect 4898 32884 4970 32936
rect 5022 32884 5094 32936
rect 5146 32884 5218 32936
rect 5270 32884 7139 32936
rect 7191 32884 7263 32936
rect 7315 32884 7387 32936
rect 7439 32884 7625 32936
rect 7677 32884 7749 32936
rect 7801 32884 7873 32936
rect 7925 32884 9794 32936
rect 9846 32884 9918 32936
rect 9970 32884 10042 32936
rect 10094 32884 10166 32936
rect 10218 32884 12066 32936
rect 12118 32884 12190 32936
rect 12242 32884 12314 32936
rect 12366 32884 12438 32936
rect 12490 32884 13202 32936
rect 13254 32884 13326 32936
rect 13378 32884 13450 32936
rect 13502 32884 13574 32936
rect 13626 32900 14352 32936
rect 14404 32900 14460 32952
rect 14512 32900 14568 32952
rect 13626 32884 14619 32900
rect 445 32844 14619 32884
rect 496 32792 552 32844
rect 604 32792 660 32844
rect 712 32812 14352 32844
rect 712 32792 1438 32812
rect 445 32760 1438 32792
rect 1490 32760 1562 32812
rect 1614 32760 1686 32812
rect 1738 32760 1810 32812
rect 1862 32760 2574 32812
rect 2626 32760 2698 32812
rect 2750 32760 2822 32812
rect 2874 32760 2946 32812
rect 2998 32760 4846 32812
rect 4898 32760 4970 32812
rect 5022 32760 5094 32812
rect 5146 32760 5218 32812
rect 5270 32760 7139 32812
rect 7191 32760 7263 32812
rect 7315 32760 7387 32812
rect 7439 32760 7625 32812
rect 7677 32760 7749 32812
rect 7801 32760 7873 32812
rect 7925 32760 9794 32812
rect 9846 32760 9918 32812
rect 9970 32760 10042 32812
rect 10094 32760 10166 32812
rect 10218 32760 12066 32812
rect 12118 32760 12190 32812
rect 12242 32760 12314 32812
rect 12366 32760 12438 32812
rect 12490 32760 13202 32812
rect 13254 32760 13326 32812
rect 13378 32760 13450 32812
rect 13502 32760 13574 32812
rect 13626 32792 14352 32812
rect 14404 32792 14460 32844
rect 14512 32792 14568 32844
rect 13626 32760 14619 32792
rect 445 32710 14619 32760
rect 445 29410 456 32710
rect 920 32639 3836 32650
rect 920 32593 931 32639
rect 3825 32593 3836 32639
rect 920 32584 978 32593
rect 1030 32584 1102 32593
rect 1154 32584 1226 32593
rect 1278 32584 3729 32593
rect 920 32582 3729 32584
rect 660 32523 860 32560
rect 660 29597 803 32523
rect 849 29597 860 32523
rect 660 29410 860 29597
rect 920 32512 1920 32582
rect 920 32460 978 32512
rect 1030 32460 1102 32512
rect 1154 32460 1226 32512
rect 1278 32460 1920 32512
rect 920 32388 1920 32460
rect 920 32336 978 32388
rect 1030 32336 1102 32388
rect 1154 32336 1226 32388
rect 1278 32336 1920 32388
rect 920 32264 1920 32336
rect 920 32212 978 32264
rect 1030 32212 1102 32264
rect 1154 32212 1226 32264
rect 1278 32212 1920 32264
rect 920 32140 1920 32212
rect 920 32088 978 32140
rect 1030 32088 1102 32140
rect 1154 32088 1226 32140
rect 1278 32088 1920 32140
rect 920 32016 1920 32088
rect 920 31964 978 32016
rect 1030 31964 1102 32016
rect 1154 31964 1226 32016
rect 1278 31964 1920 32016
rect 920 31892 1920 31964
rect 920 31840 978 31892
rect 1030 31840 1102 31892
rect 1154 31840 1226 31892
rect 1278 31840 1920 31892
rect 920 31768 1920 31840
rect 920 31716 978 31768
rect 1030 31716 1102 31768
rect 1154 31716 1226 31768
rect 1278 31716 1920 31768
rect 920 31644 1920 31716
rect 920 31592 978 31644
rect 1030 31592 1102 31644
rect 1154 31592 1226 31644
rect 1278 31592 1920 31644
rect 920 31520 1920 31592
rect 920 31468 978 31520
rect 1030 31468 1102 31520
rect 1154 31468 1226 31520
rect 1278 31468 1920 31520
rect 920 31396 1920 31468
rect 920 31344 978 31396
rect 1030 31344 1102 31396
rect 1154 31344 1226 31396
rect 1278 31344 1920 31396
rect 920 31272 1920 31344
rect 920 31220 978 31272
rect 1030 31220 1102 31272
rect 1154 31220 1226 31272
rect 1278 31220 1920 31272
rect 920 31148 1920 31220
rect 920 31096 978 31148
rect 1030 31096 1102 31148
rect 1154 31096 1226 31148
rect 1278 31096 1920 31148
rect 920 31024 1920 31096
rect 920 30972 978 31024
rect 1030 30972 1102 31024
rect 1154 30972 1226 31024
rect 1278 30972 1920 31024
rect 920 30900 1920 30972
rect 920 30848 978 30900
rect 1030 30848 1102 30900
rect 1154 30848 1226 30900
rect 1278 30848 1920 30900
rect 920 30776 1920 30848
rect 920 30724 978 30776
rect 1030 30724 1102 30776
rect 1154 30724 1226 30776
rect 1278 30724 1920 30776
rect 920 30652 1920 30724
rect 920 30600 978 30652
rect 1030 30600 1102 30652
rect 1154 30600 1226 30652
rect 1278 30600 1920 30652
rect 920 30528 1920 30600
rect 920 30476 978 30528
rect 1030 30476 1102 30528
rect 1154 30476 1226 30528
rect 1278 30476 1920 30528
rect 920 30404 1920 30476
rect 920 30352 978 30404
rect 1030 30352 1102 30404
rect 1154 30352 1226 30404
rect 1278 30352 1920 30404
rect 920 30280 1920 30352
rect 920 30228 978 30280
rect 1030 30228 1102 30280
rect 1154 30228 1226 30280
rect 1278 30228 1920 30280
rect 920 30156 1920 30228
rect 920 30104 978 30156
rect 1030 30104 1102 30156
rect 1154 30104 1226 30156
rect 1278 30104 1920 30156
rect 920 30032 1920 30104
rect 920 29980 978 30032
rect 1030 29980 1102 30032
rect 1154 29980 1226 30032
rect 1278 29980 1920 30032
rect 920 29908 1920 29980
rect 920 29856 978 29908
rect 1030 29856 1102 29908
rect 1154 29856 1226 29908
rect 1278 29856 1920 29908
rect 920 29784 1920 29856
rect 920 29732 978 29784
rect 1030 29732 1102 29784
rect 1154 29732 1226 29784
rect 1278 29732 1920 29784
rect 920 29660 1920 29732
rect 920 29608 978 29660
rect 1030 29608 1102 29660
rect 1154 29608 1226 29660
rect 1278 29608 1920 29660
rect 920 29538 1920 29608
rect 2836 32546 3729 32582
rect 3781 32546 3836 32593
rect 4356 32639 7272 32650
rect 4356 32593 4367 32639
rect 7261 32593 7272 32639
rect 4356 32582 6335 32593
rect 2836 32490 3836 32546
rect 2836 32438 3729 32490
rect 3781 32438 3836 32490
rect 2836 32382 3836 32438
rect 2836 32330 3729 32382
rect 3781 32330 3836 32382
rect 2836 32274 3836 32330
rect 2836 32222 3729 32274
rect 3781 32222 3836 32274
rect 2836 32166 3836 32222
rect 2836 32114 3729 32166
rect 3781 32114 3836 32166
rect 2836 32058 3836 32114
rect 2836 32006 3729 32058
rect 3781 32006 3836 32058
rect 2836 31950 3836 32006
rect 2836 31898 3729 31950
rect 3781 31898 3836 31950
rect 2836 31842 3836 31898
rect 2836 31790 3729 31842
rect 3781 31790 3836 31842
rect 2836 31734 3836 31790
rect 2836 31682 3729 31734
rect 3781 31682 3836 31734
rect 2836 31626 3836 31682
rect 2836 31574 3729 31626
rect 3781 31574 3836 31626
rect 2836 31518 3836 31574
rect 2836 31466 3729 31518
rect 3781 31466 3836 31518
rect 2836 31410 3836 31466
rect 2836 31358 3729 31410
rect 3781 31358 3836 31410
rect 2836 31302 3836 31358
rect 2836 31250 3729 31302
rect 3781 31250 3836 31302
rect 2836 31194 3836 31250
rect 2836 31142 3729 31194
rect 3781 31142 3836 31194
rect 2836 31086 3836 31142
rect 2836 31034 3729 31086
rect 3781 31034 3836 31086
rect 2836 30978 3836 31034
rect 2836 30926 3729 30978
rect 3781 30926 3836 30978
rect 2836 30870 3836 30926
rect 2836 30818 3729 30870
rect 3781 30818 3836 30870
rect 2836 30762 3836 30818
rect 2836 30710 3729 30762
rect 3781 30710 3836 30762
rect 2836 30654 3836 30710
rect 2836 30602 3729 30654
rect 3781 30602 3836 30654
rect 2836 30546 3836 30602
rect 2836 30494 3729 30546
rect 3781 30494 3836 30546
rect 2836 30438 3836 30494
rect 2836 30386 3729 30438
rect 3781 30386 3836 30438
rect 2836 30330 3836 30386
rect 2836 30278 3729 30330
rect 3781 30278 3836 30330
rect 2836 30222 3836 30278
rect 2836 30170 3729 30222
rect 3781 30170 3836 30222
rect 2836 30114 3836 30170
rect 2836 30062 3729 30114
rect 3781 30062 3836 30114
rect 2836 30006 3836 30062
rect 2836 29954 3729 30006
rect 3781 29954 3836 30006
rect 2836 29898 3836 29954
rect 2836 29846 3729 29898
rect 3781 29846 3836 29898
rect 2836 29790 3836 29846
rect 2836 29738 3729 29790
rect 3781 29738 3836 29790
rect 2836 29682 3836 29738
rect 2836 29630 3729 29682
rect 3781 29630 3836 29682
rect 2836 29574 3836 29630
rect 2836 29538 3729 29574
rect 920 29536 3729 29538
rect 920 29527 978 29536
rect 1030 29527 1102 29536
rect 1154 29527 1226 29536
rect 1278 29527 3729 29536
rect 3781 29527 3836 29574
rect 920 29481 931 29527
rect 3825 29481 3836 29527
rect 920 29470 3836 29481
rect 3896 32523 4296 32560
rect 3896 29597 3907 32523
rect 3953 29597 4239 32523
rect 4285 29597 4296 32523
rect 3896 29410 4296 29597
rect 4356 29538 5356 32582
rect 6272 32546 6335 32582
rect 6387 32546 7272 32593
rect 7792 32639 10708 32650
rect 7792 32593 7803 32639
rect 10697 32593 10708 32639
rect 6272 32490 7272 32546
rect 6272 32438 6335 32490
rect 6387 32438 7272 32490
rect 6272 32382 7272 32438
rect 6272 32330 6335 32382
rect 6387 32330 7272 32382
rect 6272 32274 7272 32330
rect 6272 32222 6335 32274
rect 6387 32222 7272 32274
rect 6272 32166 7272 32222
rect 6272 32114 6335 32166
rect 6387 32114 7272 32166
rect 6272 32058 7272 32114
rect 6272 32006 6335 32058
rect 6387 32006 7272 32058
rect 6272 31950 7272 32006
rect 6272 31898 6335 31950
rect 6387 31898 7272 31950
rect 6272 31842 7272 31898
rect 6272 31790 6335 31842
rect 6387 31790 7272 31842
rect 6272 31734 7272 31790
rect 6272 31682 6335 31734
rect 6387 31682 7272 31734
rect 6272 31626 7272 31682
rect 6272 31574 6335 31626
rect 6387 31574 7272 31626
rect 6272 31518 7272 31574
rect 6272 31466 6335 31518
rect 6387 31466 7272 31518
rect 6272 31410 7272 31466
rect 6272 31358 6335 31410
rect 6387 31358 7272 31410
rect 6272 31302 7272 31358
rect 6272 31250 6335 31302
rect 6387 31250 7272 31302
rect 6272 31194 7272 31250
rect 6272 31142 6335 31194
rect 6387 31142 7272 31194
rect 6272 31086 7272 31142
rect 6272 31034 6335 31086
rect 6387 31034 7272 31086
rect 6272 30978 7272 31034
rect 6272 30926 6335 30978
rect 6387 30926 7272 30978
rect 6272 30870 7272 30926
rect 6272 30818 6335 30870
rect 6387 30818 7272 30870
rect 6272 30762 7272 30818
rect 6272 30710 6335 30762
rect 6387 30710 7272 30762
rect 6272 30654 7272 30710
rect 6272 30602 6335 30654
rect 6387 30602 7272 30654
rect 6272 30546 7272 30602
rect 6272 30494 6335 30546
rect 6387 30494 7272 30546
rect 6272 30438 7272 30494
rect 6272 30386 6335 30438
rect 6387 30386 7272 30438
rect 6272 30330 7272 30386
rect 6272 30278 6335 30330
rect 6387 30278 7272 30330
rect 6272 30222 7272 30278
rect 6272 30170 6335 30222
rect 6387 30170 7272 30222
rect 6272 30114 7272 30170
rect 6272 30062 6335 30114
rect 6387 30062 7272 30114
rect 6272 30006 7272 30062
rect 6272 29954 6335 30006
rect 6387 29954 7272 30006
rect 6272 29898 7272 29954
rect 6272 29846 6335 29898
rect 6387 29846 7272 29898
rect 6272 29790 7272 29846
rect 6272 29738 6335 29790
rect 6387 29738 7272 29790
rect 6272 29682 7272 29738
rect 6272 29630 6335 29682
rect 6387 29630 7272 29682
rect 6272 29574 7272 29630
rect 6272 29538 6335 29574
rect 4356 29527 6335 29538
rect 6387 29527 7272 29574
rect 4356 29481 4367 29527
rect 7261 29481 7272 29527
rect 4356 29470 7272 29481
rect 7332 32544 7732 32560
rect 7332 32523 7388 32544
rect 7332 29597 7343 32523
rect 7440 32492 7624 32544
rect 7676 32523 7732 32544
rect 7389 32436 7675 32492
rect 7440 32384 7624 32436
rect 7389 32328 7675 32384
rect 7440 32276 7624 32328
rect 7389 32220 7675 32276
rect 7440 32168 7624 32220
rect 7389 32112 7675 32168
rect 7440 32060 7624 32112
rect 7389 32004 7675 32060
rect 7440 31952 7624 32004
rect 7389 31896 7675 31952
rect 7440 31844 7624 31896
rect 7389 31788 7675 31844
rect 7440 31736 7624 31788
rect 7389 31680 7675 31736
rect 7440 31628 7624 31680
rect 7389 31572 7675 31628
rect 7440 31520 7624 31572
rect 7389 31464 7675 31520
rect 7440 31412 7624 31464
rect 7389 31356 7675 31412
rect 7440 31304 7624 31356
rect 7389 31248 7675 31304
rect 7440 31196 7624 31248
rect 7389 31140 7675 31196
rect 7440 31088 7624 31140
rect 7389 31032 7675 31088
rect 7440 30980 7624 31032
rect 7389 30924 7675 30980
rect 7440 30872 7624 30924
rect 7389 30816 7675 30872
rect 7440 30764 7624 30816
rect 7389 30708 7675 30764
rect 7440 30656 7624 30708
rect 7389 30600 7675 30656
rect 7440 30548 7624 30600
rect 7389 30492 7675 30548
rect 7440 30440 7624 30492
rect 7389 30384 7675 30440
rect 7440 30332 7624 30384
rect 7389 30276 7675 30332
rect 7440 30224 7624 30276
rect 7389 30168 7675 30224
rect 7440 30116 7624 30168
rect 7389 30060 7675 30116
rect 7440 30008 7624 30060
rect 7389 29952 7675 30008
rect 7440 29900 7624 29952
rect 7389 29844 7675 29900
rect 7440 29792 7624 29844
rect 7389 29736 7675 29792
rect 7440 29684 7624 29736
rect 7389 29628 7675 29684
rect 7332 29576 7388 29597
rect 7440 29576 7624 29628
rect 7721 29597 7732 32523
rect 7676 29576 7732 29597
rect 7332 29410 7732 29576
rect 7792 32546 8677 32593
rect 8729 32582 10708 32593
rect 8729 32546 8792 32582
rect 7792 32490 8792 32546
rect 7792 32438 8677 32490
rect 8729 32438 8792 32490
rect 7792 32382 8792 32438
rect 7792 32330 8677 32382
rect 8729 32330 8792 32382
rect 7792 32274 8792 32330
rect 7792 32222 8677 32274
rect 8729 32222 8792 32274
rect 7792 32166 8792 32222
rect 7792 32114 8677 32166
rect 8729 32114 8792 32166
rect 7792 32058 8792 32114
rect 7792 32006 8677 32058
rect 8729 32006 8792 32058
rect 7792 31950 8792 32006
rect 7792 31898 8677 31950
rect 8729 31898 8792 31950
rect 7792 31842 8792 31898
rect 7792 31790 8677 31842
rect 8729 31790 8792 31842
rect 7792 31734 8792 31790
rect 7792 31682 8677 31734
rect 8729 31682 8792 31734
rect 7792 31626 8792 31682
rect 7792 31574 8677 31626
rect 8729 31574 8792 31626
rect 7792 31518 8792 31574
rect 7792 31466 8677 31518
rect 8729 31466 8792 31518
rect 7792 31410 8792 31466
rect 7792 31358 8677 31410
rect 8729 31358 8792 31410
rect 7792 31302 8792 31358
rect 7792 31250 8677 31302
rect 8729 31250 8792 31302
rect 7792 31194 8792 31250
rect 7792 31142 8677 31194
rect 8729 31142 8792 31194
rect 7792 31086 8792 31142
rect 7792 31034 8677 31086
rect 8729 31034 8792 31086
rect 7792 30978 8792 31034
rect 7792 30926 8677 30978
rect 8729 30926 8792 30978
rect 7792 30870 8792 30926
rect 7792 30818 8677 30870
rect 8729 30818 8792 30870
rect 7792 30762 8792 30818
rect 7792 30710 8677 30762
rect 8729 30710 8792 30762
rect 7792 30654 8792 30710
rect 7792 30602 8677 30654
rect 8729 30602 8792 30654
rect 7792 30546 8792 30602
rect 7792 30494 8677 30546
rect 8729 30494 8792 30546
rect 7792 30438 8792 30494
rect 7792 30386 8677 30438
rect 8729 30386 8792 30438
rect 7792 30330 8792 30386
rect 7792 30278 8677 30330
rect 8729 30278 8792 30330
rect 7792 30222 8792 30278
rect 7792 30170 8677 30222
rect 8729 30170 8792 30222
rect 7792 30114 8792 30170
rect 7792 30062 8677 30114
rect 8729 30062 8792 30114
rect 7792 30006 8792 30062
rect 7792 29954 8677 30006
rect 8729 29954 8792 30006
rect 7792 29898 8792 29954
rect 7792 29846 8677 29898
rect 8729 29846 8792 29898
rect 7792 29790 8792 29846
rect 7792 29738 8677 29790
rect 8729 29738 8792 29790
rect 7792 29682 8792 29738
rect 7792 29630 8677 29682
rect 8729 29630 8792 29682
rect 7792 29574 8792 29630
rect 7792 29527 8677 29574
rect 8729 29538 8792 29574
rect 9708 29538 10708 32582
rect 11228 32639 14144 32650
rect 11228 32593 11239 32639
rect 14133 32593 14144 32639
rect 8729 29527 10708 29538
rect 7792 29481 7803 29527
rect 10697 29481 10708 29527
rect 7792 29470 10708 29481
rect 10768 32523 11168 32560
rect 10768 29597 10779 32523
rect 10825 29597 11111 32523
rect 11157 29597 11168 32523
rect 10768 29410 11168 29597
rect 11228 32546 11283 32593
rect 11335 32584 13786 32593
rect 13838 32584 13910 32593
rect 13962 32584 14034 32593
rect 14086 32584 14144 32593
rect 11335 32582 14144 32584
rect 11335 32546 12228 32582
rect 11228 32490 12228 32546
rect 11228 32438 11283 32490
rect 11335 32438 12228 32490
rect 11228 32382 12228 32438
rect 11228 32330 11283 32382
rect 11335 32330 12228 32382
rect 11228 32274 12228 32330
rect 11228 32222 11283 32274
rect 11335 32222 12228 32274
rect 11228 32166 12228 32222
rect 11228 32114 11283 32166
rect 11335 32114 12228 32166
rect 11228 32058 12228 32114
rect 11228 32006 11283 32058
rect 11335 32006 12228 32058
rect 11228 31950 12228 32006
rect 11228 31898 11283 31950
rect 11335 31898 12228 31950
rect 11228 31842 12228 31898
rect 11228 31790 11283 31842
rect 11335 31790 12228 31842
rect 11228 31734 12228 31790
rect 11228 31682 11283 31734
rect 11335 31682 12228 31734
rect 11228 31626 12228 31682
rect 11228 31574 11283 31626
rect 11335 31574 12228 31626
rect 11228 31518 12228 31574
rect 11228 31466 11283 31518
rect 11335 31466 12228 31518
rect 11228 31410 12228 31466
rect 11228 31358 11283 31410
rect 11335 31358 12228 31410
rect 11228 31302 12228 31358
rect 11228 31250 11283 31302
rect 11335 31250 12228 31302
rect 11228 31194 12228 31250
rect 11228 31142 11283 31194
rect 11335 31142 12228 31194
rect 11228 31086 12228 31142
rect 11228 31034 11283 31086
rect 11335 31034 12228 31086
rect 11228 30978 12228 31034
rect 11228 30926 11283 30978
rect 11335 30926 12228 30978
rect 11228 30870 12228 30926
rect 11228 30818 11283 30870
rect 11335 30818 12228 30870
rect 11228 30762 12228 30818
rect 11228 30710 11283 30762
rect 11335 30710 12228 30762
rect 11228 30654 12228 30710
rect 11228 30602 11283 30654
rect 11335 30602 12228 30654
rect 11228 30546 12228 30602
rect 11228 30494 11283 30546
rect 11335 30494 12228 30546
rect 11228 30438 12228 30494
rect 11228 30386 11283 30438
rect 11335 30386 12228 30438
rect 11228 30330 12228 30386
rect 11228 30278 11283 30330
rect 11335 30278 12228 30330
rect 11228 30222 12228 30278
rect 11228 30170 11283 30222
rect 11335 30170 12228 30222
rect 11228 30114 12228 30170
rect 11228 30062 11283 30114
rect 11335 30062 12228 30114
rect 11228 30006 12228 30062
rect 11228 29954 11283 30006
rect 11335 29954 12228 30006
rect 11228 29898 12228 29954
rect 11228 29846 11283 29898
rect 11335 29846 12228 29898
rect 11228 29790 12228 29846
rect 11228 29738 11283 29790
rect 11335 29738 12228 29790
rect 11228 29682 12228 29738
rect 11228 29630 11283 29682
rect 11335 29630 12228 29682
rect 11228 29574 12228 29630
rect 11228 29527 11283 29574
rect 11335 29538 12228 29574
rect 13144 32512 14144 32582
rect 13144 32460 13786 32512
rect 13838 32460 13910 32512
rect 13962 32460 14034 32512
rect 14086 32460 14144 32512
rect 13144 32388 14144 32460
rect 13144 32336 13786 32388
rect 13838 32336 13910 32388
rect 13962 32336 14034 32388
rect 14086 32336 14144 32388
rect 13144 32264 14144 32336
rect 13144 32212 13786 32264
rect 13838 32212 13910 32264
rect 13962 32212 14034 32264
rect 14086 32212 14144 32264
rect 13144 32140 14144 32212
rect 13144 32088 13786 32140
rect 13838 32088 13910 32140
rect 13962 32088 14034 32140
rect 14086 32088 14144 32140
rect 13144 32016 14144 32088
rect 13144 31964 13786 32016
rect 13838 31964 13910 32016
rect 13962 31964 14034 32016
rect 14086 31964 14144 32016
rect 13144 31892 14144 31964
rect 13144 31840 13786 31892
rect 13838 31840 13910 31892
rect 13962 31840 14034 31892
rect 14086 31840 14144 31892
rect 13144 31768 14144 31840
rect 13144 31716 13786 31768
rect 13838 31716 13910 31768
rect 13962 31716 14034 31768
rect 14086 31716 14144 31768
rect 13144 31644 14144 31716
rect 13144 31592 13786 31644
rect 13838 31592 13910 31644
rect 13962 31592 14034 31644
rect 14086 31592 14144 31644
rect 13144 31520 14144 31592
rect 13144 31468 13786 31520
rect 13838 31468 13910 31520
rect 13962 31468 14034 31520
rect 14086 31468 14144 31520
rect 13144 31396 14144 31468
rect 13144 31344 13786 31396
rect 13838 31344 13910 31396
rect 13962 31344 14034 31396
rect 14086 31344 14144 31396
rect 13144 31272 14144 31344
rect 13144 31220 13786 31272
rect 13838 31220 13910 31272
rect 13962 31220 14034 31272
rect 14086 31220 14144 31272
rect 13144 31148 14144 31220
rect 13144 31096 13786 31148
rect 13838 31096 13910 31148
rect 13962 31096 14034 31148
rect 14086 31096 14144 31148
rect 13144 31024 14144 31096
rect 13144 30972 13786 31024
rect 13838 30972 13910 31024
rect 13962 30972 14034 31024
rect 14086 30972 14144 31024
rect 13144 30900 14144 30972
rect 13144 30848 13786 30900
rect 13838 30848 13910 30900
rect 13962 30848 14034 30900
rect 14086 30848 14144 30900
rect 13144 30776 14144 30848
rect 13144 30724 13786 30776
rect 13838 30724 13910 30776
rect 13962 30724 14034 30776
rect 14086 30724 14144 30776
rect 13144 30652 14144 30724
rect 13144 30600 13786 30652
rect 13838 30600 13910 30652
rect 13962 30600 14034 30652
rect 14086 30600 14144 30652
rect 13144 30528 14144 30600
rect 13144 30476 13786 30528
rect 13838 30476 13910 30528
rect 13962 30476 14034 30528
rect 14086 30476 14144 30528
rect 13144 30404 14144 30476
rect 13144 30352 13786 30404
rect 13838 30352 13910 30404
rect 13962 30352 14034 30404
rect 14086 30352 14144 30404
rect 13144 30280 14144 30352
rect 13144 30228 13786 30280
rect 13838 30228 13910 30280
rect 13962 30228 14034 30280
rect 14086 30228 14144 30280
rect 13144 30156 14144 30228
rect 13144 30104 13786 30156
rect 13838 30104 13910 30156
rect 13962 30104 14034 30156
rect 14086 30104 14144 30156
rect 13144 30032 14144 30104
rect 13144 29980 13786 30032
rect 13838 29980 13910 30032
rect 13962 29980 14034 30032
rect 14086 29980 14144 30032
rect 13144 29908 14144 29980
rect 13144 29856 13786 29908
rect 13838 29856 13910 29908
rect 13962 29856 14034 29908
rect 14086 29856 14144 29908
rect 13144 29784 14144 29856
rect 13144 29732 13786 29784
rect 13838 29732 13910 29784
rect 13962 29732 14034 29784
rect 14086 29732 14144 29784
rect 13144 29660 14144 29732
rect 13144 29608 13786 29660
rect 13838 29608 13910 29660
rect 13962 29608 14034 29660
rect 14086 29608 14144 29660
rect 13144 29538 14144 29608
rect 11335 29536 14144 29538
rect 11335 29527 13786 29536
rect 13838 29527 13910 29536
rect 13962 29527 14034 29536
rect 14086 29527 14144 29536
rect 11228 29481 11239 29527
rect 14133 29481 14144 29527
rect 11228 29470 14144 29481
rect 14204 32523 14404 32560
rect 14204 29597 14215 32523
rect 14261 29597 14404 32523
rect 14204 29410 14404 29597
rect 14608 29410 14619 32710
rect 445 29360 14619 29410
rect 445 29328 1438 29360
rect 496 29276 552 29328
rect 604 29276 660 29328
rect 712 29308 1438 29328
rect 1490 29308 1562 29360
rect 1614 29308 1686 29360
rect 1738 29308 1810 29360
rect 1862 29308 2574 29360
rect 2626 29308 2698 29360
rect 2750 29308 2822 29360
rect 2874 29308 2946 29360
rect 2998 29308 4846 29360
rect 4898 29308 4970 29360
rect 5022 29308 5094 29360
rect 5146 29308 5218 29360
rect 5270 29308 7139 29360
rect 7191 29308 7263 29360
rect 7315 29308 7387 29360
rect 7439 29308 7625 29360
rect 7677 29308 7749 29360
rect 7801 29308 7873 29360
rect 7925 29308 9794 29360
rect 9846 29308 9918 29360
rect 9970 29308 10042 29360
rect 10094 29308 10166 29360
rect 10218 29308 12066 29360
rect 12118 29308 12190 29360
rect 12242 29308 12314 29360
rect 12366 29308 12438 29360
rect 12490 29308 13202 29360
rect 13254 29308 13326 29360
rect 13378 29308 13450 29360
rect 13502 29308 13574 29360
rect 13626 29328 14619 29360
rect 13626 29308 14352 29328
rect 712 29276 14352 29308
rect 14404 29276 14460 29328
rect 14512 29276 14568 29328
rect 445 29236 14619 29276
rect 445 29220 1438 29236
rect 496 29168 552 29220
rect 604 29168 660 29220
rect 712 29184 1438 29220
rect 1490 29184 1562 29236
rect 1614 29184 1686 29236
rect 1738 29184 1810 29236
rect 1862 29184 2574 29236
rect 2626 29184 2698 29236
rect 2750 29184 2822 29236
rect 2874 29184 2946 29236
rect 2998 29184 4846 29236
rect 4898 29184 4970 29236
rect 5022 29184 5094 29236
rect 5146 29184 5218 29236
rect 5270 29184 7139 29236
rect 7191 29184 7263 29236
rect 7315 29184 7387 29236
rect 7439 29184 7625 29236
rect 7677 29184 7749 29236
rect 7801 29184 7873 29236
rect 7925 29184 9794 29236
rect 9846 29184 9918 29236
rect 9970 29184 10042 29236
rect 10094 29184 10166 29236
rect 10218 29184 12066 29236
rect 12118 29184 12190 29236
rect 12242 29184 12314 29236
rect 12366 29184 12438 29236
rect 12490 29184 13202 29236
rect 13254 29184 13326 29236
rect 13378 29184 13450 29236
rect 13502 29184 13574 29236
rect 13626 29220 14619 29236
rect 13626 29184 14352 29220
rect 712 29168 14352 29184
rect 14404 29168 14460 29220
rect 14512 29168 14568 29220
rect 445 29112 14619 29168
rect 496 29060 552 29112
rect 604 29109 660 29112
rect 712 29109 1438 29112
rect 1490 29109 1562 29112
rect 1614 29109 1686 29112
rect 1738 29109 1810 29112
rect 1862 29109 2574 29112
rect 2626 29109 2698 29112
rect 2750 29109 2822 29112
rect 2874 29109 2946 29112
rect 2998 29109 4846 29112
rect 4898 29109 4970 29112
rect 5022 29109 5094 29112
rect 5146 29109 5218 29112
rect 5270 29109 7139 29112
rect 7191 29109 7263 29112
rect 7315 29109 7387 29112
rect 7439 29109 7625 29112
rect 7677 29109 7749 29112
rect 7801 29109 7873 29112
rect 7925 29109 9794 29112
rect 9846 29109 9918 29112
rect 9970 29109 10042 29112
rect 10094 29109 10166 29112
rect 10218 29109 12066 29112
rect 12118 29109 12190 29112
rect 12242 29109 12314 29112
rect 12366 29109 12438 29112
rect 12490 29109 13202 29112
rect 13254 29109 13326 29112
rect 13378 29109 13450 29112
rect 13502 29109 13574 29112
rect 13626 29109 14352 29112
rect 14404 29109 14460 29112
rect 604 29060 660 29063
rect 712 29060 1438 29063
rect 1490 29060 1562 29063
rect 1614 29060 1686 29063
rect 1738 29060 1810 29063
rect 1862 29060 2574 29063
rect 2626 29060 2698 29063
rect 2750 29060 2822 29063
rect 2874 29060 2946 29063
rect 2998 29060 4846 29063
rect 4898 29060 4970 29063
rect 5022 29060 5094 29063
rect 5146 29060 5218 29063
rect 5270 29060 7139 29063
rect 7191 29060 7263 29063
rect 7315 29060 7387 29063
rect 7439 29060 7625 29063
rect 7677 29060 7749 29063
rect 7801 29060 7873 29063
rect 7925 29060 9794 29063
rect 9846 29060 9918 29063
rect 9970 29060 10042 29063
rect 10094 29060 10166 29063
rect 10218 29060 12066 29063
rect 12118 29060 12190 29063
rect 12242 29060 12314 29063
rect 12366 29060 12438 29063
rect 12490 29060 13202 29063
rect 13254 29060 13326 29063
rect 13378 29060 13450 29063
rect 13502 29060 13574 29063
rect 13626 29060 14352 29063
rect 14404 29060 14460 29063
rect 14512 29060 14568 29112
rect 445 29004 14619 29060
rect 496 28952 552 29004
rect 604 28952 660 29004
rect 712 28988 14352 29004
rect 712 28952 1438 28988
rect 445 28936 1438 28952
rect 1490 28936 1562 28988
rect 1614 28936 1686 28988
rect 1738 28936 1810 28988
rect 1862 28936 2574 28988
rect 2626 28936 2698 28988
rect 2750 28936 2822 28988
rect 2874 28936 2946 28988
rect 2998 28936 4846 28988
rect 4898 28936 4970 28988
rect 5022 28936 5094 28988
rect 5146 28936 5218 28988
rect 5270 28936 7139 28988
rect 7191 28936 7263 28988
rect 7315 28936 7387 28988
rect 7439 28936 7625 28988
rect 7677 28936 7749 28988
rect 7801 28936 7873 28988
rect 7925 28936 9794 28988
rect 9846 28936 9918 28988
rect 9970 28936 10042 28988
rect 10094 28936 10166 28988
rect 10218 28936 12066 28988
rect 12118 28936 12190 28988
rect 12242 28936 12314 28988
rect 12366 28936 12438 28988
rect 12490 28936 13202 28988
rect 13254 28936 13326 28988
rect 13378 28936 13450 28988
rect 13502 28936 13574 28988
rect 13626 28952 14352 28988
rect 14404 28952 14460 29004
rect 14512 28952 14568 29004
rect 13626 28936 14619 28952
rect 445 28896 14619 28936
rect 496 28844 552 28896
rect 604 28844 660 28896
rect 712 28864 14352 28896
rect 712 28844 1438 28864
rect 445 28812 1438 28844
rect 1490 28812 1562 28864
rect 1614 28812 1686 28864
rect 1738 28812 1810 28864
rect 1862 28812 2574 28864
rect 2626 28812 2698 28864
rect 2750 28812 2822 28864
rect 2874 28812 2946 28864
rect 2998 28812 4846 28864
rect 4898 28812 4970 28864
rect 5022 28812 5094 28864
rect 5146 28812 5218 28864
rect 5270 28812 7139 28864
rect 7191 28812 7263 28864
rect 7315 28812 7387 28864
rect 7439 28812 7625 28864
rect 7677 28812 7749 28864
rect 7801 28812 7873 28864
rect 7925 28812 9794 28864
rect 9846 28812 9918 28864
rect 9970 28812 10042 28864
rect 10094 28812 10166 28864
rect 10218 28812 12066 28864
rect 12118 28812 12190 28864
rect 12242 28812 12314 28864
rect 12366 28812 12438 28864
rect 12490 28812 13202 28864
rect 13254 28812 13326 28864
rect 13378 28812 13450 28864
rect 13502 28812 13574 28864
rect 13626 28844 14352 28864
rect 14404 28844 14460 28896
rect 14512 28844 14568 28896
rect 13626 28812 14619 28844
rect 445 28762 14619 28812
rect 445 25462 456 28762
rect 920 28691 3836 28702
rect 920 28645 931 28691
rect 3825 28645 3836 28691
rect 920 28636 978 28645
rect 1030 28636 1102 28645
rect 1154 28636 1226 28645
rect 1278 28636 3729 28645
rect 920 28634 3729 28636
rect 660 28575 860 28612
rect 660 25649 803 28575
rect 849 25649 860 28575
rect 660 25462 860 25649
rect 920 28564 1920 28634
rect 920 28512 978 28564
rect 1030 28512 1102 28564
rect 1154 28512 1226 28564
rect 1278 28512 1920 28564
rect 920 28440 1920 28512
rect 920 28388 978 28440
rect 1030 28388 1102 28440
rect 1154 28388 1226 28440
rect 1278 28388 1920 28440
rect 920 28316 1920 28388
rect 920 28264 978 28316
rect 1030 28264 1102 28316
rect 1154 28264 1226 28316
rect 1278 28264 1920 28316
rect 920 28192 1920 28264
rect 920 28140 978 28192
rect 1030 28140 1102 28192
rect 1154 28140 1226 28192
rect 1278 28140 1920 28192
rect 920 28068 1920 28140
rect 920 28016 978 28068
rect 1030 28016 1102 28068
rect 1154 28016 1226 28068
rect 1278 28016 1920 28068
rect 920 27944 1920 28016
rect 920 27892 978 27944
rect 1030 27892 1102 27944
rect 1154 27892 1226 27944
rect 1278 27892 1920 27944
rect 920 27820 1920 27892
rect 920 27768 978 27820
rect 1030 27768 1102 27820
rect 1154 27768 1226 27820
rect 1278 27768 1920 27820
rect 920 27696 1920 27768
rect 920 27644 978 27696
rect 1030 27644 1102 27696
rect 1154 27644 1226 27696
rect 1278 27644 1920 27696
rect 920 27572 1920 27644
rect 920 27520 978 27572
rect 1030 27520 1102 27572
rect 1154 27520 1226 27572
rect 1278 27520 1920 27572
rect 920 27448 1920 27520
rect 920 27396 978 27448
rect 1030 27396 1102 27448
rect 1154 27396 1226 27448
rect 1278 27396 1920 27448
rect 920 27324 1920 27396
rect 920 27272 978 27324
rect 1030 27272 1102 27324
rect 1154 27272 1226 27324
rect 1278 27272 1920 27324
rect 920 27200 1920 27272
rect 920 27148 978 27200
rect 1030 27148 1102 27200
rect 1154 27148 1226 27200
rect 1278 27148 1920 27200
rect 920 27076 1920 27148
rect 920 27024 978 27076
rect 1030 27024 1102 27076
rect 1154 27024 1226 27076
rect 1278 27024 1920 27076
rect 920 26952 1920 27024
rect 920 26900 978 26952
rect 1030 26900 1102 26952
rect 1154 26900 1226 26952
rect 1278 26900 1920 26952
rect 920 26828 1920 26900
rect 920 26776 978 26828
rect 1030 26776 1102 26828
rect 1154 26776 1226 26828
rect 1278 26776 1920 26828
rect 920 26704 1920 26776
rect 920 26652 978 26704
rect 1030 26652 1102 26704
rect 1154 26652 1226 26704
rect 1278 26652 1920 26704
rect 920 26580 1920 26652
rect 920 26528 978 26580
rect 1030 26528 1102 26580
rect 1154 26528 1226 26580
rect 1278 26528 1920 26580
rect 920 26456 1920 26528
rect 920 26404 978 26456
rect 1030 26404 1102 26456
rect 1154 26404 1226 26456
rect 1278 26404 1920 26456
rect 920 26332 1920 26404
rect 920 26280 978 26332
rect 1030 26280 1102 26332
rect 1154 26280 1226 26332
rect 1278 26280 1920 26332
rect 920 26208 1920 26280
rect 920 26156 978 26208
rect 1030 26156 1102 26208
rect 1154 26156 1226 26208
rect 1278 26156 1920 26208
rect 920 26084 1920 26156
rect 920 26032 978 26084
rect 1030 26032 1102 26084
rect 1154 26032 1226 26084
rect 1278 26032 1920 26084
rect 920 25960 1920 26032
rect 920 25908 978 25960
rect 1030 25908 1102 25960
rect 1154 25908 1226 25960
rect 1278 25908 1920 25960
rect 920 25836 1920 25908
rect 920 25784 978 25836
rect 1030 25784 1102 25836
rect 1154 25784 1226 25836
rect 1278 25784 1920 25836
rect 920 25712 1920 25784
rect 920 25660 978 25712
rect 1030 25660 1102 25712
rect 1154 25660 1226 25712
rect 1278 25660 1920 25712
rect 920 25590 1920 25660
rect 2836 28598 3729 28634
rect 3781 28598 3836 28645
rect 4356 28691 7272 28702
rect 4356 28645 4367 28691
rect 7261 28645 7272 28691
rect 4356 28634 6335 28645
rect 2836 28542 3836 28598
rect 2836 28490 3729 28542
rect 3781 28490 3836 28542
rect 2836 28434 3836 28490
rect 2836 28382 3729 28434
rect 3781 28382 3836 28434
rect 2836 28326 3836 28382
rect 2836 28274 3729 28326
rect 3781 28274 3836 28326
rect 2836 28218 3836 28274
rect 2836 28166 3729 28218
rect 3781 28166 3836 28218
rect 2836 28110 3836 28166
rect 2836 28058 3729 28110
rect 3781 28058 3836 28110
rect 2836 28002 3836 28058
rect 2836 27950 3729 28002
rect 3781 27950 3836 28002
rect 2836 27894 3836 27950
rect 2836 27842 3729 27894
rect 3781 27842 3836 27894
rect 2836 27786 3836 27842
rect 2836 27734 3729 27786
rect 3781 27734 3836 27786
rect 2836 27678 3836 27734
rect 2836 27626 3729 27678
rect 3781 27626 3836 27678
rect 2836 27570 3836 27626
rect 2836 27518 3729 27570
rect 3781 27518 3836 27570
rect 2836 27462 3836 27518
rect 2836 27410 3729 27462
rect 3781 27410 3836 27462
rect 2836 27354 3836 27410
rect 2836 27302 3729 27354
rect 3781 27302 3836 27354
rect 2836 27246 3836 27302
rect 2836 27194 3729 27246
rect 3781 27194 3836 27246
rect 2836 27138 3836 27194
rect 2836 27086 3729 27138
rect 3781 27086 3836 27138
rect 2836 27030 3836 27086
rect 2836 26978 3729 27030
rect 3781 26978 3836 27030
rect 2836 26922 3836 26978
rect 2836 26870 3729 26922
rect 3781 26870 3836 26922
rect 2836 26814 3836 26870
rect 2836 26762 3729 26814
rect 3781 26762 3836 26814
rect 2836 26706 3836 26762
rect 2836 26654 3729 26706
rect 3781 26654 3836 26706
rect 2836 26598 3836 26654
rect 2836 26546 3729 26598
rect 3781 26546 3836 26598
rect 2836 26490 3836 26546
rect 2836 26438 3729 26490
rect 3781 26438 3836 26490
rect 2836 26382 3836 26438
rect 2836 26330 3729 26382
rect 3781 26330 3836 26382
rect 2836 26274 3836 26330
rect 2836 26222 3729 26274
rect 3781 26222 3836 26274
rect 2836 26166 3836 26222
rect 2836 26114 3729 26166
rect 3781 26114 3836 26166
rect 2836 26058 3836 26114
rect 2836 26006 3729 26058
rect 3781 26006 3836 26058
rect 2836 25950 3836 26006
rect 2836 25898 3729 25950
rect 3781 25898 3836 25950
rect 2836 25842 3836 25898
rect 2836 25790 3729 25842
rect 3781 25790 3836 25842
rect 2836 25734 3836 25790
rect 2836 25682 3729 25734
rect 3781 25682 3836 25734
rect 2836 25626 3836 25682
rect 2836 25590 3729 25626
rect 920 25588 3729 25590
rect 920 25579 978 25588
rect 1030 25579 1102 25588
rect 1154 25579 1226 25588
rect 1278 25579 3729 25588
rect 3781 25579 3836 25626
rect 920 25533 931 25579
rect 3825 25533 3836 25579
rect 920 25522 3836 25533
rect 3896 28575 4296 28612
rect 3896 25649 3907 28575
rect 3953 25649 4239 28575
rect 4285 25649 4296 28575
rect 3896 25462 4296 25649
rect 4356 25590 5356 28634
rect 6272 28598 6335 28634
rect 6387 28598 7272 28645
rect 7792 28691 10708 28702
rect 7792 28645 7803 28691
rect 10697 28645 10708 28691
rect 6272 28542 7272 28598
rect 6272 28490 6335 28542
rect 6387 28490 7272 28542
rect 6272 28434 7272 28490
rect 6272 28382 6335 28434
rect 6387 28382 7272 28434
rect 6272 28326 7272 28382
rect 6272 28274 6335 28326
rect 6387 28274 7272 28326
rect 6272 28218 7272 28274
rect 6272 28166 6335 28218
rect 6387 28166 7272 28218
rect 6272 28110 7272 28166
rect 6272 28058 6335 28110
rect 6387 28058 7272 28110
rect 6272 28002 7272 28058
rect 6272 27950 6335 28002
rect 6387 27950 7272 28002
rect 6272 27894 7272 27950
rect 6272 27842 6335 27894
rect 6387 27842 7272 27894
rect 6272 27786 7272 27842
rect 6272 27734 6335 27786
rect 6387 27734 7272 27786
rect 6272 27678 7272 27734
rect 6272 27626 6335 27678
rect 6387 27626 7272 27678
rect 6272 27570 7272 27626
rect 6272 27518 6335 27570
rect 6387 27518 7272 27570
rect 6272 27462 7272 27518
rect 6272 27410 6335 27462
rect 6387 27410 7272 27462
rect 6272 27354 7272 27410
rect 6272 27302 6335 27354
rect 6387 27302 7272 27354
rect 6272 27246 7272 27302
rect 6272 27194 6335 27246
rect 6387 27194 7272 27246
rect 6272 27138 7272 27194
rect 6272 27086 6335 27138
rect 6387 27086 7272 27138
rect 6272 27030 7272 27086
rect 6272 26978 6335 27030
rect 6387 26978 7272 27030
rect 6272 26922 7272 26978
rect 6272 26870 6335 26922
rect 6387 26870 7272 26922
rect 6272 26814 7272 26870
rect 6272 26762 6335 26814
rect 6387 26762 7272 26814
rect 6272 26706 7272 26762
rect 6272 26654 6335 26706
rect 6387 26654 7272 26706
rect 6272 26598 7272 26654
rect 6272 26546 6335 26598
rect 6387 26546 7272 26598
rect 6272 26490 7272 26546
rect 6272 26438 6335 26490
rect 6387 26438 7272 26490
rect 6272 26382 7272 26438
rect 6272 26330 6335 26382
rect 6387 26330 7272 26382
rect 6272 26274 7272 26330
rect 6272 26222 6335 26274
rect 6387 26222 7272 26274
rect 6272 26166 7272 26222
rect 6272 26114 6335 26166
rect 6387 26114 7272 26166
rect 6272 26058 7272 26114
rect 6272 26006 6335 26058
rect 6387 26006 7272 26058
rect 6272 25950 7272 26006
rect 6272 25898 6335 25950
rect 6387 25898 7272 25950
rect 6272 25842 7272 25898
rect 6272 25790 6335 25842
rect 6387 25790 7272 25842
rect 6272 25734 7272 25790
rect 6272 25682 6335 25734
rect 6387 25682 7272 25734
rect 6272 25626 7272 25682
rect 6272 25590 6335 25626
rect 4356 25579 6335 25590
rect 6387 25579 7272 25626
rect 4356 25533 4367 25579
rect 7261 25533 7272 25579
rect 4356 25522 7272 25533
rect 7332 28596 7732 28612
rect 7332 28575 7388 28596
rect 7332 25649 7343 28575
rect 7440 28544 7624 28596
rect 7676 28575 7732 28596
rect 7389 28488 7675 28544
rect 7440 28436 7624 28488
rect 7389 28380 7675 28436
rect 7440 28328 7624 28380
rect 7389 28272 7675 28328
rect 7440 28220 7624 28272
rect 7389 28164 7675 28220
rect 7440 28112 7624 28164
rect 7389 28056 7675 28112
rect 7440 28004 7624 28056
rect 7389 27948 7675 28004
rect 7440 27896 7624 27948
rect 7389 27840 7675 27896
rect 7440 27788 7624 27840
rect 7389 27732 7675 27788
rect 7440 27680 7624 27732
rect 7389 27624 7675 27680
rect 7440 27572 7624 27624
rect 7389 27516 7675 27572
rect 7440 27464 7624 27516
rect 7389 27408 7675 27464
rect 7440 27356 7624 27408
rect 7389 27300 7675 27356
rect 7440 27248 7624 27300
rect 7389 27192 7675 27248
rect 7440 27140 7624 27192
rect 7389 27084 7675 27140
rect 7440 27032 7624 27084
rect 7389 26976 7675 27032
rect 7440 26924 7624 26976
rect 7389 26868 7675 26924
rect 7440 26816 7624 26868
rect 7389 26760 7675 26816
rect 7440 26708 7624 26760
rect 7389 26652 7675 26708
rect 7440 26600 7624 26652
rect 7389 26544 7675 26600
rect 7440 26492 7624 26544
rect 7389 26436 7675 26492
rect 7440 26384 7624 26436
rect 7389 26328 7675 26384
rect 7440 26276 7624 26328
rect 7389 26220 7675 26276
rect 7440 26168 7624 26220
rect 7389 26112 7675 26168
rect 7440 26060 7624 26112
rect 7389 26004 7675 26060
rect 7440 25952 7624 26004
rect 7389 25896 7675 25952
rect 7440 25844 7624 25896
rect 7389 25788 7675 25844
rect 7440 25736 7624 25788
rect 7389 25680 7675 25736
rect 7332 25628 7388 25649
rect 7440 25628 7624 25680
rect 7721 25649 7732 28575
rect 7676 25628 7732 25649
rect 7332 25462 7732 25628
rect 7792 28598 8677 28645
rect 8729 28634 10708 28645
rect 8729 28598 8792 28634
rect 7792 28542 8792 28598
rect 7792 28490 8677 28542
rect 8729 28490 8792 28542
rect 7792 28434 8792 28490
rect 7792 28382 8677 28434
rect 8729 28382 8792 28434
rect 7792 28326 8792 28382
rect 7792 28274 8677 28326
rect 8729 28274 8792 28326
rect 7792 28218 8792 28274
rect 7792 28166 8677 28218
rect 8729 28166 8792 28218
rect 7792 28110 8792 28166
rect 7792 28058 8677 28110
rect 8729 28058 8792 28110
rect 7792 28002 8792 28058
rect 7792 27950 8677 28002
rect 8729 27950 8792 28002
rect 7792 27894 8792 27950
rect 7792 27842 8677 27894
rect 8729 27842 8792 27894
rect 7792 27786 8792 27842
rect 7792 27734 8677 27786
rect 8729 27734 8792 27786
rect 7792 27678 8792 27734
rect 7792 27626 8677 27678
rect 8729 27626 8792 27678
rect 7792 27570 8792 27626
rect 7792 27518 8677 27570
rect 8729 27518 8792 27570
rect 7792 27462 8792 27518
rect 7792 27410 8677 27462
rect 8729 27410 8792 27462
rect 7792 27354 8792 27410
rect 7792 27302 8677 27354
rect 8729 27302 8792 27354
rect 7792 27246 8792 27302
rect 7792 27194 8677 27246
rect 8729 27194 8792 27246
rect 7792 27138 8792 27194
rect 7792 27086 8677 27138
rect 8729 27086 8792 27138
rect 7792 27030 8792 27086
rect 7792 26978 8677 27030
rect 8729 26978 8792 27030
rect 7792 26922 8792 26978
rect 7792 26870 8677 26922
rect 8729 26870 8792 26922
rect 7792 26814 8792 26870
rect 7792 26762 8677 26814
rect 8729 26762 8792 26814
rect 7792 26706 8792 26762
rect 7792 26654 8677 26706
rect 8729 26654 8792 26706
rect 7792 26598 8792 26654
rect 7792 26546 8677 26598
rect 8729 26546 8792 26598
rect 7792 26490 8792 26546
rect 7792 26438 8677 26490
rect 8729 26438 8792 26490
rect 7792 26382 8792 26438
rect 7792 26330 8677 26382
rect 8729 26330 8792 26382
rect 7792 26274 8792 26330
rect 7792 26222 8677 26274
rect 8729 26222 8792 26274
rect 7792 26166 8792 26222
rect 7792 26114 8677 26166
rect 8729 26114 8792 26166
rect 7792 26058 8792 26114
rect 7792 26006 8677 26058
rect 8729 26006 8792 26058
rect 7792 25950 8792 26006
rect 7792 25898 8677 25950
rect 8729 25898 8792 25950
rect 7792 25842 8792 25898
rect 7792 25790 8677 25842
rect 8729 25790 8792 25842
rect 7792 25734 8792 25790
rect 7792 25682 8677 25734
rect 8729 25682 8792 25734
rect 7792 25626 8792 25682
rect 7792 25579 8677 25626
rect 8729 25590 8792 25626
rect 9708 25590 10708 28634
rect 11228 28691 14144 28702
rect 11228 28645 11239 28691
rect 14133 28645 14144 28691
rect 8729 25579 10708 25590
rect 7792 25533 7803 25579
rect 10697 25533 10708 25579
rect 7792 25522 10708 25533
rect 10768 28575 11168 28612
rect 10768 25649 10779 28575
rect 10825 25649 11111 28575
rect 11157 25649 11168 28575
rect 10768 25462 11168 25649
rect 11228 28598 11283 28645
rect 11335 28636 13786 28645
rect 13838 28636 13910 28645
rect 13962 28636 14034 28645
rect 14086 28636 14144 28645
rect 11335 28634 14144 28636
rect 11335 28598 12228 28634
rect 11228 28542 12228 28598
rect 11228 28490 11283 28542
rect 11335 28490 12228 28542
rect 11228 28434 12228 28490
rect 11228 28382 11283 28434
rect 11335 28382 12228 28434
rect 11228 28326 12228 28382
rect 11228 28274 11283 28326
rect 11335 28274 12228 28326
rect 11228 28218 12228 28274
rect 11228 28166 11283 28218
rect 11335 28166 12228 28218
rect 11228 28110 12228 28166
rect 11228 28058 11283 28110
rect 11335 28058 12228 28110
rect 11228 28002 12228 28058
rect 11228 27950 11283 28002
rect 11335 27950 12228 28002
rect 11228 27894 12228 27950
rect 11228 27842 11283 27894
rect 11335 27842 12228 27894
rect 11228 27786 12228 27842
rect 11228 27734 11283 27786
rect 11335 27734 12228 27786
rect 11228 27678 12228 27734
rect 11228 27626 11283 27678
rect 11335 27626 12228 27678
rect 11228 27570 12228 27626
rect 11228 27518 11283 27570
rect 11335 27518 12228 27570
rect 11228 27462 12228 27518
rect 11228 27410 11283 27462
rect 11335 27410 12228 27462
rect 11228 27354 12228 27410
rect 11228 27302 11283 27354
rect 11335 27302 12228 27354
rect 11228 27246 12228 27302
rect 11228 27194 11283 27246
rect 11335 27194 12228 27246
rect 11228 27138 12228 27194
rect 11228 27086 11283 27138
rect 11335 27086 12228 27138
rect 11228 27030 12228 27086
rect 11228 26978 11283 27030
rect 11335 26978 12228 27030
rect 11228 26922 12228 26978
rect 11228 26870 11283 26922
rect 11335 26870 12228 26922
rect 11228 26814 12228 26870
rect 11228 26762 11283 26814
rect 11335 26762 12228 26814
rect 11228 26706 12228 26762
rect 11228 26654 11283 26706
rect 11335 26654 12228 26706
rect 11228 26598 12228 26654
rect 11228 26546 11283 26598
rect 11335 26546 12228 26598
rect 11228 26490 12228 26546
rect 11228 26438 11283 26490
rect 11335 26438 12228 26490
rect 11228 26382 12228 26438
rect 11228 26330 11283 26382
rect 11335 26330 12228 26382
rect 11228 26274 12228 26330
rect 11228 26222 11283 26274
rect 11335 26222 12228 26274
rect 11228 26166 12228 26222
rect 11228 26114 11283 26166
rect 11335 26114 12228 26166
rect 11228 26058 12228 26114
rect 11228 26006 11283 26058
rect 11335 26006 12228 26058
rect 11228 25950 12228 26006
rect 11228 25898 11283 25950
rect 11335 25898 12228 25950
rect 11228 25842 12228 25898
rect 11228 25790 11283 25842
rect 11335 25790 12228 25842
rect 11228 25734 12228 25790
rect 11228 25682 11283 25734
rect 11335 25682 12228 25734
rect 11228 25626 12228 25682
rect 11228 25579 11283 25626
rect 11335 25590 12228 25626
rect 13144 28564 14144 28634
rect 13144 28512 13786 28564
rect 13838 28512 13910 28564
rect 13962 28512 14034 28564
rect 14086 28512 14144 28564
rect 13144 28440 14144 28512
rect 13144 28388 13786 28440
rect 13838 28388 13910 28440
rect 13962 28388 14034 28440
rect 14086 28388 14144 28440
rect 13144 28316 14144 28388
rect 13144 28264 13786 28316
rect 13838 28264 13910 28316
rect 13962 28264 14034 28316
rect 14086 28264 14144 28316
rect 13144 28192 14144 28264
rect 13144 28140 13786 28192
rect 13838 28140 13910 28192
rect 13962 28140 14034 28192
rect 14086 28140 14144 28192
rect 13144 28068 14144 28140
rect 13144 28016 13786 28068
rect 13838 28016 13910 28068
rect 13962 28016 14034 28068
rect 14086 28016 14144 28068
rect 13144 27944 14144 28016
rect 13144 27892 13786 27944
rect 13838 27892 13910 27944
rect 13962 27892 14034 27944
rect 14086 27892 14144 27944
rect 13144 27820 14144 27892
rect 13144 27768 13786 27820
rect 13838 27768 13910 27820
rect 13962 27768 14034 27820
rect 14086 27768 14144 27820
rect 13144 27696 14144 27768
rect 13144 27644 13786 27696
rect 13838 27644 13910 27696
rect 13962 27644 14034 27696
rect 14086 27644 14144 27696
rect 13144 27572 14144 27644
rect 13144 27520 13786 27572
rect 13838 27520 13910 27572
rect 13962 27520 14034 27572
rect 14086 27520 14144 27572
rect 13144 27448 14144 27520
rect 13144 27396 13786 27448
rect 13838 27396 13910 27448
rect 13962 27396 14034 27448
rect 14086 27396 14144 27448
rect 13144 27324 14144 27396
rect 13144 27272 13786 27324
rect 13838 27272 13910 27324
rect 13962 27272 14034 27324
rect 14086 27272 14144 27324
rect 13144 27200 14144 27272
rect 13144 27148 13786 27200
rect 13838 27148 13910 27200
rect 13962 27148 14034 27200
rect 14086 27148 14144 27200
rect 13144 27076 14144 27148
rect 13144 27024 13786 27076
rect 13838 27024 13910 27076
rect 13962 27024 14034 27076
rect 14086 27024 14144 27076
rect 13144 26952 14144 27024
rect 13144 26900 13786 26952
rect 13838 26900 13910 26952
rect 13962 26900 14034 26952
rect 14086 26900 14144 26952
rect 13144 26828 14144 26900
rect 13144 26776 13786 26828
rect 13838 26776 13910 26828
rect 13962 26776 14034 26828
rect 14086 26776 14144 26828
rect 13144 26704 14144 26776
rect 13144 26652 13786 26704
rect 13838 26652 13910 26704
rect 13962 26652 14034 26704
rect 14086 26652 14144 26704
rect 13144 26580 14144 26652
rect 13144 26528 13786 26580
rect 13838 26528 13910 26580
rect 13962 26528 14034 26580
rect 14086 26528 14144 26580
rect 13144 26456 14144 26528
rect 13144 26404 13786 26456
rect 13838 26404 13910 26456
rect 13962 26404 14034 26456
rect 14086 26404 14144 26456
rect 13144 26332 14144 26404
rect 13144 26280 13786 26332
rect 13838 26280 13910 26332
rect 13962 26280 14034 26332
rect 14086 26280 14144 26332
rect 13144 26208 14144 26280
rect 13144 26156 13786 26208
rect 13838 26156 13910 26208
rect 13962 26156 14034 26208
rect 14086 26156 14144 26208
rect 13144 26084 14144 26156
rect 13144 26032 13786 26084
rect 13838 26032 13910 26084
rect 13962 26032 14034 26084
rect 14086 26032 14144 26084
rect 13144 25960 14144 26032
rect 13144 25908 13786 25960
rect 13838 25908 13910 25960
rect 13962 25908 14034 25960
rect 14086 25908 14144 25960
rect 13144 25836 14144 25908
rect 13144 25784 13786 25836
rect 13838 25784 13910 25836
rect 13962 25784 14034 25836
rect 14086 25784 14144 25836
rect 13144 25712 14144 25784
rect 13144 25660 13786 25712
rect 13838 25660 13910 25712
rect 13962 25660 14034 25712
rect 14086 25660 14144 25712
rect 13144 25590 14144 25660
rect 11335 25588 14144 25590
rect 11335 25579 13786 25588
rect 13838 25579 13910 25588
rect 13962 25579 14034 25588
rect 14086 25579 14144 25588
rect 11228 25533 11239 25579
rect 14133 25533 14144 25579
rect 11228 25522 14144 25533
rect 14204 28575 14404 28612
rect 14204 25649 14215 28575
rect 14261 25649 14404 28575
rect 14204 25462 14404 25649
rect 14608 25462 14619 28762
rect 445 25412 14619 25462
rect 445 25380 1438 25412
rect 496 25328 552 25380
rect 604 25328 660 25380
rect 712 25360 1438 25380
rect 1490 25360 1562 25412
rect 1614 25360 1686 25412
rect 1738 25360 1810 25412
rect 1862 25360 2574 25412
rect 2626 25360 2698 25412
rect 2750 25360 2822 25412
rect 2874 25360 2946 25412
rect 2998 25360 4846 25412
rect 4898 25360 4970 25412
rect 5022 25360 5094 25412
rect 5146 25360 5218 25412
rect 5270 25360 7139 25412
rect 7191 25360 7263 25412
rect 7315 25360 7387 25412
rect 7439 25360 7625 25412
rect 7677 25360 7749 25412
rect 7801 25360 7873 25412
rect 7925 25360 9794 25412
rect 9846 25360 9918 25412
rect 9970 25360 10042 25412
rect 10094 25360 10166 25412
rect 10218 25360 12066 25412
rect 12118 25360 12190 25412
rect 12242 25360 12314 25412
rect 12366 25360 12438 25412
rect 12490 25360 13202 25412
rect 13254 25360 13326 25412
rect 13378 25360 13450 25412
rect 13502 25360 13574 25412
rect 13626 25380 14619 25412
rect 13626 25360 14352 25380
rect 712 25328 14352 25360
rect 14404 25328 14460 25380
rect 14512 25328 14568 25380
rect 445 25288 14619 25328
rect 445 25272 1438 25288
rect 496 25220 552 25272
rect 604 25220 660 25272
rect 712 25236 1438 25272
rect 1490 25236 1562 25288
rect 1614 25236 1686 25288
rect 1738 25236 1810 25288
rect 1862 25236 2574 25288
rect 2626 25236 2698 25288
rect 2750 25236 2822 25288
rect 2874 25236 2946 25288
rect 2998 25236 4846 25288
rect 4898 25236 4970 25288
rect 5022 25236 5094 25288
rect 5146 25236 5218 25288
rect 5270 25236 7139 25288
rect 7191 25236 7263 25288
rect 7315 25236 7387 25288
rect 7439 25236 7625 25288
rect 7677 25236 7749 25288
rect 7801 25236 7873 25288
rect 7925 25236 9794 25288
rect 9846 25236 9918 25288
rect 9970 25236 10042 25288
rect 10094 25236 10166 25288
rect 10218 25236 12066 25288
rect 12118 25236 12190 25288
rect 12242 25236 12314 25288
rect 12366 25236 12438 25288
rect 12490 25236 13202 25288
rect 13254 25236 13326 25288
rect 13378 25236 13450 25288
rect 13502 25236 13574 25288
rect 13626 25272 14619 25288
rect 13626 25236 14352 25272
rect 712 25220 14352 25236
rect 14404 25220 14460 25272
rect 14512 25220 14568 25272
rect 445 25164 14619 25220
rect 496 25112 552 25164
rect 604 25161 660 25164
rect 712 25161 1438 25164
rect 1490 25161 1562 25164
rect 1614 25161 1686 25164
rect 1738 25161 1810 25164
rect 1862 25161 2574 25164
rect 2626 25161 2698 25164
rect 2750 25161 2822 25164
rect 2874 25161 2946 25164
rect 2998 25161 4846 25164
rect 4898 25161 4970 25164
rect 5022 25161 5094 25164
rect 5146 25161 5218 25164
rect 5270 25161 7139 25164
rect 7191 25161 7263 25164
rect 7315 25161 7387 25164
rect 7439 25161 7625 25164
rect 7677 25161 7749 25164
rect 7801 25161 7873 25164
rect 7925 25161 9794 25164
rect 9846 25161 9918 25164
rect 9970 25161 10042 25164
rect 10094 25161 10166 25164
rect 10218 25161 12066 25164
rect 12118 25161 12190 25164
rect 12242 25161 12314 25164
rect 12366 25161 12438 25164
rect 12490 25161 13202 25164
rect 13254 25161 13326 25164
rect 13378 25161 13450 25164
rect 13502 25161 13574 25164
rect 13626 25161 14352 25164
rect 14404 25161 14460 25164
rect 604 25112 660 25115
rect 712 25112 1438 25115
rect 1490 25112 1562 25115
rect 1614 25112 1686 25115
rect 1738 25112 1810 25115
rect 1862 25112 2574 25115
rect 2626 25112 2698 25115
rect 2750 25112 2822 25115
rect 2874 25112 2946 25115
rect 2998 25112 4846 25115
rect 4898 25112 4970 25115
rect 5022 25112 5094 25115
rect 5146 25112 5218 25115
rect 5270 25112 7139 25115
rect 7191 25112 7263 25115
rect 7315 25112 7387 25115
rect 7439 25112 7625 25115
rect 7677 25112 7749 25115
rect 7801 25112 7873 25115
rect 7925 25112 9794 25115
rect 9846 25112 9918 25115
rect 9970 25112 10042 25115
rect 10094 25112 10166 25115
rect 10218 25112 12066 25115
rect 12118 25112 12190 25115
rect 12242 25112 12314 25115
rect 12366 25112 12438 25115
rect 12490 25112 13202 25115
rect 13254 25112 13326 25115
rect 13378 25112 13450 25115
rect 13502 25112 13574 25115
rect 13626 25112 14352 25115
rect 14404 25112 14460 25115
rect 14512 25112 14568 25164
rect 445 25056 14619 25112
rect 496 25004 552 25056
rect 604 25004 660 25056
rect 712 25040 14352 25056
rect 712 25004 1438 25040
rect 445 24988 1438 25004
rect 1490 24988 1562 25040
rect 1614 24988 1686 25040
rect 1738 24988 1810 25040
rect 1862 24988 2574 25040
rect 2626 24988 2698 25040
rect 2750 24988 2822 25040
rect 2874 24988 2946 25040
rect 2998 24988 4846 25040
rect 4898 24988 4970 25040
rect 5022 24988 5094 25040
rect 5146 24988 5218 25040
rect 5270 24988 7139 25040
rect 7191 24988 7263 25040
rect 7315 24988 7387 25040
rect 7439 24988 7625 25040
rect 7677 24988 7749 25040
rect 7801 24988 7873 25040
rect 7925 24988 9794 25040
rect 9846 24988 9918 25040
rect 9970 24988 10042 25040
rect 10094 24988 10166 25040
rect 10218 24988 12066 25040
rect 12118 24988 12190 25040
rect 12242 24988 12314 25040
rect 12366 24988 12438 25040
rect 12490 24988 13202 25040
rect 13254 24988 13326 25040
rect 13378 24988 13450 25040
rect 13502 24988 13574 25040
rect 13626 25004 14352 25040
rect 14404 25004 14460 25056
rect 14512 25004 14568 25056
rect 13626 24988 14619 25004
rect 445 24948 14619 24988
rect 496 24896 552 24948
rect 604 24896 660 24948
rect 712 24916 14352 24948
rect 712 24896 1438 24916
rect 445 24864 1438 24896
rect 1490 24864 1562 24916
rect 1614 24864 1686 24916
rect 1738 24864 1810 24916
rect 1862 24864 2574 24916
rect 2626 24864 2698 24916
rect 2750 24864 2822 24916
rect 2874 24864 2946 24916
rect 2998 24864 4846 24916
rect 4898 24864 4970 24916
rect 5022 24864 5094 24916
rect 5146 24864 5218 24916
rect 5270 24864 7139 24916
rect 7191 24864 7263 24916
rect 7315 24864 7387 24916
rect 7439 24864 7625 24916
rect 7677 24864 7749 24916
rect 7801 24864 7873 24916
rect 7925 24864 9794 24916
rect 9846 24864 9918 24916
rect 9970 24864 10042 24916
rect 10094 24864 10166 24916
rect 10218 24864 12066 24916
rect 12118 24864 12190 24916
rect 12242 24864 12314 24916
rect 12366 24864 12438 24916
rect 12490 24864 13202 24916
rect 13254 24864 13326 24916
rect 13378 24864 13450 24916
rect 13502 24864 13574 24916
rect 13626 24896 14352 24916
rect 14404 24896 14460 24948
rect 14512 24896 14568 24948
rect 13626 24864 14619 24896
rect 445 24814 14619 24864
rect 445 21514 456 24814
rect 920 24743 3836 24754
rect 920 24697 931 24743
rect 3825 24697 3836 24743
rect 920 24688 978 24697
rect 1030 24688 1102 24697
rect 1154 24688 1226 24697
rect 1278 24688 3729 24697
rect 920 24686 3729 24688
rect 660 24627 860 24664
rect 660 21701 803 24627
rect 849 21701 860 24627
rect 660 21514 860 21701
rect 920 24616 1920 24686
rect 920 24564 978 24616
rect 1030 24564 1102 24616
rect 1154 24564 1226 24616
rect 1278 24564 1920 24616
rect 920 24492 1920 24564
rect 920 24440 978 24492
rect 1030 24440 1102 24492
rect 1154 24440 1226 24492
rect 1278 24440 1920 24492
rect 920 24368 1920 24440
rect 920 24316 978 24368
rect 1030 24316 1102 24368
rect 1154 24316 1226 24368
rect 1278 24316 1920 24368
rect 920 24244 1920 24316
rect 920 24192 978 24244
rect 1030 24192 1102 24244
rect 1154 24192 1226 24244
rect 1278 24192 1920 24244
rect 920 24120 1920 24192
rect 920 24068 978 24120
rect 1030 24068 1102 24120
rect 1154 24068 1226 24120
rect 1278 24068 1920 24120
rect 920 23996 1920 24068
rect 920 23944 978 23996
rect 1030 23944 1102 23996
rect 1154 23944 1226 23996
rect 1278 23944 1920 23996
rect 920 23872 1920 23944
rect 920 23820 978 23872
rect 1030 23820 1102 23872
rect 1154 23820 1226 23872
rect 1278 23820 1920 23872
rect 920 23748 1920 23820
rect 920 23696 978 23748
rect 1030 23696 1102 23748
rect 1154 23696 1226 23748
rect 1278 23696 1920 23748
rect 920 23624 1920 23696
rect 920 23572 978 23624
rect 1030 23572 1102 23624
rect 1154 23572 1226 23624
rect 1278 23572 1920 23624
rect 920 23500 1920 23572
rect 920 23448 978 23500
rect 1030 23448 1102 23500
rect 1154 23448 1226 23500
rect 1278 23448 1920 23500
rect 920 23376 1920 23448
rect 920 23324 978 23376
rect 1030 23324 1102 23376
rect 1154 23324 1226 23376
rect 1278 23324 1920 23376
rect 920 23252 1920 23324
rect 920 23200 978 23252
rect 1030 23200 1102 23252
rect 1154 23200 1226 23252
rect 1278 23200 1920 23252
rect 920 23128 1920 23200
rect 920 23076 978 23128
rect 1030 23076 1102 23128
rect 1154 23076 1226 23128
rect 1278 23076 1920 23128
rect 920 23004 1920 23076
rect 920 22952 978 23004
rect 1030 22952 1102 23004
rect 1154 22952 1226 23004
rect 1278 22952 1920 23004
rect 920 22880 1920 22952
rect 920 22828 978 22880
rect 1030 22828 1102 22880
rect 1154 22828 1226 22880
rect 1278 22828 1920 22880
rect 920 22756 1920 22828
rect 920 22704 978 22756
rect 1030 22704 1102 22756
rect 1154 22704 1226 22756
rect 1278 22704 1920 22756
rect 920 22632 1920 22704
rect 920 22580 978 22632
rect 1030 22580 1102 22632
rect 1154 22580 1226 22632
rect 1278 22580 1920 22632
rect 920 22508 1920 22580
rect 920 22456 978 22508
rect 1030 22456 1102 22508
rect 1154 22456 1226 22508
rect 1278 22456 1920 22508
rect 920 22384 1920 22456
rect 920 22332 978 22384
rect 1030 22332 1102 22384
rect 1154 22332 1226 22384
rect 1278 22332 1920 22384
rect 920 22260 1920 22332
rect 920 22208 978 22260
rect 1030 22208 1102 22260
rect 1154 22208 1226 22260
rect 1278 22208 1920 22260
rect 920 22136 1920 22208
rect 920 22084 978 22136
rect 1030 22084 1102 22136
rect 1154 22084 1226 22136
rect 1278 22084 1920 22136
rect 920 22012 1920 22084
rect 920 21960 978 22012
rect 1030 21960 1102 22012
rect 1154 21960 1226 22012
rect 1278 21960 1920 22012
rect 920 21888 1920 21960
rect 920 21836 978 21888
rect 1030 21836 1102 21888
rect 1154 21836 1226 21888
rect 1278 21836 1920 21888
rect 920 21764 1920 21836
rect 920 21712 978 21764
rect 1030 21712 1102 21764
rect 1154 21712 1226 21764
rect 1278 21712 1920 21764
rect 920 21642 1920 21712
rect 2836 24650 3729 24686
rect 3781 24650 3836 24697
rect 4356 24743 7272 24754
rect 4356 24697 4367 24743
rect 7261 24697 7272 24743
rect 4356 24686 6335 24697
rect 2836 24594 3836 24650
rect 2836 24542 3729 24594
rect 3781 24542 3836 24594
rect 2836 24486 3836 24542
rect 2836 24434 3729 24486
rect 3781 24434 3836 24486
rect 2836 24378 3836 24434
rect 2836 24326 3729 24378
rect 3781 24326 3836 24378
rect 2836 24270 3836 24326
rect 2836 24218 3729 24270
rect 3781 24218 3836 24270
rect 2836 24162 3836 24218
rect 2836 24110 3729 24162
rect 3781 24110 3836 24162
rect 2836 24054 3836 24110
rect 2836 24002 3729 24054
rect 3781 24002 3836 24054
rect 2836 23946 3836 24002
rect 2836 23894 3729 23946
rect 3781 23894 3836 23946
rect 2836 23838 3836 23894
rect 2836 23786 3729 23838
rect 3781 23786 3836 23838
rect 2836 23730 3836 23786
rect 2836 23678 3729 23730
rect 3781 23678 3836 23730
rect 2836 23622 3836 23678
rect 2836 23570 3729 23622
rect 3781 23570 3836 23622
rect 2836 23514 3836 23570
rect 2836 23462 3729 23514
rect 3781 23462 3836 23514
rect 2836 23406 3836 23462
rect 2836 23354 3729 23406
rect 3781 23354 3836 23406
rect 2836 23298 3836 23354
rect 2836 23246 3729 23298
rect 3781 23246 3836 23298
rect 2836 23190 3836 23246
rect 2836 23138 3729 23190
rect 3781 23138 3836 23190
rect 2836 23082 3836 23138
rect 2836 23030 3729 23082
rect 3781 23030 3836 23082
rect 2836 22974 3836 23030
rect 2836 22922 3729 22974
rect 3781 22922 3836 22974
rect 2836 22866 3836 22922
rect 2836 22814 3729 22866
rect 3781 22814 3836 22866
rect 2836 22758 3836 22814
rect 2836 22706 3729 22758
rect 3781 22706 3836 22758
rect 2836 22650 3836 22706
rect 2836 22598 3729 22650
rect 3781 22598 3836 22650
rect 2836 22542 3836 22598
rect 2836 22490 3729 22542
rect 3781 22490 3836 22542
rect 2836 22434 3836 22490
rect 2836 22382 3729 22434
rect 3781 22382 3836 22434
rect 2836 22326 3836 22382
rect 2836 22274 3729 22326
rect 3781 22274 3836 22326
rect 2836 22218 3836 22274
rect 2836 22166 3729 22218
rect 3781 22166 3836 22218
rect 2836 22110 3836 22166
rect 2836 22058 3729 22110
rect 3781 22058 3836 22110
rect 2836 22002 3836 22058
rect 2836 21950 3729 22002
rect 3781 21950 3836 22002
rect 2836 21894 3836 21950
rect 2836 21842 3729 21894
rect 3781 21842 3836 21894
rect 2836 21786 3836 21842
rect 2836 21734 3729 21786
rect 3781 21734 3836 21786
rect 2836 21678 3836 21734
rect 2836 21642 3729 21678
rect 920 21640 3729 21642
rect 920 21631 978 21640
rect 1030 21631 1102 21640
rect 1154 21631 1226 21640
rect 1278 21631 3729 21640
rect 3781 21631 3836 21678
rect 920 21585 931 21631
rect 3825 21585 3836 21631
rect 920 21574 3836 21585
rect 3896 24627 4296 24664
rect 3896 21701 3907 24627
rect 3953 21701 4239 24627
rect 4285 21701 4296 24627
rect 3896 21514 4296 21701
rect 4356 21642 5356 24686
rect 6272 24650 6335 24686
rect 6387 24650 7272 24697
rect 7792 24743 10708 24754
rect 7792 24697 7803 24743
rect 10697 24697 10708 24743
rect 6272 24594 7272 24650
rect 6272 24542 6335 24594
rect 6387 24542 7272 24594
rect 6272 24486 7272 24542
rect 6272 24434 6335 24486
rect 6387 24434 7272 24486
rect 6272 24378 7272 24434
rect 6272 24326 6335 24378
rect 6387 24326 7272 24378
rect 6272 24270 7272 24326
rect 6272 24218 6335 24270
rect 6387 24218 7272 24270
rect 6272 24162 7272 24218
rect 6272 24110 6335 24162
rect 6387 24110 7272 24162
rect 6272 24054 7272 24110
rect 6272 24002 6335 24054
rect 6387 24002 7272 24054
rect 6272 23946 7272 24002
rect 6272 23894 6335 23946
rect 6387 23894 7272 23946
rect 6272 23838 7272 23894
rect 6272 23786 6335 23838
rect 6387 23786 7272 23838
rect 6272 23730 7272 23786
rect 6272 23678 6335 23730
rect 6387 23678 7272 23730
rect 6272 23622 7272 23678
rect 6272 23570 6335 23622
rect 6387 23570 7272 23622
rect 6272 23514 7272 23570
rect 6272 23462 6335 23514
rect 6387 23462 7272 23514
rect 6272 23406 7272 23462
rect 6272 23354 6335 23406
rect 6387 23354 7272 23406
rect 6272 23298 7272 23354
rect 6272 23246 6335 23298
rect 6387 23246 7272 23298
rect 6272 23190 7272 23246
rect 6272 23138 6335 23190
rect 6387 23138 7272 23190
rect 6272 23082 7272 23138
rect 6272 23030 6335 23082
rect 6387 23030 7272 23082
rect 6272 22974 7272 23030
rect 6272 22922 6335 22974
rect 6387 22922 7272 22974
rect 6272 22866 7272 22922
rect 6272 22814 6335 22866
rect 6387 22814 7272 22866
rect 6272 22758 7272 22814
rect 6272 22706 6335 22758
rect 6387 22706 7272 22758
rect 6272 22650 7272 22706
rect 6272 22598 6335 22650
rect 6387 22598 7272 22650
rect 6272 22542 7272 22598
rect 6272 22490 6335 22542
rect 6387 22490 7272 22542
rect 6272 22434 7272 22490
rect 6272 22382 6335 22434
rect 6387 22382 7272 22434
rect 6272 22326 7272 22382
rect 6272 22274 6335 22326
rect 6387 22274 7272 22326
rect 6272 22218 7272 22274
rect 6272 22166 6335 22218
rect 6387 22166 7272 22218
rect 6272 22110 7272 22166
rect 6272 22058 6335 22110
rect 6387 22058 7272 22110
rect 6272 22002 7272 22058
rect 6272 21950 6335 22002
rect 6387 21950 7272 22002
rect 6272 21894 7272 21950
rect 6272 21842 6335 21894
rect 6387 21842 7272 21894
rect 6272 21786 7272 21842
rect 6272 21734 6335 21786
rect 6387 21734 7272 21786
rect 6272 21678 7272 21734
rect 6272 21642 6335 21678
rect 4356 21631 6335 21642
rect 6387 21631 7272 21678
rect 4356 21585 4367 21631
rect 7261 21585 7272 21631
rect 4356 21574 7272 21585
rect 7332 24648 7732 24664
rect 7332 24627 7388 24648
rect 7332 21701 7343 24627
rect 7440 24596 7624 24648
rect 7676 24627 7732 24648
rect 7389 24540 7675 24596
rect 7440 24488 7624 24540
rect 7389 24432 7675 24488
rect 7440 24380 7624 24432
rect 7389 24324 7675 24380
rect 7440 24272 7624 24324
rect 7389 24216 7675 24272
rect 7440 24164 7624 24216
rect 7389 24108 7675 24164
rect 7440 24056 7624 24108
rect 7389 24000 7675 24056
rect 7440 23948 7624 24000
rect 7389 23892 7675 23948
rect 7440 23840 7624 23892
rect 7389 23784 7675 23840
rect 7440 23732 7624 23784
rect 7389 23676 7675 23732
rect 7440 23624 7624 23676
rect 7389 23568 7675 23624
rect 7440 23516 7624 23568
rect 7389 23460 7675 23516
rect 7440 23408 7624 23460
rect 7389 23352 7675 23408
rect 7440 23300 7624 23352
rect 7389 23244 7675 23300
rect 7440 23192 7624 23244
rect 7389 23136 7675 23192
rect 7440 23084 7624 23136
rect 7389 23028 7675 23084
rect 7440 22976 7624 23028
rect 7389 22920 7675 22976
rect 7440 22868 7624 22920
rect 7389 22812 7675 22868
rect 7440 22760 7624 22812
rect 7389 22704 7675 22760
rect 7440 22652 7624 22704
rect 7389 22596 7675 22652
rect 7440 22544 7624 22596
rect 7389 22488 7675 22544
rect 7440 22436 7624 22488
rect 7389 22380 7675 22436
rect 7440 22328 7624 22380
rect 7389 22272 7675 22328
rect 7440 22220 7624 22272
rect 7389 22164 7675 22220
rect 7440 22112 7624 22164
rect 7389 22056 7675 22112
rect 7440 22004 7624 22056
rect 7389 21948 7675 22004
rect 7440 21896 7624 21948
rect 7389 21840 7675 21896
rect 7440 21788 7624 21840
rect 7389 21732 7675 21788
rect 7332 21680 7388 21701
rect 7440 21680 7624 21732
rect 7721 21701 7732 24627
rect 7676 21680 7732 21701
rect 7332 21514 7732 21680
rect 7792 24650 8677 24697
rect 8729 24686 10708 24697
rect 8729 24650 8792 24686
rect 7792 24594 8792 24650
rect 7792 24542 8677 24594
rect 8729 24542 8792 24594
rect 7792 24486 8792 24542
rect 7792 24434 8677 24486
rect 8729 24434 8792 24486
rect 7792 24378 8792 24434
rect 7792 24326 8677 24378
rect 8729 24326 8792 24378
rect 7792 24270 8792 24326
rect 7792 24218 8677 24270
rect 8729 24218 8792 24270
rect 7792 24162 8792 24218
rect 7792 24110 8677 24162
rect 8729 24110 8792 24162
rect 7792 24054 8792 24110
rect 7792 24002 8677 24054
rect 8729 24002 8792 24054
rect 7792 23946 8792 24002
rect 7792 23894 8677 23946
rect 8729 23894 8792 23946
rect 7792 23838 8792 23894
rect 7792 23786 8677 23838
rect 8729 23786 8792 23838
rect 7792 23730 8792 23786
rect 7792 23678 8677 23730
rect 8729 23678 8792 23730
rect 7792 23622 8792 23678
rect 7792 23570 8677 23622
rect 8729 23570 8792 23622
rect 7792 23514 8792 23570
rect 7792 23462 8677 23514
rect 8729 23462 8792 23514
rect 7792 23406 8792 23462
rect 7792 23354 8677 23406
rect 8729 23354 8792 23406
rect 7792 23298 8792 23354
rect 7792 23246 8677 23298
rect 8729 23246 8792 23298
rect 7792 23190 8792 23246
rect 7792 23138 8677 23190
rect 8729 23138 8792 23190
rect 7792 23082 8792 23138
rect 7792 23030 8677 23082
rect 8729 23030 8792 23082
rect 7792 22974 8792 23030
rect 7792 22922 8677 22974
rect 8729 22922 8792 22974
rect 7792 22866 8792 22922
rect 7792 22814 8677 22866
rect 8729 22814 8792 22866
rect 7792 22758 8792 22814
rect 7792 22706 8677 22758
rect 8729 22706 8792 22758
rect 7792 22650 8792 22706
rect 7792 22598 8677 22650
rect 8729 22598 8792 22650
rect 7792 22542 8792 22598
rect 7792 22490 8677 22542
rect 8729 22490 8792 22542
rect 7792 22434 8792 22490
rect 7792 22382 8677 22434
rect 8729 22382 8792 22434
rect 7792 22326 8792 22382
rect 7792 22274 8677 22326
rect 8729 22274 8792 22326
rect 7792 22218 8792 22274
rect 7792 22166 8677 22218
rect 8729 22166 8792 22218
rect 7792 22110 8792 22166
rect 7792 22058 8677 22110
rect 8729 22058 8792 22110
rect 7792 22002 8792 22058
rect 7792 21950 8677 22002
rect 8729 21950 8792 22002
rect 7792 21894 8792 21950
rect 7792 21842 8677 21894
rect 8729 21842 8792 21894
rect 7792 21786 8792 21842
rect 7792 21734 8677 21786
rect 8729 21734 8792 21786
rect 7792 21678 8792 21734
rect 7792 21631 8677 21678
rect 8729 21642 8792 21678
rect 9708 21642 10708 24686
rect 11228 24743 14144 24754
rect 11228 24697 11239 24743
rect 14133 24697 14144 24743
rect 8729 21631 10708 21642
rect 7792 21585 7803 21631
rect 10697 21585 10708 21631
rect 7792 21574 10708 21585
rect 10768 24627 11168 24664
rect 10768 21701 10779 24627
rect 10825 21701 11111 24627
rect 11157 21701 11168 24627
rect 10768 21514 11168 21701
rect 11228 24650 11283 24697
rect 11335 24688 13786 24697
rect 13838 24688 13910 24697
rect 13962 24688 14034 24697
rect 14086 24688 14144 24697
rect 11335 24686 14144 24688
rect 11335 24650 12228 24686
rect 11228 24594 12228 24650
rect 11228 24542 11283 24594
rect 11335 24542 12228 24594
rect 11228 24486 12228 24542
rect 11228 24434 11283 24486
rect 11335 24434 12228 24486
rect 11228 24378 12228 24434
rect 11228 24326 11283 24378
rect 11335 24326 12228 24378
rect 11228 24270 12228 24326
rect 11228 24218 11283 24270
rect 11335 24218 12228 24270
rect 11228 24162 12228 24218
rect 11228 24110 11283 24162
rect 11335 24110 12228 24162
rect 11228 24054 12228 24110
rect 11228 24002 11283 24054
rect 11335 24002 12228 24054
rect 11228 23946 12228 24002
rect 11228 23894 11283 23946
rect 11335 23894 12228 23946
rect 11228 23838 12228 23894
rect 11228 23786 11283 23838
rect 11335 23786 12228 23838
rect 11228 23730 12228 23786
rect 11228 23678 11283 23730
rect 11335 23678 12228 23730
rect 11228 23622 12228 23678
rect 11228 23570 11283 23622
rect 11335 23570 12228 23622
rect 11228 23514 12228 23570
rect 11228 23462 11283 23514
rect 11335 23462 12228 23514
rect 11228 23406 12228 23462
rect 11228 23354 11283 23406
rect 11335 23354 12228 23406
rect 11228 23298 12228 23354
rect 11228 23246 11283 23298
rect 11335 23246 12228 23298
rect 11228 23190 12228 23246
rect 11228 23138 11283 23190
rect 11335 23138 12228 23190
rect 11228 23082 12228 23138
rect 11228 23030 11283 23082
rect 11335 23030 12228 23082
rect 11228 22974 12228 23030
rect 11228 22922 11283 22974
rect 11335 22922 12228 22974
rect 11228 22866 12228 22922
rect 11228 22814 11283 22866
rect 11335 22814 12228 22866
rect 11228 22758 12228 22814
rect 11228 22706 11283 22758
rect 11335 22706 12228 22758
rect 11228 22650 12228 22706
rect 11228 22598 11283 22650
rect 11335 22598 12228 22650
rect 11228 22542 12228 22598
rect 11228 22490 11283 22542
rect 11335 22490 12228 22542
rect 11228 22434 12228 22490
rect 11228 22382 11283 22434
rect 11335 22382 12228 22434
rect 11228 22326 12228 22382
rect 11228 22274 11283 22326
rect 11335 22274 12228 22326
rect 11228 22218 12228 22274
rect 11228 22166 11283 22218
rect 11335 22166 12228 22218
rect 11228 22110 12228 22166
rect 11228 22058 11283 22110
rect 11335 22058 12228 22110
rect 11228 22002 12228 22058
rect 11228 21950 11283 22002
rect 11335 21950 12228 22002
rect 11228 21894 12228 21950
rect 11228 21842 11283 21894
rect 11335 21842 12228 21894
rect 11228 21786 12228 21842
rect 11228 21734 11283 21786
rect 11335 21734 12228 21786
rect 11228 21678 12228 21734
rect 11228 21631 11283 21678
rect 11335 21642 12228 21678
rect 13144 24616 14144 24686
rect 13144 24564 13786 24616
rect 13838 24564 13910 24616
rect 13962 24564 14034 24616
rect 14086 24564 14144 24616
rect 13144 24492 14144 24564
rect 13144 24440 13786 24492
rect 13838 24440 13910 24492
rect 13962 24440 14034 24492
rect 14086 24440 14144 24492
rect 13144 24368 14144 24440
rect 13144 24316 13786 24368
rect 13838 24316 13910 24368
rect 13962 24316 14034 24368
rect 14086 24316 14144 24368
rect 13144 24244 14144 24316
rect 13144 24192 13786 24244
rect 13838 24192 13910 24244
rect 13962 24192 14034 24244
rect 14086 24192 14144 24244
rect 13144 24120 14144 24192
rect 13144 24068 13786 24120
rect 13838 24068 13910 24120
rect 13962 24068 14034 24120
rect 14086 24068 14144 24120
rect 13144 23996 14144 24068
rect 13144 23944 13786 23996
rect 13838 23944 13910 23996
rect 13962 23944 14034 23996
rect 14086 23944 14144 23996
rect 13144 23872 14144 23944
rect 13144 23820 13786 23872
rect 13838 23820 13910 23872
rect 13962 23820 14034 23872
rect 14086 23820 14144 23872
rect 13144 23748 14144 23820
rect 13144 23696 13786 23748
rect 13838 23696 13910 23748
rect 13962 23696 14034 23748
rect 14086 23696 14144 23748
rect 13144 23624 14144 23696
rect 13144 23572 13786 23624
rect 13838 23572 13910 23624
rect 13962 23572 14034 23624
rect 14086 23572 14144 23624
rect 13144 23500 14144 23572
rect 13144 23448 13786 23500
rect 13838 23448 13910 23500
rect 13962 23448 14034 23500
rect 14086 23448 14144 23500
rect 13144 23376 14144 23448
rect 13144 23324 13786 23376
rect 13838 23324 13910 23376
rect 13962 23324 14034 23376
rect 14086 23324 14144 23376
rect 13144 23252 14144 23324
rect 13144 23200 13786 23252
rect 13838 23200 13910 23252
rect 13962 23200 14034 23252
rect 14086 23200 14144 23252
rect 13144 23128 14144 23200
rect 13144 23076 13786 23128
rect 13838 23076 13910 23128
rect 13962 23076 14034 23128
rect 14086 23076 14144 23128
rect 13144 23004 14144 23076
rect 13144 22952 13786 23004
rect 13838 22952 13910 23004
rect 13962 22952 14034 23004
rect 14086 22952 14144 23004
rect 13144 22880 14144 22952
rect 13144 22828 13786 22880
rect 13838 22828 13910 22880
rect 13962 22828 14034 22880
rect 14086 22828 14144 22880
rect 13144 22756 14144 22828
rect 13144 22704 13786 22756
rect 13838 22704 13910 22756
rect 13962 22704 14034 22756
rect 14086 22704 14144 22756
rect 13144 22632 14144 22704
rect 13144 22580 13786 22632
rect 13838 22580 13910 22632
rect 13962 22580 14034 22632
rect 14086 22580 14144 22632
rect 13144 22508 14144 22580
rect 13144 22456 13786 22508
rect 13838 22456 13910 22508
rect 13962 22456 14034 22508
rect 14086 22456 14144 22508
rect 13144 22384 14144 22456
rect 13144 22332 13786 22384
rect 13838 22332 13910 22384
rect 13962 22332 14034 22384
rect 14086 22332 14144 22384
rect 13144 22260 14144 22332
rect 13144 22208 13786 22260
rect 13838 22208 13910 22260
rect 13962 22208 14034 22260
rect 14086 22208 14144 22260
rect 13144 22136 14144 22208
rect 13144 22084 13786 22136
rect 13838 22084 13910 22136
rect 13962 22084 14034 22136
rect 14086 22084 14144 22136
rect 13144 22012 14144 22084
rect 13144 21960 13786 22012
rect 13838 21960 13910 22012
rect 13962 21960 14034 22012
rect 14086 21960 14144 22012
rect 13144 21888 14144 21960
rect 13144 21836 13786 21888
rect 13838 21836 13910 21888
rect 13962 21836 14034 21888
rect 14086 21836 14144 21888
rect 13144 21764 14144 21836
rect 13144 21712 13786 21764
rect 13838 21712 13910 21764
rect 13962 21712 14034 21764
rect 14086 21712 14144 21764
rect 13144 21642 14144 21712
rect 11335 21640 14144 21642
rect 11335 21631 13786 21640
rect 13838 21631 13910 21640
rect 13962 21631 14034 21640
rect 14086 21631 14144 21640
rect 11228 21585 11239 21631
rect 14133 21585 14144 21631
rect 11228 21574 14144 21585
rect 14204 24627 14404 24664
rect 14204 21701 14215 24627
rect 14261 21701 14404 24627
rect 14204 21514 14404 21701
rect 14608 21514 14619 24814
rect 445 21469 14619 21514
rect 496 21417 552 21469
rect 604 21417 660 21469
rect 712 21417 1408 21469
rect 1460 21417 1516 21469
rect 1568 21417 1624 21469
rect 1676 21417 1732 21469
rect 1784 21417 1840 21469
rect 1892 21417 2544 21469
rect 2596 21417 2652 21469
rect 2704 21417 2760 21469
rect 2812 21417 2868 21469
rect 2920 21417 2976 21469
rect 3028 21417 4816 21469
rect 4868 21417 4924 21469
rect 4976 21417 5032 21469
rect 5084 21417 5140 21469
rect 5192 21417 5248 21469
rect 5300 21417 7101 21469
rect 7153 21417 7209 21469
rect 7261 21417 7317 21469
rect 7369 21417 7425 21469
rect 7477 21417 7587 21469
rect 7639 21417 7695 21469
rect 7747 21417 7803 21469
rect 7855 21417 7911 21469
rect 7963 21417 9764 21469
rect 9816 21417 9872 21469
rect 9924 21417 9980 21469
rect 10032 21417 10088 21469
rect 10140 21417 10196 21469
rect 10248 21417 12036 21469
rect 12088 21417 12144 21469
rect 12196 21417 12252 21469
rect 12304 21417 12360 21469
rect 12412 21417 12468 21469
rect 12520 21417 13172 21469
rect 13224 21417 13280 21469
rect 13332 21417 13388 21469
rect 13440 21417 13496 21469
rect 13548 21417 13604 21469
rect 13656 21417 14352 21469
rect 14404 21417 14460 21469
rect 14512 21417 14568 21469
rect 445 21361 14619 21417
rect 496 21309 552 21361
rect 604 21309 660 21361
rect 712 21309 1408 21361
rect 1460 21309 1516 21361
rect 1568 21309 1624 21361
rect 1676 21309 1732 21361
rect 1784 21309 1840 21361
rect 1892 21309 2544 21361
rect 2596 21309 2652 21361
rect 2704 21309 2760 21361
rect 2812 21309 2868 21361
rect 2920 21309 2976 21361
rect 3028 21309 4816 21361
rect 4868 21309 4924 21361
rect 4976 21309 5032 21361
rect 5084 21309 5140 21361
rect 5192 21309 5248 21361
rect 5300 21309 7101 21361
rect 7153 21309 7209 21361
rect 7261 21309 7317 21361
rect 7369 21309 7425 21361
rect 7477 21309 7587 21361
rect 7639 21309 7695 21361
rect 7747 21309 7803 21361
rect 7855 21309 7911 21361
rect 7963 21309 9764 21361
rect 9816 21309 9872 21361
rect 9924 21309 9980 21361
rect 10032 21309 10088 21361
rect 10140 21309 10196 21361
rect 10248 21309 12036 21361
rect 12088 21309 12144 21361
rect 12196 21309 12252 21361
rect 12304 21309 12360 21361
rect 12412 21309 12468 21361
rect 12520 21309 13172 21361
rect 13224 21309 13280 21361
rect 13332 21309 13388 21361
rect 13440 21309 13496 21361
rect 13548 21309 13604 21361
rect 13656 21309 14352 21361
rect 14404 21309 14460 21361
rect 14512 21309 14568 21361
rect 445 21253 14619 21309
rect 496 21201 552 21253
rect 604 21213 660 21253
rect 712 21213 1408 21253
rect 1460 21213 1516 21253
rect 1568 21213 1624 21253
rect 1676 21213 1732 21253
rect 1784 21213 1840 21253
rect 1892 21213 2544 21253
rect 2596 21213 2652 21253
rect 2704 21213 2760 21253
rect 2812 21213 2868 21253
rect 2920 21213 2976 21253
rect 3028 21213 4816 21253
rect 4868 21213 4924 21253
rect 4976 21213 5032 21253
rect 5084 21213 5140 21253
rect 5192 21213 5248 21253
rect 5300 21213 7101 21253
rect 7153 21213 7209 21253
rect 7261 21213 7317 21253
rect 7369 21213 7425 21253
rect 7477 21213 7587 21253
rect 7639 21213 7695 21253
rect 7747 21213 7803 21253
rect 7855 21213 7911 21253
rect 7963 21213 9764 21253
rect 9816 21213 9872 21253
rect 9924 21213 9980 21253
rect 10032 21213 10088 21253
rect 10140 21213 10196 21253
rect 10248 21213 12036 21253
rect 12088 21213 12144 21253
rect 12196 21213 12252 21253
rect 12304 21213 12360 21253
rect 12412 21213 12468 21253
rect 12520 21213 13172 21253
rect 13224 21213 13280 21253
rect 13332 21213 13388 21253
rect 13440 21213 13496 21253
rect 13548 21213 13604 21253
rect 13656 21213 14352 21253
rect 14404 21213 14460 21253
rect 14512 21201 14568 21253
rect 445 21167 553 21201
rect 14511 21167 14619 21201
rect 14665 21167 14676 56745
rect 388 21156 14676 21167
rect 14942 52271 15064 57254
rect 14942 52219 14954 52271
rect 15006 52219 15064 52271
rect 14942 52163 15064 52219
rect 14942 52111 14954 52163
rect 15006 52111 15064 52163
rect 14942 52055 15064 52111
rect 14942 52003 14954 52055
rect 15006 52003 15064 52055
rect 14942 51947 15064 52003
rect 14942 51895 14954 51947
rect 15006 51895 15064 51947
rect 14942 51839 15064 51895
rect 14942 51787 14954 51839
rect 15006 51787 15064 51839
rect 14942 51731 15064 51787
rect 14942 51679 14954 51731
rect 15006 51679 15064 51731
rect 14942 51623 15064 51679
rect 14942 51571 14954 51623
rect 15006 51571 15064 51623
rect 14942 51515 15064 51571
rect 14942 51463 14954 51515
rect 15006 51463 15064 51515
rect 14942 51407 15064 51463
rect 14942 51355 14954 51407
rect 15006 51355 15064 51407
rect 14942 51299 15064 51355
rect 14942 51247 14954 51299
rect 15006 51247 15064 51299
rect 14942 51191 15064 51247
rect 14942 51139 14954 51191
rect 15006 51139 15064 51191
rect 14942 51083 15064 51139
rect 14942 51031 14954 51083
rect 15006 51031 15064 51083
rect 14942 50975 15064 51031
rect 14942 50923 14954 50975
rect 15006 50923 15064 50975
rect 14942 37871 15064 50923
rect 14942 37819 14954 37871
rect 15006 37819 15064 37871
rect 14942 37763 15064 37819
rect 14942 37711 14954 37763
rect 15006 37711 15064 37763
rect 14942 37655 15064 37711
rect 14942 37603 14954 37655
rect 15006 37603 15064 37655
rect 14942 37547 15064 37603
rect 14942 37495 14954 37547
rect 15006 37495 15064 37547
rect 14942 37439 15064 37495
rect 14942 37387 14954 37439
rect 15006 37387 15064 37439
rect 14942 37331 15064 37387
rect 14942 37279 14954 37331
rect 15006 37279 15064 37331
rect 14942 37223 15064 37279
rect 14942 37171 14954 37223
rect 15006 37171 15064 37223
rect 14942 37115 15064 37171
rect 14942 37063 14954 37115
rect 15006 37063 15064 37115
rect 14942 37007 15064 37063
rect 14942 36955 14954 37007
rect 15006 36955 15064 37007
rect 14942 36899 15064 36955
rect 14942 36847 14954 36899
rect 15006 36847 15064 36899
rect 14942 36791 15064 36847
rect 14942 36739 14954 36791
rect 15006 36739 15064 36791
rect 14942 36683 15064 36739
rect 14942 36631 14954 36683
rect 15006 36631 15064 36683
rect 14942 36575 15064 36631
rect 14942 36523 14954 36575
rect 15006 36523 15064 36575
rect 2494 20619 12570 20630
rect 0 20357 1068 20368
rect 0 19368 311 20357
rect 0 19168 122 19368
rect 300 19168 311 19368
rect 0 18168 311 19168
rect 0 17968 122 18168
rect 300 17968 311 18168
rect 0 16968 311 17968
rect 0 16768 122 16968
rect 300 16768 311 16968
rect 0 15768 311 16768
rect 0 15568 122 15768
rect 300 15568 311 15768
rect 0 14568 311 15568
rect 0 14368 122 14568
rect 300 14368 311 14568
rect 0 13368 311 14368
rect 0 13168 122 13368
rect 300 13168 311 13368
rect 0 12168 311 13168
rect 0 11968 122 12168
rect 300 11968 311 12168
rect 0 10968 311 11968
rect 0 10768 122 10968
rect 300 10768 311 10968
rect 0 9768 311 10768
rect 0 9100 122 9768
rect 300 9100 311 9768
rect 0 8100 311 9100
rect 0 7900 122 8100
rect 300 7900 311 8100
rect 0 6900 311 7900
rect 0 6700 122 6900
rect 300 6700 311 6900
rect 0 5700 311 6700
rect 0 5500 122 5700
rect 300 5500 311 5700
rect 0 4500 311 5500
rect 0 4300 122 4500
rect 300 4300 311 4500
rect 0 3300 311 4300
rect 0 3100 122 3300
rect 300 3100 311 3300
rect 0 2100 311 3100
rect 0 1900 122 2100
rect 300 1900 311 2100
rect 0 911 311 1900
rect 1057 911 1068 20357
rect 2494 15773 2505 20619
rect 2851 20273 2959 20619
rect 12105 20273 12213 20619
rect 2851 20262 12213 20273
rect 2851 16130 2862 20262
rect 3127 19971 11937 19982
rect 3127 19925 3138 19971
rect 11926 19925 11937 19971
rect 3127 19899 4816 19925
rect 4868 19899 4924 19925
rect 4976 19899 5032 19925
rect 5084 19899 5140 19925
rect 5192 19899 5248 19925
rect 5300 19899 7101 19925
rect 7153 19899 7209 19925
rect 7261 19899 7317 19925
rect 7369 19899 7425 19925
rect 7477 19899 7587 19925
rect 7639 19899 7695 19925
rect 7747 19899 7803 19925
rect 7855 19899 7911 19925
rect 7963 19899 9764 19925
rect 9816 19899 9872 19925
rect 9924 19899 9980 19925
rect 10032 19899 10088 19925
rect 10140 19899 10196 19925
rect 10248 19899 11937 19925
rect 3127 19843 11937 19899
rect 3127 19817 4816 19843
rect 4868 19817 4924 19843
rect 4976 19817 5032 19843
rect 5084 19817 5140 19843
rect 5192 19817 5248 19843
rect 5300 19817 7101 19843
rect 7153 19817 7209 19843
rect 7261 19817 7317 19843
rect 7369 19817 7425 19843
rect 7477 19817 7587 19843
rect 7639 19817 7695 19843
rect 7747 19817 7803 19843
rect 7855 19817 7911 19843
rect 7963 19817 9764 19843
rect 9816 19817 9872 19843
rect 9924 19817 9980 19843
rect 10032 19817 10088 19843
rect 10140 19817 10196 19843
rect 10248 19817 11937 19843
rect 3127 16575 3138 19817
rect 3184 19809 3467 19817
rect 3184 19199 3292 19809
rect 3338 19771 3467 19809
rect 11597 19809 11880 19817
rect 11597 19771 11726 19809
rect 3338 19760 11726 19771
rect 3338 19256 3349 19760
rect 3532 19591 11532 19604
rect 3532 19545 3545 19591
rect 11519 19545 11532 19591
rect 3532 19532 3680 19545
rect 3732 19532 3788 19545
rect 3840 19532 3896 19545
rect 3948 19532 4004 19545
rect 4056 19532 4112 19545
rect 4164 19532 5952 19545
rect 6004 19532 6060 19545
rect 6112 19532 6168 19545
rect 6220 19532 6276 19545
rect 6328 19532 6384 19545
rect 6436 19532 8628 19545
rect 8680 19532 8736 19545
rect 8788 19532 8844 19545
rect 8896 19532 8952 19545
rect 9004 19532 9060 19545
rect 9112 19532 10900 19545
rect 10952 19532 11008 19545
rect 11060 19532 11116 19545
rect 11168 19532 11224 19545
rect 11276 19532 11332 19545
rect 11384 19532 11532 19545
rect 3532 19476 11532 19532
rect 3532 19463 3680 19476
rect 3732 19463 3788 19476
rect 3840 19463 3896 19476
rect 3948 19463 4004 19476
rect 4056 19463 4112 19476
rect 4164 19463 5952 19476
rect 6004 19463 6060 19476
rect 6112 19463 6168 19476
rect 6220 19463 6276 19476
rect 6328 19463 6384 19476
rect 6436 19463 8628 19476
rect 8680 19463 8736 19476
rect 8788 19463 8844 19476
rect 8896 19463 8952 19476
rect 9004 19463 9060 19476
rect 9112 19463 10900 19476
rect 10952 19463 11008 19476
rect 11060 19463 11116 19476
rect 11168 19463 11224 19476
rect 11276 19463 11332 19476
rect 11384 19463 11532 19476
rect 3532 19417 3545 19463
rect 11519 19417 11532 19463
rect 3532 19404 11532 19417
rect 11715 19256 11726 19760
rect 3338 19245 11726 19256
rect 3338 19199 3467 19245
rect 11597 19199 11726 19245
rect 11772 19199 11880 19809
rect 3184 19150 4816 19199
rect 4868 19150 4924 19199
rect 4976 19150 5032 19199
rect 5084 19150 5140 19199
rect 5192 19150 5248 19199
rect 5300 19150 7101 19199
rect 7153 19150 7209 19199
rect 7261 19150 7317 19199
rect 7369 19150 7425 19199
rect 7477 19150 7587 19199
rect 7639 19150 7695 19199
rect 7747 19150 7803 19199
rect 7855 19150 7911 19199
rect 7963 19150 9764 19199
rect 9816 19150 9872 19199
rect 9924 19150 9980 19199
rect 10032 19150 10088 19199
rect 10140 19150 10196 19199
rect 10248 19150 11880 19199
rect 3184 19094 11880 19150
rect 3184 19091 4816 19094
rect 4868 19091 4924 19094
rect 4976 19091 5032 19094
rect 5084 19091 5140 19094
rect 5192 19091 5248 19094
rect 5300 19091 7101 19094
rect 7153 19091 7209 19094
rect 7261 19091 7317 19094
rect 7369 19091 7425 19094
rect 7477 19091 7587 19094
rect 7639 19091 7695 19094
rect 7747 19091 7803 19094
rect 7855 19091 7911 19094
rect 7963 19091 9764 19094
rect 9816 19091 9872 19094
rect 9924 19091 9980 19094
rect 10032 19091 10088 19094
rect 10140 19091 10196 19094
rect 10248 19091 11880 19094
rect 3184 19045 3326 19091
rect 11738 19045 11880 19091
rect 3184 19042 4816 19045
rect 4868 19042 4924 19045
rect 4976 19042 5032 19045
rect 5084 19042 5140 19045
rect 5192 19042 5248 19045
rect 5300 19042 7101 19045
rect 7153 19042 7209 19045
rect 7261 19042 7317 19045
rect 7369 19042 7425 19045
rect 7477 19042 7587 19045
rect 7639 19042 7695 19045
rect 7747 19042 7803 19045
rect 7855 19042 7911 19045
rect 7963 19042 9764 19045
rect 9816 19042 9872 19045
rect 9924 19042 9980 19045
rect 10032 19042 10088 19045
rect 10140 19042 10196 19045
rect 10248 19042 11880 19045
rect 3184 18986 11880 19042
rect 3184 18937 4816 18986
rect 4868 18937 4924 18986
rect 4976 18937 5032 18986
rect 5084 18937 5140 18986
rect 5192 18937 5248 18986
rect 5300 18937 7101 18986
rect 7153 18937 7209 18986
rect 7261 18937 7317 18986
rect 7369 18937 7425 18986
rect 7477 18937 7587 18986
rect 7639 18937 7695 18986
rect 7747 18937 7803 18986
rect 7855 18937 7911 18986
rect 7963 18937 9764 18986
rect 9816 18937 9872 18986
rect 9924 18937 9980 18986
rect 10032 18937 10088 18986
rect 10140 18937 10196 18986
rect 10248 18937 11880 18986
rect 3184 18327 3292 18937
rect 3338 18891 3467 18937
rect 11597 18891 11726 18937
rect 3338 18880 11726 18891
rect 3338 18384 3349 18880
rect 3532 18719 11532 18732
rect 3532 18673 3545 18719
rect 11519 18673 11532 18719
rect 3532 18660 3680 18673
rect 3732 18660 3788 18673
rect 3840 18660 3896 18673
rect 3948 18660 4004 18673
rect 4056 18660 4112 18673
rect 4164 18660 5952 18673
rect 6004 18660 6060 18673
rect 6112 18660 6168 18673
rect 6220 18660 6276 18673
rect 6328 18660 6384 18673
rect 6436 18660 8628 18673
rect 8680 18660 8736 18673
rect 8788 18660 8844 18673
rect 8896 18660 8952 18673
rect 9004 18660 9060 18673
rect 9112 18660 10900 18673
rect 10952 18660 11008 18673
rect 11060 18660 11116 18673
rect 11168 18660 11224 18673
rect 11276 18660 11332 18673
rect 11384 18660 11532 18673
rect 3532 18604 11532 18660
rect 3532 18591 3680 18604
rect 3732 18591 3788 18604
rect 3840 18591 3896 18604
rect 3948 18591 4004 18604
rect 4056 18591 4112 18604
rect 4164 18591 5952 18604
rect 6004 18591 6060 18604
rect 6112 18591 6168 18604
rect 6220 18591 6276 18604
rect 6328 18591 6384 18604
rect 6436 18591 8628 18604
rect 8680 18591 8736 18604
rect 8788 18591 8844 18604
rect 8896 18591 8952 18604
rect 9004 18591 9060 18604
rect 9112 18591 10900 18604
rect 10952 18591 11008 18604
rect 11060 18591 11116 18604
rect 11168 18591 11224 18604
rect 11276 18591 11332 18604
rect 11384 18591 11532 18604
rect 3532 18545 3545 18591
rect 11519 18545 11532 18591
rect 3532 18532 11532 18545
rect 11715 18384 11726 18880
rect 3338 18373 11726 18384
rect 3338 18327 3467 18373
rect 11597 18327 11726 18373
rect 11772 18327 11880 18937
rect 3184 18278 4816 18327
rect 4868 18278 4924 18327
rect 4976 18278 5032 18327
rect 5084 18278 5140 18327
rect 5192 18278 5248 18327
rect 5300 18278 7101 18327
rect 7153 18278 7209 18327
rect 7261 18278 7317 18327
rect 7369 18278 7425 18327
rect 7477 18278 7587 18327
rect 7639 18278 7695 18327
rect 7747 18278 7803 18327
rect 7855 18278 7911 18327
rect 7963 18278 9764 18327
rect 9816 18278 9872 18327
rect 9924 18278 9980 18327
rect 10032 18278 10088 18327
rect 10140 18278 10196 18327
rect 10248 18278 11880 18327
rect 3184 18222 11880 18278
rect 3184 18219 4816 18222
rect 4868 18219 4924 18222
rect 4976 18219 5032 18222
rect 5084 18219 5140 18222
rect 5192 18219 5248 18222
rect 5300 18219 7101 18222
rect 7153 18219 7209 18222
rect 7261 18219 7317 18222
rect 7369 18219 7425 18222
rect 7477 18219 7587 18222
rect 7639 18219 7695 18222
rect 7747 18219 7803 18222
rect 7855 18219 7911 18222
rect 7963 18219 9764 18222
rect 9816 18219 9872 18222
rect 9924 18219 9980 18222
rect 10032 18219 10088 18222
rect 10140 18219 10196 18222
rect 10248 18219 11880 18222
rect 3184 18173 3326 18219
rect 11738 18173 11880 18219
rect 3184 18170 4816 18173
rect 4868 18170 4924 18173
rect 4976 18170 5032 18173
rect 5084 18170 5140 18173
rect 5192 18170 5248 18173
rect 5300 18170 7101 18173
rect 7153 18170 7209 18173
rect 7261 18170 7317 18173
rect 7369 18170 7425 18173
rect 7477 18170 7587 18173
rect 7639 18170 7695 18173
rect 7747 18170 7803 18173
rect 7855 18170 7911 18173
rect 7963 18170 9764 18173
rect 9816 18170 9872 18173
rect 9924 18170 9980 18173
rect 10032 18170 10088 18173
rect 10140 18170 10196 18173
rect 10248 18170 11880 18173
rect 3184 18114 11880 18170
rect 3184 18065 4816 18114
rect 4868 18065 4924 18114
rect 4976 18065 5032 18114
rect 5084 18065 5140 18114
rect 5192 18065 5248 18114
rect 5300 18065 7101 18114
rect 7153 18065 7209 18114
rect 7261 18065 7317 18114
rect 7369 18065 7425 18114
rect 7477 18065 7587 18114
rect 7639 18065 7695 18114
rect 7747 18065 7803 18114
rect 7855 18065 7911 18114
rect 7963 18065 9764 18114
rect 9816 18065 9872 18114
rect 9924 18065 9980 18114
rect 10032 18065 10088 18114
rect 10140 18065 10196 18114
rect 10248 18065 11880 18114
rect 3184 17455 3292 18065
rect 3338 18019 3467 18065
rect 11597 18019 11726 18065
rect 3338 18008 11726 18019
rect 3338 17512 3349 18008
rect 3532 17847 11532 17860
rect 3532 17801 3545 17847
rect 11519 17801 11532 17847
rect 3532 17788 3680 17801
rect 3732 17788 3788 17801
rect 3840 17788 3896 17801
rect 3948 17788 4004 17801
rect 4056 17788 4112 17801
rect 4164 17788 5952 17801
rect 6004 17788 6060 17801
rect 6112 17788 6168 17801
rect 6220 17788 6276 17801
rect 6328 17788 6384 17801
rect 6436 17788 8628 17801
rect 8680 17788 8736 17801
rect 8788 17788 8844 17801
rect 8896 17788 8952 17801
rect 9004 17788 9060 17801
rect 9112 17788 10900 17801
rect 10952 17788 11008 17801
rect 11060 17788 11116 17801
rect 11168 17788 11224 17801
rect 11276 17788 11332 17801
rect 11384 17788 11532 17801
rect 3532 17732 11532 17788
rect 3532 17719 3680 17732
rect 3732 17719 3788 17732
rect 3840 17719 3896 17732
rect 3948 17719 4004 17732
rect 4056 17719 4112 17732
rect 4164 17719 5952 17732
rect 6004 17719 6060 17732
rect 6112 17719 6168 17732
rect 6220 17719 6276 17732
rect 6328 17719 6384 17732
rect 6436 17719 8628 17732
rect 8680 17719 8736 17732
rect 8788 17719 8844 17732
rect 8896 17719 8952 17732
rect 9004 17719 9060 17732
rect 9112 17719 10900 17732
rect 10952 17719 11008 17732
rect 11060 17719 11116 17732
rect 11168 17719 11224 17732
rect 11276 17719 11332 17732
rect 11384 17719 11532 17732
rect 3532 17673 3545 17719
rect 11519 17673 11532 17719
rect 3532 17660 11532 17673
rect 11715 17512 11726 18008
rect 3338 17501 11726 17512
rect 3338 17455 3467 17501
rect 11597 17455 11726 17501
rect 11772 17455 11880 18065
rect 3184 17406 4816 17455
rect 4868 17406 4924 17455
rect 4976 17406 5032 17455
rect 5084 17406 5140 17455
rect 5192 17406 5248 17455
rect 5300 17406 7101 17455
rect 7153 17406 7209 17455
rect 7261 17406 7317 17455
rect 7369 17406 7425 17455
rect 7477 17406 7587 17455
rect 7639 17406 7695 17455
rect 7747 17406 7803 17455
rect 7855 17406 7911 17455
rect 7963 17406 9764 17455
rect 9816 17406 9872 17455
rect 9924 17406 9980 17455
rect 10032 17406 10088 17455
rect 10140 17406 10196 17455
rect 10248 17406 11880 17455
rect 3184 17350 11880 17406
rect 3184 17347 4816 17350
rect 4868 17347 4924 17350
rect 4976 17347 5032 17350
rect 5084 17347 5140 17350
rect 5192 17347 5248 17350
rect 5300 17347 7101 17350
rect 7153 17347 7209 17350
rect 7261 17347 7317 17350
rect 7369 17347 7425 17350
rect 7477 17347 7587 17350
rect 7639 17347 7695 17350
rect 7747 17347 7803 17350
rect 7855 17347 7911 17350
rect 7963 17347 9764 17350
rect 9816 17347 9872 17350
rect 9924 17347 9980 17350
rect 10032 17347 10088 17350
rect 10140 17347 10196 17350
rect 10248 17347 11880 17350
rect 3184 17301 3326 17347
rect 11738 17301 11880 17347
rect 3184 17298 4816 17301
rect 4868 17298 4924 17301
rect 4976 17298 5032 17301
rect 5084 17298 5140 17301
rect 5192 17298 5248 17301
rect 5300 17298 7101 17301
rect 7153 17298 7209 17301
rect 7261 17298 7317 17301
rect 7369 17298 7425 17301
rect 7477 17298 7587 17301
rect 7639 17298 7695 17301
rect 7747 17298 7803 17301
rect 7855 17298 7911 17301
rect 7963 17298 9764 17301
rect 9816 17298 9872 17301
rect 9924 17298 9980 17301
rect 10032 17298 10088 17301
rect 10140 17298 10196 17301
rect 10248 17298 11880 17301
rect 3184 17242 11880 17298
rect 3184 17193 4816 17242
rect 4868 17193 4924 17242
rect 4976 17193 5032 17242
rect 5084 17193 5140 17242
rect 5192 17193 5248 17242
rect 5300 17193 7101 17242
rect 7153 17193 7209 17242
rect 7261 17193 7317 17242
rect 7369 17193 7425 17242
rect 7477 17193 7587 17242
rect 7639 17193 7695 17242
rect 7747 17193 7803 17242
rect 7855 17193 7911 17242
rect 7963 17193 9764 17242
rect 9816 17193 9872 17242
rect 9924 17193 9980 17242
rect 10032 17193 10088 17242
rect 10140 17193 10196 17242
rect 10248 17193 11880 17242
rect 3184 16583 3292 17193
rect 3338 17147 3467 17193
rect 11597 17147 11726 17193
rect 3338 17136 11726 17147
rect 3338 16632 3349 17136
rect 3532 16975 11532 16988
rect 3532 16929 3545 16975
rect 11519 16929 11532 16975
rect 3532 16916 3680 16929
rect 3732 16916 3788 16929
rect 3840 16916 3896 16929
rect 3948 16916 4004 16929
rect 4056 16916 4112 16929
rect 4164 16916 5952 16929
rect 6004 16916 6060 16929
rect 6112 16916 6168 16929
rect 6220 16916 6276 16929
rect 6328 16916 6384 16929
rect 6436 16916 8628 16929
rect 8680 16916 8736 16929
rect 8788 16916 8844 16929
rect 8896 16916 8952 16929
rect 9004 16916 9060 16929
rect 9112 16916 10900 16929
rect 10952 16916 11008 16929
rect 11060 16916 11116 16929
rect 11168 16916 11224 16929
rect 11276 16916 11332 16929
rect 11384 16916 11532 16929
rect 3532 16860 11532 16916
rect 3532 16847 3680 16860
rect 3732 16847 3788 16860
rect 3840 16847 3896 16860
rect 3948 16847 4004 16860
rect 4056 16847 4112 16860
rect 4164 16847 5952 16860
rect 6004 16847 6060 16860
rect 6112 16847 6168 16860
rect 6220 16847 6276 16860
rect 6328 16847 6384 16860
rect 6436 16847 8628 16860
rect 8680 16847 8736 16860
rect 8788 16847 8844 16860
rect 8896 16847 8952 16860
rect 9004 16847 9060 16860
rect 9112 16847 10900 16860
rect 10952 16847 11008 16860
rect 11060 16847 11116 16860
rect 11168 16847 11224 16860
rect 11276 16847 11332 16860
rect 11384 16847 11532 16860
rect 3532 16801 3545 16847
rect 11519 16801 11532 16847
rect 3532 16788 11532 16801
rect 11715 16632 11726 17136
rect 3338 16621 11726 16632
rect 3338 16583 3467 16621
rect 3184 16575 3467 16583
rect 11597 16583 11726 16621
rect 11772 16583 11880 17193
rect 11597 16575 11880 16583
rect 11926 16575 11937 19817
rect 3127 16549 4816 16575
rect 4868 16549 4924 16575
rect 4976 16549 5032 16575
rect 5084 16549 5140 16575
rect 5192 16549 5248 16575
rect 5300 16549 7101 16575
rect 7153 16549 7209 16575
rect 7261 16549 7317 16575
rect 7369 16549 7425 16575
rect 7477 16549 7587 16575
rect 7639 16549 7695 16575
rect 7747 16549 7803 16575
rect 7855 16549 7911 16575
rect 7963 16549 9764 16575
rect 9816 16549 9872 16575
rect 9924 16549 9980 16575
rect 10032 16549 10088 16575
rect 10140 16549 10196 16575
rect 10248 16549 11937 16575
rect 3127 16493 11937 16549
rect 3127 16467 4816 16493
rect 4868 16467 4924 16493
rect 4976 16467 5032 16493
rect 5084 16467 5140 16493
rect 5192 16467 5248 16493
rect 5300 16467 7101 16493
rect 7153 16467 7209 16493
rect 7261 16467 7317 16493
rect 7369 16467 7425 16493
rect 7477 16467 7587 16493
rect 7639 16467 7695 16493
rect 7747 16467 7803 16493
rect 7855 16467 7911 16493
rect 7963 16467 9764 16493
rect 9816 16467 9872 16493
rect 9924 16467 9980 16493
rect 10032 16467 10088 16493
rect 10140 16467 10196 16493
rect 10248 16467 11937 16493
rect 3127 16421 3138 16467
rect 11926 16421 11937 16467
rect 3127 16410 11937 16421
rect 12202 16130 12213 20262
rect 2851 16119 12213 16130
rect 2851 15773 2959 16119
rect 12105 15773 12213 16119
rect 12559 15773 12570 20619
rect 14942 20368 15064 36523
rect 2494 15762 12570 15773
rect 13996 20357 15064 20368
rect 0 900 1068 911
rect 13996 911 14007 20357
rect 14753 19368 15064 20357
rect 14753 19168 14764 19368
rect 14942 19168 15064 19368
rect 14753 18168 15064 19168
rect 14753 17968 14764 18168
rect 14942 17968 15064 18168
rect 14753 16968 15064 17968
rect 14753 16768 14764 16968
rect 14942 16768 15064 16968
rect 14753 15768 15064 16768
rect 14753 15568 14764 15768
rect 14942 15568 15064 15768
rect 14753 14568 15064 15568
rect 14753 14368 14764 14568
rect 14942 14368 15064 14568
rect 14753 13368 15064 14368
rect 14753 13168 14764 13368
rect 14942 13168 15064 13368
rect 14753 12168 15064 13168
rect 14753 11968 14764 12168
rect 14942 11968 15064 12168
rect 14753 10968 15064 11968
rect 14753 10768 14764 10968
rect 14942 10768 15064 10968
rect 14753 9768 15064 10768
rect 14753 9100 14764 9768
rect 14942 9100 15064 9768
rect 14753 8100 15064 9100
rect 14753 7900 14764 8100
rect 14942 7900 15064 8100
rect 14753 6900 15064 7900
rect 14753 6700 14764 6900
rect 14942 6700 15064 6900
rect 14753 5700 15064 6700
rect 14753 5500 14764 5700
rect 14942 5500 15064 5700
rect 14753 4500 15064 5500
rect 14753 4300 14764 4500
rect 14942 4300 15064 4500
rect 14753 3300 15064 4300
rect 14753 3100 14764 3300
rect 14942 3100 15064 3300
rect 14753 2100 15064 3100
rect 14753 1900 14764 2100
rect 14942 1900 15064 2100
rect 14753 911 15064 1900
rect 13996 900 15064 911
rect 0 405 122 900
rect 14942 405 15064 900
<< via1 >>
rect 58 52219 110 52271
rect 58 52111 110 52163
rect 58 52003 110 52055
rect 58 51895 110 51947
rect 58 51787 110 51839
rect 58 51679 110 51731
rect 58 51571 110 51623
rect 58 51463 110 51515
rect 58 51355 110 51407
rect 58 51247 110 51299
rect 58 51139 110 51191
rect 58 51031 110 51083
rect 58 50923 110 50975
rect 58 37819 110 37871
rect 58 37711 110 37763
rect 58 37603 110 37655
rect 58 37495 110 37547
rect 58 37387 110 37439
rect 58 37279 110 37331
rect 58 37171 110 37223
rect 58 37063 110 37115
rect 58 36955 110 37007
rect 58 36847 110 36899
rect 58 36739 110 36791
rect 58 36631 110 36683
rect 58 36523 110 36575
rect 444 56659 445 56711
rect 445 56659 496 56711
rect 552 56699 553 56711
rect 553 56699 604 56711
rect 660 56699 712 56711
rect 1408 56699 1460 56711
rect 1516 56699 1568 56711
rect 1624 56699 1676 56711
rect 1732 56699 1784 56711
rect 1840 56699 1892 56711
rect 2544 56699 2596 56711
rect 2652 56699 2704 56711
rect 2760 56699 2812 56711
rect 2868 56699 2920 56711
rect 2976 56699 3028 56711
rect 4816 56699 4868 56711
rect 4924 56699 4976 56711
rect 5032 56699 5084 56711
rect 5140 56699 5192 56711
rect 5248 56699 5300 56711
rect 7101 56699 7153 56711
rect 7209 56699 7261 56711
rect 7317 56699 7369 56711
rect 7425 56699 7477 56711
rect 7587 56699 7639 56711
rect 7695 56699 7747 56711
rect 7803 56699 7855 56711
rect 7911 56699 7963 56711
rect 9764 56699 9816 56711
rect 9872 56699 9924 56711
rect 9980 56699 10032 56711
rect 10088 56699 10140 56711
rect 10196 56699 10248 56711
rect 12036 56699 12088 56711
rect 12144 56699 12196 56711
rect 12252 56699 12304 56711
rect 12360 56699 12412 56711
rect 12468 56699 12520 56711
rect 13172 56699 13224 56711
rect 13280 56699 13332 56711
rect 13388 56699 13440 56711
rect 13496 56699 13548 56711
rect 13604 56699 13656 56711
rect 14352 56699 14404 56711
rect 14460 56699 14511 56711
rect 14511 56699 14512 56711
rect 552 56659 604 56699
rect 660 56659 712 56699
rect 1408 56659 1460 56699
rect 1516 56659 1568 56699
rect 1624 56659 1676 56699
rect 1732 56659 1784 56699
rect 1840 56659 1892 56699
rect 2544 56659 2596 56699
rect 2652 56659 2704 56699
rect 2760 56659 2812 56699
rect 2868 56659 2920 56699
rect 2976 56659 3028 56699
rect 4816 56659 4868 56699
rect 4924 56659 4976 56699
rect 5032 56659 5084 56699
rect 5140 56659 5192 56699
rect 5248 56659 5300 56699
rect 7101 56659 7153 56699
rect 7209 56659 7261 56699
rect 7317 56659 7369 56699
rect 7425 56659 7477 56699
rect 7587 56659 7639 56699
rect 7695 56659 7747 56699
rect 7803 56659 7855 56699
rect 7911 56659 7963 56699
rect 9764 56659 9816 56699
rect 9872 56659 9924 56699
rect 9980 56659 10032 56699
rect 10088 56659 10140 56699
rect 10196 56659 10248 56699
rect 12036 56659 12088 56699
rect 12144 56659 12196 56699
rect 12252 56659 12304 56699
rect 12360 56659 12412 56699
rect 12468 56659 12520 56699
rect 13172 56659 13224 56699
rect 13280 56659 13332 56699
rect 13388 56659 13440 56699
rect 13496 56659 13548 56699
rect 13604 56659 13656 56699
rect 14352 56659 14404 56699
rect 14460 56659 14512 56699
rect 14568 56659 14619 56711
rect 14619 56659 14620 56711
rect 444 56551 445 56603
rect 445 56551 496 56603
rect 552 56551 604 56603
rect 660 56551 712 56603
rect 1408 56551 1460 56603
rect 1516 56551 1568 56603
rect 1624 56551 1676 56603
rect 1732 56551 1784 56603
rect 1840 56551 1892 56603
rect 2544 56551 2596 56603
rect 2652 56551 2704 56603
rect 2760 56551 2812 56603
rect 2868 56551 2920 56603
rect 2976 56551 3028 56603
rect 4816 56551 4868 56603
rect 4924 56551 4976 56603
rect 5032 56551 5084 56603
rect 5140 56551 5192 56603
rect 5248 56551 5300 56603
rect 7101 56551 7153 56603
rect 7209 56551 7261 56603
rect 7317 56551 7369 56603
rect 7425 56551 7477 56603
rect 7587 56551 7639 56603
rect 7695 56551 7747 56603
rect 7803 56551 7855 56603
rect 7911 56551 7963 56603
rect 9764 56551 9816 56603
rect 9872 56551 9924 56603
rect 9980 56551 10032 56603
rect 10088 56551 10140 56603
rect 10196 56551 10248 56603
rect 12036 56551 12088 56603
rect 12144 56551 12196 56603
rect 12252 56551 12304 56603
rect 12360 56551 12412 56603
rect 12468 56551 12520 56603
rect 13172 56551 13224 56603
rect 13280 56551 13332 56603
rect 13388 56551 13440 56603
rect 13496 56551 13548 56603
rect 13604 56551 13656 56603
rect 14352 56551 14404 56603
rect 14460 56551 14512 56603
rect 14568 56551 14619 56603
rect 14619 56551 14620 56603
rect 444 56443 445 56495
rect 445 56443 496 56495
rect 552 56443 604 56495
rect 660 56443 712 56495
rect 1408 56443 1460 56495
rect 1516 56443 1568 56495
rect 1624 56443 1676 56495
rect 1732 56443 1784 56495
rect 1840 56443 1892 56495
rect 2544 56443 2596 56495
rect 2652 56443 2704 56495
rect 2760 56443 2812 56495
rect 2868 56443 2920 56495
rect 2976 56443 3028 56495
rect 4816 56443 4868 56495
rect 4924 56443 4976 56495
rect 5032 56443 5084 56495
rect 5140 56443 5192 56495
rect 5248 56443 5300 56495
rect 7101 56443 7153 56495
rect 7209 56443 7261 56495
rect 7317 56443 7369 56495
rect 7425 56443 7477 56495
rect 7587 56443 7639 56495
rect 7695 56443 7747 56495
rect 7803 56443 7855 56495
rect 7911 56443 7963 56495
rect 9764 56443 9816 56495
rect 9872 56443 9924 56495
rect 9980 56443 10032 56495
rect 10088 56443 10140 56495
rect 10196 56443 10248 56495
rect 12036 56443 12088 56495
rect 12144 56443 12196 56495
rect 12252 56443 12304 56495
rect 12360 56443 12412 56495
rect 12468 56443 12520 56495
rect 13172 56443 13224 56495
rect 13280 56443 13332 56495
rect 13388 56443 13440 56495
rect 13496 56443 13548 56495
rect 13604 56443 13656 56495
rect 14352 56443 14404 56495
rect 14460 56443 14512 56495
rect 14568 56443 14619 56495
rect 14619 56443 14620 56495
rect 978 56281 1030 56324
rect 1102 56281 1154 56324
rect 1226 56281 1278 56324
rect 3729 56281 3781 56286
rect 978 56272 1030 56281
rect 1102 56272 1154 56281
rect 1226 56272 1278 56281
rect 978 56148 1030 56200
rect 1102 56148 1154 56200
rect 1226 56148 1278 56200
rect 978 56024 1030 56076
rect 1102 56024 1154 56076
rect 1226 56024 1278 56076
rect 978 55900 1030 55952
rect 1102 55900 1154 55952
rect 1226 55900 1278 55952
rect 978 55776 1030 55828
rect 1102 55776 1154 55828
rect 1226 55776 1278 55828
rect 978 55652 1030 55704
rect 1102 55652 1154 55704
rect 1226 55652 1278 55704
rect 978 55528 1030 55580
rect 1102 55528 1154 55580
rect 1226 55528 1278 55580
rect 978 55404 1030 55456
rect 1102 55404 1154 55456
rect 1226 55404 1278 55456
rect 978 55280 1030 55332
rect 1102 55280 1154 55332
rect 1226 55280 1278 55332
rect 978 55156 1030 55208
rect 1102 55156 1154 55208
rect 1226 55156 1278 55208
rect 978 55032 1030 55084
rect 1102 55032 1154 55084
rect 1226 55032 1278 55084
rect 978 54908 1030 54960
rect 1102 54908 1154 54960
rect 1226 54908 1278 54960
rect 978 54784 1030 54836
rect 1102 54784 1154 54836
rect 1226 54784 1278 54836
rect 978 54660 1030 54712
rect 1102 54660 1154 54712
rect 1226 54660 1278 54712
rect 978 54536 1030 54588
rect 1102 54536 1154 54588
rect 1226 54536 1278 54588
rect 978 54412 1030 54464
rect 1102 54412 1154 54464
rect 1226 54412 1278 54464
rect 978 54288 1030 54340
rect 1102 54288 1154 54340
rect 1226 54288 1278 54340
rect 978 54164 1030 54216
rect 1102 54164 1154 54216
rect 1226 54164 1278 54216
rect 978 54040 1030 54092
rect 1102 54040 1154 54092
rect 1226 54040 1278 54092
rect 978 53916 1030 53968
rect 1102 53916 1154 53968
rect 1226 53916 1278 53968
rect 978 53792 1030 53844
rect 1102 53792 1154 53844
rect 1226 53792 1278 53844
rect 978 53668 1030 53720
rect 1102 53668 1154 53720
rect 1226 53668 1278 53720
rect 978 53544 1030 53596
rect 1102 53544 1154 53596
rect 1226 53544 1278 53596
rect 978 53420 1030 53472
rect 1102 53420 1154 53472
rect 1226 53420 1278 53472
rect 978 53296 1030 53348
rect 1102 53296 1154 53348
rect 1226 53296 1278 53348
rect 3729 56234 3781 56281
rect 6335 56281 6387 56286
rect 3729 56126 3781 56178
rect 3729 56018 3781 56070
rect 3729 55910 3781 55962
rect 3729 55802 3781 55854
rect 3729 55694 3781 55746
rect 3729 55586 3781 55638
rect 3729 55478 3781 55530
rect 3729 55370 3781 55422
rect 3729 55262 3781 55314
rect 3729 55154 3781 55206
rect 3729 55046 3781 55098
rect 3729 54938 3781 54990
rect 3729 54830 3781 54882
rect 3729 54722 3781 54774
rect 3729 54614 3781 54666
rect 3729 54506 3781 54558
rect 3729 54398 3781 54450
rect 3729 54290 3781 54342
rect 3729 54182 3781 54234
rect 3729 54074 3781 54126
rect 3729 53966 3781 54018
rect 3729 53858 3781 53910
rect 3729 53750 3781 53802
rect 3729 53642 3781 53694
rect 3729 53534 3781 53586
rect 3729 53426 3781 53478
rect 3729 53318 3781 53370
rect 978 53215 1030 53224
rect 1102 53215 1154 53224
rect 1226 53215 1278 53224
rect 3729 53215 3781 53262
rect 978 53172 1030 53215
rect 1102 53172 1154 53215
rect 1226 53172 1278 53215
rect 3729 53210 3781 53215
rect 6335 56234 6387 56281
rect 8677 56281 8729 56286
rect 6335 56126 6387 56178
rect 6335 56018 6387 56070
rect 6335 55910 6387 55962
rect 6335 55802 6387 55854
rect 6335 55694 6387 55746
rect 6335 55586 6387 55638
rect 6335 55478 6387 55530
rect 6335 55370 6387 55422
rect 6335 55262 6387 55314
rect 6335 55154 6387 55206
rect 6335 55046 6387 55098
rect 6335 54938 6387 54990
rect 6335 54830 6387 54882
rect 6335 54722 6387 54774
rect 6335 54614 6387 54666
rect 6335 54506 6387 54558
rect 6335 54398 6387 54450
rect 6335 54290 6387 54342
rect 6335 54182 6387 54234
rect 6335 54074 6387 54126
rect 6335 53966 6387 54018
rect 6335 53858 6387 53910
rect 6335 53750 6387 53802
rect 6335 53642 6387 53694
rect 6335 53534 6387 53586
rect 6335 53426 6387 53478
rect 6335 53318 6387 53370
rect 6335 53215 6387 53262
rect 6335 53210 6387 53215
rect 7388 56211 7440 56232
rect 7388 56180 7389 56211
rect 7389 56180 7440 56211
rect 7624 56211 7676 56232
rect 7624 56180 7675 56211
rect 7675 56180 7676 56211
rect 7388 56072 7389 56124
rect 7389 56072 7440 56124
rect 7624 56072 7675 56124
rect 7675 56072 7676 56124
rect 7388 55964 7389 56016
rect 7389 55964 7440 56016
rect 7624 55964 7675 56016
rect 7675 55964 7676 56016
rect 7388 55856 7389 55908
rect 7389 55856 7440 55908
rect 7624 55856 7675 55908
rect 7675 55856 7676 55908
rect 7388 55748 7389 55800
rect 7389 55748 7440 55800
rect 7624 55748 7675 55800
rect 7675 55748 7676 55800
rect 7388 55640 7389 55692
rect 7389 55640 7440 55692
rect 7624 55640 7675 55692
rect 7675 55640 7676 55692
rect 7388 55532 7389 55584
rect 7389 55532 7440 55584
rect 7624 55532 7675 55584
rect 7675 55532 7676 55584
rect 7388 55424 7389 55476
rect 7389 55424 7440 55476
rect 7624 55424 7675 55476
rect 7675 55424 7676 55476
rect 7388 55316 7389 55368
rect 7389 55316 7440 55368
rect 7624 55316 7675 55368
rect 7675 55316 7676 55368
rect 7388 55208 7389 55260
rect 7389 55208 7440 55260
rect 7624 55208 7675 55260
rect 7675 55208 7676 55260
rect 7388 55100 7389 55152
rect 7389 55100 7440 55152
rect 7624 55100 7675 55152
rect 7675 55100 7676 55152
rect 7388 54992 7389 55044
rect 7389 54992 7440 55044
rect 7624 54992 7675 55044
rect 7675 54992 7676 55044
rect 7388 54884 7389 54936
rect 7389 54884 7440 54936
rect 7624 54884 7675 54936
rect 7675 54884 7676 54936
rect 7388 54776 7389 54828
rect 7389 54776 7440 54828
rect 7624 54776 7675 54828
rect 7675 54776 7676 54828
rect 7388 54668 7389 54720
rect 7389 54668 7440 54720
rect 7624 54668 7675 54720
rect 7675 54668 7676 54720
rect 7388 54560 7389 54612
rect 7389 54560 7440 54612
rect 7624 54560 7675 54612
rect 7675 54560 7676 54612
rect 7388 54452 7389 54504
rect 7389 54452 7440 54504
rect 7624 54452 7675 54504
rect 7675 54452 7676 54504
rect 7388 54344 7389 54396
rect 7389 54344 7440 54396
rect 7624 54344 7675 54396
rect 7675 54344 7676 54396
rect 7388 54236 7389 54288
rect 7389 54236 7440 54288
rect 7624 54236 7675 54288
rect 7675 54236 7676 54288
rect 7388 54128 7389 54180
rect 7389 54128 7440 54180
rect 7624 54128 7675 54180
rect 7675 54128 7676 54180
rect 7388 54020 7389 54072
rect 7389 54020 7440 54072
rect 7624 54020 7675 54072
rect 7675 54020 7676 54072
rect 7388 53912 7389 53964
rect 7389 53912 7440 53964
rect 7624 53912 7675 53964
rect 7675 53912 7676 53964
rect 7388 53804 7389 53856
rect 7389 53804 7440 53856
rect 7624 53804 7675 53856
rect 7675 53804 7676 53856
rect 7388 53696 7389 53748
rect 7389 53696 7440 53748
rect 7624 53696 7675 53748
rect 7675 53696 7676 53748
rect 7388 53588 7389 53640
rect 7389 53588 7440 53640
rect 7624 53588 7675 53640
rect 7675 53588 7676 53640
rect 7388 53480 7389 53532
rect 7389 53480 7440 53532
rect 7624 53480 7675 53532
rect 7675 53480 7676 53532
rect 7388 53372 7389 53424
rect 7389 53372 7440 53424
rect 7624 53372 7675 53424
rect 7675 53372 7676 53424
rect 7388 53285 7389 53316
rect 7389 53285 7440 53316
rect 7388 53264 7440 53285
rect 7624 53285 7675 53316
rect 7675 53285 7676 53316
rect 7624 53264 7676 53285
rect 8677 56234 8729 56281
rect 8677 56126 8729 56178
rect 8677 56018 8729 56070
rect 8677 55910 8729 55962
rect 8677 55802 8729 55854
rect 8677 55694 8729 55746
rect 8677 55586 8729 55638
rect 8677 55478 8729 55530
rect 8677 55370 8729 55422
rect 8677 55262 8729 55314
rect 8677 55154 8729 55206
rect 8677 55046 8729 55098
rect 8677 54938 8729 54990
rect 8677 54830 8729 54882
rect 8677 54722 8729 54774
rect 8677 54614 8729 54666
rect 8677 54506 8729 54558
rect 8677 54398 8729 54450
rect 8677 54290 8729 54342
rect 8677 54182 8729 54234
rect 8677 54074 8729 54126
rect 8677 53966 8729 54018
rect 8677 53858 8729 53910
rect 8677 53750 8729 53802
rect 8677 53642 8729 53694
rect 8677 53534 8729 53586
rect 8677 53426 8729 53478
rect 8677 53318 8729 53370
rect 8677 53215 8729 53262
rect 11283 56281 11335 56286
rect 13786 56281 13838 56324
rect 13910 56281 13962 56324
rect 14034 56281 14086 56324
rect 8677 53210 8729 53215
rect 11283 56234 11335 56281
rect 13786 56272 13838 56281
rect 13910 56272 13962 56281
rect 14034 56272 14086 56281
rect 11283 56126 11335 56178
rect 11283 56018 11335 56070
rect 11283 55910 11335 55962
rect 11283 55802 11335 55854
rect 11283 55694 11335 55746
rect 11283 55586 11335 55638
rect 11283 55478 11335 55530
rect 11283 55370 11335 55422
rect 11283 55262 11335 55314
rect 11283 55154 11335 55206
rect 11283 55046 11335 55098
rect 11283 54938 11335 54990
rect 11283 54830 11335 54882
rect 11283 54722 11335 54774
rect 11283 54614 11335 54666
rect 11283 54506 11335 54558
rect 11283 54398 11335 54450
rect 11283 54290 11335 54342
rect 11283 54182 11335 54234
rect 11283 54074 11335 54126
rect 11283 53966 11335 54018
rect 11283 53858 11335 53910
rect 11283 53750 11335 53802
rect 11283 53642 11335 53694
rect 11283 53534 11335 53586
rect 11283 53426 11335 53478
rect 11283 53318 11335 53370
rect 11283 53215 11335 53262
rect 13786 56148 13838 56200
rect 13910 56148 13962 56200
rect 14034 56148 14086 56200
rect 13786 56024 13838 56076
rect 13910 56024 13962 56076
rect 14034 56024 14086 56076
rect 13786 55900 13838 55952
rect 13910 55900 13962 55952
rect 14034 55900 14086 55952
rect 13786 55776 13838 55828
rect 13910 55776 13962 55828
rect 14034 55776 14086 55828
rect 13786 55652 13838 55704
rect 13910 55652 13962 55704
rect 14034 55652 14086 55704
rect 13786 55528 13838 55580
rect 13910 55528 13962 55580
rect 14034 55528 14086 55580
rect 13786 55404 13838 55456
rect 13910 55404 13962 55456
rect 14034 55404 14086 55456
rect 13786 55280 13838 55332
rect 13910 55280 13962 55332
rect 14034 55280 14086 55332
rect 13786 55156 13838 55208
rect 13910 55156 13962 55208
rect 14034 55156 14086 55208
rect 13786 55032 13838 55084
rect 13910 55032 13962 55084
rect 14034 55032 14086 55084
rect 13786 54908 13838 54960
rect 13910 54908 13962 54960
rect 14034 54908 14086 54960
rect 13786 54784 13838 54836
rect 13910 54784 13962 54836
rect 14034 54784 14086 54836
rect 13786 54660 13838 54712
rect 13910 54660 13962 54712
rect 14034 54660 14086 54712
rect 13786 54536 13838 54588
rect 13910 54536 13962 54588
rect 14034 54536 14086 54588
rect 13786 54412 13838 54464
rect 13910 54412 13962 54464
rect 14034 54412 14086 54464
rect 13786 54288 13838 54340
rect 13910 54288 13962 54340
rect 14034 54288 14086 54340
rect 13786 54164 13838 54216
rect 13910 54164 13962 54216
rect 14034 54164 14086 54216
rect 13786 54040 13838 54092
rect 13910 54040 13962 54092
rect 14034 54040 14086 54092
rect 13786 53916 13838 53968
rect 13910 53916 13962 53968
rect 14034 53916 14086 53968
rect 13786 53792 13838 53844
rect 13910 53792 13962 53844
rect 14034 53792 14086 53844
rect 13786 53668 13838 53720
rect 13910 53668 13962 53720
rect 14034 53668 14086 53720
rect 13786 53544 13838 53596
rect 13910 53544 13962 53596
rect 14034 53544 14086 53596
rect 13786 53420 13838 53472
rect 13910 53420 13962 53472
rect 14034 53420 14086 53472
rect 13786 53296 13838 53348
rect 13910 53296 13962 53348
rect 14034 53296 14086 53348
rect 13786 53215 13838 53224
rect 13910 53215 13962 53224
rect 14034 53215 14086 53224
rect 11283 53210 11335 53215
rect 13786 53172 13838 53215
rect 13910 53172 13962 53215
rect 14034 53172 14086 53215
rect 444 52964 445 53016
rect 445 52964 496 53016
rect 552 52964 604 53016
rect 660 52964 712 53016
rect 1438 52996 1490 53048
rect 1562 52996 1614 53048
rect 1686 52996 1738 53048
rect 1810 52996 1862 53048
rect 2574 52996 2626 53048
rect 2698 52996 2750 53048
rect 2822 52996 2874 53048
rect 2946 52996 2998 53048
rect 4846 52996 4898 53048
rect 4970 52996 5022 53048
rect 5094 52996 5146 53048
rect 5218 52996 5270 53048
rect 7139 52996 7191 53048
rect 7263 52996 7315 53048
rect 7387 52996 7439 53048
rect 7625 52996 7677 53048
rect 7749 52996 7801 53048
rect 7873 52996 7925 53048
rect 9794 52996 9846 53048
rect 9918 52996 9970 53048
rect 10042 52996 10094 53048
rect 10166 52996 10218 53048
rect 12066 52996 12118 53048
rect 12190 52996 12242 53048
rect 12314 52996 12366 53048
rect 12438 52996 12490 53048
rect 13202 52996 13254 53048
rect 13326 52996 13378 53048
rect 13450 52996 13502 53048
rect 13574 52996 13626 53048
rect 14352 52964 14404 53016
rect 14460 52964 14512 53016
rect 14568 52964 14619 53016
rect 14619 52964 14620 53016
rect 444 52856 445 52908
rect 445 52856 496 52908
rect 552 52856 604 52908
rect 660 52856 712 52908
rect 1438 52872 1490 52924
rect 1562 52872 1614 52924
rect 1686 52872 1738 52924
rect 1810 52872 1862 52924
rect 2574 52872 2626 52924
rect 2698 52872 2750 52924
rect 2822 52872 2874 52924
rect 2946 52872 2998 52924
rect 4846 52872 4898 52924
rect 4970 52872 5022 52924
rect 5094 52872 5146 52924
rect 5218 52872 5270 52924
rect 7139 52872 7191 52924
rect 7263 52872 7315 52924
rect 7387 52872 7439 52924
rect 7625 52872 7677 52924
rect 7749 52872 7801 52924
rect 7873 52872 7925 52924
rect 9794 52872 9846 52924
rect 9918 52872 9970 52924
rect 10042 52872 10094 52924
rect 10166 52872 10218 52924
rect 12066 52872 12118 52924
rect 12190 52872 12242 52924
rect 12314 52872 12366 52924
rect 12438 52872 12490 52924
rect 13202 52872 13254 52924
rect 13326 52872 13378 52924
rect 13450 52872 13502 52924
rect 13574 52872 13626 52924
rect 14352 52856 14404 52908
rect 14460 52856 14512 52908
rect 14568 52856 14619 52908
rect 14619 52856 14620 52908
rect 444 52748 445 52800
rect 445 52748 496 52800
rect 552 52797 604 52800
rect 660 52797 712 52800
rect 1438 52797 1490 52800
rect 1562 52797 1614 52800
rect 1686 52797 1738 52800
rect 1810 52797 1862 52800
rect 2574 52797 2626 52800
rect 2698 52797 2750 52800
rect 2822 52797 2874 52800
rect 2946 52797 2998 52800
rect 4846 52797 4898 52800
rect 4970 52797 5022 52800
rect 5094 52797 5146 52800
rect 5218 52797 5270 52800
rect 7139 52797 7191 52800
rect 7263 52797 7315 52800
rect 7387 52797 7439 52800
rect 7625 52797 7677 52800
rect 7749 52797 7801 52800
rect 7873 52797 7925 52800
rect 9794 52797 9846 52800
rect 9918 52797 9970 52800
rect 10042 52797 10094 52800
rect 10166 52797 10218 52800
rect 12066 52797 12118 52800
rect 12190 52797 12242 52800
rect 12314 52797 12366 52800
rect 12438 52797 12490 52800
rect 13202 52797 13254 52800
rect 13326 52797 13378 52800
rect 13450 52797 13502 52800
rect 13574 52797 13626 52800
rect 14352 52797 14404 52800
rect 14460 52797 14512 52800
rect 552 52751 553 52797
rect 553 52751 604 52797
rect 660 52751 712 52797
rect 1438 52751 1490 52797
rect 1562 52751 1614 52797
rect 1686 52751 1738 52797
rect 1810 52751 1862 52797
rect 2574 52751 2626 52797
rect 2698 52751 2750 52797
rect 2822 52751 2874 52797
rect 2946 52751 2998 52797
rect 4846 52751 4898 52797
rect 4970 52751 5022 52797
rect 5094 52751 5146 52797
rect 5218 52751 5270 52797
rect 7139 52751 7191 52797
rect 7263 52751 7315 52797
rect 7387 52751 7439 52797
rect 7625 52751 7677 52797
rect 7749 52751 7801 52797
rect 7873 52751 7925 52797
rect 9794 52751 9846 52797
rect 9918 52751 9970 52797
rect 10042 52751 10094 52797
rect 10166 52751 10218 52797
rect 12066 52751 12118 52797
rect 12190 52751 12242 52797
rect 12314 52751 12366 52797
rect 12438 52751 12490 52797
rect 13202 52751 13254 52797
rect 13326 52751 13378 52797
rect 13450 52751 13502 52797
rect 13574 52751 13626 52797
rect 14352 52751 14404 52797
rect 14460 52751 14511 52797
rect 14511 52751 14512 52797
rect 552 52748 604 52751
rect 660 52748 712 52751
rect 1438 52748 1490 52751
rect 1562 52748 1614 52751
rect 1686 52748 1738 52751
rect 1810 52748 1862 52751
rect 2574 52748 2626 52751
rect 2698 52748 2750 52751
rect 2822 52748 2874 52751
rect 2946 52748 2998 52751
rect 4846 52748 4898 52751
rect 4970 52748 5022 52751
rect 5094 52748 5146 52751
rect 5218 52748 5270 52751
rect 7139 52748 7191 52751
rect 7263 52748 7315 52751
rect 7387 52748 7439 52751
rect 7625 52748 7677 52751
rect 7749 52748 7801 52751
rect 7873 52748 7925 52751
rect 9794 52748 9846 52751
rect 9918 52748 9970 52751
rect 10042 52748 10094 52751
rect 10166 52748 10218 52751
rect 12066 52748 12118 52751
rect 12190 52748 12242 52751
rect 12314 52748 12366 52751
rect 12438 52748 12490 52751
rect 13202 52748 13254 52751
rect 13326 52748 13378 52751
rect 13450 52748 13502 52751
rect 13574 52748 13626 52751
rect 14352 52748 14404 52751
rect 14460 52748 14512 52751
rect 14568 52748 14619 52800
rect 14619 52748 14620 52800
rect 444 52640 445 52692
rect 445 52640 496 52692
rect 552 52640 604 52692
rect 660 52640 712 52692
rect 1438 52624 1490 52676
rect 1562 52624 1614 52676
rect 1686 52624 1738 52676
rect 1810 52624 1862 52676
rect 2574 52624 2626 52676
rect 2698 52624 2750 52676
rect 2822 52624 2874 52676
rect 2946 52624 2998 52676
rect 4846 52624 4898 52676
rect 4970 52624 5022 52676
rect 5094 52624 5146 52676
rect 5218 52624 5270 52676
rect 7139 52624 7191 52676
rect 7263 52624 7315 52676
rect 7387 52624 7439 52676
rect 7625 52624 7677 52676
rect 7749 52624 7801 52676
rect 7873 52624 7925 52676
rect 9794 52624 9846 52676
rect 9918 52624 9970 52676
rect 10042 52624 10094 52676
rect 10166 52624 10218 52676
rect 12066 52624 12118 52676
rect 12190 52624 12242 52676
rect 12314 52624 12366 52676
rect 12438 52624 12490 52676
rect 13202 52624 13254 52676
rect 13326 52624 13378 52676
rect 13450 52624 13502 52676
rect 13574 52624 13626 52676
rect 14352 52640 14404 52692
rect 14460 52640 14512 52692
rect 14568 52640 14619 52692
rect 14619 52640 14620 52692
rect 444 52532 445 52584
rect 445 52532 496 52584
rect 552 52532 604 52584
rect 660 52532 712 52584
rect 1438 52500 1490 52552
rect 1562 52500 1614 52552
rect 1686 52500 1738 52552
rect 1810 52500 1862 52552
rect 2574 52500 2626 52552
rect 2698 52500 2750 52552
rect 2822 52500 2874 52552
rect 2946 52500 2998 52552
rect 4846 52500 4898 52552
rect 4970 52500 5022 52552
rect 5094 52500 5146 52552
rect 5218 52500 5270 52552
rect 7139 52500 7191 52552
rect 7263 52500 7315 52552
rect 7387 52500 7439 52552
rect 7625 52500 7677 52552
rect 7749 52500 7801 52552
rect 7873 52500 7925 52552
rect 9794 52500 9846 52552
rect 9918 52500 9970 52552
rect 10042 52500 10094 52552
rect 10166 52500 10218 52552
rect 12066 52500 12118 52552
rect 12190 52500 12242 52552
rect 12314 52500 12366 52552
rect 12438 52500 12490 52552
rect 13202 52500 13254 52552
rect 13326 52500 13378 52552
rect 13450 52500 13502 52552
rect 13574 52500 13626 52552
rect 14352 52532 14404 52584
rect 14460 52532 14512 52584
rect 14568 52532 14619 52584
rect 14619 52532 14620 52584
rect 1148 52333 1200 52376
rect 1272 52333 1324 52376
rect 3729 52333 3781 52338
rect 1148 52324 1200 52333
rect 1272 52324 1324 52333
rect 1148 52200 1200 52252
rect 1272 52200 1324 52252
rect 1148 52076 1200 52128
rect 1272 52076 1324 52128
rect 1148 51952 1200 52004
rect 1272 51952 1324 52004
rect 1148 51828 1200 51880
rect 1272 51828 1324 51880
rect 1148 51704 1200 51756
rect 1272 51704 1324 51756
rect 1148 51580 1200 51632
rect 1272 51580 1324 51632
rect 1148 51456 1200 51508
rect 1272 51456 1324 51508
rect 1148 51332 1200 51384
rect 1272 51332 1324 51384
rect 1148 51208 1200 51260
rect 1272 51208 1324 51260
rect 1148 51084 1200 51136
rect 1272 51084 1324 51136
rect 1148 50960 1200 51012
rect 1272 50960 1324 51012
rect 1148 50836 1200 50888
rect 1272 50836 1324 50888
rect 1148 50712 1200 50764
rect 1272 50712 1324 50764
rect 1148 50588 1200 50640
rect 1272 50588 1324 50640
rect 1148 50464 1200 50516
rect 1272 50464 1324 50516
rect 1148 50340 1200 50392
rect 1272 50340 1324 50392
rect 1148 50216 1200 50268
rect 1272 50216 1324 50268
rect 1148 50092 1200 50144
rect 1272 50092 1324 50144
rect 1148 49968 1200 50020
rect 1272 49968 1324 50020
rect 1148 49844 1200 49896
rect 1272 49844 1324 49896
rect 1148 49720 1200 49772
rect 1272 49720 1324 49772
rect 1148 49596 1200 49648
rect 1272 49596 1324 49648
rect 1148 49472 1200 49524
rect 1272 49472 1324 49524
rect 1148 49348 1200 49400
rect 1272 49348 1324 49400
rect 3729 52286 3781 52333
rect 6335 52333 6387 52338
rect 3729 52178 3781 52230
rect 3729 52070 3781 52122
rect 3729 51962 3781 52014
rect 3729 51854 3781 51906
rect 3729 51746 3781 51798
rect 3729 51638 3781 51690
rect 3729 51530 3781 51582
rect 3729 51422 3781 51474
rect 3729 51314 3781 51366
rect 3729 51206 3781 51258
rect 3729 51098 3781 51150
rect 3729 50990 3781 51042
rect 3729 50882 3781 50934
rect 3729 50774 3781 50826
rect 3729 50666 3781 50718
rect 3729 50558 3781 50610
rect 3729 50450 3781 50502
rect 3729 50342 3781 50394
rect 3729 50234 3781 50286
rect 3729 50126 3781 50178
rect 3729 50018 3781 50070
rect 3729 49910 3781 49962
rect 3729 49802 3781 49854
rect 3729 49694 3781 49746
rect 3729 49586 3781 49638
rect 3729 49478 3781 49530
rect 3729 49370 3781 49422
rect 1148 49267 1200 49276
rect 1272 49267 1324 49276
rect 3729 49267 3781 49314
rect 1148 49224 1200 49267
rect 1272 49224 1324 49267
rect 3729 49262 3781 49267
rect 6335 52286 6387 52333
rect 8677 52333 8729 52338
rect 6335 52178 6387 52230
rect 6335 52070 6387 52122
rect 6335 51962 6387 52014
rect 6335 51854 6387 51906
rect 6335 51746 6387 51798
rect 6335 51638 6387 51690
rect 6335 51530 6387 51582
rect 6335 51422 6387 51474
rect 6335 51314 6387 51366
rect 6335 51206 6387 51258
rect 6335 51098 6387 51150
rect 6335 50990 6387 51042
rect 6335 50882 6387 50934
rect 6335 50774 6387 50826
rect 6335 50666 6387 50718
rect 6335 50558 6387 50610
rect 6335 50450 6387 50502
rect 6335 50342 6387 50394
rect 6335 50234 6387 50286
rect 6335 50126 6387 50178
rect 6335 50018 6387 50070
rect 6335 49910 6387 49962
rect 6335 49802 6387 49854
rect 6335 49694 6387 49746
rect 6335 49586 6387 49638
rect 6335 49478 6387 49530
rect 6335 49370 6387 49422
rect 6335 49267 6387 49314
rect 6335 49262 6387 49267
rect 7388 52263 7440 52284
rect 7388 52232 7389 52263
rect 7389 52232 7440 52263
rect 7624 52263 7676 52284
rect 7624 52232 7675 52263
rect 7675 52232 7676 52263
rect 7388 52124 7389 52176
rect 7389 52124 7440 52176
rect 7624 52124 7675 52176
rect 7675 52124 7676 52176
rect 7388 52016 7389 52068
rect 7389 52016 7440 52068
rect 7624 52016 7675 52068
rect 7675 52016 7676 52068
rect 7388 51908 7389 51960
rect 7389 51908 7440 51960
rect 7624 51908 7675 51960
rect 7675 51908 7676 51960
rect 7388 51800 7389 51852
rect 7389 51800 7440 51852
rect 7624 51800 7675 51852
rect 7675 51800 7676 51852
rect 7388 51692 7389 51744
rect 7389 51692 7440 51744
rect 7624 51692 7675 51744
rect 7675 51692 7676 51744
rect 7388 51584 7389 51636
rect 7389 51584 7440 51636
rect 7624 51584 7675 51636
rect 7675 51584 7676 51636
rect 7388 51476 7389 51528
rect 7389 51476 7440 51528
rect 7624 51476 7675 51528
rect 7675 51476 7676 51528
rect 7388 51368 7389 51420
rect 7389 51368 7440 51420
rect 7624 51368 7675 51420
rect 7675 51368 7676 51420
rect 7388 51260 7389 51312
rect 7389 51260 7440 51312
rect 7624 51260 7675 51312
rect 7675 51260 7676 51312
rect 7388 51152 7389 51204
rect 7389 51152 7440 51204
rect 7624 51152 7675 51204
rect 7675 51152 7676 51204
rect 7388 51044 7389 51096
rect 7389 51044 7440 51096
rect 7624 51044 7675 51096
rect 7675 51044 7676 51096
rect 7388 50936 7389 50988
rect 7389 50936 7440 50988
rect 7624 50936 7675 50988
rect 7675 50936 7676 50988
rect 7388 50828 7389 50880
rect 7389 50828 7440 50880
rect 7624 50828 7675 50880
rect 7675 50828 7676 50880
rect 7388 50720 7389 50772
rect 7389 50720 7440 50772
rect 7624 50720 7675 50772
rect 7675 50720 7676 50772
rect 7388 50612 7389 50664
rect 7389 50612 7440 50664
rect 7624 50612 7675 50664
rect 7675 50612 7676 50664
rect 7388 50504 7389 50556
rect 7389 50504 7440 50556
rect 7624 50504 7675 50556
rect 7675 50504 7676 50556
rect 7388 50396 7389 50448
rect 7389 50396 7440 50448
rect 7624 50396 7675 50448
rect 7675 50396 7676 50448
rect 7388 50288 7389 50340
rect 7389 50288 7440 50340
rect 7624 50288 7675 50340
rect 7675 50288 7676 50340
rect 7388 50180 7389 50232
rect 7389 50180 7440 50232
rect 7624 50180 7675 50232
rect 7675 50180 7676 50232
rect 7388 50072 7389 50124
rect 7389 50072 7440 50124
rect 7624 50072 7675 50124
rect 7675 50072 7676 50124
rect 7388 49964 7389 50016
rect 7389 49964 7440 50016
rect 7624 49964 7675 50016
rect 7675 49964 7676 50016
rect 7388 49856 7389 49908
rect 7389 49856 7440 49908
rect 7624 49856 7675 49908
rect 7675 49856 7676 49908
rect 7388 49748 7389 49800
rect 7389 49748 7440 49800
rect 7624 49748 7675 49800
rect 7675 49748 7676 49800
rect 7388 49640 7389 49692
rect 7389 49640 7440 49692
rect 7624 49640 7675 49692
rect 7675 49640 7676 49692
rect 7388 49532 7389 49584
rect 7389 49532 7440 49584
rect 7624 49532 7675 49584
rect 7675 49532 7676 49584
rect 7388 49424 7389 49476
rect 7389 49424 7440 49476
rect 7624 49424 7675 49476
rect 7675 49424 7676 49476
rect 7388 49337 7389 49368
rect 7389 49337 7440 49368
rect 7388 49316 7440 49337
rect 7624 49337 7675 49368
rect 7675 49337 7676 49368
rect 7624 49316 7676 49337
rect 8677 52286 8729 52333
rect 8677 52178 8729 52230
rect 8677 52070 8729 52122
rect 8677 51962 8729 52014
rect 8677 51854 8729 51906
rect 8677 51746 8729 51798
rect 8677 51638 8729 51690
rect 8677 51530 8729 51582
rect 8677 51422 8729 51474
rect 8677 51314 8729 51366
rect 8677 51206 8729 51258
rect 8677 51098 8729 51150
rect 8677 50990 8729 51042
rect 8677 50882 8729 50934
rect 8677 50774 8729 50826
rect 8677 50666 8729 50718
rect 8677 50558 8729 50610
rect 8677 50450 8729 50502
rect 8677 50342 8729 50394
rect 8677 50234 8729 50286
rect 8677 50126 8729 50178
rect 8677 50018 8729 50070
rect 8677 49910 8729 49962
rect 8677 49802 8729 49854
rect 8677 49694 8729 49746
rect 8677 49586 8729 49638
rect 8677 49478 8729 49530
rect 8677 49370 8729 49422
rect 8677 49267 8729 49314
rect 11283 52333 11335 52338
rect 13786 52333 13838 52376
rect 13910 52333 13962 52376
rect 14034 52333 14086 52376
rect 8677 49262 8729 49267
rect 11283 52286 11335 52333
rect 13786 52324 13838 52333
rect 13910 52324 13962 52333
rect 14034 52324 14086 52333
rect 11283 52178 11335 52230
rect 11283 52070 11335 52122
rect 11283 51962 11335 52014
rect 11283 51854 11335 51906
rect 11283 51746 11335 51798
rect 11283 51638 11335 51690
rect 11283 51530 11335 51582
rect 11283 51422 11335 51474
rect 11283 51314 11335 51366
rect 11283 51206 11335 51258
rect 11283 51098 11335 51150
rect 11283 50990 11335 51042
rect 11283 50882 11335 50934
rect 11283 50774 11335 50826
rect 11283 50666 11335 50718
rect 11283 50558 11335 50610
rect 11283 50450 11335 50502
rect 11283 50342 11335 50394
rect 11283 50234 11335 50286
rect 11283 50126 11335 50178
rect 11283 50018 11335 50070
rect 11283 49910 11335 49962
rect 11283 49802 11335 49854
rect 11283 49694 11335 49746
rect 11283 49586 11335 49638
rect 11283 49478 11335 49530
rect 11283 49370 11335 49422
rect 11283 49267 11335 49314
rect 13786 52200 13838 52252
rect 13910 52200 13962 52252
rect 14034 52200 14086 52252
rect 13786 52076 13838 52128
rect 13910 52076 13962 52128
rect 14034 52076 14086 52128
rect 13786 51952 13838 52004
rect 13910 51952 13962 52004
rect 14034 51952 14086 52004
rect 13786 51828 13838 51880
rect 13910 51828 13962 51880
rect 14034 51828 14086 51880
rect 13786 51704 13838 51756
rect 13910 51704 13962 51756
rect 14034 51704 14086 51756
rect 13786 51580 13838 51632
rect 13910 51580 13962 51632
rect 14034 51580 14086 51632
rect 13786 51456 13838 51508
rect 13910 51456 13962 51508
rect 14034 51456 14086 51508
rect 13786 51332 13838 51384
rect 13910 51332 13962 51384
rect 14034 51332 14086 51384
rect 13786 51208 13838 51260
rect 13910 51208 13962 51260
rect 14034 51208 14086 51260
rect 13786 51084 13838 51136
rect 13910 51084 13962 51136
rect 14034 51084 14086 51136
rect 13786 50960 13838 51012
rect 13910 50960 13962 51012
rect 14034 50960 14086 51012
rect 13786 50836 13838 50888
rect 13910 50836 13962 50888
rect 14034 50836 14086 50888
rect 13786 50712 13838 50764
rect 13910 50712 13962 50764
rect 14034 50712 14086 50764
rect 13786 50588 13838 50640
rect 13910 50588 13962 50640
rect 14034 50588 14086 50640
rect 13786 50464 13838 50516
rect 13910 50464 13962 50516
rect 14034 50464 14086 50516
rect 13786 50340 13838 50392
rect 13910 50340 13962 50392
rect 14034 50340 14086 50392
rect 13786 50216 13838 50268
rect 13910 50216 13962 50268
rect 14034 50216 14086 50268
rect 13786 50092 13838 50144
rect 13910 50092 13962 50144
rect 14034 50092 14086 50144
rect 13786 49968 13838 50020
rect 13910 49968 13962 50020
rect 14034 49968 14086 50020
rect 13786 49844 13838 49896
rect 13910 49844 13962 49896
rect 14034 49844 14086 49896
rect 13786 49720 13838 49772
rect 13910 49720 13962 49772
rect 14034 49720 14086 49772
rect 13786 49596 13838 49648
rect 13910 49596 13962 49648
rect 14034 49596 14086 49648
rect 13786 49472 13838 49524
rect 13910 49472 13962 49524
rect 14034 49472 14086 49524
rect 13786 49348 13838 49400
rect 13910 49348 13962 49400
rect 14034 49348 14086 49400
rect 13786 49267 13838 49276
rect 13910 49267 13962 49276
rect 14034 49267 14086 49276
rect 11283 49262 11335 49267
rect 13786 49224 13838 49267
rect 13910 49224 13962 49267
rect 14034 49224 14086 49267
rect 444 49016 445 49068
rect 445 49016 496 49068
rect 552 49016 604 49068
rect 660 49016 712 49068
rect 1438 49048 1490 49100
rect 1562 49048 1614 49100
rect 1686 49048 1738 49100
rect 1810 49048 1862 49100
rect 2574 49048 2626 49100
rect 2698 49048 2750 49100
rect 2822 49048 2874 49100
rect 2946 49048 2998 49100
rect 4846 49048 4898 49100
rect 4970 49048 5022 49100
rect 5094 49048 5146 49100
rect 5218 49048 5270 49100
rect 7139 49048 7191 49100
rect 7263 49048 7315 49100
rect 7387 49048 7439 49100
rect 7625 49048 7677 49100
rect 7749 49048 7801 49100
rect 7873 49048 7925 49100
rect 9794 49048 9846 49100
rect 9918 49048 9970 49100
rect 10042 49048 10094 49100
rect 10166 49048 10218 49100
rect 12066 49048 12118 49100
rect 12190 49048 12242 49100
rect 12314 49048 12366 49100
rect 12438 49048 12490 49100
rect 13480 49048 13532 49100
rect 13604 49048 13656 49100
rect 14352 49016 14404 49068
rect 14460 49016 14512 49068
rect 14568 49016 14619 49068
rect 14619 49016 14620 49068
rect 444 48908 445 48960
rect 445 48908 496 48960
rect 552 48908 604 48960
rect 660 48908 712 48960
rect 1438 48924 1490 48976
rect 1562 48924 1614 48976
rect 1686 48924 1738 48976
rect 1810 48924 1862 48976
rect 2574 48924 2626 48976
rect 2698 48924 2750 48976
rect 2822 48924 2874 48976
rect 2946 48924 2998 48976
rect 4846 48924 4898 48976
rect 4970 48924 5022 48976
rect 5094 48924 5146 48976
rect 5218 48924 5270 48976
rect 7139 48924 7191 48976
rect 7263 48924 7315 48976
rect 7387 48924 7439 48976
rect 7625 48924 7677 48976
rect 7749 48924 7801 48976
rect 7873 48924 7925 48976
rect 9794 48924 9846 48976
rect 9918 48924 9970 48976
rect 10042 48924 10094 48976
rect 10166 48924 10218 48976
rect 12066 48924 12118 48976
rect 12190 48924 12242 48976
rect 12314 48924 12366 48976
rect 12438 48924 12490 48976
rect 13480 48924 13532 48976
rect 13604 48924 13656 48976
rect 14352 48908 14404 48960
rect 14460 48908 14512 48960
rect 14568 48908 14619 48960
rect 14619 48908 14620 48960
rect 444 48800 445 48852
rect 445 48800 496 48852
rect 552 48849 604 48852
rect 660 48849 712 48852
rect 1438 48849 1490 48852
rect 1562 48849 1614 48852
rect 1686 48849 1738 48852
rect 1810 48849 1862 48852
rect 2574 48849 2626 48852
rect 2698 48849 2750 48852
rect 2822 48849 2874 48852
rect 2946 48849 2998 48852
rect 4846 48849 4898 48852
rect 4970 48849 5022 48852
rect 5094 48849 5146 48852
rect 5218 48849 5270 48852
rect 7139 48849 7191 48852
rect 7263 48849 7315 48852
rect 7387 48849 7439 48852
rect 7625 48849 7677 48852
rect 7749 48849 7801 48852
rect 7873 48849 7925 48852
rect 9794 48849 9846 48852
rect 9918 48849 9970 48852
rect 10042 48849 10094 48852
rect 10166 48849 10218 48852
rect 12066 48849 12118 48852
rect 12190 48849 12242 48852
rect 12314 48849 12366 48852
rect 12438 48849 12490 48852
rect 13480 48849 13532 48852
rect 13604 48849 13656 48852
rect 14352 48849 14404 48852
rect 14460 48849 14512 48852
rect 552 48803 553 48849
rect 553 48803 604 48849
rect 660 48803 712 48849
rect 1438 48803 1490 48849
rect 1562 48803 1614 48849
rect 1686 48803 1738 48849
rect 1810 48803 1862 48849
rect 2574 48803 2626 48849
rect 2698 48803 2750 48849
rect 2822 48803 2874 48849
rect 2946 48803 2998 48849
rect 4846 48803 4898 48849
rect 4970 48803 5022 48849
rect 5094 48803 5146 48849
rect 5218 48803 5270 48849
rect 7139 48803 7191 48849
rect 7263 48803 7315 48849
rect 7387 48803 7439 48849
rect 7625 48803 7677 48849
rect 7749 48803 7801 48849
rect 7873 48803 7925 48849
rect 9794 48803 9846 48849
rect 9918 48803 9970 48849
rect 10042 48803 10094 48849
rect 10166 48803 10218 48849
rect 12066 48803 12118 48849
rect 12190 48803 12242 48849
rect 12314 48803 12366 48849
rect 12438 48803 12490 48849
rect 13480 48803 13532 48849
rect 13604 48803 13656 48849
rect 14352 48803 14404 48849
rect 14460 48803 14511 48849
rect 14511 48803 14512 48849
rect 552 48800 604 48803
rect 660 48800 712 48803
rect 1438 48800 1490 48803
rect 1562 48800 1614 48803
rect 1686 48800 1738 48803
rect 1810 48800 1862 48803
rect 2574 48800 2626 48803
rect 2698 48800 2750 48803
rect 2822 48800 2874 48803
rect 2946 48800 2998 48803
rect 4846 48800 4898 48803
rect 4970 48800 5022 48803
rect 5094 48800 5146 48803
rect 5218 48800 5270 48803
rect 7139 48800 7191 48803
rect 7263 48800 7315 48803
rect 7387 48800 7439 48803
rect 7625 48800 7677 48803
rect 7749 48800 7801 48803
rect 7873 48800 7925 48803
rect 9794 48800 9846 48803
rect 9918 48800 9970 48803
rect 10042 48800 10094 48803
rect 10166 48800 10218 48803
rect 12066 48800 12118 48803
rect 12190 48800 12242 48803
rect 12314 48800 12366 48803
rect 12438 48800 12490 48803
rect 13480 48800 13532 48803
rect 13604 48800 13656 48803
rect 14352 48800 14404 48803
rect 14460 48800 14512 48803
rect 14568 48800 14619 48852
rect 14619 48800 14620 48852
rect 444 48692 445 48744
rect 445 48692 496 48744
rect 552 48692 604 48744
rect 660 48692 712 48744
rect 1438 48676 1490 48728
rect 1562 48676 1614 48728
rect 1686 48676 1738 48728
rect 1810 48676 1862 48728
rect 2574 48676 2626 48728
rect 2698 48676 2750 48728
rect 2822 48676 2874 48728
rect 2946 48676 2998 48728
rect 4846 48676 4898 48728
rect 4970 48676 5022 48728
rect 5094 48676 5146 48728
rect 5218 48676 5270 48728
rect 7139 48676 7191 48728
rect 7263 48676 7315 48728
rect 7387 48676 7439 48728
rect 7625 48676 7677 48728
rect 7749 48676 7801 48728
rect 7873 48676 7925 48728
rect 9794 48676 9846 48728
rect 9918 48676 9970 48728
rect 10042 48676 10094 48728
rect 10166 48676 10218 48728
rect 12066 48676 12118 48728
rect 12190 48676 12242 48728
rect 12314 48676 12366 48728
rect 12438 48676 12490 48728
rect 13480 48676 13532 48728
rect 13604 48676 13656 48728
rect 14352 48692 14404 48744
rect 14460 48692 14512 48744
rect 14568 48692 14619 48744
rect 14619 48692 14620 48744
rect 444 48584 445 48636
rect 445 48584 496 48636
rect 552 48584 604 48636
rect 660 48584 712 48636
rect 1438 48552 1490 48604
rect 1562 48552 1614 48604
rect 1686 48552 1738 48604
rect 1810 48552 1862 48604
rect 2574 48552 2626 48604
rect 2698 48552 2750 48604
rect 2822 48552 2874 48604
rect 2946 48552 2998 48604
rect 4846 48552 4898 48604
rect 4970 48552 5022 48604
rect 5094 48552 5146 48604
rect 5218 48552 5270 48604
rect 7139 48552 7191 48604
rect 7263 48552 7315 48604
rect 7387 48552 7439 48604
rect 7625 48552 7677 48604
rect 7749 48552 7801 48604
rect 7873 48552 7925 48604
rect 9794 48552 9846 48604
rect 9918 48552 9970 48604
rect 10042 48552 10094 48604
rect 10166 48552 10218 48604
rect 12066 48552 12118 48604
rect 12190 48552 12242 48604
rect 12314 48552 12366 48604
rect 12438 48552 12490 48604
rect 13480 48552 13532 48604
rect 13604 48552 13656 48604
rect 14352 48584 14404 48636
rect 14460 48584 14512 48636
rect 14568 48584 14619 48636
rect 14619 48584 14620 48636
rect 1148 48385 1200 48428
rect 1272 48385 1324 48428
rect 3729 48385 3781 48390
rect 1148 48376 1200 48385
rect 1272 48376 1324 48385
rect 1148 48252 1200 48304
rect 1272 48252 1324 48304
rect 1148 48128 1200 48180
rect 1272 48128 1324 48180
rect 1148 48004 1200 48056
rect 1272 48004 1324 48056
rect 1148 47880 1200 47932
rect 1272 47880 1324 47932
rect 1148 47756 1200 47808
rect 1272 47756 1324 47808
rect 1148 47632 1200 47684
rect 1272 47632 1324 47684
rect 1148 47508 1200 47560
rect 1272 47508 1324 47560
rect 1148 47384 1200 47436
rect 1272 47384 1324 47436
rect 1148 47260 1200 47312
rect 1272 47260 1324 47312
rect 1148 47136 1200 47188
rect 1272 47136 1324 47188
rect 1148 47012 1200 47064
rect 1272 47012 1324 47064
rect 1148 46888 1200 46940
rect 1272 46888 1324 46940
rect 1148 46764 1200 46816
rect 1272 46764 1324 46816
rect 1148 46640 1200 46692
rect 1272 46640 1324 46692
rect 1148 46516 1200 46568
rect 1272 46516 1324 46568
rect 1148 46392 1200 46444
rect 1272 46392 1324 46444
rect 1148 46268 1200 46320
rect 1272 46268 1324 46320
rect 1148 46144 1200 46196
rect 1272 46144 1324 46196
rect 1148 46020 1200 46072
rect 1272 46020 1324 46072
rect 1148 45896 1200 45948
rect 1272 45896 1324 45948
rect 1148 45772 1200 45824
rect 1272 45772 1324 45824
rect 1148 45648 1200 45700
rect 1272 45648 1324 45700
rect 1148 45524 1200 45576
rect 1272 45524 1324 45576
rect 1148 45400 1200 45452
rect 1272 45400 1324 45452
rect 3729 48338 3781 48385
rect 6335 48385 6387 48390
rect 3729 48230 3781 48282
rect 3729 48122 3781 48174
rect 3729 48014 3781 48066
rect 3729 47906 3781 47958
rect 3729 47798 3781 47850
rect 3729 47690 3781 47742
rect 3729 47582 3781 47634
rect 3729 47474 3781 47526
rect 3729 47366 3781 47418
rect 3729 47258 3781 47310
rect 3729 47150 3781 47202
rect 3729 47042 3781 47094
rect 3729 46934 3781 46986
rect 3729 46826 3781 46878
rect 3729 46718 3781 46770
rect 3729 46610 3781 46662
rect 3729 46502 3781 46554
rect 3729 46394 3781 46446
rect 3729 46286 3781 46338
rect 3729 46178 3781 46230
rect 3729 46070 3781 46122
rect 3729 45962 3781 46014
rect 3729 45854 3781 45906
rect 3729 45746 3781 45798
rect 3729 45638 3781 45690
rect 3729 45530 3781 45582
rect 3729 45422 3781 45474
rect 1148 45319 1200 45328
rect 1272 45319 1324 45328
rect 3729 45319 3781 45366
rect 1148 45276 1200 45319
rect 1272 45276 1324 45319
rect 3729 45314 3781 45319
rect 6335 48338 6387 48385
rect 8677 48385 8729 48390
rect 6335 48230 6387 48282
rect 6335 48122 6387 48174
rect 6335 48014 6387 48066
rect 6335 47906 6387 47958
rect 6335 47798 6387 47850
rect 6335 47690 6387 47742
rect 6335 47582 6387 47634
rect 6335 47474 6387 47526
rect 6335 47366 6387 47418
rect 6335 47258 6387 47310
rect 6335 47150 6387 47202
rect 6335 47042 6387 47094
rect 6335 46934 6387 46986
rect 6335 46826 6387 46878
rect 6335 46718 6387 46770
rect 6335 46610 6387 46662
rect 6335 46502 6387 46554
rect 6335 46394 6387 46446
rect 6335 46286 6387 46338
rect 6335 46178 6387 46230
rect 6335 46070 6387 46122
rect 6335 45962 6387 46014
rect 6335 45854 6387 45906
rect 6335 45746 6387 45798
rect 6335 45638 6387 45690
rect 6335 45530 6387 45582
rect 6335 45422 6387 45474
rect 6335 45319 6387 45366
rect 6335 45314 6387 45319
rect 7388 48315 7440 48336
rect 7388 48284 7389 48315
rect 7389 48284 7440 48315
rect 7624 48315 7676 48336
rect 7624 48284 7675 48315
rect 7675 48284 7676 48315
rect 7388 48176 7389 48228
rect 7389 48176 7440 48228
rect 7624 48176 7675 48228
rect 7675 48176 7676 48228
rect 7388 48068 7389 48120
rect 7389 48068 7440 48120
rect 7624 48068 7675 48120
rect 7675 48068 7676 48120
rect 7388 47960 7389 48012
rect 7389 47960 7440 48012
rect 7624 47960 7675 48012
rect 7675 47960 7676 48012
rect 7388 47852 7389 47904
rect 7389 47852 7440 47904
rect 7624 47852 7675 47904
rect 7675 47852 7676 47904
rect 7388 47744 7389 47796
rect 7389 47744 7440 47796
rect 7624 47744 7675 47796
rect 7675 47744 7676 47796
rect 7388 47636 7389 47688
rect 7389 47636 7440 47688
rect 7624 47636 7675 47688
rect 7675 47636 7676 47688
rect 7388 47528 7389 47580
rect 7389 47528 7440 47580
rect 7624 47528 7675 47580
rect 7675 47528 7676 47580
rect 7388 47420 7389 47472
rect 7389 47420 7440 47472
rect 7624 47420 7675 47472
rect 7675 47420 7676 47472
rect 7388 47312 7389 47364
rect 7389 47312 7440 47364
rect 7624 47312 7675 47364
rect 7675 47312 7676 47364
rect 7388 47204 7389 47256
rect 7389 47204 7440 47256
rect 7624 47204 7675 47256
rect 7675 47204 7676 47256
rect 7388 47096 7389 47148
rect 7389 47096 7440 47148
rect 7624 47096 7675 47148
rect 7675 47096 7676 47148
rect 7388 46988 7389 47040
rect 7389 46988 7440 47040
rect 7624 46988 7675 47040
rect 7675 46988 7676 47040
rect 7388 46880 7389 46932
rect 7389 46880 7440 46932
rect 7624 46880 7675 46932
rect 7675 46880 7676 46932
rect 7388 46772 7389 46824
rect 7389 46772 7440 46824
rect 7624 46772 7675 46824
rect 7675 46772 7676 46824
rect 7388 46664 7389 46716
rect 7389 46664 7440 46716
rect 7624 46664 7675 46716
rect 7675 46664 7676 46716
rect 7388 46556 7389 46608
rect 7389 46556 7440 46608
rect 7624 46556 7675 46608
rect 7675 46556 7676 46608
rect 7388 46448 7389 46500
rect 7389 46448 7440 46500
rect 7624 46448 7675 46500
rect 7675 46448 7676 46500
rect 7388 46340 7389 46392
rect 7389 46340 7440 46392
rect 7624 46340 7675 46392
rect 7675 46340 7676 46392
rect 7388 46232 7389 46284
rect 7389 46232 7440 46284
rect 7624 46232 7675 46284
rect 7675 46232 7676 46284
rect 7388 46124 7389 46176
rect 7389 46124 7440 46176
rect 7624 46124 7675 46176
rect 7675 46124 7676 46176
rect 7388 46016 7389 46068
rect 7389 46016 7440 46068
rect 7624 46016 7675 46068
rect 7675 46016 7676 46068
rect 7388 45908 7389 45960
rect 7389 45908 7440 45960
rect 7624 45908 7675 45960
rect 7675 45908 7676 45960
rect 7388 45800 7389 45852
rect 7389 45800 7440 45852
rect 7624 45800 7675 45852
rect 7675 45800 7676 45852
rect 7388 45692 7389 45744
rect 7389 45692 7440 45744
rect 7624 45692 7675 45744
rect 7675 45692 7676 45744
rect 7388 45584 7389 45636
rect 7389 45584 7440 45636
rect 7624 45584 7675 45636
rect 7675 45584 7676 45636
rect 7388 45476 7389 45528
rect 7389 45476 7440 45528
rect 7624 45476 7675 45528
rect 7675 45476 7676 45528
rect 7388 45389 7389 45420
rect 7389 45389 7440 45420
rect 7388 45368 7440 45389
rect 7624 45389 7675 45420
rect 7675 45389 7676 45420
rect 7624 45368 7676 45389
rect 8677 48338 8729 48385
rect 8677 48230 8729 48282
rect 8677 48122 8729 48174
rect 8677 48014 8729 48066
rect 8677 47906 8729 47958
rect 8677 47798 8729 47850
rect 8677 47690 8729 47742
rect 8677 47582 8729 47634
rect 8677 47474 8729 47526
rect 8677 47366 8729 47418
rect 8677 47258 8729 47310
rect 8677 47150 8729 47202
rect 8677 47042 8729 47094
rect 8677 46934 8729 46986
rect 8677 46826 8729 46878
rect 8677 46718 8729 46770
rect 8677 46610 8729 46662
rect 8677 46502 8729 46554
rect 8677 46394 8729 46446
rect 8677 46286 8729 46338
rect 8677 46178 8729 46230
rect 8677 46070 8729 46122
rect 8677 45962 8729 46014
rect 8677 45854 8729 45906
rect 8677 45746 8729 45798
rect 8677 45638 8729 45690
rect 8677 45530 8729 45582
rect 8677 45422 8729 45474
rect 8677 45319 8729 45366
rect 11283 48385 11335 48390
rect 13786 48385 13838 48428
rect 13910 48385 13962 48428
rect 14034 48385 14086 48428
rect 8677 45314 8729 45319
rect 11283 48338 11335 48385
rect 13786 48376 13838 48385
rect 13910 48376 13962 48385
rect 14034 48376 14086 48385
rect 11283 48230 11335 48282
rect 11283 48122 11335 48174
rect 11283 48014 11335 48066
rect 11283 47906 11335 47958
rect 11283 47798 11335 47850
rect 11283 47690 11335 47742
rect 11283 47582 11335 47634
rect 11283 47474 11335 47526
rect 11283 47366 11335 47418
rect 11283 47258 11335 47310
rect 11283 47150 11335 47202
rect 11283 47042 11335 47094
rect 11283 46934 11335 46986
rect 11283 46826 11335 46878
rect 11283 46718 11335 46770
rect 11283 46610 11335 46662
rect 11283 46502 11335 46554
rect 11283 46394 11335 46446
rect 11283 46286 11335 46338
rect 11283 46178 11335 46230
rect 11283 46070 11335 46122
rect 11283 45962 11335 46014
rect 11283 45854 11335 45906
rect 11283 45746 11335 45798
rect 11283 45638 11335 45690
rect 11283 45530 11335 45582
rect 11283 45422 11335 45474
rect 11283 45319 11335 45366
rect 13786 48252 13838 48304
rect 13910 48252 13962 48304
rect 14034 48252 14086 48304
rect 13786 48128 13838 48180
rect 13910 48128 13962 48180
rect 14034 48128 14086 48180
rect 13786 48004 13838 48056
rect 13910 48004 13962 48056
rect 14034 48004 14086 48056
rect 13786 47880 13838 47932
rect 13910 47880 13962 47932
rect 14034 47880 14086 47932
rect 13786 47756 13838 47808
rect 13910 47756 13962 47808
rect 14034 47756 14086 47808
rect 13786 47632 13838 47684
rect 13910 47632 13962 47684
rect 14034 47632 14086 47684
rect 13786 47508 13838 47560
rect 13910 47508 13962 47560
rect 14034 47508 14086 47560
rect 13786 47384 13838 47436
rect 13910 47384 13962 47436
rect 14034 47384 14086 47436
rect 13786 47260 13838 47312
rect 13910 47260 13962 47312
rect 14034 47260 14086 47312
rect 13786 47136 13838 47188
rect 13910 47136 13962 47188
rect 14034 47136 14086 47188
rect 13786 47012 13838 47064
rect 13910 47012 13962 47064
rect 14034 47012 14086 47064
rect 13786 46888 13838 46940
rect 13910 46888 13962 46940
rect 14034 46888 14086 46940
rect 13786 46764 13838 46816
rect 13910 46764 13962 46816
rect 14034 46764 14086 46816
rect 13786 46640 13838 46692
rect 13910 46640 13962 46692
rect 14034 46640 14086 46692
rect 13786 46516 13838 46568
rect 13910 46516 13962 46568
rect 14034 46516 14086 46568
rect 13786 46392 13838 46444
rect 13910 46392 13962 46444
rect 14034 46392 14086 46444
rect 13786 46268 13838 46320
rect 13910 46268 13962 46320
rect 14034 46268 14086 46320
rect 13786 46144 13838 46196
rect 13910 46144 13962 46196
rect 14034 46144 14086 46196
rect 13786 46020 13838 46072
rect 13910 46020 13962 46072
rect 14034 46020 14086 46072
rect 13786 45896 13838 45948
rect 13910 45896 13962 45948
rect 14034 45896 14086 45948
rect 13786 45772 13838 45824
rect 13910 45772 13962 45824
rect 14034 45772 14086 45824
rect 13786 45648 13838 45700
rect 13910 45648 13962 45700
rect 14034 45648 14086 45700
rect 13786 45524 13838 45576
rect 13910 45524 13962 45576
rect 14034 45524 14086 45576
rect 13786 45400 13838 45452
rect 13910 45400 13962 45452
rect 14034 45400 14086 45452
rect 13786 45319 13838 45328
rect 13910 45319 13962 45328
rect 14034 45319 14086 45328
rect 11283 45314 11335 45319
rect 13786 45276 13838 45319
rect 13910 45276 13962 45319
rect 14034 45276 14086 45319
rect 444 45068 445 45120
rect 445 45068 496 45120
rect 552 45068 604 45120
rect 660 45068 712 45120
rect 1438 45100 1490 45152
rect 1562 45100 1614 45152
rect 1686 45100 1738 45152
rect 1810 45100 1862 45152
rect 2574 45100 2626 45152
rect 2698 45100 2750 45152
rect 2822 45100 2874 45152
rect 2946 45100 2998 45152
rect 4846 45100 4898 45152
rect 4970 45100 5022 45152
rect 5094 45100 5146 45152
rect 5218 45100 5270 45152
rect 7139 45100 7191 45152
rect 7263 45100 7315 45152
rect 7387 45100 7439 45152
rect 7625 45100 7677 45152
rect 7749 45100 7801 45152
rect 7873 45100 7925 45152
rect 9794 45100 9846 45152
rect 9918 45100 9970 45152
rect 10042 45100 10094 45152
rect 10166 45100 10218 45152
rect 12066 45100 12118 45152
rect 12190 45100 12242 45152
rect 12314 45100 12366 45152
rect 12438 45100 12490 45152
rect 13480 45100 13532 45152
rect 13604 45100 13656 45152
rect 14352 45068 14404 45120
rect 14460 45068 14512 45120
rect 14568 45068 14619 45120
rect 14619 45068 14620 45120
rect 444 44960 445 45012
rect 445 44960 496 45012
rect 552 44960 604 45012
rect 660 44960 712 45012
rect 1438 44976 1490 45028
rect 1562 44976 1614 45028
rect 1686 44976 1738 45028
rect 1810 44976 1862 45028
rect 2574 44976 2626 45028
rect 2698 44976 2750 45028
rect 2822 44976 2874 45028
rect 2946 44976 2998 45028
rect 4846 44976 4898 45028
rect 4970 44976 5022 45028
rect 5094 44976 5146 45028
rect 5218 44976 5270 45028
rect 7139 44976 7191 45028
rect 7263 44976 7315 45028
rect 7387 44976 7439 45028
rect 7625 44976 7677 45028
rect 7749 44976 7801 45028
rect 7873 44976 7925 45028
rect 9794 44976 9846 45028
rect 9918 44976 9970 45028
rect 10042 44976 10094 45028
rect 10166 44976 10218 45028
rect 12066 44976 12118 45028
rect 12190 44976 12242 45028
rect 12314 44976 12366 45028
rect 12438 44976 12490 45028
rect 13480 44976 13532 45028
rect 13604 44976 13656 45028
rect 14352 44960 14404 45012
rect 14460 44960 14512 45012
rect 14568 44960 14619 45012
rect 14619 44960 14620 45012
rect 444 44852 445 44904
rect 445 44852 496 44904
rect 552 44901 604 44904
rect 660 44901 712 44904
rect 1438 44901 1490 44904
rect 1562 44901 1614 44904
rect 1686 44901 1738 44904
rect 1810 44901 1862 44904
rect 2574 44901 2626 44904
rect 2698 44901 2750 44904
rect 2822 44901 2874 44904
rect 2946 44901 2998 44904
rect 4846 44901 4898 44904
rect 4970 44901 5022 44904
rect 5094 44901 5146 44904
rect 5218 44901 5270 44904
rect 7139 44901 7191 44904
rect 7263 44901 7315 44904
rect 7387 44901 7439 44904
rect 7625 44901 7677 44904
rect 7749 44901 7801 44904
rect 7873 44901 7925 44904
rect 9794 44901 9846 44904
rect 9918 44901 9970 44904
rect 10042 44901 10094 44904
rect 10166 44901 10218 44904
rect 12066 44901 12118 44904
rect 12190 44901 12242 44904
rect 12314 44901 12366 44904
rect 12438 44901 12490 44904
rect 13480 44901 13532 44904
rect 13604 44901 13656 44904
rect 14352 44901 14404 44904
rect 14460 44901 14512 44904
rect 552 44855 553 44901
rect 553 44855 604 44901
rect 660 44855 712 44901
rect 1438 44855 1490 44901
rect 1562 44855 1614 44901
rect 1686 44855 1738 44901
rect 1810 44855 1862 44901
rect 2574 44855 2626 44901
rect 2698 44855 2750 44901
rect 2822 44855 2874 44901
rect 2946 44855 2998 44901
rect 4846 44855 4898 44901
rect 4970 44855 5022 44901
rect 5094 44855 5146 44901
rect 5218 44855 5270 44901
rect 7139 44855 7191 44901
rect 7263 44855 7315 44901
rect 7387 44855 7439 44901
rect 7625 44855 7677 44901
rect 7749 44855 7801 44901
rect 7873 44855 7925 44901
rect 9794 44855 9846 44901
rect 9918 44855 9970 44901
rect 10042 44855 10094 44901
rect 10166 44855 10218 44901
rect 12066 44855 12118 44901
rect 12190 44855 12242 44901
rect 12314 44855 12366 44901
rect 12438 44855 12490 44901
rect 13480 44855 13532 44901
rect 13604 44855 13656 44901
rect 14352 44855 14404 44901
rect 14460 44855 14511 44901
rect 14511 44855 14512 44901
rect 552 44852 604 44855
rect 660 44852 712 44855
rect 1438 44852 1490 44855
rect 1562 44852 1614 44855
rect 1686 44852 1738 44855
rect 1810 44852 1862 44855
rect 2574 44852 2626 44855
rect 2698 44852 2750 44855
rect 2822 44852 2874 44855
rect 2946 44852 2998 44855
rect 4846 44852 4898 44855
rect 4970 44852 5022 44855
rect 5094 44852 5146 44855
rect 5218 44852 5270 44855
rect 7139 44852 7191 44855
rect 7263 44852 7315 44855
rect 7387 44852 7439 44855
rect 7625 44852 7677 44855
rect 7749 44852 7801 44855
rect 7873 44852 7925 44855
rect 9794 44852 9846 44855
rect 9918 44852 9970 44855
rect 10042 44852 10094 44855
rect 10166 44852 10218 44855
rect 12066 44852 12118 44855
rect 12190 44852 12242 44855
rect 12314 44852 12366 44855
rect 12438 44852 12490 44855
rect 13480 44852 13532 44855
rect 13604 44852 13656 44855
rect 14352 44852 14404 44855
rect 14460 44852 14512 44855
rect 14568 44852 14619 44904
rect 14619 44852 14620 44904
rect 444 44744 445 44796
rect 445 44744 496 44796
rect 552 44744 604 44796
rect 660 44744 712 44796
rect 1438 44728 1490 44780
rect 1562 44728 1614 44780
rect 1686 44728 1738 44780
rect 1810 44728 1862 44780
rect 2574 44728 2626 44780
rect 2698 44728 2750 44780
rect 2822 44728 2874 44780
rect 2946 44728 2998 44780
rect 4846 44728 4898 44780
rect 4970 44728 5022 44780
rect 5094 44728 5146 44780
rect 5218 44728 5270 44780
rect 7139 44728 7191 44780
rect 7263 44728 7315 44780
rect 7387 44728 7439 44780
rect 7625 44728 7677 44780
rect 7749 44728 7801 44780
rect 7873 44728 7925 44780
rect 9794 44728 9846 44780
rect 9918 44728 9970 44780
rect 10042 44728 10094 44780
rect 10166 44728 10218 44780
rect 12066 44728 12118 44780
rect 12190 44728 12242 44780
rect 12314 44728 12366 44780
rect 12438 44728 12490 44780
rect 13480 44728 13532 44780
rect 13604 44728 13656 44780
rect 14352 44744 14404 44796
rect 14460 44744 14512 44796
rect 14568 44744 14619 44796
rect 14619 44744 14620 44796
rect 444 44636 445 44688
rect 445 44636 496 44688
rect 552 44636 604 44688
rect 660 44636 712 44688
rect 1438 44604 1490 44656
rect 1562 44604 1614 44656
rect 1686 44604 1738 44656
rect 1810 44604 1862 44656
rect 2574 44604 2626 44656
rect 2698 44604 2750 44656
rect 2822 44604 2874 44656
rect 2946 44604 2998 44656
rect 4846 44604 4898 44656
rect 4970 44604 5022 44656
rect 5094 44604 5146 44656
rect 5218 44604 5270 44656
rect 7139 44604 7191 44656
rect 7263 44604 7315 44656
rect 7387 44604 7439 44656
rect 7625 44604 7677 44656
rect 7749 44604 7801 44656
rect 7873 44604 7925 44656
rect 9794 44604 9846 44656
rect 9918 44604 9970 44656
rect 10042 44604 10094 44656
rect 10166 44604 10218 44656
rect 12066 44604 12118 44656
rect 12190 44604 12242 44656
rect 12314 44604 12366 44656
rect 12438 44604 12490 44656
rect 13480 44604 13532 44656
rect 13604 44604 13656 44656
rect 14352 44636 14404 44688
rect 14460 44636 14512 44688
rect 14568 44636 14619 44688
rect 14619 44636 14620 44688
rect 1148 44437 1200 44480
rect 1272 44437 1324 44480
rect 3729 44437 3781 44442
rect 1148 44428 1200 44437
rect 1272 44428 1324 44437
rect 1148 44304 1200 44356
rect 1272 44304 1324 44356
rect 1148 44180 1200 44232
rect 1272 44180 1324 44232
rect 1148 44056 1200 44108
rect 1272 44056 1324 44108
rect 1148 43932 1200 43984
rect 1272 43932 1324 43984
rect 1148 43808 1200 43860
rect 1272 43808 1324 43860
rect 1148 43684 1200 43736
rect 1272 43684 1324 43736
rect 1148 43560 1200 43612
rect 1272 43560 1324 43612
rect 1148 43436 1200 43488
rect 1272 43436 1324 43488
rect 1148 43312 1200 43364
rect 1272 43312 1324 43364
rect 1148 43188 1200 43240
rect 1272 43188 1324 43240
rect 1148 43064 1200 43116
rect 1272 43064 1324 43116
rect 1148 42940 1200 42992
rect 1272 42940 1324 42992
rect 1148 42816 1200 42868
rect 1272 42816 1324 42868
rect 1148 42692 1200 42744
rect 1272 42692 1324 42744
rect 1148 42568 1200 42620
rect 1272 42568 1324 42620
rect 1148 42444 1200 42496
rect 1272 42444 1324 42496
rect 1148 42320 1200 42372
rect 1272 42320 1324 42372
rect 1148 42196 1200 42248
rect 1272 42196 1324 42248
rect 1148 42072 1200 42124
rect 1272 42072 1324 42124
rect 1148 41948 1200 42000
rect 1272 41948 1324 42000
rect 1148 41824 1200 41876
rect 1272 41824 1324 41876
rect 1148 41700 1200 41752
rect 1272 41700 1324 41752
rect 1148 41576 1200 41628
rect 1272 41576 1324 41628
rect 1148 41452 1200 41504
rect 1272 41452 1324 41504
rect 3729 44390 3781 44437
rect 6335 44437 6387 44442
rect 3729 44282 3781 44334
rect 3729 44174 3781 44226
rect 3729 44066 3781 44118
rect 3729 43958 3781 44010
rect 3729 43850 3781 43902
rect 3729 43742 3781 43794
rect 3729 43634 3781 43686
rect 3729 43526 3781 43578
rect 3729 43418 3781 43470
rect 3729 43310 3781 43362
rect 3729 43202 3781 43254
rect 3729 43094 3781 43146
rect 3729 42986 3781 43038
rect 3729 42878 3781 42930
rect 3729 42770 3781 42822
rect 3729 42662 3781 42714
rect 3729 42554 3781 42606
rect 3729 42446 3781 42498
rect 3729 42338 3781 42390
rect 3729 42230 3781 42282
rect 3729 42122 3781 42174
rect 3729 42014 3781 42066
rect 3729 41906 3781 41958
rect 3729 41798 3781 41850
rect 3729 41690 3781 41742
rect 3729 41582 3781 41634
rect 3729 41474 3781 41526
rect 1148 41371 1200 41380
rect 1272 41371 1324 41380
rect 3729 41371 3781 41418
rect 1148 41328 1200 41371
rect 1272 41328 1324 41371
rect 3729 41366 3781 41371
rect 6335 44390 6387 44437
rect 8677 44437 8729 44442
rect 6335 44282 6387 44334
rect 6335 44174 6387 44226
rect 6335 44066 6387 44118
rect 6335 43958 6387 44010
rect 6335 43850 6387 43902
rect 6335 43742 6387 43794
rect 6335 43634 6387 43686
rect 6335 43526 6387 43578
rect 6335 43418 6387 43470
rect 6335 43310 6387 43362
rect 6335 43202 6387 43254
rect 6335 43094 6387 43146
rect 6335 42986 6387 43038
rect 6335 42878 6387 42930
rect 6335 42770 6387 42822
rect 6335 42662 6387 42714
rect 6335 42554 6387 42606
rect 6335 42446 6387 42498
rect 6335 42338 6387 42390
rect 6335 42230 6387 42282
rect 6335 42122 6387 42174
rect 6335 42014 6387 42066
rect 6335 41906 6387 41958
rect 6335 41798 6387 41850
rect 6335 41690 6387 41742
rect 6335 41582 6387 41634
rect 6335 41474 6387 41526
rect 6335 41371 6387 41418
rect 6335 41366 6387 41371
rect 7388 44367 7440 44388
rect 7388 44336 7389 44367
rect 7389 44336 7440 44367
rect 7624 44367 7676 44388
rect 7624 44336 7675 44367
rect 7675 44336 7676 44367
rect 7388 44228 7389 44280
rect 7389 44228 7440 44280
rect 7624 44228 7675 44280
rect 7675 44228 7676 44280
rect 7388 44120 7389 44172
rect 7389 44120 7440 44172
rect 7624 44120 7675 44172
rect 7675 44120 7676 44172
rect 7388 44012 7389 44064
rect 7389 44012 7440 44064
rect 7624 44012 7675 44064
rect 7675 44012 7676 44064
rect 7388 43904 7389 43956
rect 7389 43904 7440 43956
rect 7624 43904 7675 43956
rect 7675 43904 7676 43956
rect 7388 43796 7389 43848
rect 7389 43796 7440 43848
rect 7624 43796 7675 43848
rect 7675 43796 7676 43848
rect 7388 43688 7389 43740
rect 7389 43688 7440 43740
rect 7624 43688 7675 43740
rect 7675 43688 7676 43740
rect 7388 43580 7389 43632
rect 7389 43580 7440 43632
rect 7624 43580 7675 43632
rect 7675 43580 7676 43632
rect 7388 43472 7389 43524
rect 7389 43472 7440 43524
rect 7624 43472 7675 43524
rect 7675 43472 7676 43524
rect 7388 43364 7389 43416
rect 7389 43364 7440 43416
rect 7624 43364 7675 43416
rect 7675 43364 7676 43416
rect 7388 43256 7389 43308
rect 7389 43256 7440 43308
rect 7624 43256 7675 43308
rect 7675 43256 7676 43308
rect 7388 43148 7389 43200
rect 7389 43148 7440 43200
rect 7624 43148 7675 43200
rect 7675 43148 7676 43200
rect 7388 43040 7389 43092
rect 7389 43040 7440 43092
rect 7624 43040 7675 43092
rect 7675 43040 7676 43092
rect 7388 42932 7389 42984
rect 7389 42932 7440 42984
rect 7624 42932 7675 42984
rect 7675 42932 7676 42984
rect 7388 42824 7389 42876
rect 7389 42824 7440 42876
rect 7624 42824 7675 42876
rect 7675 42824 7676 42876
rect 7388 42716 7389 42768
rect 7389 42716 7440 42768
rect 7624 42716 7675 42768
rect 7675 42716 7676 42768
rect 7388 42608 7389 42660
rect 7389 42608 7440 42660
rect 7624 42608 7675 42660
rect 7675 42608 7676 42660
rect 7388 42500 7389 42552
rect 7389 42500 7440 42552
rect 7624 42500 7675 42552
rect 7675 42500 7676 42552
rect 7388 42392 7389 42444
rect 7389 42392 7440 42444
rect 7624 42392 7675 42444
rect 7675 42392 7676 42444
rect 7388 42284 7389 42336
rect 7389 42284 7440 42336
rect 7624 42284 7675 42336
rect 7675 42284 7676 42336
rect 7388 42176 7389 42228
rect 7389 42176 7440 42228
rect 7624 42176 7675 42228
rect 7675 42176 7676 42228
rect 7388 42068 7389 42120
rect 7389 42068 7440 42120
rect 7624 42068 7675 42120
rect 7675 42068 7676 42120
rect 7388 41960 7389 42012
rect 7389 41960 7440 42012
rect 7624 41960 7675 42012
rect 7675 41960 7676 42012
rect 7388 41852 7389 41904
rect 7389 41852 7440 41904
rect 7624 41852 7675 41904
rect 7675 41852 7676 41904
rect 7388 41744 7389 41796
rect 7389 41744 7440 41796
rect 7624 41744 7675 41796
rect 7675 41744 7676 41796
rect 7388 41636 7389 41688
rect 7389 41636 7440 41688
rect 7624 41636 7675 41688
rect 7675 41636 7676 41688
rect 7388 41528 7389 41580
rect 7389 41528 7440 41580
rect 7624 41528 7675 41580
rect 7675 41528 7676 41580
rect 7388 41441 7389 41472
rect 7389 41441 7440 41472
rect 7388 41420 7440 41441
rect 7624 41441 7675 41472
rect 7675 41441 7676 41472
rect 7624 41420 7676 41441
rect 8677 44390 8729 44437
rect 8677 44282 8729 44334
rect 8677 44174 8729 44226
rect 8677 44066 8729 44118
rect 8677 43958 8729 44010
rect 8677 43850 8729 43902
rect 8677 43742 8729 43794
rect 8677 43634 8729 43686
rect 8677 43526 8729 43578
rect 8677 43418 8729 43470
rect 8677 43310 8729 43362
rect 8677 43202 8729 43254
rect 8677 43094 8729 43146
rect 8677 42986 8729 43038
rect 8677 42878 8729 42930
rect 8677 42770 8729 42822
rect 8677 42662 8729 42714
rect 8677 42554 8729 42606
rect 8677 42446 8729 42498
rect 8677 42338 8729 42390
rect 8677 42230 8729 42282
rect 8677 42122 8729 42174
rect 8677 42014 8729 42066
rect 8677 41906 8729 41958
rect 8677 41798 8729 41850
rect 8677 41690 8729 41742
rect 8677 41582 8729 41634
rect 8677 41474 8729 41526
rect 8677 41371 8729 41418
rect 11283 44437 11335 44442
rect 13786 44437 13838 44480
rect 13910 44437 13962 44480
rect 14034 44437 14086 44480
rect 8677 41366 8729 41371
rect 11283 44390 11335 44437
rect 13786 44428 13838 44437
rect 13910 44428 13962 44437
rect 14034 44428 14086 44437
rect 11283 44282 11335 44334
rect 11283 44174 11335 44226
rect 11283 44066 11335 44118
rect 11283 43958 11335 44010
rect 11283 43850 11335 43902
rect 11283 43742 11335 43794
rect 11283 43634 11335 43686
rect 11283 43526 11335 43578
rect 11283 43418 11335 43470
rect 11283 43310 11335 43362
rect 11283 43202 11335 43254
rect 11283 43094 11335 43146
rect 11283 42986 11335 43038
rect 11283 42878 11335 42930
rect 11283 42770 11335 42822
rect 11283 42662 11335 42714
rect 11283 42554 11335 42606
rect 11283 42446 11335 42498
rect 11283 42338 11335 42390
rect 11283 42230 11335 42282
rect 11283 42122 11335 42174
rect 11283 42014 11335 42066
rect 11283 41906 11335 41958
rect 11283 41798 11335 41850
rect 11283 41690 11335 41742
rect 11283 41582 11335 41634
rect 11283 41474 11335 41526
rect 11283 41371 11335 41418
rect 13786 44304 13838 44356
rect 13910 44304 13962 44356
rect 14034 44304 14086 44356
rect 13786 44180 13838 44232
rect 13910 44180 13962 44232
rect 14034 44180 14086 44232
rect 13786 44056 13838 44108
rect 13910 44056 13962 44108
rect 14034 44056 14086 44108
rect 13786 43932 13838 43984
rect 13910 43932 13962 43984
rect 14034 43932 14086 43984
rect 13786 43808 13838 43860
rect 13910 43808 13962 43860
rect 14034 43808 14086 43860
rect 13786 43684 13838 43736
rect 13910 43684 13962 43736
rect 14034 43684 14086 43736
rect 13786 43560 13838 43612
rect 13910 43560 13962 43612
rect 14034 43560 14086 43612
rect 13786 43436 13838 43488
rect 13910 43436 13962 43488
rect 14034 43436 14086 43488
rect 13786 43312 13838 43364
rect 13910 43312 13962 43364
rect 14034 43312 14086 43364
rect 13786 43188 13838 43240
rect 13910 43188 13962 43240
rect 14034 43188 14086 43240
rect 13786 43064 13838 43116
rect 13910 43064 13962 43116
rect 14034 43064 14086 43116
rect 13786 42940 13838 42992
rect 13910 42940 13962 42992
rect 14034 42940 14086 42992
rect 13786 42816 13838 42868
rect 13910 42816 13962 42868
rect 14034 42816 14086 42868
rect 13786 42692 13838 42744
rect 13910 42692 13962 42744
rect 14034 42692 14086 42744
rect 13786 42568 13838 42620
rect 13910 42568 13962 42620
rect 14034 42568 14086 42620
rect 13786 42444 13838 42496
rect 13910 42444 13962 42496
rect 14034 42444 14086 42496
rect 13786 42320 13838 42372
rect 13910 42320 13962 42372
rect 14034 42320 14086 42372
rect 13786 42196 13838 42248
rect 13910 42196 13962 42248
rect 14034 42196 14086 42248
rect 13786 42072 13838 42124
rect 13910 42072 13962 42124
rect 14034 42072 14086 42124
rect 13786 41948 13838 42000
rect 13910 41948 13962 42000
rect 14034 41948 14086 42000
rect 13786 41824 13838 41876
rect 13910 41824 13962 41876
rect 14034 41824 14086 41876
rect 13786 41700 13838 41752
rect 13910 41700 13962 41752
rect 14034 41700 14086 41752
rect 13786 41576 13838 41628
rect 13910 41576 13962 41628
rect 14034 41576 14086 41628
rect 13786 41452 13838 41504
rect 13910 41452 13962 41504
rect 14034 41452 14086 41504
rect 13786 41371 13838 41380
rect 13910 41371 13962 41380
rect 14034 41371 14086 41380
rect 11283 41366 11335 41371
rect 13786 41328 13838 41371
rect 13910 41328 13962 41371
rect 14034 41328 14086 41371
rect 444 41120 445 41172
rect 445 41120 496 41172
rect 552 41120 604 41172
rect 660 41120 712 41172
rect 1438 41152 1490 41204
rect 1562 41152 1614 41204
rect 1686 41152 1738 41204
rect 1810 41152 1862 41204
rect 2574 41152 2626 41204
rect 2698 41152 2750 41204
rect 2822 41152 2874 41204
rect 2946 41152 2998 41204
rect 4846 41152 4898 41204
rect 4970 41152 5022 41204
rect 5094 41152 5146 41204
rect 5218 41152 5270 41204
rect 7139 41152 7191 41204
rect 7263 41152 7315 41204
rect 7387 41152 7439 41204
rect 7625 41152 7677 41204
rect 7749 41152 7801 41204
rect 7873 41152 7925 41204
rect 9794 41152 9846 41204
rect 9918 41152 9970 41204
rect 10042 41152 10094 41204
rect 10166 41152 10218 41204
rect 12066 41152 12118 41204
rect 12190 41152 12242 41204
rect 12314 41152 12366 41204
rect 12438 41152 12490 41204
rect 13480 41152 13532 41204
rect 13604 41152 13656 41204
rect 14352 41120 14404 41172
rect 14460 41120 14512 41172
rect 14568 41120 14619 41172
rect 14619 41120 14620 41172
rect 444 41012 445 41064
rect 445 41012 496 41064
rect 552 41012 604 41064
rect 660 41012 712 41064
rect 1438 41028 1490 41080
rect 1562 41028 1614 41080
rect 1686 41028 1738 41080
rect 1810 41028 1862 41080
rect 2574 41028 2626 41080
rect 2698 41028 2750 41080
rect 2822 41028 2874 41080
rect 2946 41028 2998 41080
rect 4846 41028 4898 41080
rect 4970 41028 5022 41080
rect 5094 41028 5146 41080
rect 5218 41028 5270 41080
rect 7139 41028 7191 41080
rect 7263 41028 7315 41080
rect 7387 41028 7439 41080
rect 7625 41028 7677 41080
rect 7749 41028 7801 41080
rect 7873 41028 7925 41080
rect 9794 41028 9846 41080
rect 9918 41028 9970 41080
rect 10042 41028 10094 41080
rect 10166 41028 10218 41080
rect 12066 41028 12118 41080
rect 12190 41028 12242 41080
rect 12314 41028 12366 41080
rect 12438 41028 12490 41080
rect 13480 41028 13532 41080
rect 13604 41028 13656 41080
rect 14352 41012 14404 41064
rect 14460 41012 14512 41064
rect 14568 41012 14619 41064
rect 14619 41012 14620 41064
rect 444 40904 445 40956
rect 445 40904 496 40956
rect 552 40953 604 40956
rect 660 40953 712 40956
rect 1438 40953 1490 40956
rect 1562 40953 1614 40956
rect 1686 40953 1738 40956
rect 1810 40953 1862 40956
rect 2574 40953 2626 40956
rect 2698 40953 2750 40956
rect 2822 40953 2874 40956
rect 2946 40953 2998 40956
rect 4846 40953 4898 40956
rect 4970 40953 5022 40956
rect 5094 40953 5146 40956
rect 5218 40953 5270 40956
rect 7139 40953 7191 40956
rect 7263 40953 7315 40956
rect 7387 40953 7439 40956
rect 7625 40953 7677 40956
rect 7749 40953 7801 40956
rect 7873 40953 7925 40956
rect 9794 40953 9846 40956
rect 9918 40953 9970 40956
rect 10042 40953 10094 40956
rect 10166 40953 10218 40956
rect 12066 40953 12118 40956
rect 12190 40953 12242 40956
rect 12314 40953 12366 40956
rect 12438 40953 12490 40956
rect 13480 40953 13532 40956
rect 13604 40953 13656 40956
rect 14352 40953 14404 40956
rect 14460 40953 14512 40956
rect 552 40907 553 40953
rect 553 40907 604 40953
rect 660 40907 712 40953
rect 1438 40907 1490 40953
rect 1562 40907 1614 40953
rect 1686 40907 1738 40953
rect 1810 40907 1862 40953
rect 2574 40907 2626 40953
rect 2698 40907 2750 40953
rect 2822 40907 2874 40953
rect 2946 40907 2998 40953
rect 4846 40907 4898 40953
rect 4970 40907 5022 40953
rect 5094 40907 5146 40953
rect 5218 40907 5270 40953
rect 7139 40907 7191 40953
rect 7263 40907 7315 40953
rect 7387 40907 7439 40953
rect 7625 40907 7677 40953
rect 7749 40907 7801 40953
rect 7873 40907 7925 40953
rect 9794 40907 9846 40953
rect 9918 40907 9970 40953
rect 10042 40907 10094 40953
rect 10166 40907 10218 40953
rect 12066 40907 12118 40953
rect 12190 40907 12242 40953
rect 12314 40907 12366 40953
rect 12438 40907 12490 40953
rect 13480 40907 13532 40953
rect 13604 40907 13656 40953
rect 14352 40907 14404 40953
rect 14460 40907 14511 40953
rect 14511 40907 14512 40953
rect 552 40904 604 40907
rect 660 40904 712 40907
rect 1438 40904 1490 40907
rect 1562 40904 1614 40907
rect 1686 40904 1738 40907
rect 1810 40904 1862 40907
rect 2574 40904 2626 40907
rect 2698 40904 2750 40907
rect 2822 40904 2874 40907
rect 2946 40904 2998 40907
rect 4846 40904 4898 40907
rect 4970 40904 5022 40907
rect 5094 40904 5146 40907
rect 5218 40904 5270 40907
rect 7139 40904 7191 40907
rect 7263 40904 7315 40907
rect 7387 40904 7439 40907
rect 7625 40904 7677 40907
rect 7749 40904 7801 40907
rect 7873 40904 7925 40907
rect 9794 40904 9846 40907
rect 9918 40904 9970 40907
rect 10042 40904 10094 40907
rect 10166 40904 10218 40907
rect 12066 40904 12118 40907
rect 12190 40904 12242 40907
rect 12314 40904 12366 40907
rect 12438 40904 12490 40907
rect 13480 40904 13532 40907
rect 13604 40904 13656 40907
rect 14352 40904 14404 40907
rect 14460 40904 14512 40907
rect 14568 40904 14619 40956
rect 14619 40904 14620 40956
rect 444 40796 445 40848
rect 445 40796 496 40848
rect 552 40796 604 40848
rect 660 40796 712 40848
rect 1438 40780 1490 40832
rect 1562 40780 1614 40832
rect 1686 40780 1738 40832
rect 1810 40780 1862 40832
rect 2574 40780 2626 40832
rect 2698 40780 2750 40832
rect 2822 40780 2874 40832
rect 2946 40780 2998 40832
rect 4846 40780 4898 40832
rect 4970 40780 5022 40832
rect 5094 40780 5146 40832
rect 5218 40780 5270 40832
rect 7139 40780 7191 40832
rect 7263 40780 7315 40832
rect 7387 40780 7439 40832
rect 7625 40780 7677 40832
rect 7749 40780 7801 40832
rect 7873 40780 7925 40832
rect 9794 40780 9846 40832
rect 9918 40780 9970 40832
rect 10042 40780 10094 40832
rect 10166 40780 10218 40832
rect 12066 40780 12118 40832
rect 12190 40780 12242 40832
rect 12314 40780 12366 40832
rect 12438 40780 12490 40832
rect 13480 40780 13532 40832
rect 13604 40780 13656 40832
rect 14352 40796 14404 40848
rect 14460 40796 14512 40848
rect 14568 40796 14619 40848
rect 14619 40796 14620 40848
rect 444 40688 445 40740
rect 445 40688 496 40740
rect 552 40688 604 40740
rect 660 40688 712 40740
rect 1438 40656 1490 40708
rect 1562 40656 1614 40708
rect 1686 40656 1738 40708
rect 1810 40656 1862 40708
rect 2574 40656 2626 40708
rect 2698 40656 2750 40708
rect 2822 40656 2874 40708
rect 2946 40656 2998 40708
rect 4846 40656 4898 40708
rect 4970 40656 5022 40708
rect 5094 40656 5146 40708
rect 5218 40656 5270 40708
rect 7139 40656 7191 40708
rect 7263 40656 7315 40708
rect 7387 40656 7439 40708
rect 7625 40656 7677 40708
rect 7749 40656 7801 40708
rect 7873 40656 7925 40708
rect 9794 40656 9846 40708
rect 9918 40656 9970 40708
rect 10042 40656 10094 40708
rect 10166 40656 10218 40708
rect 12066 40656 12118 40708
rect 12190 40656 12242 40708
rect 12314 40656 12366 40708
rect 12438 40656 12490 40708
rect 13480 40656 13532 40708
rect 13604 40656 13656 40708
rect 14352 40688 14404 40740
rect 14460 40688 14512 40740
rect 14568 40688 14619 40740
rect 14619 40688 14620 40740
rect 1148 40489 1200 40532
rect 1272 40489 1324 40532
rect 3729 40489 3781 40494
rect 1148 40480 1200 40489
rect 1272 40480 1324 40489
rect 1148 40356 1200 40408
rect 1272 40356 1324 40408
rect 1148 40232 1200 40284
rect 1272 40232 1324 40284
rect 1148 40108 1200 40160
rect 1272 40108 1324 40160
rect 1148 39984 1200 40036
rect 1272 39984 1324 40036
rect 1148 39860 1200 39912
rect 1272 39860 1324 39912
rect 1148 39736 1200 39788
rect 1272 39736 1324 39788
rect 1148 39612 1200 39664
rect 1272 39612 1324 39664
rect 1148 39488 1200 39540
rect 1272 39488 1324 39540
rect 1148 39364 1200 39416
rect 1272 39364 1324 39416
rect 1148 39240 1200 39292
rect 1272 39240 1324 39292
rect 1148 39116 1200 39168
rect 1272 39116 1324 39168
rect 1148 38992 1200 39044
rect 1272 38992 1324 39044
rect 1148 38868 1200 38920
rect 1272 38868 1324 38920
rect 1148 38744 1200 38796
rect 1272 38744 1324 38796
rect 1148 38620 1200 38672
rect 1272 38620 1324 38672
rect 1148 38496 1200 38548
rect 1272 38496 1324 38548
rect 1148 38372 1200 38424
rect 1272 38372 1324 38424
rect 1148 38248 1200 38300
rect 1272 38248 1324 38300
rect 1148 38124 1200 38176
rect 1272 38124 1324 38176
rect 1148 38000 1200 38052
rect 1272 38000 1324 38052
rect 1148 37876 1200 37928
rect 1272 37876 1324 37928
rect 1148 37752 1200 37804
rect 1272 37752 1324 37804
rect 1148 37628 1200 37680
rect 1272 37628 1324 37680
rect 1148 37504 1200 37556
rect 1272 37504 1324 37556
rect 3729 40442 3781 40489
rect 6335 40489 6387 40494
rect 3729 40334 3781 40386
rect 3729 40226 3781 40278
rect 3729 40118 3781 40170
rect 3729 40010 3781 40062
rect 3729 39902 3781 39954
rect 3729 39794 3781 39846
rect 3729 39686 3781 39738
rect 3729 39578 3781 39630
rect 3729 39470 3781 39522
rect 3729 39362 3781 39414
rect 3729 39254 3781 39306
rect 3729 39146 3781 39198
rect 3729 39038 3781 39090
rect 3729 38930 3781 38982
rect 3729 38822 3781 38874
rect 3729 38714 3781 38766
rect 3729 38606 3781 38658
rect 3729 38498 3781 38550
rect 3729 38390 3781 38442
rect 3729 38282 3781 38334
rect 3729 38174 3781 38226
rect 3729 38066 3781 38118
rect 3729 37958 3781 38010
rect 3729 37850 3781 37902
rect 3729 37742 3781 37794
rect 3729 37634 3781 37686
rect 3729 37526 3781 37578
rect 1148 37423 1200 37432
rect 1272 37423 1324 37432
rect 3729 37423 3781 37470
rect 1148 37380 1200 37423
rect 1272 37380 1324 37423
rect 3729 37418 3781 37423
rect 6335 40442 6387 40489
rect 8677 40489 8729 40494
rect 6335 40334 6387 40386
rect 6335 40226 6387 40278
rect 6335 40118 6387 40170
rect 6335 40010 6387 40062
rect 6335 39902 6387 39954
rect 6335 39794 6387 39846
rect 6335 39686 6387 39738
rect 6335 39578 6387 39630
rect 6335 39470 6387 39522
rect 6335 39362 6387 39414
rect 6335 39254 6387 39306
rect 6335 39146 6387 39198
rect 6335 39038 6387 39090
rect 6335 38930 6387 38982
rect 6335 38822 6387 38874
rect 6335 38714 6387 38766
rect 6335 38606 6387 38658
rect 6335 38498 6387 38550
rect 6335 38390 6387 38442
rect 6335 38282 6387 38334
rect 6335 38174 6387 38226
rect 6335 38066 6387 38118
rect 6335 37958 6387 38010
rect 6335 37850 6387 37902
rect 6335 37742 6387 37794
rect 6335 37634 6387 37686
rect 6335 37526 6387 37578
rect 6335 37423 6387 37470
rect 6335 37418 6387 37423
rect 7388 40419 7440 40440
rect 7388 40388 7389 40419
rect 7389 40388 7440 40419
rect 7624 40419 7676 40440
rect 7624 40388 7675 40419
rect 7675 40388 7676 40419
rect 7388 40280 7389 40332
rect 7389 40280 7440 40332
rect 7624 40280 7675 40332
rect 7675 40280 7676 40332
rect 7388 40172 7389 40224
rect 7389 40172 7440 40224
rect 7624 40172 7675 40224
rect 7675 40172 7676 40224
rect 7388 40064 7389 40116
rect 7389 40064 7440 40116
rect 7624 40064 7675 40116
rect 7675 40064 7676 40116
rect 7388 39956 7389 40008
rect 7389 39956 7440 40008
rect 7624 39956 7675 40008
rect 7675 39956 7676 40008
rect 7388 39848 7389 39900
rect 7389 39848 7440 39900
rect 7624 39848 7675 39900
rect 7675 39848 7676 39900
rect 7388 39740 7389 39792
rect 7389 39740 7440 39792
rect 7624 39740 7675 39792
rect 7675 39740 7676 39792
rect 7388 39632 7389 39684
rect 7389 39632 7440 39684
rect 7624 39632 7675 39684
rect 7675 39632 7676 39684
rect 7388 39524 7389 39576
rect 7389 39524 7440 39576
rect 7624 39524 7675 39576
rect 7675 39524 7676 39576
rect 7388 39416 7389 39468
rect 7389 39416 7440 39468
rect 7624 39416 7675 39468
rect 7675 39416 7676 39468
rect 7388 39308 7389 39360
rect 7389 39308 7440 39360
rect 7624 39308 7675 39360
rect 7675 39308 7676 39360
rect 7388 39200 7389 39252
rect 7389 39200 7440 39252
rect 7624 39200 7675 39252
rect 7675 39200 7676 39252
rect 7388 39092 7389 39144
rect 7389 39092 7440 39144
rect 7624 39092 7675 39144
rect 7675 39092 7676 39144
rect 7388 38984 7389 39036
rect 7389 38984 7440 39036
rect 7624 38984 7675 39036
rect 7675 38984 7676 39036
rect 7388 38876 7389 38928
rect 7389 38876 7440 38928
rect 7624 38876 7675 38928
rect 7675 38876 7676 38928
rect 7388 38768 7389 38820
rect 7389 38768 7440 38820
rect 7624 38768 7675 38820
rect 7675 38768 7676 38820
rect 7388 38660 7389 38712
rect 7389 38660 7440 38712
rect 7624 38660 7675 38712
rect 7675 38660 7676 38712
rect 7388 38552 7389 38604
rect 7389 38552 7440 38604
rect 7624 38552 7675 38604
rect 7675 38552 7676 38604
rect 7388 38444 7389 38496
rect 7389 38444 7440 38496
rect 7624 38444 7675 38496
rect 7675 38444 7676 38496
rect 7388 38336 7389 38388
rect 7389 38336 7440 38388
rect 7624 38336 7675 38388
rect 7675 38336 7676 38388
rect 7388 38228 7389 38280
rect 7389 38228 7440 38280
rect 7624 38228 7675 38280
rect 7675 38228 7676 38280
rect 7388 38120 7389 38172
rect 7389 38120 7440 38172
rect 7624 38120 7675 38172
rect 7675 38120 7676 38172
rect 7388 38012 7389 38064
rect 7389 38012 7440 38064
rect 7624 38012 7675 38064
rect 7675 38012 7676 38064
rect 7388 37904 7389 37956
rect 7389 37904 7440 37956
rect 7624 37904 7675 37956
rect 7675 37904 7676 37956
rect 7388 37796 7389 37848
rect 7389 37796 7440 37848
rect 7624 37796 7675 37848
rect 7675 37796 7676 37848
rect 7388 37688 7389 37740
rect 7389 37688 7440 37740
rect 7624 37688 7675 37740
rect 7675 37688 7676 37740
rect 7388 37580 7389 37632
rect 7389 37580 7440 37632
rect 7624 37580 7675 37632
rect 7675 37580 7676 37632
rect 7388 37493 7389 37524
rect 7389 37493 7440 37524
rect 7388 37472 7440 37493
rect 7624 37493 7675 37524
rect 7675 37493 7676 37524
rect 7624 37472 7676 37493
rect 8677 40442 8729 40489
rect 8677 40334 8729 40386
rect 8677 40226 8729 40278
rect 8677 40118 8729 40170
rect 8677 40010 8729 40062
rect 8677 39902 8729 39954
rect 8677 39794 8729 39846
rect 8677 39686 8729 39738
rect 8677 39578 8729 39630
rect 8677 39470 8729 39522
rect 8677 39362 8729 39414
rect 8677 39254 8729 39306
rect 8677 39146 8729 39198
rect 8677 39038 8729 39090
rect 8677 38930 8729 38982
rect 8677 38822 8729 38874
rect 8677 38714 8729 38766
rect 8677 38606 8729 38658
rect 8677 38498 8729 38550
rect 8677 38390 8729 38442
rect 8677 38282 8729 38334
rect 8677 38174 8729 38226
rect 8677 38066 8729 38118
rect 8677 37958 8729 38010
rect 8677 37850 8729 37902
rect 8677 37742 8729 37794
rect 8677 37634 8729 37686
rect 8677 37526 8729 37578
rect 8677 37423 8729 37470
rect 11283 40489 11335 40494
rect 13786 40489 13838 40532
rect 13910 40489 13962 40532
rect 14034 40489 14086 40532
rect 8677 37418 8729 37423
rect 11283 40442 11335 40489
rect 13786 40480 13838 40489
rect 13910 40480 13962 40489
rect 14034 40480 14086 40489
rect 11283 40334 11335 40386
rect 11283 40226 11335 40278
rect 11283 40118 11335 40170
rect 11283 40010 11335 40062
rect 11283 39902 11335 39954
rect 11283 39794 11335 39846
rect 11283 39686 11335 39738
rect 11283 39578 11335 39630
rect 11283 39470 11335 39522
rect 11283 39362 11335 39414
rect 11283 39254 11335 39306
rect 11283 39146 11335 39198
rect 11283 39038 11335 39090
rect 11283 38930 11335 38982
rect 11283 38822 11335 38874
rect 11283 38714 11335 38766
rect 11283 38606 11335 38658
rect 11283 38498 11335 38550
rect 11283 38390 11335 38442
rect 11283 38282 11335 38334
rect 11283 38174 11335 38226
rect 11283 38066 11335 38118
rect 11283 37958 11335 38010
rect 11283 37850 11335 37902
rect 11283 37742 11335 37794
rect 11283 37634 11335 37686
rect 11283 37526 11335 37578
rect 11283 37423 11335 37470
rect 13786 40356 13838 40408
rect 13910 40356 13962 40408
rect 14034 40356 14086 40408
rect 13786 40232 13838 40284
rect 13910 40232 13962 40284
rect 14034 40232 14086 40284
rect 13786 40108 13838 40160
rect 13910 40108 13962 40160
rect 14034 40108 14086 40160
rect 13786 39984 13838 40036
rect 13910 39984 13962 40036
rect 14034 39984 14086 40036
rect 13786 39860 13838 39912
rect 13910 39860 13962 39912
rect 14034 39860 14086 39912
rect 13786 39736 13838 39788
rect 13910 39736 13962 39788
rect 14034 39736 14086 39788
rect 13786 39612 13838 39664
rect 13910 39612 13962 39664
rect 14034 39612 14086 39664
rect 13786 39488 13838 39540
rect 13910 39488 13962 39540
rect 14034 39488 14086 39540
rect 13786 39364 13838 39416
rect 13910 39364 13962 39416
rect 14034 39364 14086 39416
rect 13786 39240 13838 39292
rect 13910 39240 13962 39292
rect 14034 39240 14086 39292
rect 13786 39116 13838 39168
rect 13910 39116 13962 39168
rect 14034 39116 14086 39168
rect 13786 38992 13838 39044
rect 13910 38992 13962 39044
rect 14034 38992 14086 39044
rect 13786 38868 13838 38920
rect 13910 38868 13962 38920
rect 14034 38868 14086 38920
rect 13786 38744 13838 38796
rect 13910 38744 13962 38796
rect 14034 38744 14086 38796
rect 13786 38620 13838 38672
rect 13910 38620 13962 38672
rect 14034 38620 14086 38672
rect 13786 38496 13838 38548
rect 13910 38496 13962 38548
rect 14034 38496 14086 38548
rect 13786 38372 13838 38424
rect 13910 38372 13962 38424
rect 14034 38372 14086 38424
rect 13786 38248 13838 38300
rect 13910 38248 13962 38300
rect 14034 38248 14086 38300
rect 13786 38124 13838 38176
rect 13910 38124 13962 38176
rect 14034 38124 14086 38176
rect 13786 38000 13838 38052
rect 13910 38000 13962 38052
rect 14034 38000 14086 38052
rect 13786 37876 13838 37928
rect 13910 37876 13962 37928
rect 14034 37876 14086 37928
rect 13786 37752 13838 37804
rect 13910 37752 13962 37804
rect 14034 37752 14086 37804
rect 13786 37628 13838 37680
rect 13910 37628 13962 37680
rect 14034 37628 14086 37680
rect 13786 37504 13838 37556
rect 13910 37504 13962 37556
rect 14034 37504 14086 37556
rect 13786 37423 13838 37432
rect 13910 37423 13962 37432
rect 14034 37423 14086 37432
rect 11283 37418 11335 37423
rect 13786 37380 13838 37423
rect 13910 37380 13962 37423
rect 14034 37380 14086 37423
rect 444 37172 445 37224
rect 445 37172 496 37224
rect 552 37172 604 37224
rect 660 37172 712 37224
rect 1438 37204 1490 37256
rect 1562 37204 1614 37256
rect 1686 37204 1738 37256
rect 1810 37204 1862 37256
rect 2574 37204 2626 37256
rect 2698 37204 2750 37256
rect 2822 37204 2874 37256
rect 2946 37204 2998 37256
rect 4846 37204 4898 37256
rect 4970 37204 5022 37256
rect 5094 37204 5146 37256
rect 5218 37204 5270 37256
rect 7139 37204 7191 37256
rect 7263 37204 7315 37256
rect 7387 37204 7439 37256
rect 7625 37204 7677 37256
rect 7749 37204 7801 37256
rect 7873 37204 7925 37256
rect 9794 37204 9846 37256
rect 9918 37204 9970 37256
rect 10042 37204 10094 37256
rect 10166 37204 10218 37256
rect 12066 37204 12118 37256
rect 12190 37204 12242 37256
rect 12314 37204 12366 37256
rect 12438 37204 12490 37256
rect 13480 37204 13532 37256
rect 13604 37204 13656 37256
rect 14352 37172 14404 37224
rect 14460 37172 14512 37224
rect 14568 37172 14619 37224
rect 14619 37172 14620 37224
rect 444 37064 445 37116
rect 445 37064 496 37116
rect 552 37064 604 37116
rect 660 37064 712 37116
rect 1438 37080 1490 37132
rect 1562 37080 1614 37132
rect 1686 37080 1738 37132
rect 1810 37080 1862 37132
rect 2574 37080 2626 37132
rect 2698 37080 2750 37132
rect 2822 37080 2874 37132
rect 2946 37080 2998 37132
rect 4846 37080 4898 37132
rect 4970 37080 5022 37132
rect 5094 37080 5146 37132
rect 5218 37080 5270 37132
rect 7139 37080 7191 37132
rect 7263 37080 7315 37132
rect 7387 37080 7439 37132
rect 7625 37080 7677 37132
rect 7749 37080 7801 37132
rect 7873 37080 7925 37132
rect 9794 37080 9846 37132
rect 9918 37080 9970 37132
rect 10042 37080 10094 37132
rect 10166 37080 10218 37132
rect 12066 37080 12118 37132
rect 12190 37080 12242 37132
rect 12314 37080 12366 37132
rect 12438 37080 12490 37132
rect 13480 37080 13532 37132
rect 13604 37080 13656 37132
rect 14352 37064 14404 37116
rect 14460 37064 14512 37116
rect 14568 37064 14619 37116
rect 14619 37064 14620 37116
rect 444 36956 445 37008
rect 445 36956 496 37008
rect 552 37005 604 37008
rect 660 37005 712 37008
rect 1438 37005 1490 37008
rect 1562 37005 1614 37008
rect 1686 37005 1738 37008
rect 1810 37005 1862 37008
rect 2574 37005 2626 37008
rect 2698 37005 2750 37008
rect 2822 37005 2874 37008
rect 2946 37005 2998 37008
rect 4846 37005 4898 37008
rect 4970 37005 5022 37008
rect 5094 37005 5146 37008
rect 5218 37005 5270 37008
rect 7139 37005 7191 37008
rect 7263 37005 7315 37008
rect 7387 37005 7439 37008
rect 7625 37005 7677 37008
rect 7749 37005 7801 37008
rect 7873 37005 7925 37008
rect 9794 37005 9846 37008
rect 9918 37005 9970 37008
rect 10042 37005 10094 37008
rect 10166 37005 10218 37008
rect 12066 37005 12118 37008
rect 12190 37005 12242 37008
rect 12314 37005 12366 37008
rect 12438 37005 12490 37008
rect 13480 37005 13532 37008
rect 13604 37005 13656 37008
rect 14352 37005 14404 37008
rect 14460 37005 14512 37008
rect 552 36959 553 37005
rect 553 36959 604 37005
rect 660 36959 712 37005
rect 1438 36959 1490 37005
rect 1562 36959 1614 37005
rect 1686 36959 1738 37005
rect 1810 36959 1862 37005
rect 2574 36959 2626 37005
rect 2698 36959 2750 37005
rect 2822 36959 2874 37005
rect 2946 36959 2998 37005
rect 4846 36959 4898 37005
rect 4970 36959 5022 37005
rect 5094 36959 5146 37005
rect 5218 36959 5270 37005
rect 7139 36959 7191 37005
rect 7263 36959 7315 37005
rect 7387 36959 7439 37005
rect 7625 36959 7677 37005
rect 7749 36959 7801 37005
rect 7873 36959 7925 37005
rect 9794 36959 9846 37005
rect 9918 36959 9970 37005
rect 10042 36959 10094 37005
rect 10166 36959 10218 37005
rect 12066 36959 12118 37005
rect 12190 36959 12242 37005
rect 12314 36959 12366 37005
rect 12438 36959 12490 37005
rect 13480 36959 13532 37005
rect 13604 36959 13656 37005
rect 14352 36959 14404 37005
rect 14460 36959 14511 37005
rect 14511 36959 14512 37005
rect 552 36956 604 36959
rect 660 36956 712 36959
rect 1438 36956 1490 36959
rect 1562 36956 1614 36959
rect 1686 36956 1738 36959
rect 1810 36956 1862 36959
rect 2574 36956 2626 36959
rect 2698 36956 2750 36959
rect 2822 36956 2874 36959
rect 2946 36956 2998 36959
rect 4846 36956 4898 36959
rect 4970 36956 5022 36959
rect 5094 36956 5146 36959
rect 5218 36956 5270 36959
rect 7139 36956 7191 36959
rect 7263 36956 7315 36959
rect 7387 36956 7439 36959
rect 7625 36956 7677 36959
rect 7749 36956 7801 36959
rect 7873 36956 7925 36959
rect 9794 36956 9846 36959
rect 9918 36956 9970 36959
rect 10042 36956 10094 36959
rect 10166 36956 10218 36959
rect 12066 36956 12118 36959
rect 12190 36956 12242 36959
rect 12314 36956 12366 36959
rect 12438 36956 12490 36959
rect 13480 36956 13532 36959
rect 13604 36956 13656 36959
rect 14352 36956 14404 36959
rect 14460 36956 14512 36959
rect 14568 36956 14619 37008
rect 14619 36956 14620 37008
rect 444 36848 445 36900
rect 445 36848 496 36900
rect 552 36848 604 36900
rect 660 36848 712 36900
rect 1438 36832 1490 36884
rect 1562 36832 1614 36884
rect 1686 36832 1738 36884
rect 1810 36832 1862 36884
rect 2574 36832 2626 36884
rect 2698 36832 2750 36884
rect 2822 36832 2874 36884
rect 2946 36832 2998 36884
rect 4846 36832 4898 36884
rect 4970 36832 5022 36884
rect 5094 36832 5146 36884
rect 5218 36832 5270 36884
rect 7139 36832 7191 36884
rect 7263 36832 7315 36884
rect 7387 36832 7439 36884
rect 7625 36832 7677 36884
rect 7749 36832 7801 36884
rect 7873 36832 7925 36884
rect 9794 36832 9846 36884
rect 9918 36832 9970 36884
rect 10042 36832 10094 36884
rect 10166 36832 10218 36884
rect 12066 36832 12118 36884
rect 12190 36832 12242 36884
rect 12314 36832 12366 36884
rect 12438 36832 12490 36884
rect 13480 36832 13532 36884
rect 13604 36832 13656 36884
rect 14352 36848 14404 36900
rect 14460 36848 14512 36900
rect 14568 36848 14619 36900
rect 14619 36848 14620 36900
rect 444 36740 445 36792
rect 445 36740 496 36792
rect 552 36740 604 36792
rect 660 36740 712 36792
rect 1438 36708 1490 36760
rect 1562 36708 1614 36760
rect 1686 36708 1738 36760
rect 1810 36708 1862 36760
rect 2574 36708 2626 36760
rect 2698 36708 2750 36760
rect 2822 36708 2874 36760
rect 2946 36708 2998 36760
rect 4846 36708 4898 36760
rect 4970 36708 5022 36760
rect 5094 36708 5146 36760
rect 5218 36708 5270 36760
rect 7139 36708 7191 36760
rect 7263 36708 7315 36760
rect 7387 36708 7439 36760
rect 7625 36708 7677 36760
rect 7749 36708 7801 36760
rect 7873 36708 7925 36760
rect 9794 36708 9846 36760
rect 9918 36708 9970 36760
rect 10042 36708 10094 36760
rect 10166 36708 10218 36760
rect 12066 36708 12118 36760
rect 12190 36708 12242 36760
rect 12314 36708 12366 36760
rect 12438 36708 12490 36760
rect 13480 36708 13532 36760
rect 13604 36708 13656 36760
rect 14352 36740 14404 36792
rect 14460 36740 14512 36792
rect 14568 36740 14619 36792
rect 14619 36740 14620 36792
rect 978 36541 1030 36584
rect 1102 36541 1154 36584
rect 1226 36541 1278 36584
rect 3729 36541 3781 36546
rect 978 36532 1030 36541
rect 1102 36532 1154 36541
rect 1226 36532 1278 36541
rect 978 36408 1030 36460
rect 1102 36408 1154 36460
rect 1226 36408 1278 36460
rect 978 36284 1030 36336
rect 1102 36284 1154 36336
rect 1226 36284 1278 36336
rect 978 36160 1030 36212
rect 1102 36160 1154 36212
rect 1226 36160 1278 36212
rect 978 36036 1030 36088
rect 1102 36036 1154 36088
rect 1226 36036 1278 36088
rect 978 35912 1030 35964
rect 1102 35912 1154 35964
rect 1226 35912 1278 35964
rect 978 35788 1030 35840
rect 1102 35788 1154 35840
rect 1226 35788 1278 35840
rect 978 35664 1030 35716
rect 1102 35664 1154 35716
rect 1226 35664 1278 35716
rect 978 35540 1030 35592
rect 1102 35540 1154 35592
rect 1226 35540 1278 35592
rect 978 35416 1030 35468
rect 1102 35416 1154 35468
rect 1226 35416 1278 35468
rect 978 35292 1030 35344
rect 1102 35292 1154 35344
rect 1226 35292 1278 35344
rect 978 35168 1030 35220
rect 1102 35168 1154 35220
rect 1226 35168 1278 35220
rect 978 35044 1030 35096
rect 1102 35044 1154 35096
rect 1226 35044 1278 35096
rect 978 34920 1030 34972
rect 1102 34920 1154 34972
rect 1226 34920 1278 34972
rect 978 34796 1030 34848
rect 1102 34796 1154 34848
rect 1226 34796 1278 34848
rect 978 34672 1030 34724
rect 1102 34672 1154 34724
rect 1226 34672 1278 34724
rect 978 34548 1030 34600
rect 1102 34548 1154 34600
rect 1226 34548 1278 34600
rect 978 34424 1030 34476
rect 1102 34424 1154 34476
rect 1226 34424 1278 34476
rect 978 34300 1030 34352
rect 1102 34300 1154 34352
rect 1226 34300 1278 34352
rect 978 34176 1030 34228
rect 1102 34176 1154 34228
rect 1226 34176 1278 34228
rect 978 34052 1030 34104
rect 1102 34052 1154 34104
rect 1226 34052 1278 34104
rect 978 33928 1030 33980
rect 1102 33928 1154 33980
rect 1226 33928 1278 33980
rect 978 33804 1030 33856
rect 1102 33804 1154 33856
rect 1226 33804 1278 33856
rect 978 33680 1030 33732
rect 1102 33680 1154 33732
rect 1226 33680 1278 33732
rect 978 33556 1030 33608
rect 1102 33556 1154 33608
rect 1226 33556 1278 33608
rect 3729 36494 3781 36541
rect 6335 36541 6387 36546
rect 3729 36386 3781 36438
rect 3729 36278 3781 36330
rect 3729 36170 3781 36222
rect 3729 36062 3781 36114
rect 3729 35954 3781 36006
rect 3729 35846 3781 35898
rect 3729 35738 3781 35790
rect 3729 35630 3781 35682
rect 3729 35522 3781 35574
rect 3729 35414 3781 35466
rect 3729 35306 3781 35358
rect 3729 35198 3781 35250
rect 3729 35090 3781 35142
rect 3729 34982 3781 35034
rect 3729 34874 3781 34926
rect 3729 34766 3781 34818
rect 3729 34658 3781 34710
rect 3729 34550 3781 34602
rect 3729 34442 3781 34494
rect 3729 34334 3781 34386
rect 3729 34226 3781 34278
rect 3729 34118 3781 34170
rect 3729 34010 3781 34062
rect 3729 33902 3781 33954
rect 3729 33794 3781 33846
rect 3729 33686 3781 33738
rect 3729 33578 3781 33630
rect 978 33475 1030 33484
rect 1102 33475 1154 33484
rect 1226 33475 1278 33484
rect 3729 33475 3781 33522
rect 978 33432 1030 33475
rect 1102 33432 1154 33475
rect 1226 33432 1278 33475
rect 3729 33470 3781 33475
rect 6335 36494 6387 36541
rect 8677 36541 8729 36546
rect 6335 36386 6387 36438
rect 6335 36278 6387 36330
rect 6335 36170 6387 36222
rect 6335 36062 6387 36114
rect 6335 35954 6387 36006
rect 6335 35846 6387 35898
rect 6335 35738 6387 35790
rect 6335 35630 6387 35682
rect 6335 35522 6387 35574
rect 6335 35414 6387 35466
rect 6335 35306 6387 35358
rect 6335 35198 6387 35250
rect 6335 35090 6387 35142
rect 6335 34982 6387 35034
rect 6335 34874 6387 34926
rect 6335 34766 6387 34818
rect 6335 34658 6387 34710
rect 6335 34550 6387 34602
rect 6335 34442 6387 34494
rect 6335 34334 6387 34386
rect 6335 34226 6387 34278
rect 6335 34118 6387 34170
rect 6335 34010 6387 34062
rect 6335 33902 6387 33954
rect 6335 33794 6387 33846
rect 6335 33686 6387 33738
rect 6335 33578 6387 33630
rect 6335 33475 6387 33522
rect 6335 33470 6387 33475
rect 7388 36471 7440 36492
rect 7388 36440 7389 36471
rect 7389 36440 7440 36471
rect 7624 36471 7676 36492
rect 7624 36440 7675 36471
rect 7675 36440 7676 36471
rect 7388 36332 7389 36384
rect 7389 36332 7440 36384
rect 7624 36332 7675 36384
rect 7675 36332 7676 36384
rect 7388 36224 7389 36276
rect 7389 36224 7440 36276
rect 7624 36224 7675 36276
rect 7675 36224 7676 36276
rect 7388 36116 7389 36168
rect 7389 36116 7440 36168
rect 7624 36116 7675 36168
rect 7675 36116 7676 36168
rect 7388 36008 7389 36060
rect 7389 36008 7440 36060
rect 7624 36008 7675 36060
rect 7675 36008 7676 36060
rect 7388 35900 7389 35952
rect 7389 35900 7440 35952
rect 7624 35900 7675 35952
rect 7675 35900 7676 35952
rect 7388 35792 7389 35844
rect 7389 35792 7440 35844
rect 7624 35792 7675 35844
rect 7675 35792 7676 35844
rect 7388 35684 7389 35736
rect 7389 35684 7440 35736
rect 7624 35684 7675 35736
rect 7675 35684 7676 35736
rect 7388 35576 7389 35628
rect 7389 35576 7440 35628
rect 7624 35576 7675 35628
rect 7675 35576 7676 35628
rect 7388 35468 7389 35520
rect 7389 35468 7440 35520
rect 7624 35468 7675 35520
rect 7675 35468 7676 35520
rect 7388 35360 7389 35412
rect 7389 35360 7440 35412
rect 7624 35360 7675 35412
rect 7675 35360 7676 35412
rect 7388 35252 7389 35304
rect 7389 35252 7440 35304
rect 7624 35252 7675 35304
rect 7675 35252 7676 35304
rect 7388 35144 7389 35196
rect 7389 35144 7440 35196
rect 7624 35144 7675 35196
rect 7675 35144 7676 35196
rect 7388 35036 7389 35088
rect 7389 35036 7440 35088
rect 7624 35036 7675 35088
rect 7675 35036 7676 35088
rect 7388 34928 7389 34980
rect 7389 34928 7440 34980
rect 7624 34928 7675 34980
rect 7675 34928 7676 34980
rect 7388 34820 7389 34872
rect 7389 34820 7440 34872
rect 7624 34820 7675 34872
rect 7675 34820 7676 34872
rect 7388 34712 7389 34764
rect 7389 34712 7440 34764
rect 7624 34712 7675 34764
rect 7675 34712 7676 34764
rect 7388 34604 7389 34656
rect 7389 34604 7440 34656
rect 7624 34604 7675 34656
rect 7675 34604 7676 34656
rect 7388 34496 7389 34548
rect 7389 34496 7440 34548
rect 7624 34496 7675 34548
rect 7675 34496 7676 34548
rect 7388 34388 7389 34440
rect 7389 34388 7440 34440
rect 7624 34388 7675 34440
rect 7675 34388 7676 34440
rect 7388 34280 7389 34332
rect 7389 34280 7440 34332
rect 7624 34280 7675 34332
rect 7675 34280 7676 34332
rect 7388 34172 7389 34224
rect 7389 34172 7440 34224
rect 7624 34172 7675 34224
rect 7675 34172 7676 34224
rect 7388 34064 7389 34116
rect 7389 34064 7440 34116
rect 7624 34064 7675 34116
rect 7675 34064 7676 34116
rect 7388 33956 7389 34008
rect 7389 33956 7440 34008
rect 7624 33956 7675 34008
rect 7675 33956 7676 34008
rect 7388 33848 7389 33900
rect 7389 33848 7440 33900
rect 7624 33848 7675 33900
rect 7675 33848 7676 33900
rect 7388 33740 7389 33792
rect 7389 33740 7440 33792
rect 7624 33740 7675 33792
rect 7675 33740 7676 33792
rect 7388 33632 7389 33684
rect 7389 33632 7440 33684
rect 7624 33632 7675 33684
rect 7675 33632 7676 33684
rect 7388 33545 7389 33576
rect 7389 33545 7440 33576
rect 7388 33524 7440 33545
rect 7624 33545 7675 33576
rect 7675 33545 7676 33576
rect 7624 33524 7676 33545
rect 8677 36494 8729 36541
rect 8677 36386 8729 36438
rect 8677 36278 8729 36330
rect 8677 36170 8729 36222
rect 8677 36062 8729 36114
rect 8677 35954 8729 36006
rect 8677 35846 8729 35898
rect 8677 35738 8729 35790
rect 8677 35630 8729 35682
rect 8677 35522 8729 35574
rect 8677 35414 8729 35466
rect 8677 35306 8729 35358
rect 8677 35198 8729 35250
rect 8677 35090 8729 35142
rect 8677 34982 8729 35034
rect 8677 34874 8729 34926
rect 8677 34766 8729 34818
rect 8677 34658 8729 34710
rect 8677 34550 8729 34602
rect 8677 34442 8729 34494
rect 8677 34334 8729 34386
rect 8677 34226 8729 34278
rect 8677 34118 8729 34170
rect 8677 34010 8729 34062
rect 8677 33902 8729 33954
rect 8677 33794 8729 33846
rect 8677 33686 8729 33738
rect 8677 33578 8729 33630
rect 8677 33475 8729 33522
rect 11283 36541 11335 36546
rect 13786 36541 13838 36584
rect 13910 36541 13962 36584
rect 14034 36541 14086 36584
rect 8677 33470 8729 33475
rect 11283 36494 11335 36541
rect 13786 36532 13838 36541
rect 13910 36532 13962 36541
rect 14034 36532 14086 36541
rect 11283 36386 11335 36438
rect 11283 36278 11335 36330
rect 11283 36170 11335 36222
rect 11283 36062 11335 36114
rect 11283 35954 11335 36006
rect 11283 35846 11335 35898
rect 11283 35738 11335 35790
rect 11283 35630 11335 35682
rect 11283 35522 11335 35574
rect 11283 35414 11335 35466
rect 11283 35306 11335 35358
rect 11283 35198 11335 35250
rect 11283 35090 11335 35142
rect 11283 34982 11335 35034
rect 11283 34874 11335 34926
rect 11283 34766 11335 34818
rect 11283 34658 11335 34710
rect 11283 34550 11335 34602
rect 11283 34442 11335 34494
rect 11283 34334 11335 34386
rect 11283 34226 11335 34278
rect 11283 34118 11335 34170
rect 11283 34010 11335 34062
rect 11283 33902 11335 33954
rect 11283 33794 11335 33846
rect 11283 33686 11335 33738
rect 11283 33578 11335 33630
rect 11283 33475 11335 33522
rect 13786 36408 13838 36460
rect 13910 36408 13962 36460
rect 14034 36408 14086 36460
rect 13786 36284 13838 36336
rect 13910 36284 13962 36336
rect 14034 36284 14086 36336
rect 13786 36160 13838 36212
rect 13910 36160 13962 36212
rect 14034 36160 14086 36212
rect 13786 36036 13838 36088
rect 13910 36036 13962 36088
rect 14034 36036 14086 36088
rect 13786 35912 13838 35964
rect 13910 35912 13962 35964
rect 14034 35912 14086 35964
rect 13786 35788 13838 35840
rect 13910 35788 13962 35840
rect 14034 35788 14086 35840
rect 13786 35664 13838 35716
rect 13910 35664 13962 35716
rect 14034 35664 14086 35716
rect 13786 35540 13838 35592
rect 13910 35540 13962 35592
rect 14034 35540 14086 35592
rect 13786 35416 13838 35468
rect 13910 35416 13962 35468
rect 14034 35416 14086 35468
rect 13786 35292 13838 35344
rect 13910 35292 13962 35344
rect 14034 35292 14086 35344
rect 13786 35168 13838 35220
rect 13910 35168 13962 35220
rect 14034 35168 14086 35220
rect 13786 35044 13838 35096
rect 13910 35044 13962 35096
rect 14034 35044 14086 35096
rect 13786 34920 13838 34972
rect 13910 34920 13962 34972
rect 14034 34920 14086 34972
rect 13786 34796 13838 34848
rect 13910 34796 13962 34848
rect 14034 34796 14086 34848
rect 13786 34672 13838 34724
rect 13910 34672 13962 34724
rect 14034 34672 14086 34724
rect 13786 34548 13838 34600
rect 13910 34548 13962 34600
rect 14034 34548 14086 34600
rect 13786 34424 13838 34476
rect 13910 34424 13962 34476
rect 14034 34424 14086 34476
rect 13786 34300 13838 34352
rect 13910 34300 13962 34352
rect 14034 34300 14086 34352
rect 13786 34176 13838 34228
rect 13910 34176 13962 34228
rect 14034 34176 14086 34228
rect 13786 34052 13838 34104
rect 13910 34052 13962 34104
rect 14034 34052 14086 34104
rect 13786 33928 13838 33980
rect 13910 33928 13962 33980
rect 14034 33928 14086 33980
rect 13786 33804 13838 33856
rect 13910 33804 13962 33856
rect 14034 33804 14086 33856
rect 13786 33680 13838 33732
rect 13910 33680 13962 33732
rect 14034 33680 14086 33732
rect 13786 33556 13838 33608
rect 13910 33556 13962 33608
rect 14034 33556 14086 33608
rect 13786 33475 13838 33484
rect 13910 33475 13962 33484
rect 14034 33475 14086 33484
rect 11283 33470 11335 33475
rect 13786 33432 13838 33475
rect 13910 33432 13962 33475
rect 14034 33432 14086 33475
rect 444 33224 445 33276
rect 445 33224 496 33276
rect 552 33224 604 33276
rect 660 33224 712 33276
rect 1438 33256 1490 33308
rect 1562 33256 1614 33308
rect 1686 33256 1738 33308
rect 1810 33256 1862 33308
rect 2574 33256 2626 33308
rect 2698 33256 2750 33308
rect 2822 33256 2874 33308
rect 2946 33256 2998 33308
rect 4846 33256 4898 33308
rect 4970 33256 5022 33308
rect 5094 33256 5146 33308
rect 5218 33256 5270 33308
rect 7139 33256 7191 33308
rect 7263 33256 7315 33308
rect 7387 33256 7439 33308
rect 7625 33256 7677 33308
rect 7749 33256 7801 33308
rect 7873 33256 7925 33308
rect 9794 33256 9846 33308
rect 9918 33256 9970 33308
rect 10042 33256 10094 33308
rect 10166 33256 10218 33308
rect 12066 33256 12118 33308
rect 12190 33256 12242 33308
rect 12314 33256 12366 33308
rect 12438 33256 12490 33308
rect 13202 33256 13254 33308
rect 13326 33256 13378 33308
rect 13450 33256 13502 33308
rect 13574 33256 13626 33308
rect 14352 33224 14404 33276
rect 14460 33224 14512 33276
rect 14568 33224 14619 33276
rect 14619 33224 14620 33276
rect 444 33116 445 33168
rect 445 33116 496 33168
rect 552 33116 604 33168
rect 660 33116 712 33168
rect 1438 33132 1490 33184
rect 1562 33132 1614 33184
rect 1686 33132 1738 33184
rect 1810 33132 1862 33184
rect 2574 33132 2626 33184
rect 2698 33132 2750 33184
rect 2822 33132 2874 33184
rect 2946 33132 2998 33184
rect 4846 33132 4898 33184
rect 4970 33132 5022 33184
rect 5094 33132 5146 33184
rect 5218 33132 5270 33184
rect 7139 33132 7191 33184
rect 7263 33132 7315 33184
rect 7387 33132 7439 33184
rect 7625 33132 7677 33184
rect 7749 33132 7801 33184
rect 7873 33132 7925 33184
rect 9794 33132 9846 33184
rect 9918 33132 9970 33184
rect 10042 33132 10094 33184
rect 10166 33132 10218 33184
rect 12066 33132 12118 33184
rect 12190 33132 12242 33184
rect 12314 33132 12366 33184
rect 12438 33132 12490 33184
rect 13202 33132 13254 33184
rect 13326 33132 13378 33184
rect 13450 33132 13502 33184
rect 13574 33132 13626 33184
rect 14352 33116 14404 33168
rect 14460 33116 14512 33168
rect 14568 33116 14619 33168
rect 14619 33116 14620 33168
rect 444 33008 445 33060
rect 445 33008 496 33060
rect 552 33057 604 33060
rect 660 33057 712 33060
rect 1438 33057 1490 33060
rect 1562 33057 1614 33060
rect 1686 33057 1738 33060
rect 1810 33057 1862 33060
rect 2574 33057 2626 33060
rect 2698 33057 2750 33060
rect 2822 33057 2874 33060
rect 2946 33057 2998 33060
rect 4846 33057 4898 33060
rect 4970 33057 5022 33060
rect 5094 33057 5146 33060
rect 5218 33057 5270 33060
rect 7139 33057 7191 33060
rect 7263 33057 7315 33060
rect 7387 33057 7439 33060
rect 7625 33057 7677 33060
rect 7749 33057 7801 33060
rect 7873 33057 7925 33060
rect 9794 33057 9846 33060
rect 9918 33057 9970 33060
rect 10042 33057 10094 33060
rect 10166 33057 10218 33060
rect 12066 33057 12118 33060
rect 12190 33057 12242 33060
rect 12314 33057 12366 33060
rect 12438 33057 12490 33060
rect 13202 33057 13254 33060
rect 13326 33057 13378 33060
rect 13450 33057 13502 33060
rect 13574 33057 13626 33060
rect 14352 33057 14404 33060
rect 14460 33057 14512 33060
rect 552 33011 553 33057
rect 553 33011 604 33057
rect 660 33011 712 33057
rect 1438 33011 1490 33057
rect 1562 33011 1614 33057
rect 1686 33011 1738 33057
rect 1810 33011 1862 33057
rect 2574 33011 2626 33057
rect 2698 33011 2750 33057
rect 2822 33011 2874 33057
rect 2946 33011 2998 33057
rect 4846 33011 4898 33057
rect 4970 33011 5022 33057
rect 5094 33011 5146 33057
rect 5218 33011 5270 33057
rect 7139 33011 7191 33057
rect 7263 33011 7315 33057
rect 7387 33011 7439 33057
rect 7625 33011 7677 33057
rect 7749 33011 7801 33057
rect 7873 33011 7925 33057
rect 9794 33011 9846 33057
rect 9918 33011 9970 33057
rect 10042 33011 10094 33057
rect 10166 33011 10218 33057
rect 12066 33011 12118 33057
rect 12190 33011 12242 33057
rect 12314 33011 12366 33057
rect 12438 33011 12490 33057
rect 13202 33011 13254 33057
rect 13326 33011 13378 33057
rect 13450 33011 13502 33057
rect 13574 33011 13626 33057
rect 14352 33011 14404 33057
rect 14460 33011 14511 33057
rect 14511 33011 14512 33057
rect 552 33008 604 33011
rect 660 33008 712 33011
rect 1438 33008 1490 33011
rect 1562 33008 1614 33011
rect 1686 33008 1738 33011
rect 1810 33008 1862 33011
rect 2574 33008 2626 33011
rect 2698 33008 2750 33011
rect 2822 33008 2874 33011
rect 2946 33008 2998 33011
rect 4846 33008 4898 33011
rect 4970 33008 5022 33011
rect 5094 33008 5146 33011
rect 5218 33008 5270 33011
rect 7139 33008 7191 33011
rect 7263 33008 7315 33011
rect 7387 33008 7439 33011
rect 7625 33008 7677 33011
rect 7749 33008 7801 33011
rect 7873 33008 7925 33011
rect 9794 33008 9846 33011
rect 9918 33008 9970 33011
rect 10042 33008 10094 33011
rect 10166 33008 10218 33011
rect 12066 33008 12118 33011
rect 12190 33008 12242 33011
rect 12314 33008 12366 33011
rect 12438 33008 12490 33011
rect 13202 33008 13254 33011
rect 13326 33008 13378 33011
rect 13450 33008 13502 33011
rect 13574 33008 13626 33011
rect 14352 33008 14404 33011
rect 14460 33008 14512 33011
rect 14568 33008 14619 33060
rect 14619 33008 14620 33060
rect 444 32900 445 32952
rect 445 32900 496 32952
rect 552 32900 604 32952
rect 660 32900 712 32952
rect 1438 32884 1490 32936
rect 1562 32884 1614 32936
rect 1686 32884 1738 32936
rect 1810 32884 1862 32936
rect 2574 32884 2626 32936
rect 2698 32884 2750 32936
rect 2822 32884 2874 32936
rect 2946 32884 2998 32936
rect 4846 32884 4898 32936
rect 4970 32884 5022 32936
rect 5094 32884 5146 32936
rect 5218 32884 5270 32936
rect 7139 32884 7191 32936
rect 7263 32884 7315 32936
rect 7387 32884 7439 32936
rect 7625 32884 7677 32936
rect 7749 32884 7801 32936
rect 7873 32884 7925 32936
rect 9794 32884 9846 32936
rect 9918 32884 9970 32936
rect 10042 32884 10094 32936
rect 10166 32884 10218 32936
rect 12066 32884 12118 32936
rect 12190 32884 12242 32936
rect 12314 32884 12366 32936
rect 12438 32884 12490 32936
rect 13202 32884 13254 32936
rect 13326 32884 13378 32936
rect 13450 32884 13502 32936
rect 13574 32884 13626 32936
rect 14352 32900 14404 32952
rect 14460 32900 14512 32952
rect 14568 32900 14619 32952
rect 14619 32900 14620 32952
rect 444 32792 445 32844
rect 445 32792 496 32844
rect 552 32792 604 32844
rect 660 32792 712 32844
rect 1438 32760 1490 32812
rect 1562 32760 1614 32812
rect 1686 32760 1738 32812
rect 1810 32760 1862 32812
rect 2574 32760 2626 32812
rect 2698 32760 2750 32812
rect 2822 32760 2874 32812
rect 2946 32760 2998 32812
rect 4846 32760 4898 32812
rect 4970 32760 5022 32812
rect 5094 32760 5146 32812
rect 5218 32760 5270 32812
rect 7139 32760 7191 32812
rect 7263 32760 7315 32812
rect 7387 32760 7439 32812
rect 7625 32760 7677 32812
rect 7749 32760 7801 32812
rect 7873 32760 7925 32812
rect 9794 32760 9846 32812
rect 9918 32760 9970 32812
rect 10042 32760 10094 32812
rect 10166 32760 10218 32812
rect 12066 32760 12118 32812
rect 12190 32760 12242 32812
rect 12314 32760 12366 32812
rect 12438 32760 12490 32812
rect 13202 32760 13254 32812
rect 13326 32760 13378 32812
rect 13450 32760 13502 32812
rect 13574 32760 13626 32812
rect 14352 32792 14404 32844
rect 14460 32792 14512 32844
rect 14568 32792 14619 32844
rect 14619 32792 14620 32844
rect 978 32593 1030 32636
rect 1102 32593 1154 32636
rect 1226 32593 1278 32636
rect 3729 32593 3781 32598
rect 978 32584 1030 32593
rect 1102 32584 1154 32593
rect 1226 32584 1278 32593
rect 978 32460 1030 32512
rect 1102 32460 1154 32512
rect 1226 32460 1278 32512
rect 978 32336 1030 32388
rect 1102 32336 1154 32388
rect 1226 32336 1278 32388
rect 978 32212 1030 32264
rect 1102 32212 1154 32264
rect 1226 32212 1278 32264
rect 978 32088 1030 32140
rect 1102 32088 1154 32140
rect 1226 32088 1278 32140
rect 978 31964 1030 32016
rect 1102 31964 1154 32016
rect 1226 31964 1278 32016
rect 978 31840 1030 31892
rect 1102 31840 1154 31892
rect 1226 31840 1278 31892
rect 978 31716 1030 31768
rect 1102 31716 1154 31768
rect 1226 31716 1278 31768
rect 978 31592 1030 31644
rect 1102 31592 1154 31644
rect 1226 31592 1278 31644
rect 978 31468 1030 31520
rect 1102 31468 1154 31520
rect 1226 31468 1278 31520
rect 978 31344 1030 31396
rect 1102 31344 1154 31396
rect 1226 31344 1278 31396
rect 978 31220 1030 31272
rect 1102 31220 1154 31272
rect 1226 31220 1278 31272
rect 978 31096 1030 31148
rect 1102 31096 1154 31148
rect 1226 31096 1278 31148
rect 978 30972 1030 31024
rect 1102 30972 1154 31024
rect 1226 30972 1278 31024
rect 978 30848 1030 30900
rect 1102 30848 1154 30900
rect 1226 30848 1278 30900
rect 978 30724 1030 30776
rect 1102 30724 1154 30776
rect 1226 30724 1278 30776
rect 978 30600 1030 30652
rect 1102 30600 1154 30652
rect 1226 30600 1278 30652
rect 978 30476 1030 30528
rect 1102 30476 1154 30528
rect 1226 30476 1278 30528
rect 978 30352 1030 30404
rect 1102 30352 1154 30404
rect 1226 30352 1278 30404
rect 978 30228 1030 30280
rect 1102 30228 1154 30280
rect 1226 30228 1278 30280
rect 978 30104 1030 30156
rect 1102 30104 1154 30156
rect 1226 30104 1278 30156
rect 978 29980 1030 30032
rect 1102 29980 1154 30032
rect 1226 29980 1278 30032
rect 978 29856 1030 29908
rect 1102 29856 1154 29908
rect 1226 29856 1278 29908
rect 978 29732 1030 29784
rect 1102 29732 1154 29784
rect 1226 29732 1278 29784
rect 978 29608 1030 29660
rect 1102 29608 1154 29660
rect 1226 29608 1278 29660
rect 3729 32546 3781 32593
rect 6335 32593 6387 32598
rect 3729 32438 3781 32490
rect 3729 32330 3781 32382
rect 3729 32222 3781 32274
rect 3729 32114 3781 32166
rect 3729 32006 3781 32058
rect 3729 31898 3781 31950
rect 3729 31790 3781 31842
rect 3729 31682 3781 31734
rect 3729 31574 3781 31626
rect 3729 31466 3781 31518
rect 3729 31358 3781 31410
rect 3729 31250 3781 31302
rect 3729 31142 3781 31194
rect 3729 31034 3781 31086
rect 3729 30926 3781 30978
rect 3729 30818 3781 30870
rect 3729 30710 3781 30762
rect 3729 30602 3781 30654
rect 3729 30494 3781 30546
rect 3729 30386 3781 30438
rect 3729 30278 3781 30330
rect 3729 30170 3781 30222
rect 3729 30062 3781 30114
rect 3729 29954 3781 30006
rect 3729 29846 3781 29898
rect 3729 29738 3781 29790
rect 3729 29630 3781 29682
rect 978 29527 1030 29536
rect 1102 29527 1154 29536
rect 1226 29527 1278 29536
rect 3729 29527 3781 29574
rect 978 29484 1030 29527
rect 1102 29484 1154 29527
rect 1226 29484 1278 29527
rect 3729 29522 3781 29527
rect 6335 32546 6387 32593
rect 8677 32593 8729 32598
rect 6335 32438 6387 32490
rect 6335 32330 6387 32382
rect 6335 32222 6387 32274
rect 6335 32114 6387 32166
rect 6335 32006 6387 32058
rect 6335 31898 6387 31950
rect 6335 31790 6387 31842
rect 6335 31682 6387 31734
rect 6335 31574 6387 31626
rect 6335 31466 6387 31518
rect 6335 31358 6387 31410
rect 6335 31250 6387 31302
rect 6335 31142 6387 31194
rect 6335 31034 6387 31086
rect 6335 30926 6387 30978
rect 6335 30818 6387 30870
rect 6335 30710 6387 30762
rect 6335 30602 6387 30654
rect 6335 30494 6387 30546
rect 6335 30386 6387 30438
rect 6335 30278 6387 30330
rect 6335 30170 6387 30222
rect 6335 30062 6387 30114
rect 6335 29954 6387 30006
rect 6335 29846 6387 29898
rect 6335 29738 6387 29790
rect 6335 29630 6387 29682
rect 6335 29527 6387 29574
rect 6335 29522 6387 29527
rect 7388 32523 7440 32544
rect 7388 32492 7389 32523
rect 7389 32492 7440 32523
rect 7624 32523 7676 32544
rect 7624 32492 7675 32523
rect 7675 32492 7676 32523
rect 7388 32384 7389 32436
rect 7389 32384 7440 32436
rect 7624 32384 7675 32436
rect 7675 32384 7676 32436
rect 7388 32276 7389 32328
rect 7389 32276 7440 32328
rect 7624 32276 7675 32328
rect 7675 32276 7676 32328
rect 7388 32168 7389 32220
rect 7389 32168 7440 32220
rect 7624 32168 7675 32220
rect 7675 32168 7676 32220
rect 7388 32060 7389 32112
rect 7389 32060 7440 32112
rect 7624 32060 7675 32112
rect 7675 32060 7676 32112
rect 7388 31952 7389 32004
rect 7389 31952 7440 32004
rect 7624 31952 7675 32004
rect 7675 31952 7676 32004
rect 7388 31844 7389 31896
rect 7389 31844 7440 31896
rect 7624 31844 7675 31896
rect 7675 31844 7676 31896
rect 7388 31736 7389 31788
rect 7389 31736 7440 31788
rect 7624 31736 7675 31788
rect 7675 31736 7676 31788
rect 7388 31628 7389 31680
rect 7389 31628 7440 31680
rect 7624 31628 7675 31680
rect 7675 31628 7676 31680
rect 7388 31520 7389 31572
rect 7389 31520 7440 31572
rect 7624 31520 7675 31572
rect 7675 31520 7676 31572
rect 7388 31412 7389 31464
rect 7389 31412 7440 31464
rect 7624 31412 7675 31464
rect 7675 31412 7676 31464
rect 7388 31304 7389 31356
rect 7389 31304 7440 31356
rect 7624 31304 7675 31356
rect 7675 31304 7676 31356
rect 7388 31196 7389 31248
rect 7389 31196 7440 31248
rect 7624 31196 7675 31248
rect 7675 31196 7676 31248
rect 7388 31088 7389 31140
rect 7389 31088 7440 31140
rect 7624 31088 7675 31140
rect 7675 31088 7676 31140
rect 7388 30980 7389 31032
rect 7389 30980 7440 31032
rect 7624 30980 7675 31032
rect 7675 30980 7676 31032
rect 7388 30872 7389 30924
rect 7389 30872 7440 30924
rect 7624 30872 7675 30924
rect 7675 30872 7676 30924
rect 7388 30764 7389 30816
rect 7389 30764 7440 30816
rect 7624 30764 7675 30816
rect 7675 30764 7676 30816
rect 7388 30656 7389 30708
rect 7389 30656 7440 30708
rect 7624 30656 7675 30708
rect 7675 30656 7676 30708
rect 7388 30548 7389 30600
rect 7389 30548 7440 30600
rect 7624 30548 7675 30600
rect 7675 30548 7676 30600
rect 7388 30440 7389 30492
rect 7389 30440 7440 30492
rect 7624 30440 7675 30492
rect 7675 30440 7676 30492
rect 7388 30332 7389 30384
rect 7389 30332 7440 30384
rect 7624 30332 7675 30384
rect 7675 30332 7676 30384
rect 7388 30224 7389 30276
rect 7389 30224 7440 30276
rect 7624 30224 7675 30276
rect 7675 30224 7676 30276
rect 7388 30116 7389 30168
rect 7389 30116 7440 30168
rect 7624 30116 7675 30168
rect 7675 30116 7676 30168
rect 7388 30008 7389 30060
rect 7389 30008 7440 30060
rect 7624 30008 7675 30060
rect 7675 30008 7676 30060
rect 7388 29900 7389 29952
rect 7389 29900 7440 29952
rect 7624 29900 7675 29952
rect 7675 29900 7676 29952
rect 7388 29792 7389 29844
rect 7389 29792 7440 29844
rect 7624 29792 7675 29844
rect 7675 29792 7676 29844
rect 7388 29684 7389 29736
rect 7389 29684 7440 29736
rect 7624 29684 7675 29736
rect 7675 29684 7676 29736
rect 7388 29597 7389 29628
rect 7389 29597 7440 29628
rect 7388 29576 7440 29597
rect 7624 29597 7675 29628
rect 7675 29597 7676 29628
rect 7624 29576 7676 29597
rect 8677 32546 8729 32593
rect 8677 32438 8729 32490
rect 8677 32330 8729 32382
rect 8677 32222 8729 32274
rect 8677 32114 8729 32166
rect 8677 32006 8729 32058
rect 8677 31898 8729 31950
rect 8677 31790 8729 31842
rect 8677 31682 8729 31734
rect 8677 31574 8729 31626
rect 8677 31466 8729 31518
rect 8677 31358 8729 31410
rect 8677 31250 8729 31302
rect 8677 31142 8729 31194
rect 8677 31034 8729 31086
rect 8677 30926 8729 30978
rect 8677 30818 8729 30870
rect 8677 30710 8729 30762
rect 8677 30602 8729 30654
rect 8677 30494 8729 30546
rect 8677 30386 8729 30438
rect 8677 30278 8729 30330
rect 8677 30170 8729 30222
rect 8677 30062 8729 30114
rect 8677 29954 8729 30006
rect 8677 29846 8729 29898
rect 8677 29738 8729 29790
rect 8677 29630 8729 29682
rect 8677 29527 8729 29574
rect 11283 32593 11335 32598
rect 13786 32593 13838 32636
rect 13910 32593 13962 32636
rect 14034 32593 14086 32636
rect 8677 29522 8729 29527
rect 11283 32546 11335 32593
rect 13786 32584 13838 32593
rect 13910 32584 13962 32593
rect 14034 32584 14086 32593
rect 11283 32438 11335 32490
rect 11283 32330 11335 32382
rect 11283 32222 11335 32274
rect 11283 32114 11335 32166
rect 11283 32006 11335 32058
rect 11283 31898 11335 31950
rect 11283 31790 11335 31842
rect 11283 31682 11335 31734
rect 11283 31574 11335 31626
rect 11283 31466 11335 31518
rect 11283 31358 11335 31410
rect 11283 31250 11335 31302
rect 11283 31142 11335 31194
rect 11283 31034 11335 31086
rect 11283 30926 11335 30978
rect 11283 30818 11335 30870
rect 11283 30710 11335 30762
rect 11283 30602 11335 30654
rect 11283 30494 11335 30546
rect 11283 30386 11335 30438
rect 11283 30278 11335 30330
rect 11283 30170 11335 30222
rect 11283 30062 11335 30114
rect 11283 29954 11335 30006
rect 11283 29846 11335 29898
rect 11283 29738 11335 29790
rect 11283 29630 11335 29682
rect 11283 29527 11335 29574
rect 13786 32460 13838 32512
rect 13910 32460 13962 32512
rect 14034 32460 14086 32512
rect 13786 32336 13838 32388
rect 13910 32336 13962 32388
rect 14034 32336 14086 32388
rect 13786 32212 13838 32264
rect 13910 32212 13962 32264
rect 14034 32212 14086 32264
rect 13786 32088 13838 32140
rect 13910 32088 13962 32140
rect 14034 32088 14086 32140
rect 13786 31964 13838 32016
rect 13910 31964 13962 32016
rect 14034 31964 14086 32016
rect 13786 31840 13838 31892
rect 13910 31840 13962 31892
rect 14034 31840 14086 31892
rect 13786 31716 13838 31768
rect 13910 31716 13962 31768
rect 14034 31716 14086 31768
rect 13786 31592 13838 31644
rect 13910 31592 13962 31644
rect 14034 31592 14086 31644
rect 13786 31468 13838 31520
rect 13910 31468 13962 31520
rect 14034 31468 14086 31520
rect 13786 31344 13838 31396
rect 13910 31344 13962 31396
rect 14034 31344 14086 31396
rect 13786 31220 13838 31272
rect 13910 31220 13962 31272
rect 14034 31220 14086 31272
rect 13786 31096 13838 31148
rect 13910 31096 13962 31148
rect 14034 31096 14086 31148
rect 13786 30972 13838 31024
rect 13910 30972 13962 31024
rect 14034 30972 14086 31024
rect 13786 30848 13838 30900
rect 13910 30848 13962 30900
rect 14034 30848 14086 30900
rect 13786 30724 13838 30776
rect 13910 30724 13962 30776
rect 14034 30724 14086 30776
rect 13786 30600 13838 30652
rect 13910 30600 13962 30652
rect 14034 30600 14086 30652
rect 13786 30476 13838 30528
rect 13910 30476 13962 30528
rect 14034 30476 14086 30528
rect 13786 30352 13838 30404
rect 13910 30352 13962 30404
rect 14034 30352 14086 30404
rect 13786 30228 13838 30280
rect 13910 30228 13962 30280
rect 14034 30228 14086 30280
rect 13786 30104 13838 30156
rect 13910 30104 13962 30156
rect 14034 30104 14086 30156
rect 13786 29980 13838 30032
rect 13910 29980 13962 30032
rect 14034 29980 14086 30032
rect 13786 29856 13838 29908
rect 13910 29856 13962 29908
rect 14034 29856 14086 29908
rect 13786 29732 13838 29784
rect 13910 29732 13962 29784
rect 14034 29732 14086 29784
rect 13786 29608 13838 29660
rect 13910 29608 13962 29660
rect 14034 29608 14086 29660
rect 13786 29527 13838 29536
rect 13910 29527 13962 29536
rect 14034 29527 14086 29536
rect 11283 29522 11335 29527
rect 13786 29484 13838 29527
rect 13910 29484 13962 29527
rect 14034 29484 14086 29527
rect 444 29276 445 29328
rect 445 29276 496 29328
rect 552 29276 604 29328
rect 660 29276 712 29328
rect 1438 29308 1490 29360
rect 1562 29308 1614 29360
rect 1686 29308 1738 29360
rect 1810 29308 1862 29360
rect 2574 29308 2626 29360
rect 2698 29308 2750 29360
rect 2822 29308 2874 29360
rect 2946 29308 2998 29360
rect 4846 29308 4898 29360
rect 4970 29308 5022 29360
rect 5094 29308 5146 29360
rect 5218 29308 5270 29360
rect 7139 29308 7191 29360
rect 7263 29308 7315 29360
rect 7387 29308 7439 29360
rect 7625 29308 7677 29360
rect 7749 29308 7801 29360
rect 7873 29308 7925 29360
rect 9794 29308 9846 29360
rect 9918 29308 9970 29360
rect 10042 29308 10094 29360
rect 10166 29308 10218 29360
rect 12066 29308 12118 29360
rect 12190 29308 12242 29360
rect 12314 29308 12366 29360
rect 12438 29308 12490 29360
rect 13202 29308 13254 29360
rect 13326 29308 13378 29360
rect 13450 29308 13502 29360
rect 13574 29308 13626 29360
rect 14352 29276 14404 29328
rect 14460 29276 14512 29328
rect 14568 29276 14619 29328
rect 14619 29276 14620 29328
rect 444 29168 445 29220
rect 445 29168 496 29220
rect 552 29168 604 29220
rect 660 29168 712 29220
rect 1438 29184 1490 29236
rect 1562 29184 1614 29236
rect 1686 29184 1738 29236
rect 1810 29184 1862 29236
rect 2574 29184 2626 29236
rect 2698 29184 2750 29236
rect 2822 29184 2874 29236
rect 2946 29184 2998 29236
rect 4846 29184 4898 29236
rect 4970 29184 5022 29236
rect 5094 29184 5146 29236
rect 5218 29184 5270 29236
rect 7139 29184 7191 29236
rect 7263 29184 7315 29236
rect 7387 29184 7439 29236
rect 7625 29184 7677 29236
rect 7749 29184 7801 29236
rect 7873 29184 7925 29236
rect 9794 29184 9846 29236
rect 9918 29184 9970 29236
rect 10042 29184 10094 29236
rect 10166 29184 10218 29236
rect 12066 29184 12118 29236
rect 12190 29184 12242 29236
rect 12314 29184 12366 29236
rect 12438 29184 12490 29236
rect 13202 29184 13254 29236
rect 13326 29184 13378 29236
rect 13450 29184 13502 29236
rect 13574 29184 13626 29236
rect 14352 29168 14404 29220
rect 14460 29168 14512 29220
rect 14568 29168 14619 29220
rect 14619 29168 14620 29220
rect 444 29060 445 29112
rect 445 29060 496 29112
rect 552 29109 604 29112
rect 660 29109 712 29112
rect 1438 29109 1490 29112
rect 1562 29109 1614 29112
rect 1686 29109 1738 29112
rect 1810 29109 1862 29112
rect 2574 29109 2626 29112
rect 2698 29109 2750 29112
rect 2822 29109 2874 29112
rect 2946 29109 2998 29112
rect 4846 29109 4898 29112
rect 4970 29109 5022 29112
rect 5094 29109 5146 29112
rect 5218 29109 5270 29112
rect 7139 29109 7191 29112
rect 7263 29109 7315 29112
rect 7387 29109 7439 29112
rect 7625 29109 7677 29112
rect 7749 29109 7801 29112
rect 7873 29109 7925 29112
rect 9794 29109 9846 29112
rect 9918 29109 9970 29112
rect 10042 29109 10094 29112
rect 10166 29109 10218 29112
rect 12066 29109 12118 29112
rect 12190 29109 12242 29112
rect 12314 29109 12366 29112
rect 12438 29109 12490 29112
rect 13202 29109 13254 29112
rect 13326 29109 13378 29112
rect 13450 29109 13502 29112
rect 13574 29109 13626 29112
rect 14352 29109 14404 29112
rect 14460 29109 14512 29112
rect 552 29063 553 29109
rect 553 29063 604 29109
rect 660 29063 712 29109
rect 1438 29063 1490 29109
rect 1562 29063 1614 29109
rect 1686 29063 1738 29109
rect 1810 29063 1862 29109
rect 2574 29063 2626 29109
rect 2698 29063 2750 29109
rect 2822 29063 2874 29109
rect 2946 29063 2998 29109
rect 4846 29063 4898 29109
rect 4970 29063 5022 29109
rect 5094 29063 5146 29109
rect 5218 29063 5270 29109
rect 7139 29063 7191 29109
rect 7263 29063 7315 29109
rect 7387 29063 7439 29109
rect 7625 29063 7677 29109
rect 7749 29063 7801 29109
rect 7873 29063 7925 29109
rect 9794 29063 9846 29109
rect 9918 29063 9970 29109
rect 10042 29063 10094 29109
rect 10166 29063 10218 29109
rect 12066 29063 12118 29109
rect 12190 29063 12242 29109
rect 12314 29063 12366 29109
rect 12438 29063 12490 29109
rect 13202 29063 13254 29109
rect 13326 29063 13378 29109
rect 13450 29063 13502 29109
rect 13574 29063 13626 29109
rect 14352 29063 14404 29109
rect 14460 29063 14511 29109
rect 14511 29063 14512 29109
rect 552 29060 604 29063
rect 660 29060 712 29063
rect 1438 29060 1490 29063
rect 1562 29060 1614 29063
rect 1686 29060 1738 29063
rect 1810 29060 1862 29063
rect 2574 29060 2626 29063
rect 2698 29060 2750 29063
rect 2822 29060 2874 29063
rect 2946 29060 2998 29063
rect 4846 29060 4898 29063
rect 4970 29060 5022 29063
rect 5094 29060 5146 29063
rect 5218 29060 5270 29063
rect 7139 29060 7191 29063
rect 7263 29060 7315 29063
rect 7387 29060 7439 29063
rect 7625 29060 7677 29063
rect 7749 29060 7801 29063
rect 7873 29060 7925 29063
rect 9794 29060 9846 29063
rect 9918 29060 9970 29063
rect 10042 29060 10094 29063
rect 10166 29060 10218 29063
rect 12066 29060 12118 29063
rect 12190 29060 12242 29063
rect 12314 29060 12366 29063
rect 12438 29060 12490 29063
rect 13202 29060 13254 29063
rect 13326 29060 13378 29063
rect 13450 29060 13502 29063
rect 13574 29060 13626 29063
rect 14352 29060 14404 29063
rect 14460 29060 14512 29063
rect 14568 29060 14619 29112
rect 14619 29060 14620 29112
rect 444 28952 445 29004
rect 445 28952 496 29004
rect 552 28952 604 29004
rect 660 28952 712 29004
rect 1438 28936 1490 28988
rect 1562 28936 1614 28988
rect 1686 28936 1738 28988
rect 1810 28936 1862 28988
rect 2574 28936 2626 28988
rect 2698 28936 2750 28988
rect 2822 28936 2874 28988
rect 2946 28936 2998 28988
rect 4846 28936 4898 28988
rect 4970 28936 5022 28988
rect 5094 28936 5146 28988
rect 5218 28936 5270 28988
rect 7139 28936 7191 28988
rect 7263 28936 7315 28988
rect 7387 28936 7439 28988
rect 7625 28936 7677 28988
rect 7749 28936 7801 28988
rect 7873 28936 7925 28988
rect 9794 28936 9846 28988
rect 9918 28936 9970 28988
rect 10042 28936 10094 28988
rect 10166 28936 10218 28988
rect 12066 28936 12118 28988
rect 12190 28936 12242 28988
rect 12314 28936 12366 28988
rect 12438 28936 12490 28988
rect 13202 28936 13254 28988
rect 13326 28936 13378 28988
rect 13450 28936 13502 28988
rect 13574 28936 13626 28988
rect 14352 28952 14404 29004
rect 14460 28952 14512 29004
rect 14568 28952 14619 29004
rect 14619 28952 14620 29004
rect 444 28844 445 28896
rect 445 28844 496 28896
rect 552 28844 604 28896
rect 660 28844 712 28896
rect 1438 28812 1490 28864
rect 1562 28812 1614 28864
rect 1686 28812 1738 28864
rect 1810 28812 1862 28864
rect 2574 28812 2626 28864
rect 2698 28812 2750 28864
rect 2822 28812 2874 28864
rect 2946 28812 2998 28864
rect 4846 28812 4898 28864
rect 4970 28812 5022 28864
rect 5094 28812 5146 28864
rect 5218 28812 5270 28864
rect 7139 28812 7191 28864
rect 7263 28812 7315 28864
rect 7387 28812 7439 28864
rect 7625 28812 7677 28864
rect 7749 28812 7801 28864
rect 7873 28812 7925 28864
rect 9794 28812 9846 28864
rect 9918 28812 9970 28864
rect 10042 28812 10094 28864
rect 10166 28812 10218 28864
rect 12066 28812 12118 28864
rect 12190 28812 12242 28864
rect 12314 28812 12366 28864
rect 12438 28812 12490 28864
rect 13202 28812 13254 28864
rect 13326 28812 13378 28864
rect 13450 28812 13502 28864
rect 13574 28812 13626 28864
rect 14352 28844 14404 28896
rect 14460 28844 14512 28896
rect 14568 28844 14619 28896
rect 14619 28844 14620 28896
rect 978 28645 1030 28688
rect 1102 28645 1154 28688
rect 1226 28645 1278 28688
rect 3729 28645 3781 28650
rect 978 28636 1030 28645
rect 1102 28636 1154 28645
rect 1226 28636 1278 28645
rect 978 28512 1030 28564
rect 1102 28512 1154 28564
rect 1226 28512 1278 28564
rect 978 28388 1030 28440
rect 1102 28388 1154 28440
rect 1226 28388 1278 28440
rect 978 28264 1030 28316
rect 1102 28264 1154 28316
rect 1226 28264 1278 28316
rect 978 28140 1030 28192
rect 1102 28140 1154 28192
rect 1226 28140 1278 28192
rect 978 28016 1030 28068
rect 1102 28016 1154 28068
rect 1226 28016 1278 28068
rect 978 27892 1030 27944
rect 1102 27892 1154 27944
rect 1226 27892 1278 27944
rect 978 27768 1030 27820
rect 1102 27768 1154 27820
rect 1226 27768 1278 27820
rect 978 27644 1030 27696
rect 1102 27644 1154 27696
rect 1226 27644 1278 27696
rect 978 27520 1030 27572
rect 1102 27520 1154 27572
rect 1226 27520 1278 27572
rect 978 27396 1030 27448
rect 1102 27396 1154 27448
rect 1226 27396 1278 27448
rect 978 27272 1030 27324
rect 1102 27272 1154 27324
rect 1226 27272 1278 27324
rect 978 27148 1030 27200
rect 1102 27148 1154 27200
rect 1226 27148 1278 27200
rect 978 27024 1030 27076
rect 1102 27024 1154 27076
rect 1226 27024 1278 27076
rect 978 26900 1030 26952
rect 1102 26900 1154 26952
rect 1226 26900 1278 26952
rect 978 26776 1030 26828
rect 1102 26776 1154 26828
rect 1226 26776 1278 26828
rect 978 26652 1030 26704
rect 1102 26652 1154 26704
rect 1226 26652 1278 26704
rect 978 26528 1030 26580
rect 1102 26528 1154 26580
rect 1226 26528 1278 26580
rect 978 26404 1030 26456
rect 1102 26404 1154 26456
rect 1226 26404 1278 26456
rect 978 26280 1030 26332
rect 1102 26280 1154 26332
rect 1226 26280 1278 26332
rect 978 26156 1030 26208
rect 1102 26156 1154 26208
rect 1226 26156 1278 26208
rect 978 26032 1030 26084
rect 1102 26032 1154 26084
rect 1226 26032 1278 26084
rect 978 25908 1030 25960
rect 1102 25908 1154 25960
rect 1226 25908 1278 25960
rect 978 25784 1030 25836
rect 1102 25784 1154 25836
rect 1226 25784 1278 25836
rect 978 25660 1030 25712
rect 1102 25660 1154 25712
rect 1226 25660 1278 25712
rect 3729 28598 3781 28645
rect 6335 28645 6387 28650
rect 3729 28490 3781 28542
rect 3729 28382 3781 28434
rect 3729 28274 3781 28326
rect 3729 28166 3781 28218
rect 3729 28058 3781 28110
rect 3729 27950 3781 28002
rect 3729 27842 3781 27894
rect 3729 27734 3781 27786
rect 3729 27626 3781 27678
rect 3729 27518 3781 27570
rect 3729 27410 3781 27462
rect 3729 27302 3781 27354
rect 3729 27194 3781 27246
rect 3729 27086 3781 27138
rect 3729 26978 3781 27030
rect 3729 26870 3781 26922
rect 3729 26762 3781 26814
rect 3729 26654 3781 26706
rect 3729 26546 3781 26598
rect 3729 26438 3781 26490
rect 3729 26330 3781 26382
rect 3729 26222 3781 26274
rect 3729 26114 3781 26166
rect 3729 26006 3781 26058
rect 3729 25898 3781 25950
rect 3729 25790 3781 25842
rect 3729 25682 3781 25734
rect 978 25579 1030 25588
rect 1102 25579 1154 25588
rect 1226 25579 1278 25588
rect 3729 25579 3781 25626
rect 978 25536 1030 25579
rect 1102 25536 1154 25579
rect 1226 25536 1278 25579
rect 3729 25574 3781 25579
rect 6335 28598 6387 28645
rect 8677 28645 8729 28650
rect 6335 28490 6387 28542
rect 6335 28382 6387 28434
rect 6335 28274 6387 28326
rect 6335 28166 6387 28218
rect 6335 28058 6387 28110
rect 6335 27950 6387 28002
rect 6335 27842 6387 27894
rect 6335 27734 6387 27786
rect 6335 27626 6387 27678
rect 6335 27518 6387 27570
rect 6335 27410 6387 27462
rect 6335 27302 6387 27354
rect 6335 27194 6387 27246
rect 6335 27086 6387 27138
rect 6335 26978 6387 27030
rect 6335 26870 6387 26922
rect 6335 26762 6387 26814
rect 6335 26654 6387 26706
rect 6335 26546 6387 26598
rect 6335 26438 6387 26490
rect 6335 26330 6387 26382
rect 6335 26222 6387 26274
rect 6335 26114 6387 26166
rect 6335 26006 6387 26058
rect 6335 25898 6387 25950
rect 6335 25790 6387 25842
rect 6335 25682 6387 25734
rect 6335 25579 6387 25626
rect 6335 25574 6387 25579
rect 7388 28575 7440 28596
rect 7388 28544 7389 28575
rect 7389 28544 7440 28575
rect 7624 28575 7676 28596
rect 7624 28544 7675 28575
rect 7675 28544 7676 28575
rect 7388 28436 7389 28488
rect 7389 28436 7440 28488
rect 7624 28436 7675 28488
rect 7675 28436 7676 28488
rect 7388 28328 7389 28380
rect 7389 28328 7440 28380
rect 7624 28328 7675 28380
rect 7675 28328 7676 28380
rect 7388 28220 7389 28272
rect 7389 28220 7440 28272
rect 7624 28220 7675 28272
rect 7675 28220 7676 28272
rect 7388 28112 7389 28164
rect 7389 28112 7440 28164
rect 7624 28112 7675 28164
rect 7675 28112 7676 28164
rect 7388 28004 7389 28056
rect 7389 28004 7440 28056
rect 7624 28004 7675 28056
rect 7675 28004 7676 28056
rect 7388 27896 7389 27948
rect 7389 27896 7440 27948
rect 7624 27896 7675 27948
rect 7675 27896 7676 27948
rect 7388 27788 7389 27840
rect 7389 27788 7440 27840
rect 7624 27788 7675 27840
rect 7675 27788 7676 27840
rect 7388 27680 7389 27732
rect 7389 27680 7440 27732
rect 7624 27680 7675 27732
rect 7675 27680 7676 27732
rect 7388 27572 7389 27624
rect 7389 27572 7440 27624
rect 7624 27572 7675 27624
rect 7675 27572 7676 27624
rect 7388 27464 7389 27516
rect 7389 27464 7440 27516
rect 7624 27464 7675 27516
rect 7675 27464 7676 27516
rect 7388 27356 7389 27408
rect 7389 27356 7440 27408
rect 7624 27356 7675 27408
rect 7675 27356 7676 27408
rect 7388 27248 7389 27300
rect 7389 27248 7440 27300
rect 7624 27248 7675 27300
rect 7675 27248 7676 27300
rect 7388 27140 7389 27192
rect 7389 27140 7440 27192
rect 7624 27140 7675 27192
rect 7675 27140 7676 27192
rect 7388 27032 7389 27084
rect 7389 27032 7440 27084
rect 7624 27032 7675 27084
rect 7675 27032 7676 27084
rect 7388 26924 7389 26976
rect 7389 26924 7440 26976
rect 7624 26924 7675 26976
rect 7675 26924 7676 26976
rect 7388 26816 7389 26868
rect 7389 26816 7440 26868
rect 7624 26816 7675 26868
rect 7675 26816 7676 26868
rect 7388 26708 7389 26760
rect 7389 26708 7440 26760
rect 7624 26708 7675 26760
rect 7675 26708 7676 26760
rect 7388 26600 7389 26652
rect 7389 26600 7440 26652
rect 7624 26600 7675 26652
rect 7675 26600 7676 26652
rect 7388 26492 7389 26544
rect 7389 26492 7440 26544
rect 7624 26492 7675 26544
rect 7675 26492 7676 26544
rect 7388 26384 7389 26436
rect 7389 26384 7440 26436
rect 7624 26384 7675 26436
rect 7675 26384 7676 26436
rect 7388 26276 7389 26328
rect 7389 26276 7440 26328
rect 7624 26276 7675 26328
rect 7675 26276 7676 26328
rect 7388 26168 7389 26220
rect 7389 26168 7440 26220
rect 7624 26168 7675 26220
rect 7675 26168 7676 26220
rect 7388 26060 7389 26112
rect 7389 26060 7440 26112
rect 7624 26060 7675 26112
rect 7675 26060 7676 26112
rect 7388 25952 7389 26004
rect 7389 25952 7440 26004
rect 7624 25952 7675 26004
rect 7675 25952 7676 26004
rect 7388 25844 7389 25896
rect 7389 25844 7440 25896
rect 7624 25844 7675 25896
rect 7675 25844 7676 25896
rect 7388 25736 7389 25788
rect 7389 25736 7440 25788
rect 7624 25736 7675 25788
rect 7675 25736 7676 25788
rect 7388 25649 7389 25680
rect 7389 25649 7440 25680
rect 7388 25628 7440 25649
rect 7624 25649 7675 25680
rect 7675 25649 7676 25680
rect 7624 25628 7676 25649
rect 8677 28598 8729 28645
rect 8677 28490 8729 28542
rect 8677 28382 8729 28434
rect 8677 28274 8729 28326
rect 8677 28166 8729 28218
rect 8677 28058 8729 28110
rect 8677 27950 8729 28002
rect 8677 27842 8729 27894
rect 8677 27734 8729 27786
rect 8677 27626 8729 27678
rect 8677 27518 8729 27570
rect 8677 27410 8729 27462
rect 8677 27302 8729 27354
rect 8677 27194 8729 27246
rect 8677 27086 8729 27138
rect 8677 26978 8729 27030
rect 8677 26870 8729 26922
rect 8677 26762 8729 26814
rect 8677 26654 8729 26706
rect 8677 26546 8729 26598
rect 8677 26438 8729 26490
rect 8677 26330 8729 26382
rect 8677 26222 8729 26274
rect 8677 26114 8729 26166
rect 8677 26006 8729 26058
rect 8677 25898 8729 25950
rect 8677 25790 8729 25842
rect 8677 25682 8729 25734
rect 8677 25579 8729 25626
rect 11283 28645 11335 28650
rect 13786 28645 13838 28688
rect 13910 28645 13962 28688
rect 14034 28645 14086 28688
rect 8677 25574 8729 25579
rect 11283 28598 11335 28645
rect 13786 28636 13838 28645
rect 13910 28636 13962 28645
rect 14034 28636 14086 28645
rect 11283 28490 11335 28542
rect 11283 28382 11335 28434
rect 11283 28274 11335 28326
rect 11283 28166 11335 28218
rect 11283 28058 11335 28110
rect 11283 27950 11335 28002
rect 11283 27842 11335 27894
rect 11283 27734 11335 27786
rect 11283 27626 11335 27678
rect 11283 27518 11335 27570
rect 11283 27410 11335 27462
rect 11283 27302 11335 27354
rect 11283 27194 11335 27246
rect 11283 27086 11335 27138
rect 11283 26978 11335 27030
rect 11283 26870 11335 26922
rect 11283 26762 11335 26814
rect 11283 26654 11335 26706
rect 11283 26546 11335 26598
rect 11283 26438 11335 26490
rect 11283 26330 11335 26382
rect 11283 26222 11335 26274
rect 11283 26114 11335 26166
rect 11283 26006 11335 26058
rect 11283 25898 11335 25950
rect 11283 25790 11335 25842
rect 11283 25682 11335 25734
rect 11283 25579 11335 25626
rect 13786 28512 13838 28564
rect 13910 28512 13962 28564
rect 14034 28512 14086 28564
rect 13786 28388 13838 28440
rect 13910 28388 13962 28440
rect 14034 28388 14086 28440
rect 13786 28264 13838 28316
rect 13910 28264 13962 28316
rect 14034 28264 14086 28316
rect 13786 28140 13838 28192
rect 13910 28140 13962 28192
rect 14034 28140 14086 28192
rect 13786 28016 13838 28068
rect 13910 28016 13962 28068
rect 14034 28016 14086 28068
rect 13786 27892 13838 27944
rect 13910 27892 13962 27944
rect 14034 27892 14086 27944
rect 13786 27768 13838 27820
rect 13910 27768 13962 27820
rect 14034 27768 14086 27820
rect 13786 27644 13838 27696
rect 13910 27644 13962 27696
rect 14034 27644 14086 27696
rect 13786 27520 13838 27572
rect 13910 27520 13962 27572
rect 14034 27520 14086 27572
rect 13786 27396 13838 27448
rect 13910 27396 13962 27448
rect 14034 27396 14086 27448
rect 13786 27272 13838 27324
rect 13910 27272 13962 27324
rect 14034 27272 14086 27324
rect 13786 27148 13838 27200
rect 13910 27148 13962 27200
rect 14034 27148 14086 27200
rect 13786 27024 13838 27076
rect 13910 27024 13962 27076
rect 14034 27024 14086 27076
rect 13786 26900 13838 26952
rect 13910 26900 13962 26952
rect 14034 26900 14086 26952
rect 13786 26776 13838 26828
rect 13910 26776 13962 26828
rect 14034 26776 14086 26828
rect 13786 26652 13838 26704
rect 13910 26652 13962 26704
rect 14034 26652 14086 26704
rect 13786 26528 13838 26580
rect 13910 26528 13962 26580
rect 14034 26528 14086 26580
rect 13786 26404 13838 26456
rect 13910 26404 13962 26456
rect 14034 26404 14086 26456
rect 13786 26280 13838 26332
rect 13910 26280 13962 26332
rect 14034 26280 14086 26332
rect 13786 26156 13838 26208
rect 13910 26156 13962 26208
rect 14034 26156 14086 26208
rect 13786 26032 13838 26084
rect 13910 26032 13962 26084
rect 14034 26032 14086 26084
rect 13786 25908 13838 25960
rect 13910 25908 13962 25960
rect 14034 25908 14086 25960
rect 13786 25784 13838 25836
rect 13910 25784 13962 25836
rect 14034 25784 14086 25836
rect 13786 25660 13838 25712
rect 13910 25660 13962 25712
rect 14034 25660 14086 25712
rect 13786 25579 13838 25588
rect 13910 25579 13962 25588
rect 14034 25579 14086 25588
rect 11283 25574 11335 25579
rect 13786 25536 13838 25579
rect 13910 25536 13962 25579
rect 14034 25536 14086 25579
rect 444 25328 445 25380
rect 445 25328 496 25380
rect 552 25328 604 25380
rect 660 25328 712 25380
rect 1438 25360 1490 25412
rect 1562 25360 1614 25412
rect 1686 25360 1738 25412
rect 1810 25360 1862 25412
rect 2574 25360 2626 25412
rect 2698 25360 2750 25412
rect 2822 25360 2874 25412
rect 2946 25360 2998 25412
rect 4846 25360 4898 25412
rect 4970 25360 5022 25412
rect 5094 25360 5146 25412
rect 5218 25360 5270 25412
rect 7139 25360 7191 25412
rect 7263 25360 7315 25412
rect 7387 25360 7439 25412
rect 7625 25360 7677 25412
rect 7749 25360 7801 25412
rect 7873 25360 7925 25412
rect 9794 25360 9846 25412
rect 9918 25360 9970 25412
rect 10042 25360 10094 25412
rect 10166 25360 10218 25412
rect 12066 25360 12118 25412
rect 12190 25360 12242 25412
rect 12314 25360 12366 25412
rect 12438 25360 12490 25412
rect 13202 25360 13254 25412
rect 13326 25360 13378 25412
rect 13450 25360 13502 25412
rect 13574 25360 13626 25412
rect 14352 25328 14404 25380
rect 14460 25328 14512 25380
rect 14568 25328 14619 25380
rect 14619 25328 14620 25380
rect 444 25220 445 25272
rect 445 25220 496 25272
rect 552 25220 604 25272
rect 660 25220 712 25272
rect 1438 25236 1490 25288
rect 1562 25236 1614 25288
rect 1686 25236 1738 25288
rect 1810 25236 1862 25288
rect 2574 25236 2626 25288
rect 2698 25236 2750 25288
rect 2822 25236 2874 25288
rect 2946 25236 2998 25288
rect 4846 25236 4898 25288
rect 4970 25236 5022 25288
rect 5094 25236 5146 25288
rect 5218 25236 5270 25288
rect 7139 25236 7191 25288
rect 7263 25236 7315 25288
rect 7387 25236 7439 25288
rect 7625 25236 7677 25288
rect 7749 25236 7801 25288
rect 7873 25236 7925 25288
rect 9794 25236 9846 25288
rect 9918 25236 9970 25288
rect 10042 25236 10094 25288
rect 10166 25236 10218 25288
rect 12066 25236 12118 25288
rect 12190 25236 12242 25288
rect 12314 25236 12366 25288
rect 12438 25236 12490 25288
rect 13202 25236 13254 25288
rect 13326 25236 13378 25288
rect 13450 25236 13502 25288
rect 13574 25236 13626 25288
rect 14352 25220 14404 25272
rect 14460 25220 14512 25272
rect 14568 25220 14619 25272
rect 14619 25220 14620 25272
rect 444 25112 445 25164
rect 445 25112 496 25164
rect 552 25161 604 25164
rect 660 25161 712 25164
rect 1438 25161 1490 25164
rect 1562 25161 1614 25164
rect 1686 25161 1738 25164
rect 1810 25161 1862 25164
rect 2574 25161 2626 25164
rect 2698 25161 2750 25164
rect 2822 25161 2874 25164
rect 2946 25161 2998 25164
rect 4846 25161 4898 25164
rect 4970 25161 5022 25164
rect 5094 25161 5146 25164
rect 5218 25161 5270 25164
rect 7139 25161 7191 25164
rect 7263 25161 7315 25164
rect 7387 25161 7439 25164
rect 7625 25161 7677 25164
rect 7749 25161 7801 25164
rect 7873 25161 7925 25164
rect 9794 25161 9846 25164
rect 9918 25161 9970 25164
rect 10042 25161 10094 25164
rect 10166 25161 10218 25164
rect 12066 25161 12118 25164
rect 12190 25161 12242 25164
rect 12314 25161 12366 25164
rect 12438 25161 12490 25164
rect 13202 25161 13254 25164
rect 13326 25161 13378 25164
rect 13450 25161 13502 25164
rect 13574 25161 13626 25164
rect 14352 25161 14404 25164
rect 14460 25161 14512 25164
rect 552 25115 553 25161
rect 553 25115 604 25161
rect 660 25115 712 25161
rect 1438 25115 1490 25161
rect 1562 25115 1614 25161
rect 1686 25115 1738 25161
rect 1810 25115 1862 25161
rect 2574 25115 2626 25161
rect 2698 25115 2750 25161
rect 2822 25115 2874 25161
rect 2946 25115 2998 25161
rect 4846 25115 4898 25161
rect 4970 25115 5022 25161
rect 5094 25115 5146 25161
rect 5218 25115 5270 25161
rect 7139 25115 7191 25161
rect 7263 25115 7315 25161
rect 7387 25115 7439 25161
rect 7625 25115 7677 25161
rect 7749 25115 7801 25161
rect 7873 25115 7925 25161
rect 9794 25115 9846 25161
rect 9918 25115 9970 25161
rect 10042 25115 10094 25161
rect 10166 25115 10218 25161
rect 12066 25115 12118 25161
rect 12190 25115 12242 25161
rect 12314 25115 12366 25161
rect 12438 25115 12490 25161
rect 13202 25115 13254 25161
rect 13326 25115 13378 25161
rect 13450 25115 13502 25161
rect 13574 25115 13626 25161
rect 14352 25115 14404 25161
rect 14460 25115 14511 25161
rect 14511 25115 14512 25161
rect 552 25112 604 25115
rect 660 25112 712 25115
rect 1438 25112 1490 25115
rect 1562 25112 1614 25115
rect 1686 25112 1738 25115
rect 1810 25112 1862 25115
rect 2574 25112 2626 25115
rect 2698 25112 2750 25115
rect 2822 25112 2874 25115
rect 2946 25112 2998 25115
rect 4846 25112 4898 25115
rect 4970 25112 5022 25115
rect 5094 25112 5146 25115
rect 5218 25112 5270 25115
rect 7139 25112 7191 25115
rect 7263 25112 7315 25115
rect 7387 25112 7439 25115
rect 7625 25112 7677 25115
rect 7749 25112 7801 25115
rect 7873 25112 7925 25115
rect 9794 25112 9846 25115
rect 9918 25112 9970 25115
rect 10042 25112 10094 25115
rect 10166 25112 10218 25115
rect 12066 25112 12118 25115
rect 12190 25112 12242 25115
rect 12314 25112 12366 25115
rect 12438 25112 12490 25115
rect 13202 25112 13254 25115
rect 13326 25112 13378 25115
rect 13450 25112 13502 25115
rect 13574 25112 13626 25115
rect 14352 25112 14404 25115
rect 14460 25112 14512 25115
rect 14568 25112 14619 25164
rect 14619 25112 14620 25164
rect 444 25004 445 25056
rect 445 25004 496 25056
rect 552 25004 604 25056
rect 660 25004 712 25056
rect 1438 24988 1490 25040
rect 1562 24988 1614 25040
rect 1686 24988 1738 25040
rect 1810 24988 1862 25040
rect 2574 24988 2626 25040
rect 2698 24988 2750 25040
rect 2822 24988 2874 25040
rect 2946 24988 2998 25040
rect 4846 24988 4898 25040
rect 4970 24988 5022 25040
rect 5094 24988 5146 25040
rect 5218 24988 5270 25040
rect 7139 24988 7191 25040
rect 7263 24988 7315 25040
rect 7387 24988 7439 25040
rect 7625 24988 7677 25040
rect 7749 24988 7801 25040
rect 7873 24988 7925 25040
rect 9794 24988 9846 25040
rect 9918 24988 9970 25040
rect 10042 24988 10094 25040
rect 10166 24988 10218 25040
rect 12066 24988 12118 25040
rect 12190 24988 12242 25040
rect 12314 24988 12366 25040
rect 12438 24988 12490 25040
rect 13202 24988 13254 25040
rect 13326 24988 13378 25040
rect 13450 24988 13502 25040
rect 13574 24988 13626 25040
rect 14352 25004 14404 25056
rect 14460 25004 14512 25056
rect 14568 25004 14619 25056
rect 14619 25004 14620 25056
rect 444 24896 445 24948
rect 445 24896 496 24948
rect 552 24896 604 24948
rect 660 24896 712 24948
rect 1438 24864 1490 24916
rect 1562 24864 1614 24916
rect 1686 24864 1738 24916
rect 1810 24864 1862 24916
rect 2574 24864 2626 24916
rect 2698 24864 2750 24916
rect 2822 24864 2874 24916
rect 2946 24864 2998 24916
rect 4846 24864 4898 24916
rect 4970 24864 5022 24916
rect 5094 24864 5146 24916
rect 5218 24864 5270 24916
rect 7139 24864 7191 24916
rect 7263 24864 7315 24916
rect 7387 24864 7439 24916
rect 7625 24864 7677 24916
rect 7749 24864 7801 24916
rect 7873 24864 7925 24916
rect 9794 24864 9846 24916
rect 9918 24864 9970 24916
rect 10042 24864 10094 24916
rect 10166 24864 10218 24916
rect 12066 24864 12118 24916
rect 12190 24864 12242 24916
rect 12314 24864 12366 24916
rect 12438 24864 12490 24916
rect 13202 24864 13254 24916
rect 13326 24864 13378 24916
rect 13450 24864 13502 24916
rect 13574 24864 13626 24916
rect 14352 24896 14404 24948
rect 14460 24896 14512 24948
rect 14568 24896 14619 24948
rect 14619 24896 14620 24948
rect 978 24697 1030 24740
rect 1102 24697 1154 24740
rect 1226 24697 1278 24740
rect 3729 24697 3781 24702
rect 978 24688 1030 24697
rect 1102 24688 1154 24697
rect 1226 24688 1278 24697
rect 978 24564 1030 24616
rect 1102 24564 1154 24616
rect 1226 24564 1278 24616
rect 978 24440 1030 24492
rect 1102 24440 1154 24492
rect 1226 24440 1278 24492
rect 978 24316 1030 24368
rect 1102 24316 1154 24368
rect 1226 24316 1278 24368
rect 978 24192 1030 24244
rect 1102 24192 1154 24244
rect 1226 24192 1278 24244
rect 978 24068 1030 24120
rect 1102 24068 1154 24120
rect 1226 24068 1278 24120
rect 978 23944 1030 23996
rect 1102 23944 1154 23996
rect 1226 23944 1278 23996
rect 978 23820 1030 23872
rect 1102 23820 1154 23872
rect 1226 23820 1278 23872
rect 978 23696 1030 23748
rect 1102 23696 1154 23748
rect 1226 23696 1278 23748
rect 978 23572 1030 23624
rect 1102 23572 1154 23624
rect 1226 23572 1278 23624
rect 978 23448 1030 23500
rect 1102 23448 1154 23500
rect 1226 23448 1278 23500
rect 978 23324 1030 23376
rect 1102 23324 1154 23376
rect 1226 23324 1278 23376
rect 978 23200 1030 23252
rect 1102 23200 1154 23252
rect 1226 23200 1278 23252
rect 978 23076 1030 23128
rect 1102 23076 1154 23128
rect 1226 23076 1278 23128
rect 978 22952 1030 23004
rect 1102 22952 1154 23004
rect 1226 22952 1278 23004
rect 978 22828 1030 22880
rect 1102 22828 1154 22880
rect 1226 22828 1278 22880
rect 978 22704 1030 22756
rect 1102 22704 1154 22756
rect 1226 22704 1278 22756
rect 978 22580 1030 22632
rect 1102 22580 1154 22632
rect 1226 22580 1278 22632
rect 978 22456 1030 22508
rect 1102 22456 1154 22508
rect 1226 22456 1278 22508
rect 978 22332 1030 22384
rect 1102 22332 1154 22384
rect 1226 22332 1278 22384
rect 978 22208 1030 22260
rect 1102 22208 1154 22260
rect 1226 22208 1278 22260
rect 978 22084 1030 22136
rect 1102 22084 1154 22136
rect 1226 22084 1278 22136
rect 978 21960 1030 22012
rect 1102 21960 1154 22012
rect 1226 21960 1278 22012
rect 978 21836 1030 21888
rect 1102 21836 1154 21888
rect 1226 21836 1278 21888
rect 978 21712 1030 21764
rect 1102 21712 1154 21764
rect 1226 21712 1278 21764
rect 3729 24650 3781 24697
rect 6335 24697 6387 24702
rect 3729 24542 3781 24594
rect 3729 24434 3781 24486
rect 3729 24326 3781 24378
rect 3729 24218 3781 24270
rect 3729 24110 3781 24162
rect 3729 24002 3781 24054
rect 3729 23894 3781 23946
rect 3729 23786 3781 23838
rect 3729 23678 3781 23730
rect 3729 23570 3781 23622
rect 3729 23462 3781 23514
rect 3729 23354 3781 23406
rect 3729 23246 3781 23298
rect 3729 23138 3781 23190
rect 3729 23030 3781 23082
rect 3729 22922 3781 22974
rect 3729 22814 3781 22866
rect 3729 22706 3781 22758
rect 3729 22598 3781 22650
rect 3729 22490 3781 22542
rect 3729 22382 3781 22434
rect 3729 22274 3781 22326
rect 3729 22166 3781 22218
rect 3729 22058 3781 22110
rect 3729 21950 3781 22002
rect 3729 21842 3781 21894
rect 3729 21734 3781 21786
rect 978 21631 1030 21640
rect 1102 21631 1154 21640
rect 1226 21631 1278 21640
rect 3729 21631 3781 21678
rect 978 21588 1030 21631
rect 1102 21588 1154 21631
rect 1226 21588 1278 21631
rect 3729 21626 3781 21631
rect 6335 24650 6387 24697
rect 8677 24697 8729 24702
rect 6335 24542 6387 24594
rect 6335 24434 6387 24486
rect 6335 24326 6387 24378
rect 6335 24218 6387 24270
rect 6335 24110 6387 24162
rect 6335 24002 6387 24054
rect 6335 23894 6387 23946
rect 6335 23786 6387 23838
rect 6335 23678 6387 23730
rect 6335 23570 6387 23622
rect 6335 23462 6387 23514
rect 6335 23354 6387 23406
rect 6335 23246 6387 23298
rect 6335 23138 6387 23190
rect 6335 23030 6387 23082
rect 6335 22922 6387 22974
rect 6335 22814 6387 22866
rect 6335 22706 6387 22758
rect 6335 22598 6387 22650
rect 6335 22490 6387 22542
rect 6335 22382 6387 22434
rect 6335 22274 6387 22326
rect 6335 22166 6387 22218
rect 6335 22058 6387 22110
rect 6335 21950 6387 22002
rect 6335 21842 6387 21894
rect 6335 21734 6387 21786
rect 6335 21631 6387 21678
rect 6335 21626 6387 21631
rect 7388 24627 7440 24648
rect 7388 24596 7389 24627
rect 7389 24596 7440 24627
rect 7624 24627 7676 24648
rect 7624 24596 7675 24627
rect 7675 24596 7676 24627
rect 7388 24488 7389 24540
rect 7389 24488 7440 24540
rect 7624 24488 7675 24540
rect 7675 24488 7676 24540
rect 7388 24380 7389 24432
rect 7389 24380 7440 24432
rect 7624 24380 7675 24432
rect 7675 24380 7676 24432
rect 7388 24272 7389 24324
rect 7389 24272 7440 24324
rect 7624 24272 7675 24324
rect 7675 24272 7676 24324
rect 7388 24164 7389 24216
rect 7389 24164 7440 24216
rect 7624 24164 7675 24216
rect 7675 24164 7676 24216
rect 7388 24056 7389 24108
rect 7389 24056 7440 24108
rect 7624 24056 7675 24108
rect 7675 24056 7676 24108
rect 7388 23948 7389 24000
rect 7389 23948 7440 24000
rect 7624 23948 7675 24000
rect 7675 23948 7676 24000
rect 7388 23840 7389 23892
rect 7389 23840 7440 23892
rect 7624 23840 7675 23892
rect 7675 23840 7676 23892
rect 7388 23732 7389 23784
rect 7389 23732 7440 23784
rect 7624 23732 7675 23784
rect 7675 23732 7676 23784
rect 7388 23624 7389 23676
rect 7389 23624 7440 23676
rect 7624 23624 7675 23676
rect 7675 23624 7676 23676
rect 7388 23516 7389 23568
rect 7389 23516 7440 23568
rect 7624 23516 7675 23568
rect 7675 23516 7676 23568
rect 7388 23408 7389 23460
rect 7389 23408 7440 23460
rect 7624 23408 7675 23460
rect 7675 23408 7676 23460
rect 7388 23300 7389 23352
rect 7389 23300 7440 23352
rect 7624 23300 7675 23352
rect 7675 23300 7676 23352
rect 7388 23192 7389 23244
rect 7389 23192 7440 23244
rect 7624 23192 7675 23244
rect 7675 23192 7676 23244
rect 7388 23084 7389 23136
rect 7389 23084 7440 23136
rect 7624 23084 7675 23136
rect 7675 23084 7676 23136
rect 7388 22976 7389 23028
rect 7389 22976 7440 23028
rect 7624 22976 7675 23028
rect 7675 22976 7676 23028
rect 7388 22868 7389 22920
rect 7389 22868 7440 22920
rect 7624 22868 7675 22920
rect 7675 22868 7676 22920
rect 7388 22760 7389 22812
rect 7389 22760 7440 22812
rect 7624 22760 7675 22812
rect 7675 22760 7676 22812
rect 7388 22652 7389 22704
rect 7389 22652 7440 22704
rect 7624 22652 7675 22704
rect 7675 22652 7676 22704
rect 7388 22544 7389 22596
rect 7389 22544 7440 22596
rect 7624 22544 7675 22596
rect 7675 22544 7676 22596
rect 7388 22436 7389 22488
rect 7389 22436 7440 22488
rect 7624 22436 7675 22488
rect 7675 22436 7676 22488
rect 7388 22328 7389 22380
rect 7389 22328 7440 22380
rect 7624 22328 7675 22380
rect 7675 22328 7676 22380
rect 7388 22220 7389 22272
rect 7389 22220 7440 22272
rect 7624 22220 7675 22272
rect 7675 22220 7676 22272
rect 7388 22112 7389 22164
rect 7389 22112 7440 22164
rect 7624 22112 7675 22164
rect 7675 22112 7676 22164
rect 7388 22004 7389 22056
rect 7389 22004 7440 22056
rect 7624 22004 7675 22056
rect 7675 22004 7676 22056
rect 7388 21896 7389 21948
rect 7389 21896 7440 21948
rect 7624 21896 7675 21948
rect 7675 21896 7676 21948
rect 7388 21788 7389 21840
rect 7389 21788 7440 21840
rect 7624 21788 7675 21840
rect 7675 21788 7676 21840
rect 7388 21701 7389 21732
rect 7389 21701 7440 21732
rect 7388 21680 7440 21701
rect 7624 21701 7675 21732
rect 7675 21701 7676 21732
rect 7624 21680 7676 21701
rect 8677 24650 8729 24697
rect 8677 24542 8729 24594
rect 8677 24434 8729 24486
rect 8677 24326 8729 24378
rect 8677 24218 8729 24270
rect 8677 24110 8729 24162
rect 8677 24002 8729 24054
rect 8677 23894 8729 23946
rect 8677 23786 8729 23838
rect 8677 23678 8729 23730
rect 8677 23570 8729 23622
rect 8677 23462 8729 23514
rect 8677 23354 8729 23406
rect 8677 23246 8729 23298
rect 8677 23138 8729 23190
rect 8677 23030 8729 23082
rect 8677 22922 8729 22974
rect 8677 22814 8729 22866
rect 8677 22706 8729 22758
rect 8677 22598 8729 22650
rect 8677 22490 8729 22542
rect 8677 22382 8729 22434
rect 8677 22274 8729 22326
rect 8677 22166 8729 22218
rect 8677 22058 8729 22110
rect 8677 21950 8729 22002
rect 8677 21842 8729 21894
rect 8677 21734 8729 21786
rect 8677 21631 8729 21678
rect 11283 24697 11335 24702
rect 13786 24697 13838 24740
rect 13910 24697 13962 24740
rect 14034 24697 14086 24740
rect 8677 21626 8729 21631
rect 11283 24650 11335 24697
rect 13786 24688 13838 24697
rect 13910 24688 13962 24697
rect 14034 24688 14086 24697
rect 11283 24542 11335 24594
rect 11283 24434 11335 24486
rect 11283 24326 11335 24378
rect 11283 24218 11335 24270
rect 11283 24110 11335 24162
rect 11283 24002 11335 24054
rect 11283 23894 11335 23946
rect 11283 23786 11335 23838
rect 11283 23678 11335 23730
rect 11283 23570 11335 23622
rect 11283 23462 11335 23514
rect 11283 23354 11335 23406
rect 11283 23246 11335 23298
rect 11283 23138 11335 23190
rect 11283 23030 11335 23082
rect 11283 22922 11335 22974
rect 11283 22814 11335 22866
rect 11283 22706 11335 22758
rect 11283 22598 11335 22650
rect 11283 22490 11335 22542
rect 11283 22382 11335 22434
rect 11283 22274 11335 22326
rect 11283 22166 11335 22218
rect 11283 22058 11335 22110
rect 11283 21950 11335 22002
rect 11283 21842 11335 21894
rect 11283 21734 11335 21786
rect 11283 21631 11335 21678
rect 13786 24564 13838 24616
rect 13910 24564 13962 24616
rect 14034 24564 14086 24616
rect 13786 24440 13838 24492
rect 13910 24440 13962 24492
rect 14034 24440 14086 24492
rect 13786 24316 13838 24368
rect 13910 24316 13962 24368
rect 14034 24316 14086 24368
rect 13786 24192 13838 24244
rect 13910 24192 13962 24244
rect 14034 24192 14086 24244
rect 13786 24068 13838 24120
rect 13910 24068 13962 24120
rect 14034 24068 14086 24120
rect 13786 23944 13838 23996
rect 13910 23944 13962 23996
rect 14034 23944 14086 23996
rect 13786 23820 13838 23872
rect 13910 23820 13962 23872
rect 14034 23820 14086 23872
rect 13786 23696 13838 23748
rect 13910 23696 13962 23748
rect 14034 23696 14086 23748
rect 13786 23572 13838 23624
rect 13910 23572 13962 23624
rect 14034 23572 14086 23624
rect 13786 23448 13838 23500
rect 13910 23448 13962 23500
rect 14034 23448 14086 23500
rect 13786 23324 13838 23376
rect 13910 23324 13962 23376
rect 14034 23324 14086 23376
rect 13786 23200 13838 23252
rect 13910 23200 13962 23252
rect 14034 23200 14086 23252
rect 13786 23076 13838 23128
rect 13910 23076 13962 23128
rect 14034 23076 14086 23128
rect 13786 22952 13838 23004
rect 13910 22952 13962 23004
rect 14034 22952 14086 23004
rect 13786 22828 13838 22880
rect 13910 22828 13962 22880
rect 14034 22828 14086 22880
rect 13786 22704 13838 22756
rect 13910 22704 13962 22756
rect 14034 22704 14086 22756
rect 13786 22580 13838 22632
rect 13910 22580 13962 22632
rect 14034 22580 14086 22632
rect 13786 22456 13838 22508
rect 13910 22456 13962 22508
rect 14034 22456 14086 22508
rect 13786 22332 13838 22384
rect 13910 22332 13962 22384
rect 14034 22332 14086 22384
rect 13786 22208 13838 22260
rect 13910 22208 13962 22260
rect 14034 22208 14086 22260
rect 13786 22084 13838 22136
rect 13910 22084 13962 22136
rect 14034 22084 14086 22136
rect 13786 21960 13838 22012
rect 13910 21960 13962 22012
rect 14034 21960 14086 22012
rect 13786 21836 13838 21888
rect 13910 21836 13962 21888
rect 14034 21836 14086 21888
rect 13786 21712 13838 21764
rect 13910 21712 13962 21764
rect 14034 21712 14086 21764
rect 13786 21631 13838 21640
rect 13910 21631 13962 21640
rect 14034 21631 14086 21640
rect 11283 21626 11335 21631
rect 13786 21588 13838 21631
rect 13910 21588 13962 21631
rect 14034 21588 14086 21631
rect 444 21417 445 21469
rect 445 21417 496 21469
rect 552 21417 604 21469
rect 660 21417 712 21469
rect 1408 21417 1460 21469
rect 1516 21417 1568 21469
rect 1624 21417 1676 21469
rect 1732 21417 1784 21469
rect 1840 21417 1892 21469
rect 2544 21417 2596 21469
rect 2652 21417 2704 21469
rect 2760 21417 2812 21469
rect 2868 21417 2920 21469
rect 2976 21417 3028 21469
rect 4816 21417 4868 21469
rect 4924 21417 4976 21469
rect 5032 21417 5084 21469
rect 5140 21417 5192 21469
rect 5248 21417 5300 21469
rect 7101 21417 7153 21469
rect 7209 21417 7261 21469
rect 7317 21417 7369 21469
rect 7425 21417 7477 21469
rect 7587 21417 7639 21469
rect 7695 21417 7747 21469
rect 7803 21417 7855 21469
rect 7911 21417 7963 21469
rect 9764 21417 9816 21469
rect 9872 21417 9924 21469
rect 9980 21417 10032 21469
rect 10088 21417 10140 21469
rect 10196 21417 10248 21469
rect 12036 21417 12088 21469
rect 12144 21417 12196 21469
rect 12252 21417 12304 21469
rect 12360 21417 12412 21469
rect 12468 21417 12520 21469
rect 13172 21417 13224 21469
rect 13280 21417 13332 21469
rect 13388 21417 13440 21469
rect 13496 21417 13548 21469
rect 13604 21417 13656 21469
rect 14352 21417 14404 21469
rect 14460 21417 14512 21469
rect 14568 21417 14619 21469
rect 14619 21417 14620 21469
rect 444 21309 445 21361
rect 445 21309 496 21361
rect 552 21309 604 21361
rect 660 21309 712 21361
rect 1408 21309 1460 21361
rect 1516 21309 1568 21361
rect 1624 21309 1676 21361
rect 1732 21309 1784 21361
rect 1840 21309 1892 21361
rect 2544 21309 2596 21361
rect 2652 21309 2704 21361
rect 2760 21309 2812 21361
rect 2868 21309 2920 21361
rect 2976 21309 3028 21361
rect 4816 21309 4868 21361
rect 4924 21309 4976 21361
rect 5032 21309 5084 21361
rect 5140 21309 5192 21361
rect 5248 21309 5300 21361
rect 7101 21309 7153 21361
rect 7209 21309 7261 21361
rect 7317 21309 7369 21361
rect 7425 21309 7477 21361
rect 7587 21309 7639 21361
rect 7695 21309 7747 21361
rect 7803 21309 7855 21361
rect 7911 21309 7963 21361
rect 9764 21309 9816 21361
rect 9872 21309 9924 21361
rect 9980 21309 10032 21361
rect 10088 21309 10140 21361
rect 10196 21309 10248 21361
rect 12036 21309 12088 21361
rect 12144 21309 12196 21361
rect 12252 21309 12304 21361
rect 12360 21309 12412 21361
rect 12468 21309 12520 21361
rect 13172 21309 13224 21361
rect 13280 21309 13332 21361
rect 13388 21309 13440 21361
rect 13496 21309 13548 21361
rect 13604 21309 13656 21361
rect 14352 21309 14404 21361
rect 14460 21309 14512 21361
rect 14568 21309 14619 21361
rect 14619 21309 14620 21361
rect 444 21201 445 21253
rect 445 21201 496 21253
rect 552 21213 604 21253
rect 660 21213 712 21253
rect 1408 21213 1460 21253
rect 1516 21213 1568 21253
rect 1624 21213 1676 21253
rect 1732 21213 1784 21253
rect 1840 21213 1892 21253
rect 2544 21213 2596 21253
rect 2652 21213 2704 21253
rect 2760 21213 2812 21253
rect 2868 21213 2920 21253
rect 2976 21213 3028 21253
rect 4816 21213 4868 21253
rect 4924 21213 4976 21253
rect 5032 21213 5084 21253
rect 5140 21213 5192 21253
rect 5248 21213 5300 21253
rect 7101 21213 7153 21253
rect 7209 21213 7261 21253
rect 7317 21213 7369 21253
rect 7425 21213 7477 21253
rect 7587 21213 7639 21253
rect 7695 21213 7747 21253
rect 7803 21213 7855 21253
rect 7911 21213 7963 21253
rect 9764 21213 9816 21253
rect 9872 21213 9924 21253
rect 9980 21213 10032 21253
rect 10088 21213 10140 21253
rect 10196 21213 10248 21253
rect 12036 21213 12088 21253
rect 12144 21213 12196 21253
rect 12252 21213 12304 21253
rect 12360 21213 12412 21253
rect 12468 21213 12520 21253
rect 13172 21213 13224 21253
rect 13280 21213 13332 21253
rect 13388 21213 13440 21253
rect 13496 21213 13548 21253
rect 13604 21213 13656 21253
rect 14352 21213 14404 21253
rect 14460 21213 14512 21253
rect 552 21201 553 21213
rect 553 21201 604 21213
rect 660 21201 712 21213
rect 1408 21201 1460 21213
rect 1516 21201 1568 21213
rect 1624 21201 1676 21213
rect 1732 21201 1784 21213
rect 1840 21201 1892 21213
rect 2544 21201 2596 21213
rect 2652 21201 2704 21213
rect 2760 21201 2812 21213
rect 2868 21201 2920 21213
rect 2976 21201 3028 21213
rect 4816 21201 4868 21213
rect 4924 21201 4976 21213
rect 5032 21201 5084 21213
rect 5140 21201 5192 21213
rect 5248 21201 5300 21213
rect 7101 21201 7153 21213
rect 7209 21201 7261 21213
rect 7317 21201 7369 21213
rect 7425 21201 7477 21213
rect 7587 21201 7639 21213
rect 7695 21201 7747 21213
rect 7803 21201 7855 21213
rect 7911 21201 7963 21213
rect 9764 21201 9816 21213
rect 9872 21201 9924 21213
rect 9980 21201 10032 21213
rect 10088 21201 10140 21213
rect 10196 21201 10248 21213
rect 12036 21201 12088 21213
rect 12144 21201 12196 21213
rect 12252 21201 12304 21213
rect 12360 21201 12412 21213
rect 12468 21201 12520 21213
rect 13172 21201 13224 21213
rect 13280 21201 13332 21213
rect 13388 21201 13440 21213
rect 13496 21201 13548 21213
rect 13604 21201 13656 21213
rect 14352 21201 14404 21213
rect 14460 21201 14511 21213
rect 14511 21201 14512 21213
rect 14568 21201 14619 21253
rect 14619 21201 14620 21253
rect 14954 52219 15006 52271
rect 14954 52111 15006 52163
rect 14954 52003 15006 52055
rect 14954 51895 15006 51947
rect 14954 51787 15006 51839
rect 14954 51679 15006 51731
rect 14954 51571 15006 51623
rect 14954 51463 15006 51515
rect 14954 51355 15006 51407
rect 14954 51247 15006 51299
rect 14954 51139 15006 51191
rect 14954 51031 15006 51083
rect 14954 50923 15006 50975
rect 14954 37819 15006 37871
rect 14954 37711 15006 37763
rect 14954 37603 15006 37655
rect 14954 37495 15006 37547
rect 14954 37387 15006 37439
rect 14954 37279 15006 37331
rect 14954 37171 15006 37223
rect 14954 37063 15006 37115
rect 14954 36955 15006 37007
rect 14954 36847 15006 36899
rect 14954 36739 15006 36791
rect 14954 36631 15006 36683
rect 14954 36523 15006 36575
rect 3680 20525 3732 20577
rect 3788 20525 3840 20577
rect 3896 20525 3948 20577
rect 4004 20525 4056 20577
rect 4112 20525 4164 20577
rect 5952 20525 6004 20577
rect 6060 20525 6112 20577
rect 6168 20525 6220 20577
rect 6276 20525 6328 20577
rect 6384 20525 6436 20577
rect 8628 20525 8680 20577
rect 8736 20525 8788 20577
rect 8844 20525 8896 20577
rect 8952 20525 9004 20577
rect 9060 20525 9112 20577
rect 10900 20525 10952 20577
rect 11008 20525 11060 20577
rect 11116 20525 11168 20577
rect 11224 20525 11276 20577
rect 11332 20525 11384 20577
rect 3680 20417 3732 20469
rect 3788 20417 3840 20469
rect 3896 20417 3948 20469
rect 4004 20417 4056 20469
rect 4112 20417 4164 20469
rect 5952 20417 6004 20469
rect 6060 20417 6112 20469
rect 6168 20417 6220 20469
rect 6276 20417 6328 20469
rect 6384 20417 6436 20469
rect 8628 20417 8680 20469
rect 8736 20417 8788 20469
rect 8844 20417 8896 20469
rect 8952 20417 9004 20469
rect 9060 20417 9112 20469
rect 10900 20417 10952 20469
rect 11008 20417 11060 20469
rect 11116 20417 11168 20469
rect 11224 20417 11276 20469
rect 11332 20417 11384 20469
rect 3680 20309 3732 20361
rect 3788 20309 3840 20361
rect 3896 20309 3948 20361
rect 4004 20309 4056 20361
rect 4112 20309 4164 20361
rect 5952 20309 6004 20361
rect 6060 20309 6112 20361
rect 6168 20309 6220 20361
rect 6276 20309 6328 20361
rect 6384 20309 6436 20361
rect 8628 20309 8680 20361
rect 8736 20309 8788 20361
rect 8844 20309 8896 20361
rect 8952 20309 9004 20361
rect 9060 20309 9112 20361
rect 10900 20309 10952 20361
rect 11008 20309 11060 20361
rect 11116 20309 11168 20361
rect 11224 20309 11276 20361
rect 11332 20309 11384 20361
rect 4816 19925 4868 19951
rect 4924 19925 4976 19951
rect 5032 19925 5084 19951
rect 5140 19925 5192 19951
rect 5248 19925 5300 19951
rect 7101 19925 7153 19951
rect 7209 19925 7261 19951
rect 7317 19925 7369 19951
rect 7425 19925 7477 19951
rect 7587 19925 7639 19951
rect 7695 19925 7747 19951
rect 7803 19925 7855 19951
rect 7911 19925 7963 19951
rect 9764 19925 9816 19951
rect 9872 19925 9924 19951
rect 9980 19925 10032 19951
rect 10088 19925 10140 19951
rect 10196 19925 10248 19951
rect 4816 19899 4868 19925
rect 4924 19899 4976 19925
rect 5032 19899 5084 19925
rect 5140 19899 5192 19925
rect 5248 19899 5300 19925
rect 7101 19899 7153 19925
rect 7209 19899 7261 19925
rect 7317 19899 7369 19925
rect 7425 19899 7477 19925
rect 7587 19899 7639 19925
rect 7695 19899 7747 19925
rect 7803 19899 7855 19925
rect 7911 19899 7963 19925
rect 9764 19899 9816 19925
rect 9872 19899 9924 19925
rect 9980 19899 10032 19925
rect 10088 19899 10140 19925
rect 10196 19899 10248 19925
rect 4816 19817 4868 19843
rect 4924 19817 4976 19843
rect 5032 19817 5084 19843
rect 5140 19817 5192 19843
rect 5248 19817 5300 19843
rect 7101 19817 7153 19843
rect 7209 19817 7261 19843
rect 7317 19817 7369 19843
rect 7425 19817 7477 19843
rect 7587 19817 7639 19843
rect 7695 19817 7747 19843
rect 7803 19817 7855 19843
rect 7911 19817 7963 19843
rect 9764 19817 9816 19843
rect 9872 19817 9924 19843
rect 9980 19817 10032 19843
rect 10088 19817 10140 19843
rect 10196 19817 10248 19843
rect 4816 19791 4868 19817
rect 4924 19791 4976 19817
rect 5032 19791 5084 19817
rect 5140 19791 5192 19817
rect 5248 19791 5300 19817
rect 7101 19791 7153 19817
rect 7209 19791 7261 19817
rect 7317 19791 7369 19817
rect 7425 19791 7477 19817
rect 7587 19791 7639 19817
rect 7695 19791 7747 19817
rect 7803 19791 7855 19817
rect 7911 19791 7963 19817
rect 9764 19791 9816 19817
rect 9872 19791 9924 19817
rect 9980 19791 10032 19817
rect 10088 19791 10140 19817
rect 10196 19791 10248 19817
rect 3680 19545 3732 19584
rect 3788 19545 3840 19584
rect 3896 19545 3948 19584
rect 4004 19545 4056 19584
rect 4112 19545 4164 19584
rect 5952 19545 6004 19584
rect 6060 19545 6112 19584
rect 6168 19545 6220 19584
rect 6276 19545 6328 19584
rect 6384 19545 6436 19584
rect 8628 19545 8680 19584
rect 8736 19545 8788 19584
rect 8844 19545 8896 19584
rect 8952 19545 9004 19584
rect 9060 19545 9112 19584
rect 10900 19545 10952 19584
rect 11008 19545 11060 19584
rect 11116 19545 11168 19584
rect 11224 19545 11276 19584
rect 11332 19545 11384 19584
rect 3680 19532 3732 19545
rect 3788 19532 3840 19545
rect 3896 19532 3948 19545
rect 4004 19532 4056 19545
rect 4112 19532 4164 19545
rect 5952 19532 6004 19545
rect 6060 19532 6112 19545
rect 6168 19532 6220 19545
rect 6276 19532 6328 19545
rect 6384 19532 6436 19545
rect 8628 19532 8680 19545
rect 8736 19532 8788 19545
rect 8844 19532 8896 19545
rect 8952 19532 9004 19545
rect 9060 19532 9112 19545
rect 10900 19532 10952 19545
rect 11008 19532 11060 19545
rect 11116 19532 11168 19545
rect 11224 19532 11276 19545
rect 11332 19532 11384 19545
rect 3680 19463 3732 19476
rect 3788 19463 3840 19476
rect 3896 19463 3948 19476
rect 4004 19463 4056 19476
rect 4112 19463 4164 19476
rect 5952 19463 6004 19476
rect 6060 19463 6112 19476
rect 6168 19463 6220 19476
rect 6276 19463 6328 19476
rect 6384 19463 6436 19476
rect 8628 19463 8680 19476
rect 8736 19463 8788 19476
rect 8844 19463 8896 19476
rect 8952 19463 9004 19476
rect 9060 19463 9112 19476
rect 10900 19463 10952 19476
rect 11008 19463 11060 19476
rect 11116 19463 11168 19476
rect 11224 19463 11276 19476
rect 11332 19463 11384 19476
rect 3680 19424 3732 19463
rect 3788 19424 3840 19463
rect 3896 19424 3948 19463
rect 4004 19424 4056 19463
rect 4112 19424 4164 19463
rect 5952 19424 6004 19463
rect 6060 19424 6112 19463
rect 6168 19424 6220 19463
rect 6276 19424 6328 19463
rect 6384 19424 6436 19463
rect 8628 19424 8680 19463
rect 8736 19424 8788 19463
rect 8844 19424 8896 19463
rect 8952 19424 9004 19463
rect 9060 19424 9112 19463
rect 10900 19424 10952 19463
rect 11008 19424 11060 19463
rect 11116 19424 11168 19463
rect 11224 19424 11276 19463
rect 11332 19424 11384 19463
rect 4816 19199 4868 19202
rect 4924 19199 4976 19202
rect 5032 19199 5084 19202
rect 5140 19199 5192 19202
rect 5248 19199 5300 19202
rect 7101 19199 7153 19202
rect 7209 19199 7261 19202
rect 7317 19199 7369 19202
rect 7425 19199 7477 19202
rect 7587 19199 7639 19202
rect 7695 19199 7747 19202
rect 7803 19199 7855 19202
rect 7911 19199 7963 19202
rect 9764 19199 9816 19202
rect 9872 19199 9924 19202
rect 9980 19199 10032 19202
rect 10088 19199 10140 19202
rect 10196 19199 10248 19202
rect 4816 19150 4868 19199
rect 4924 19150 4976 19199
rect 5032 19150 5084 19199
rect 5140 19150 5192 19199
rect 5248 19150 5300 19199
rect 7101 19150 7153 19199
rect 7209 19150 7261 19199
rect 7317 19150 7369 19199
rect 7425 19150 7477 19199
rect 7587 19150 7639 19199
rect 7695 19150 7747 19199
rect 7803 19150 7855 19199
rect 7911 19150 7963 19199
rect 9764 19150 9816 19199
rect 9872 19150 9924 19199
rect 9980 19150 10032 19199
rect 10088 19150 10140 19199
rect 10196 19150 10248 19199
rect 4816 19091 4868 19094
rect 4924 19091 4976 19094
rect 5032 19091 5084 19094
rect 5140 19091 5192 19094
rect 5248 19091 5300 19094
rect 7101 19091 7153 19094
rect 7209 19091 7261 19094
rect 7317 19091 7369 19094
rect 7425 19091 7477 19094
rect 7587 19091 7639 19094
rect 7695 19091 7747 19094
rect 7803 19091 7855 19094
rect 7911 19091 7963 19094
rect 9764 19091 9816 19094
rect 9872 19091 9924 19094
rect 9980 19091 10032 19094
rect 10088 19091 10140 19094
rect 10196 19091 10248 19094
rect 4816 19045 4868 19091
rect 4924 19045 4976 19091
rect 5032 19045 5084 19091
rect 5140 19045 5192 19091
rect 5248 19045 5300 19091
rect 7101 19045 7153 19091
rect 7209 19045 7261 19091
rect 7317 19045 7369 19091
rect 7425 19045 7477 19091
rect 7587 19045 7639 19091
rect 7695 19045 7747 19091
rect 7803 19045 7855 19091
rect 7911 19045 7963 19091
rect 9764 19045 9816 19091
rect 9872 19045 9924 19091
rect 9980 19045 10032 19091
rect 10088 19045 10140 19091
rect 10196 19045 10248 19091
rect 4816 19042 4868 19045
rect 4924 19042 4976 19045
rect 5032 19042 5084 19045
rect 5140 19042 5192 19045
rect 5248 19042 5300 19045
rect 7101 19042 7153 19045
rect 7209 19042 7261 19045
rect 7317 19042 7369 19045
rect 7425 19042 7477 19045
rect 7587 19042 7639 19045
rect 7695 19042 7747 19045
rect 7803 19042 7855 19045
rect 7911 19042 7963 19045
rect 9764 19042 9816 19045
rect 9872 19042 9924 19045
rect 9980 19042 10032 19045
rect 10088 19042 10140 19045
rect 10196 19042 10248 19045
rect 4816 18937 4868 18986
rect 4924 18937 4976 18986
rect 5032 18937 5084 18986
rect 5140 18937 5192 18986
rect 5248 18937 5300 18986
rect 7101 18937 7153 18986
rect 7209 18937 7261 18986
rect 7317 18937 7369 18986
rect 7425 18937 7477 18986
rect 7587 18937 7639 18986
rect 7695 18937 7747 18986
rect 7803 18937 7855 18986
rect 7911 18937 7963 18986
rect 9764 18937 9816 18986
rect 9872 18937 9924 18986
rect 9980 18937 10032 18986
rect 10088 18937 10140 18986
rect 10196 18937 10248 18986
rect 4816 18934 4868 18937
rect 4924 18934 4976 18937
rect 5032 18934 5084 18937
rect 5140 18934 5192 18937
rect 5248 18934 5300 18937
rect 7101 18934 7153 18937
rect 7209 18934 7261 18937
rect 7317 18934 7369 18937
rect 7425 18934 7477 18937
rect 7587 18934 7639 18937
rect 7695 18934 7747 18937
rect 7803 18934 7855 18937
rect 7911 18934 7963 18937
rect 9764 18934 9816 18937
rect 9872 18934 9924 18937
rect 9980 18934 10032 18937
rect 10088 18934 10140 18937
rect 10196 18934 10248 18937
rect 3680 18673 3732 18712
rect 3788 18673 3840 18712
rect 3896 18673 3948 18712
rect 4004 18673 4056 18712
rect 4112 18673 4164 18712
rect 5952 18673 6004 18712
rect 6060 18673 6112 18712
rect 6168 18673 6220 18712
rect 6276 18673 6328 18712
rect 6384 18673 6436 18712
rect 8628 18673 8680 18712
rect 8736 18673 8788 18712
rect 8844 18673 8896 18712
rect 8952 18673 9004 18712
rect 9060 18673 9112 18712
rect 10900 18673 10952 18712
rect 11008 18673 11060 18712
rect 11116 18673 11168 18712
rect 11224 18673 11276 18712
rect 11332 18673 11384 18712
rect 3680 18660 3732 18673
rect 3788 18660 3840 18673
rect 3896 18660 3948 18673
rect 4004 18660 4056 18673
rect 4112 18660 4164 18673
rect 5952 18660 6004 18673
rect 6060 18660 6112 18673
rect 6168 18660 6220 18673
rect 6276 18660 6328 18673
rect 6384 18660 6436 18673
rect 8628 18660 8680 18673
rect 8736 18660 8788 18673
rect 8844 18660 8896 18673
rect 8952 18660 9004 18673
rect 9060 18660 9112 18673
rect 10900 18660 10952 18673
rect 11008 18660 11060 18673
rect 11116 18660 11168 18673
rect 11224 18660 11276 18673
rect 11332 18660 11384 18673
rect 3680 18591 3732 18604
rect 3788 18591 3840 18604
rect 3896 18591 3948 18604
rect 4004 18591 4056 18604
rect 4112 18591 4164 18604
rect 5952 18591 6004 18604
rect 6060 18591 6112 18604
rect 6168 18591 6220 18604
rect 6276 18591 6328 18604
rect 6384 18591 6436 18604
rect 8628 18591 8680 18604
rect 8736 18591 8788 18604
rect 8844 18591 8896 18604
rect 8952 18591 9004 18604
rect 9060 18591 9112 18604
rect 10900 18591 10952 18604
rect 11008 18591 11060 18604
rect 11116 18591 11168 18604
rect 11224 18591 11276 18604
rect 11332 18591 11384 18604
rect 3680 18552 3732 18591
rect 3788 18552 3840 18591
rect 3896 18552 3948 18591
rect 4004 18552 4056 18591
rect 4112 18552 4164 18591
rect 5952 18552 6004 18591
rect 6060 18552 6112 18591
rect 6168 18552 6220 18591
rect 6276 18552 6328 18591
rect 6384 18552 6436 18591
rect 8628 18552 8680 18591
rect 8736 18552 8788 18591
rect 8844 18552 8896 18591
rect 8952 18552 9004 18591
rect 9060 18552 9112 18591
rect 10900 18552 10952 18591
rect 11008 18552 11060 18591
rect 11116 18552 11168 18591
rect 11224 18552 11276 18591
rect 11332 18552 11384 18591
rect 4816 18327 4868 18330
rect 4924 18327 4976 18330
rect 5032 18327 5084 18330
rect 5140 18327 5192 18330
rect 5248 18327 5300 18330
rect 7101 18327 7153 18330
rect 7209 18327 7261 18330
rect 7317 18327 7369 18330
rect 7425 18327 7477 18330
rect 7587 18327 7639 18330
rect 7695 18327 7747 18330
rect 7803 18327 7855 18330
rect 7911 18327 7963 18330
rect 9764 18327 9816 18330
rect 9872 18327 9924 18330
rect 9980 18327 10032 18330
rect 10088 18327 10140 18330
rect 10196 18327 10248 18330
rect 4816 18278 4868 18327
rect 4924 18278 4976 18327
rect 5032 18278 5084 18327
rect 5140 18278 5192 18327
rect 5248 18278 5300 18327
rect 7101 18278 7153 18327
rect 7209 18278 7261 18327
rect 7317 18278 7369 18327
rect 7425 18278 7477 18327
rect 7587 18278 7639 18327
rect 7695 18278 7747 18327
rect 7803 18278 7855 18327
rect 7911 18278 7963 18327
rect 9764 18278 9816 18327
rect 9872 18278 9924 18327
rect 9980 18278 10032 18327
rect 10088 18278 10140 18327
rect 10196 18278 10248 18327
rect 4816 18219 4868 18222
rect 4924 18219 4976 18222
rect 5032 18219 5084 18222
rect 5140 18219 5192 18222
rect 5248 18219 5300 18222
rect 7101 18219 7153 18222
rect 7209 18219 7261 18222
rect 7317 18219 7369 18222
rect 7425 18219 7477 18222
rect 7587 18219 7639 18222
rect 7695 18219 7747 18222
rect 7803 18219 7855 18222
rect 7911 18219 7963 18222
rect 9764 18219 9816 18222
rect 9872 18219 9924 18222
rect 9980 18219 10032 18222
rect 10088 18219 10140 18222
rect 10196 18219 10248 18222
rect 4816 18173 4868 18219
rect 4924 18173 4976 18219
rect 5032 18173 5084 18219
rect 5140 18173 5192 18219
rect 5248 18173 5300 18219
rect 7101 18173 7153 18219
rect 7209 18173 7261 18219
rect 7317 18173 7369 18219
rect 7425 18173 7477 18219
rect 7587 18173 7639 18219
rect 7695 18173 7747 18219
rect 7803 18173 7855 18219
rect 7911 18173 7963 18219
rect 9764 18173 9816 18219
rect 9872 18173 9924 18219
rect 9980 18173 10032 18219
rect 10088 18173 10140 18219
rect 10196 18173 10248 18219
rect 4816 18170 4868 18173
rect 4924 18170 4976 18173
rect 5032 18170 5084 18173
rect 5140 18170 5192 18173
rect 5248 18170 5300 18173
rect 7101 18170 7153 18173
rect 7209 18170 7261 18173
rect 7317 18170 7369 18173
rect 7425 18170 7477 18173
rect 7587 18170 7639 18173
rect 7695 18170 7747 18173
rect 7803 18170 7855 18173
rect 7911 18170 7963 18173
rect 9764 18170 9816 18173
rect 9872 18170 9924 18173
rect 9980 18170 10032 18173
rect 10088 18170 10140 18173
rect 10196 18170 10248 18173
rect 4816 18065 4868 18114
rect 4924 18065 4976 18114
rect 5032 18065 5084 18114
rect 5140 18065 5192 18114
rect 5248 18065 5300 18114
rect 7101 18065 7153 18114
rect 7209 18065 7261 18114
rect 7317 18065 7369 18114
rect 7425 18065 7477 18114
rect 7587 18065 7639 18114
rect 7695 18065 7747 18114
rect 7803 18065 7855 18114
rect 7911 18065 7963 18114
rect 9764 18065 9816 18114
rect 9872 18065 9924 18114
rect 9980 18065 10032 18114
rect 10088 18065 10140 18114
rect 10196 18065 10248 18114
rect 4816 18062 4868 18065
rect 4924 18062 4976 18065
rect 5032 18062 5084 18065
rect 5140 18062 5192 18065
rect 5248 18062 5300 18065
rect 7101 18062 7153 18065
rect 7209 18062 7261 18065
rect 7317 18062 7369 18065
rect 7425 18062 7477 18065
rect 7587 18062 7639 18065
rect 7695 18062 7747 18065
rect 7803 18062 7855 18065
rect 7911 18062 7963 18065
rect 9764 18062 9816 18065
rect 9872 18062 9924 18065
rect 9980 18062 10032 18065
rect 10088 18062 10140 18065
rect 10196 18062 10248 18065
rect 3680 17801 3732 17840
rect 3788 17801 3840 17840
rect 3896 17801 3948 17840
rect 4004 17801 4056 17840
rect 4112 17801 4164 17840
rect 5952 17801 6004 17840
rect 6060 17801 6112 17840
rect 6168 17801 6220 17840
rect 6276 17801 6328 17840
rect 6384 17801 6436 17840
rect 8628 17801 8680 17840
rect 8736 17801 8788 17840
rect 8844 17801 8896 17840
rect 8952 17801 9004 17840
rect 9060 17801 9112 17840
rect 10900 17801 10952 17840
rect 11008 17801 11060 17840
rect 11116 17801 11168 17840
rect 11224 17801 11276 17840
rect 11332 17801 11384 17840
rect 3680 17788 3732 17801
rect 3788 17788 3840 17801
rect 3896 17788 3948 17801
rect 4004 17788 4056 17801
rect 4112 17788 4164 17801
rect 5952 17788 6004 17801
rect 6060 17788 6112 17801
rect 6168 17788 6220 17801
rect 6276 17788 6328 17801
rect 6384 17788 6436 17801
rect 8628 17788 8680 17801
rect 8736 17788 8788 17801
rect 8844 17788 8896 17801
rect 8952 17788 9004 17801
rect 9060 17788 9112 17801
rect 10900 17788 10952 17801
rect 11008 17788 11060 17801
rect 11116 17788 11168 17801
rect 11224 17788 11276 17801
rect 11332 17788 11384 17801
rect 3680 17719 3732 17732
rect 3788 17719 3840 17732
rect 3896 17719 3948 17732
rect 4004 17719 4056 17732
rect 4112 17719 4164 17732
rect 5952 17719 6004 17732
rect 6060 17719 6112 17732
rect 6168 17719 6220 17732
rect 6276 17719 6328 17732
rect 6384 17719 6436 17732
rect 8628 17719 8680 17732
rect 8736 17719 8788 17732
rect 8844 17719 8896 17732
rect 8952 17719 9004 17732
rect 9060 17719 9112 17732
rect 10900 17719 10952 17732
rect 11008 17719 11060 17732
rect 11116 17719 11168 17732
rect 11224 17719 11276 17732
rect 11332 17719 11384 17732
rect 3680 17680 3732 17719
rect 3788 17680 3840 17719
rect 3896 17680 3948 17719
rect 4004 17680 4056 17719
rect 4112 17680 4164 17719
rect 5952 17680 6004 17719
rect 6060 17680 6112 17719
rect 6168 17680 6220 17719
rect 6276 17680 6328 17719
rect 6384 17680 6436 17719
rect 8628 17680 8680 17719
rect 8736 17680 8788 17719
rect 8844 17680 8896 17719
rect 8952 17680 9004 17719
rect 9060 17680 9112 17719
rect 10900 17680 10952 17719
rect 11008 17680 11060 17719
rect 11116 17680 11168 17719
rect 11224 17680 11276 17719
rect 11332 17680 11384 17719
rect 4816 17455 4868 17458
rect 4924 17455 4976 17458
rect 5032 17455 5084 17458
rect 5140 17455 5192 17458
rect 5248 17455 5300 17458
rect 7101 17455 7153 17458
rect 7209 17455 7261 17458
rect 7317 17455 7369 17458
rect 7425 17455 7477 17458
rect 7587 17455 7639 17458
rect 7695 17455 7747 17458
rect 7803 17455 7855 17458
rect 7911 17455 7963 17458
rect 9764 17455 9816 17458
rect 9872 17455 9924 17458
rect 9980 17455 10032 17458
rect 10088 17455 10140 17458
rect 10196 17455 10248 17458
rect 4816 17406 4868 17455
rect 4924 17406 4976 17455
rect 5032 17406 5084 17455
rect 5140 17406 5192 17455
rect 5248 17406 5300 17455
rect 7101 17406 7153 17455
rect 7209 17406 7261 17455
rect 7317 17406 7369 17455
rect 7425 17406 7477 17455
rect 7587 17406 7639 17455
rect 7695 17406 7747 17455
rect 7803 17406 7855 17455
rect 7911 17406 7963 17455
rect 9764 17406 9816 17455
rect 9872 17406 9924 17455
rect 9980 17406 10032 17455
rect 10088 17406 10140 17455
rect 10196 17406 10248 17455
rect 4816 17347 4868 17350
rect 4924 17347 4976 17350
rect 5032 17347 5084 17350
rect 5140 17347 5192 17350
rect 5248 17347 5300 17350
rect 7101 17347 7153 17350
rect 7209 17347 7261 17350
rect 7317 17347 7369 17350
rect 7425 17347 7477 17350
rect 7587 17347 7639 17350
rect 7695 17347 7747 17350
rect 7803 17347 7855 17350
rect 7911 17347 7963 17350
rect 9764 17347 9816 17350
rect 9872 17347 9924 17350
rect 9980 17347 10032 17350
rect 10088 17347 10140 17350
rect 10196 17347 10248 17350
rect 4816 17301 4868 17347
rect 4924 17301 4976 17347
rect 5032 17301 5084 17347
rect 5140 17301 5192 17347
rect 5248 17301 5300 17347
rect 7101 17301 7153 17347
rect 7209 17301 7261 17347
rect 7317 17301 7369 17347
rect 7425 17301 7477 17347
rect 7587 17301 7639 17347
rect 7695 17301 7747 17347
rect 7803 17301 7855 17347
rect 7911 17301 7963 17347
rect 9764 17301 9816 17347
rect 9872 17301 9924 17347
rect 9980 17301 10032 17347
rect 10088 17301 10140 17347
rect 10196 17301 10248 17347
rect 4816 17298 4868 17301
rect 4924 17298 4976 17301
rect 5032 17298 5084 17301
rect 5140 17298 5192 17301
rect 5248 17298 5300 17301
rect 7101 17298 7153 17301
rect 7209 17298 7261 17301
rect 7317 17298 7369 17301
rect 7425 17298 7477 17301
rect 7587 17298 7639 17301
rect 7695 17298 7747 17301
rect 7803 17298 7855 17301
rect 7911 17298 7963 17301
rect 9764 17298 9816 17301
rect 9872 17298 9924 17301
rect 9980 17298 10032 17301
rect 10088 17298 10140 17301
rect 10196 17298 10248 17301
rect 4816 17193 4868 17242
rect 4924 17193 4976 17242
rect 5032 17193 5084 17242
rect 5140 17193 5192 17242
rect 5248 17193 5300 17242
rect 7101 17193 7153 17242
rect 7209 17193 7261 17242
rect 7317 17193 7369 17242
rect 7425 17193 7477 17242
rect 7587 17193 7639 17242
rect 7695 17193 7747 17242
rect 7803 17193 7855 17242
rect 7911 17193 7963 17242
rect 9764 17193 9816 17242
rect 9872 17193 9924 17242
rect 9980 17193 10032 17242
rect 10088 17193 10140 17242
rect 10196 17193 10248 17242
rect 4816 17190 4868 17193
rect 4924 17190 4976 17193
rect 5032 17190 5084 17193
rect 5140 17190 5192 17193
rect 5248 17190 5300 17193
rect 7101 17190 7153 17193
rect 7209 17190 7261 17193
rect 7317 17190 7369 17193
rect 7425 17190 7477 17193
rect 7587 17190 7639 17193
rect 7695 17190 7747 17193
rect 7803 17190 7855 17193
rect 7911 17190 7963 17193
rect 9764 17190 9816 17193
rect 9872 17190 9924 17193
rect 9980 17190 10032 17193
rect 10088 17190 10140 17193
rect 10196 17190 10248 17193
rect 3680 16929 3732 16968
rect 3788 16929 3840 16968
rect 3896 16929 3948 16968
rect 4004 16929 4056 16968
rect 4112 16929 4164 16968
rect 5952 16929 6004 16968
rect 6060 16929 6112 16968
rect 6168 16929 6220 16968
rect 6276 16929 6328 16968
rect 6384 16929 6436 16968
rect 8628 16929 8680 16968
rect 8736 16929 8788 16968
rect 8844 16929 8896 16968
rect 8952 16929 9004 16968
rect 9060 16929 9112 16968
rect 10900 16929 10952 16968
rect 11008 16929 11060 16968
rect 11116 16929 11168 16968
rect 11224 16929 11276 16968
rect 11332 16929 11384 16968
rect 3680 16916 3732 16929
rect 3788 16916 3840 16929
rect 3896 16916 3948 16929
rect 4004 16916 4056 16929
rect 4112 16916 4164 16929
rect 5952 16916 6004 16929
rect 6060 16916 6112 16929
rect 6168 16916 6220 16929
rect 6276 16916 6328 16929
rect 6384 16916 6436 16929
rect 8628 16916 8680 16929
rect 8736 16916 8788 16929
rect 8844 16916 8896 16929
rect 8952 16916 9004 16929
rect 9060 16916 9112 16929
rect 10900 16916 10952 16929
rect 11008 16916 11060 16929
rect 11116 16916 11168 16929
rect 11224 16916 11276 16929
rect 11332 16916 11384 16929
rect 3680 16847 3732 16860
rect 3788 16847 3840 16860
rect 3896 16847 3948 16860
rect 4004 16847 4056 16860
rect 4112 16847 4164 16860
rect 5952 16847 6004 16860
rect 6060 16847 6112 16860
rect 6168 16847 6220 16860
rect 6276 16847 6328 16860
rect 6384 16847 6436 16860
rect 8628 16847 8680 16860
rect 8736 16847 8788 16860
rect 8844 16847 8896 16860
rect 8952 16847 9004 16860
rect 9060 16847 9112 16860
rect 10900 16847 10952 16860
rect 11008 16847 11060 16860
rect 11116 16847 11168 16860
rect 11224 16847 11276 16860
rect 11332 16847 11384 16860
rect 3680 16808 3732 16847
rect 3788 16808 3840 16847
rect 3896 16808 3948 16847
rect 4004 16808 4056 16847
rect 4112 16808 4164 16847
rect 5952 16808 6004 16847
rect 6060 16808 6112 16847
rect 6168 16808 6220 16847
rect 6276 16808 6328 16847
rect 6384 16808 6436 16847
rect 8628 16808 8680 16847
rect 8736 16808 8788 16847
rect 8844 16808 8896 16847
rect 8952 16808 9004 16847
rect 9060 16808 9112 16847
rect 10900 16808 10952 16847
rect 11008 16808 11060 16847
rect 11116 16808 11168 16847
rect 11224 16808 11276 16847
rect 11332 16808 11384 16847
rect 4816 16575 4868 16601
rect 4924 16575 4976 16601
rect 5032 16575 5084 16601
rect 5140 16575 5192 16601
rect 5248 16575 5300 16601
rect 7101 16575 7153 16601
rect 7209 16575 7261 16601
rect 7317 16575 7369 16601
rect 7425 16575 7477 16601
rect 7587 16575 7639 16601
rect 7695 16575 7747 16601
rect 7803 16575 7855 16601
rect 7911 16575 7963 16601
rect 9764 16575 9816 16601
rect 9872 16575 9924 16601
rect 9980 16575 10032 16601
rect 10088 16575 10140 16601
rect 10196 16575 10248 16601
rect 4816 16549 4868 16575
rect 4924 16549 4976 16575
rect 5032 16549 5084 16575
rect 5140 16549 5192 16575
rect 5248 16549 5300 16575
rect 7101 16549 7153 16575
rect 7209 16549 7261 16575
rect 7317 16549 7369 16575
rect 7425 16549 7477 16575
rect 7587 16549 7639 16575
rect 7695 16549 7747 16575
rect 7803 16549 7855 16575
rect 7911 16549 7963 16575
rect 9764 16549 9816 16575
rect 9872 16549 9924 16575
rect 9980 16549 10032 16575
rect 10088 16549 10140 16575
rect 10196 16549 10248 16575
rect 4816 16467 4868 16493
rect 4924 16467 4976 16493
rect 5032 16467 5084 16493
rect 5140 16467 5192 16493
rect 5248 16467 5300 16493
rect 7101 16467 7153 16493
rect 7209 16467 7261 16493
rect 7317 16467 7369 16493
rect 7425 16467 7477 16493
rect 7587 16467 7639 16493
rect 7695 16467 7747 16493
rect 7803 16467 7855 16493
rect 7911 16467 7963 16493
rect 9764 16467 9816 16493
rect 9872 16467 9924 16493
rect 9980 16467 10032 16493
rect 10088 16467 10140 16493
rect 10196 16467 10248 16493
rect 4816 16441 4868 16467
rect 4924 16441 4976 16467
rect 5032 16441 5084 16467
rect 5140 16441 5192 16467
rect 5248 16441 5300 16467
rect 7101 16441 7153 16467
rect 7209 16441 7261 16467
rect 7317 16441 7369 16467
rect 7425 16441 7477 16467
rect 7587 16441 7639 16467
rect 7695 16441 7747 16467
rect 7803 16441 7855 16467
rect 7911 16441 7963 16467
rect 9764 16441 9816 16467
rect 9872 16441 9924 16467
rect 9980 16441 10032 16467
rect 10088 16441 10140 16467
rect 10196 16441 10248 16467
rect 3680 16031 3732 16083
rect 3788 16031 3840 16083
rect 3896 16031 3948 16083
rect 4004 16031 4056 16083
rect 4112 16031 4164 16083
rect 5952 16031 6004 16083
rect 6060 16031 6112 16083
rect 6168 16031 6220 16083
rect 6276 16031 6328 16083
rect 6384 16031 6436 16083
rect 8628 16031 8680 16083
rect 8736 16031 8788 16083
rect 8844 16031 8896 16083
rect 8952 16031 9004 16083
rect 9060 16031 9112 16083
rect 10900 16031 10952 16083
rect 11008 16031 11060 16083
rect 11116 16031 11168 16083
rect 11224 16031 11276 16083
rect 11332 16031 11384 16083
rect 3680 15923 3732 15975
rect 3788 15923 3840 15975
rect 3896 15923 3948 15975
rect 4004 15923 4056 15975
rect 4112 15923 4164 15975
rect 5952 15923 6004 15975
rect 6060 15923 6112 15975
rect 6168 15923 6220 15975
rect 6276 15923 6328 15975
rect 6384 15923 6436 15975
rect 8628 15923 8680 15975
rect 8736 15923 8788 15975
rect 8844 15923 8896 15975
rect 8952 15923 9004 15975
rect 9060 15923 9112 15975
rect 10900 15923 10952 15975
rect 11008 15923 11060 15975
rect 11116 15923 11168 15975
rect 11224 15923 11276 15975
rect 11332 15923 11384 15975
rect 3680 15815 3732 15867
rect 3788 15815 3840 15867
rect 3896 15815 3948 15867
rect 4004 15815 4056 15867
rect 4112 15815 4164 15867
rect 5952 15815 6004 15867
rect 6060 15815 6112 15867
rect 6168 15815 6220 15867
rect 6276 15815 6328 15867
rect 6384 15815 6436 15867
rect 8628 15815 8680 15867
rect 8736 15815 8788 15867
rect 8844 15815 8896 15867
rect 8952 15815 9004 15867
rect 9060 15815 9112 15867
rect 10900 15815 10952 15867
rect 11008 15815 11060 15867
rect 11116 15815 11168 15867
rect 11224 15815 11276 15867
rect 11332 15815 11384 15867
<< metal2 >>
rect 260 56922 768 56975
rect 260 56866 300 56922
rect 356 56866 424 56922
rect 480 56866 548 56922
rect 604 56866 672 56922
rect 728 56866 768 56922
rect 260 56798 768 56866
rect 260 56742 300 56798
rect 356 56742 424 56798
rect 480 56742 548 56798
rect 604 56742 672 56798
rect 728 56742 768 56798
rect 260 56711 768 56742
rect 260 56674 444 56711
rect 496 56674 552 56711
rect 260 56618 300 56674
rect 356 56618 424 56674
rect 496 56659 548 56674
rect 604 56659 660 56711
rect 712 56674 768 56711
rect 480 56618 548 56659
rect 604 56618 672 56659
rect 728 56618 768 56674
rect 260 56603 768 56618
rect 260 56551 444 56603
rect 496 56551 552 56603
rect 604 56551 660 56603
rect 712 56551 768 56603
rect 260 56550 768 56551
rect 260 56494 300 56550
rect 356 56494 424 56550
rect 480 56495 548 56550
rect 604 56495 672 56550
rect 496 56494 548 56495
rect 260 56443 444 56494
rect 496 56443 552 56494
rect 604 56443 660 56495
rect 728 56494 768 56550
rect 712 56443 768 56494
rect 260 56426 768 56443
rect 260 56370 300 56426
rect 356 56370 424 56426
rect 480 56370 548 56426
rect 604 56370 672 56426
rect 728 56370 768 56426
rect 260 56302 768 56370
rect 1396 56922 1904 56975
rect 1396 56866 1436 56922
rect 1492 56866 1560 56922
rect 1616 56866 1684 56922
rect 1740 56866 1808 56922
rect 1864 56866 1904 56922
rect 1396 56798 1904 56866
rect 1396 56742 1436 56798
rect 1492 56742 1560 56798
rect 1616 56742 1684 56798
rect 1740 56742 1808 56798
rect 1864 56742 1904 56798
rect 1396 56711 1904 56742
rect 1396 56659 1408 56711
rect 1460 56674 1516 56711
rect 1568 56674 1624 56711
rect 1492 56659 1516 56674
rect 1616 56659 1624 56674
rect 1676 56674 1732 56711
rect 1784 56674 1840 56711
rect 1676 56659 1684 56674
rect 1784 56659 1808 56674
rect 1892 56659 1904 56711
rect 1396 56618 1436 56659
rect 1492 56618 1560 56659
rect 1616 56618 1684 56659
rect 1740 56618 1808 56659
rect 1864 56618 1904 56659
rect 1396 56603 1904 56618
rect 1396 56551 1408 56603
rect 1460 56551 1516 56603
rect 1568 56551 1624 56603
rect 1676 56551 1732 56603
rect 1784 56551 1840 56603
rect 1892 56551 1904 56603
rect 1396 56550 1904 56551
rect 1396 56495 1436 56550
rect 1492 56495 1560 56550
rect 1616 56495 1684 56550
rect 1740 56495 1808 56550
rect 1864 56495 1904 56550
rect 1396 56443 1408 56495
rect 1492 56494 1516 56495
rect 1616 56494 1624 56495
rect 1460 56443 1516 56494
rect 1568 56443 1624 56494
rect 1676 56494 1684 56495
rect 1784 56494 1808 56495
rect 1676 56443 1732 56494
rect 1784 56443 1840 56494
rect 1892 56443 1904 56495
rect 1396 56426 1904 56443
rect 1396 56370 1436 56426
rect 1492 56370 1560 56426
rect 1616 56370 1684 56426
rect 1740 56370 1808 56426
rect 1864 56370 1904 56426
rect 260 56246 300 56302
rect 356 56246 424 56302
rect 480 56246 548 56302
rect 604 56246 672 56302
rect 728 56246 768 56302
rect 260 56178 768 56246
rect 260 56122 300 56178
rect 356 56122 424 56178
rect 480 56122 548 56178
rect 604 56122 672 56178
rect 728 56122 768 56178
rect 260 56054 768 56122
rect 260 55998 300 56054
rect 356 55998 424 56054
rect 480 55998 548 56054
rect 604 55998 672 56054
rect 728 55998 768 56054
rect 260 55930 768 55998
rect 260 55874 300 55930
rect 356 55874 424 55930
rect 480 55874 548 55930
rect 604 55874 672 55930
rect 728 55874 768 55930
rect 260 55806 768 55874
rect 260 55750 300 55806
rect 356 55750 424 55806
rect 480 55750 548 55806
rect 604 55750 672 55806
rect 728 55750 768 55806
rect 260 53845 768 55750
rect 966 56324 1290 56336
rect 966 56272 978 56324
rect 1030 56272 1102 56324
rect 1154 56272 1226 56324
rect 1278 56272 1290 56324
rect 966 56200 1290 56272
rect 966 56148 978 56200
rect 1030 56148 1102 56200
rect 1154 56148 1226 56200
rect 1278 56148 1290 56200
rect 966 56076 1290 56148
rect 966 56024 978 56076
rect 1030 56024 1102 56076
rect 1154 56024 1226 56076
rect 1278 56024 1290 56076
rect 966 55952 1290 56024
rect 966 55900 978 55952
rect 1030 55900 1102 55952
rect 1154 55900 1226 55952
rect 1278 55900 1290 55952
rect 966 55828 1290 55900
rect 966 55776 978 55828
rect 1030 55776 1102 55828
rect 1154 55776 1226 55828
rect 1278 55776 1290 55828
rect 966 55704 1290 55776
rect 966 55652 978 55704
rect 1030 55652 1102 55704
rect 1154 55652 1226 55704
rect 1278 55652 1290 55704
rect 966 55580 1290 55652
rect 966 55528 978 55580
rect 1030 55528 1102 55580
rect 1154 55528 1226 55580
rect 1278 55528 1290 55580
rect 966 55456 1290 55528
rect 966 55455 978 55456
rect 858 55445 978 55455
rect 1030 55445 1102 55456
rect 1154 55445 1226 55456
rect 1278 55455 1290 55456
rect 1396 56302 1904 56370
rect 1396 56246 1436 56302
rect 1492 56246 1560 56302
rect 1616 56246 1684 56302
rect 1740 56246 1808 56302
rect 1864 56246 1904 56302
rect 1396 56178 1904 56246
rect 1396 56122 1436 56178
rect 1492 56122 1560 56178
rect 1616 56122 1684 56178
rect 1740 56122 1808 56178
rect 1864 56122 1904 56178
rect 1396 56054 1904 56122
rect 1396 55998 1436 56054
rect 1492 55998 1560 56054
rect 1616 55998 1684 56054
rect 1740 55998 1808 56054
rect 1864 55998 1904 56054
rect 1396 55930 1904 55998
rect 1396 55874 1436 55930
rect 1492 55874 1560 55930
rect 1616 55874 1684 55930
rect 1740 55874 1808 55930
rect 1864 55874 1904 55930
rect 1396 55806 1904 55874
rect 1396 55750 1436 55806
rect 1492 55750 1560 55806
rect 1616 55750 1684 55806
rect 1740 55750 1808 55806
rect 1864 55750 1904 55806
rect 1278 55445 1306 55455
rect 858 55389 868 55445
rect 924 55404 978 55445
rect 1048 55404 1102 55445
rect 1172 55404 1226 55445
rect 924 55389 992 55404
rect 1048 55389 1116 55404
rect 1172 55389 1240 55404
rect 1296 55389 1306 55445
rect 858 55332 1306 55389
rect 858 55321 978 55332
rect 1030 55321 1102 55332
rect 1154 55321 1226 55332
rect 1278 55321 1306 55332
rect 858 55265 868 55321
rect 924 55280 978 55321
rect 1048 55280 1102 55321
rect 1172 55280 1226 55321
rect 924 55265 992 55280
rect 1048 55265 1116 55280
rect 1172 55265 1240 55280
rect 1296 55265 1306 55321
rect 858 55208 1306 55265
rect 858 55197 978 55208
rect 1030 55197 1102 55208
rect 1154 55197 1226 55208
rect 1278 55197 1306 55208
rect 858 55141 868 55197
rect 924 55156 978 55197
rect 1048 55156 1102 55197
rect 1172 55156 1226 55197
rect 924 55141 992 55156
rect 1048 55141 1116 55156
rect 1172 55141 1240 55156
rect 1296 55141 1306 55197
rect 858 55084 1306 55141
rect 858 55073 978 55084
rect 1030 55073 1102 55084
rect 1154 55073 1226 55084
rect 1278 55073 1306 55084
rect 858 55017 868 55073
rect 924 55032 978 55073
rect 1048 55032 1102 55073
rect 1172 55032 1226 55073
rect 924 55017 992 55032
rect 1048 55017 1116 55032
rect 1172 55017 1240 55032
rect 1296 55017 1306 55073
rect 858 54960 1306 55017
rect 858 54949 978 54960
rect 1030 54949 1102 54960
rect 1154 54949 1226 54960
rect 1278 54949 1306 54960
rect 858 54893 868 54949
rect 924 54908 978 54949
rect 1048 54908 1102 54949
rect 1172 54908 1226 54949
rect 924 54893 992 54908
rect 1048 54893 1116 54908
rect 1172 54893 1240 54908
rect 1296 54893 1306 54949
rect 858 54836 1306 54893
rect 858 54825 978 54836
rect 1030 54825 1102 54836
rect 1154 54825 1226 54836
rect 1278 54825 1306 54836
rect 858 54769 868 54825
rect 924 54784 978 54825
rect 1048 54784 1102 54825
rect 1172 54784 1226 54825
rect 924 54769 992 54784
rect 1048 54769 1116 54784
rect 1172 54769 1240 54784
rect 1296 54769 1306 54825
rect 858 54712 1306 54769
rect 858 54701 978 54712
rect 1030 54701 1102 54712
rect 1154 54701 1226 54712
rect 1278 54701 1306 54712
rect 858 54645 868 54701
rect 924 54660 978 54701
rect 1048 54660 1102 54701
rect 1172 54660 1226 54701
rect 924 54645 992 54660
rect 1048 54645 1116 54660
rect 1172 54645 1240 54660
rect 1296 54645 1306 54701
rect 858 54588 1306 54645
rect 858 54577 978 54588
rect 1030 54577 1102 54588
rect 1154 54577 1226 54588
rect 1278 54577 1306 54588
rect 858 54521 868 54577
rect 924 54536 978 54577
rect 1048 54536 1102 54577
rect 1172 54536 1226 54577
rect 924 54521 992 54536
rect 1048 54521 1116 54536
rect 1172 54521 1240 54536
rect 1296 54521 1306 54577
rect 858 54464 1306 54521
rect 858 54453 978 54464
rect 1030 54453 1102 54464
rect 1154 54453 1226 54464
rect 1278 54453 1306 54464
rect 858 54397 868 54453
rect 924 54412 978 54453
rect 1048 54412 1102 54453
rect 1172 54412 1226 54453
rect 924 54397 992 54412
rect 1048 54397 1116 54412
rect 1172 54397 1240 54412
rect 1296 54397 1306 54453
rect 858 54340 1306 54397
rect 858 54329 978 54340
rect 1030 54329 1102 54340
rect 1154 54329 1226 54340
rect 1278 54329 1306 54340
rect 858 54273 868 54329
rect 924 54288 978 54329
rect 1048 54288 1102 54329
rect 1172 54288 1226 54329
rect 924 54273 992 54288
rect 1048 54273 1116 54288
rect 1172 54273 1240 54288
rect 1296 54273 1306 54329
rect 858 54216 1306 54273
rect 858 54205 978 54216
rect 1030 54205 1102 54216
rect 1154 54205 1226 54216
rect 1278 54205 1306 54216
rect 858 54149 868 54205
rect 924 54164 978 54205
rect 1048 54164 1102 54205
rect 1172 54164 1226 54205
rect 924 54149 992 54164
rect 1048 54149 1116 54164
rect 1172 54149 1240 54164
rect 1296 54149 1306 54205
rect 858 54139 1306 54149
rect 260 53789 300 53845
rect 356 53789 424 53845
rect 480 53789 548 53845
rect 604 53789 672 53845
rect 728 53789 768 53845
rect 260 53721 768 53789
rect 260 53665 300 53721
rect 356 53665 424 53721
rect 480 53665 548 53721
rect 604 53665 672 53721
rect 728 53665 768 53721
rect 260 53597 768 53665
rect 260 53541 300 53597
rect 356 53541 424 53597
rect 480 53541 548 53597
rect 604 53541 672 53597
rect 728 53541 768 53597
rect 260 53473 768 53541
rect 260 53417 300 53473
rect 356 53417 424 53473
rect 480 53417 548 53473
rect 604 53417 672 53473
rect 728 53417 768 53473
rect 260 53349 768 53417
rect 260 53293 300 53349
rect 356 53293 424 53349
rect 480 53293 548 53349
rect 604 53293 672 53349
rect 728 53293 768 53349
rect 260 53225 768 53293
rect 260 53169 300 53225
rect 356 53169 424 53225
rect 480 53169 548 53225
rect 604 53169 672 53225
rect 728 53169 768 53225
rect 260 53101 768 53169
rect 966 54092 1290 54139
rect 966 54040 978 54092
rect 1030 54040 1102 54092
rect 1154 54040 1226 54092
rect 1278 54040 1290 54092
rect 966 53968 1290 54040
rect 966 53916 978 53968
rect 1030 53916 1102 53968
rect 1154 53916 1226 53968
rect 1278 53916 1290 53968
rect 966 53844 1290 53916
rect 966 53792 978 53844
rect 1030 53792 1102 53844
rect 1154 53792 1226 53844
rect 1278 53792 1290 53844
rect 966 53720 1290 53792
rect 966 53668 978 53720
rect 1030 53668 1102 53720
rect 1154 53668 1226 53720
rect 1278 53668 1290 53720
rect 966 53596 1290 53668
rect 966 53544 978 53596
rect 1030 53544 1102 53596
rect 1154 53544 1226 53596
rect 1278 53544 1290 53596
rect 966 53472 1290 53544
rect 966 53420 978 53472
rect 1030 53420 1102 53472
rect 1154 53420 1226 53472
rect 1278 53420 1290 53472
rect 966 53348 1290 53420
rect 966 53296 978 53348
rect 1030 53296 1102 53348
rect 1154 53296 1226 53348
rect 1278 53296 1290 53348
rect 966 53224 1290 53296
rect 966 53172 978 53224
rect 1030 53172 1102 53224
rect 1154 53172 1226 53224
rect 1278 53172 1290 53224
rect 966 53160 1290 53172
rect 1396 53845 1904 55750
rect 1396 53789 1436 53845
rect 1492 53789 1560 53845
rect 1616 53789 1684 53845
rect 1740 53789 1808 53845
rect 1864 53789 1904 53845
rect 1396 53721 1904 53789
rect 1396 53665 1436 53721
rect 1492 53665 1560 53721
rect 1616 53665 1684 53721
rect 1740 53665 1808 53721
rect 1864 53665 1904 53721
rect 1396 53597 1904 53665
rect 1396 53541 1436 53597
rect 1492 53541 1560 53597
rect 1616 53541 1684 53597
rect 1740 53541 1808 53597
rect 1864 53541 1904 53597
rect 1396 53473 1904 53541
rect 1396 53417 1436 53473
rect 1492 53417 1560 53473
rect 1616 53417 1684 53473
rect 1740 53417 1808 53473
rect 1864 53417 1904 53473
rect 1396 53349 1904 53417
rect 1396 53293 1436 53349
rect 1492 53293 1560 53349
rect 1616 53293 1684 53349
rect 1740 53293 1808 53349
rect 1864 53293 1904 53349
rect 1396 53225 1904 53293
rect 1396 53169 1436 53225
rect 1492 53169 1560 53225
rect 1616 53169 1684 53225
rect 1740 53169 1808 53225
rect 1864 53169 1904 53225
rect 260 53045 300 53101
rect 356 53045 424 53101
rect 480 53045 548 53101
rect 604 53045 672 53101
rect 728 53045 768 53101
rect 260 53016 768 53045
rect 260 52977 444 53016
rect 496 52977 552 53016
rect 260 52921 300 52977
rect 356 52921 424 52977
rect 496 52964 548 52977
rect 604 52964 660 53016
rect 712 52977 768 53016
rect 480 52921 548 52964
rect 604 52921 672 52964
rect 728 52921 768 52977
rect 260 52908 768 52921
rect 260 52856 444 52908
rect 496 52856 552 52908
rect 604 52856 660 52908
rect 712 52856 768 52908
rect 260 52853 768 52856
rect 260 52797 300 52853
rect 356 52797 424 52853
rect 480 52800 548 52853
rect 604 52800 672 52853
rect 496 52797 548 52800
rect 260 52748 444 52797
rect 496 52748 552 52797
rect 604 52748 660 52800
rect 728 52797 768 52853
rect 712 52748 768 52797
rect 260 52729 768 52748
rect 260 52673 300 52729
rect 356 52673 424 52729
rect 480 52692 548 52729
rect 604 52692 672 52729
rect 496 52673 548 52692
rect 260 52640 444 52673
rect 496 52640 552 52673
rect 604 52640 660 52692
rect 728 52673 768 52729
rect 712 52640 768 52673
rect 260 52605 768 52640
rect 260 52549 300 52605
rect 356 52549 424 52605
rect 480 52584 548 52605
rect 604 52584 672 52605
rect 496 52549 548 52584
rect 260 52532 444 52549
rect 496 52532 552 52549
rect 604 52532 660 52584
rect 728 52549 768 52605
rect 712 52532 768 52549
rect 32 52273 122 52297
rect 32 50921 56 52273
rect 112 50921 122 52273
rect 32 50897 122 50921
rect 260 49068 768 52532
rect 1136 52376 1336 53160
rect 1136 52324 1148 52376
rect 1200 52324 1272 52376
rect 1324 52324 1336 52376
rect 1136 52252 1336 52324
rect 1136 52200 1148 52252
rect 1200 52200 1272 52252
rect 1324 52200 1336 52252
rect 1136 52128 1336 52200
rect 1136 52076 1148 52128
rect 1200 52076 1272 52128
rect 1324 52076 1336 52128
rect 1136 52004 1336 52076
rect 1136 51952 1148 52004
rect 1200 51952 1272 52004
rect 1324 51952 1336 52004
rect 1136 51880 1336 51952
rect 1136 51828 1148 51880
rect 1200 51828 1272 51880
rect 1324 51828 1336 51880
rect 1136 51756 1336 51828
rect 1136 51704 1148 51756
rect 1200 51704 1272 51756
rect 1324 51704 1336 51756
rect 1136 51632 1336 51704
rect 1136 51580 1148 51632
rect 1200 51580 1272 51632
rect 1324 51580 1336 51632
rect 1136 51508 1336 51580
rect 1136 51456 1148 51508
rect 1200 51456 1272 51508
rect 1324 51456 1336 51508
rect 1136 51384 1336 51456
rect 1136 51332 1148 51384
rect 1200 51332 1272 51384
rect 1324 51332 1336 51384
rect 1136 51260 1336 51332
rect 1136 51208 1148 51260
rect 1200 51208 1272 51260
rect 1324 51208 1336 51260
rect 1136 51136 1336 51208
rect 1136 51084 1148 51136
rect 1200 51084 1272 51136
rect 1324 51084 1336 51136
rect 1136 51012 1336 51084
rect 1136 50960 1148 51012
rect 1200 50960 1272 51012
rect 1324 50960 1336 51012
rect 1136 50888 1336 50960
rect 1136 50836 1148 50888
rect 1200 50836 1272 50888
rect 1324 50836 1336 50888
rect 1136 50764 1336 50836
rect 1136 50712 1148 50764
rect 1200 50712 1272 50764
rect 1324 50712 1336 50764
rect 260 49045 444 49068
rect 496 49045 552 49068
rect 260 48989 300 49045
rect 356 48989 424 49045
rect 496 49016 548 49045
rect 604 49016 660 49068
rect 712 49045 768 49068
rect 480 48989 548 49016
rect 604 48989 672 49016
rect 728 48989 768 49045
rect 260 48960 768 48989
rect 260 48921 444 48960
rect 496 48921 552 48960
rect 260 48865 300 48921
rect 356 48865 424 48921
rect 496 48908 548 48921
rect 604 48908 660 48960
rect 712 48921 768 48960
rect 480 48865 548 48908
rect 604 48865 672 48908
rect 728 48865 768 48921
rect 260 48852 768 48865
rect 260 48800 444 48852
rect 496 48800 552 48852
rect 604 48800 660 48852
rect 712 48800 768 48852
rect 260 48797 768 48800
rect 260 48741 300 48797
rect 356 48741 424 48797
rect 480 48744 548 48797
rect 604 48744 672 48797
rect 496 48741 548 48744
rect 260 48692 444 48741
rect 496 48692 552 48741
rect 604 48692 660 48744
rect 728 48741 768 48797
rect 712 48692 768 48741
rect 260 48673 768 48692
rect 260 48617 300 48673
rect 356 48617 424 48673
rect 480 48636 548 48673
rect 604 48636 672 48673
rect 496 48617 548 48636
rect 260 48584 444 48617
rect 496 48584 552 48617
rect 604 48584 660 48636
rect 728 48617 768 48673
rect 712 48584 768 48617
rect 260 48549 768 48584
rect 260 48493 300 48549
rect 356 48493 424 48549
rect 480 48493 548 48549
rect 604 48493 672 48549
rect 728 48493 768 48549
rect 260 48425 768 48493
rect 260 48369 300 48425
rect 356 48369 424 48425
rect 480 48369 548 48425
rect 604 48369 672 48425
rect 728 48369 768 48425
rect 260 48301 768 48369
rect 260 48245 300 48301
rect 356 48245 424 48301
rect 480 48245 548 48301
rect 604 48245 672 48301
rect 728 48245 768 48301
rect 260 48177 768 48245
rect 260 48121 300 48177
rect 356 48121 424 48177
rect 480 48121 548 48177
rect 604 48121 672 48177
rect 728 48121 768 48177
rect 260 48053 768 48121
rect 260 47997 300 48053
rect 356 47997 424 48053
rect 480 47997 548 48053
rect 604 47997 672 48053
rect 728 47997 768 48053
rect 260 47929 768 47997
rect 260 47873 300 47929
rect 356 47873 424 47929
rect 480 47873 548 47929
rect 604 47873 672 47929
rect 728 47873 768 47929
rect 260 47805 768 47873
rect 260 47749 300 47805
rect 356 47749 424 47805
rect 480 47749 548 47805
rect 604 47749 672 47805
rect 728 47749 768 47805
rect 260 45845 768 47749
rect 260 45789 300 45845
rect 356 45789 424 45845
rect 480 45789 548 45845
rect 604 45789 672 45845
rect 728 45789 768 45845
rect 260 45721 768 45789
rect 260 45665 300 45721
rect 356 45665 424 45721
rect 480 45665 548 45721
rect 604 45665 672 45721
rect 728 45665 768 45721
rect 260 45597 768 45665
rect 260 45541 300 45597
rect 356 45541 424 45597
rect 480 45541 548 45597
rect 604 45541 672 45597
rect 728 45541 768 45597
rect 260 45473 768 45541
rect 260 45417 300 45473
rect 356 45417 424 45473
rect 480 45417 548 45473
rect 604 45417 672 45473
rect 728 45417 768 45473
rect 260 45349 768 45417
rect 260 45293 300 45349
rect 356 45293 424 45349
rect 480 45293 548 45349
rect 604 45293 672 45349
rect 728 45293 768 45349
rect 260 45225 768 45293
rect 260 45169 300 45225
rect 356 45169 424 45225
rect 480 45169 548 45225
rect 604 45169 672 45225
rect 728 45169 768 45225
rect 260 45120 768 45169
rect 260 45101 444 45120
rect 496 45101 552 45120
rect 260 45045 300 45101
rect 356 45045 424 45101
rect 496 45068 548 45101
rect 604 45068 660 45120
rect 712 45101 768 45120
rect 480 45045 548 45068
rect 604 45045 672 45068
rect 728 45045 768 45101
rect 260 45012 768 45045
rect 260 44977 444 45012
rect 496 44977 552 45012
rect 260 44921 300 44977
rect 356 44921 424 44977
rect 496 44960 548 44977
rect 604 44960 660 45012
rect 712 44977 768 45012
rect 480 44921 548 44960
rect 604 44921 672 44960
rect 728 44921 768 44977
rect 260 44904 768 44921
rect 260 44853 444 44904
rect 496 44853 552 44904
rect 260 44797 300 44853
rect 356 44797 424 44853
rect 496 44852 548 44853
rect 604 44852 660 44904
rect 712 44853 768 44904
rect 480 44797 548 44852
rect 604 44797 672 44852
rect 728 44797 768 44853
rect 260 44796 768 44797
rect 260 44744 444 44796
rect 496 44744 552 44796
rect 604 44744 660 44796
rect 712 44744 768 44796
rect 260 44729 768 44744
rect 260 44673 300 44729
rect 356 44673 424 44729
rect 480 44688 548 44729
rect 604 44688 672 44729
rect 496 44673 548 44688
rect 260 44636 444 44673
rect 496 44636 552 44673
rect 604 44636 660 44688
rect 728 44673 768 44729
rect 712 44636 768 44673
rect 260 44605 768 44636
rect 260 44549 300 44605
rect 356 44549 424 44605
rect 480 44549 548 44605
rect 604 44549 672 44605
rect 728 44549 768 44605
rect 260 41172 768 44549
rect 260 41120 444 41172
rect 496 41120 552 41172
rect 604 41120 660 41172
rect 712 41120 768 41172
rect 260 41064 768 41120
rect 260 41012 444 41064
rect 496 41012 552 41064
rect 604 41012 660 41064
rect 712 41012 768 41064
rect 260 40956 768 41012
rect 260 40904 444 40956
rect 496 40904 552 40956
rect 604 40904 660 40956
rect 712 40904 768 40956
rect 260 40848 768 40904
rect 260 40796 444 40848
rect 496 40796 552 40848
rect 604 40796 660 40848
rect 712 40796 768 40848
rect 260 40740 768 40796
rect 260 40688 444 40740
rect 496 40688 552 40740
rect 604 40688 660 40740
rect 712 40688 768 40740
rect 32 37873 122 37897
rect 32 36521 56 37873
rect 112 36521 122 37873
rect 32 36497 122 36521
rect 260 37224 768 40688
rect 828 50645 1028 50697
rect 828 50589 838 50645
rect 894 50589 962 50645
rect 1018 50589 1028 50645
rect 828 50521 1028 50589
rect 828 50465 838 50521
rect 894 50465 962 50521
rect 1018 50465 1028 50521
rect 828 50397 1028 50465
rect 828 50341 838 50397
rect 894 50341 962 50397
rect 1018 50341 1028 50397
rect 828 50273 1028 50341
rect 828 50217 838 50273
rect 894 50217 962 50273
rect 1018 50217 1028 50273
rect 828 50149 1028 50217
rect 828 50093 838 50149
rect 894 50093 962 50149
rect 1018 50093 1028 50149
rect 828 50025 1028 50093
rect 828 49969 838 50025
rect 894 49969 962 50025
rect 1018 49969 1028 50025
rect 828 49901 1028 49969
rect 828 49845 838 49901
rect 894 49845 962 49901
rect 1018 49845 1028 49901
rect 828 49777 1028 49845
rect 828 49721 838 49777
rect 894 49721 962 49777
rect 1018 49721 1028 49777
rect 828 49653 1028 49721
rect 828 49597 838 49653
rect 894 49597 962 49653
rect 1018 49597 1028 49653
rect 828 49529 1028 49597
rect 828 49473 838 49529
rect 894 49473 962 49529
rect 1018 49473 1028 49529
rect 828 49405 1028 49473
rect 828 49349 838 49405
rect 894 49349 962 49405
rect 1018 49349 1028 49405
rect 828 39445 1028 49349
rect 828 39389 838 39445
rect 894 39389 962 39445
rect 1018 39389 1028 39445
rect 828 39321 1028 39389
rect 828 39265 838 39321
rect 894 39265 962 39321
rect 1018 39265 1028 39321
rect 828 39197 1028 39265
rect 828 39141 838 39197
rect 894 39141 962 39197
rect 1018 39141 1028 39197
rect 828 39073 1028 39141
rect 828 39017 838 39073
rect 894 39017 962 39073
rect 1018 39017 1028 39073
rect 828 38949 1028 39017
rect 828 38893 838 38949
rect 894 38893 962 38949
rect 1018 38893 1028 38949
rect 828 38825 1028 38893
rect 828 38769 838 38825
rect 894 38769 962 38825
rect 1018 38769 1028 38825
rect 828 38701 1028 38769
rect 828 38645 838 38701
rect 894 38645 962 38701
rect 1018 38645 1028 38701
rect 828 38577 1028 38645
rect 828 38521 838 38577
rect 894 38521 962 38577
rect 1018 38521 1028 38577
rect 828 38453 1028 38521
rect 828 38397 838 38453
rect 894 38397 962 38453
rect 1018 38397 1028 38453
rect 828 38329 1028 38397
rect 828 38273 838 38329
rect 894 38273 962 38329
rect 1018 38273 1028 38329
rect 828 38205 1028 38273
rect 828 38149 838 38205
rect 894 38149 962 38205
rect 1018 38149 1028 38205
rect 828 38097 1028 38149
rect 1136 50640 1336 50712
rect 1136 50588 1148 50640
rect 1200 50588 1272 50640
rect 1324 50588 1336 50640
rect 1136 50516 1336 50588
rect 1136 50464 1148 50516
rect 1200 50464 1272 50516
rect 1324 50464 1336 50516
rect 1136 50392 1336 50464
rect 1136 50340 1148 50392
rect 1200 50340 1272 50392
rect 1324 50340 1336 50392
rect 1136 50268 1336 50340
rect 1136 50216 1148 50268
rect 1200 50216 1272 50268
rect 1324 50216 1336 50268
rect 1136 50144 1336 50216
rect 1136 50092 1148 50144
rect 1200 50092 1272 50144
rect 1324 50092 1336 50144
rect 1136 50020 1336 50092
rect 1136 49968 1148 50020
rect 1200 49968 1272 50020
rect 1324 49968 1336 50020
rect 1136 49896 1336 49968
rect 1136 49844 1148 49896
rect 1200 49844 1272 49896
rect 1324 49844 1336 49896
rect 1136 49772 1336 49844
rect 1136 49720 1148 49772
rect 1200 49720 1272 49772
rect 1324 49720 1336 49772
rect 1136 49648 1336 49720
rect 1136 49596 1148 49648
rect 1200 49596 1272 49648
rect 1324 49596 1336 49648
rect 1136 49524 1336 49596
rect 1136 49472 1148 49524
rect 1200 49472 1272 49524
rect 1324 49472 1336 49524
rect 1136 49400 1336 49472
rect 1136 49348 1148 49400
rect 1200 49348 1272 49400
rect 1324 49348 1336 49400
rect 1136 49276 1336 49348
rect 1136 49224 1148 49276
rect 1200 49224 1272 49276
rect 1324 49224 1336 49276
rect 1136 48428 1336 49224
rect 1136 48376 1148 48428
rect 1200 48376 1272 48428
rect 1324 48376 1336 48428
rect 1136 48304 1336 48376
rect 1136 48252 1148 48304
rect 1200 48252 1272 48304
rect 1324 48252 1336 48304
rect 1136 48180 1336 48252
rect 1136 48128 1148 48180
rect 1200 48128 1272 48180
rect 1324 48128 1336 48180
rect 1136 48056 1336 48128
rect 1136 48004 1148 48056
rect 1200 48004 1272 48056
rect 1324 48004 1336 48056
rect 1136 47932 1336 48004
rect 1136 47880 1148 47932
rect 1200 47880 1272 47932
rect 1324 47880 1336 47932
rect 1136 47808 1336 47880
rect 1136 47756 1148 47808
rect 1200 47756 1272 47808
rect 1324 47756 1336 47808
rect 1136 47684 1336 47756
rect 1136 47632 1148 47684
rect 1200 47632 1272 47684
rect 1324 47632 1336 47684
rect 1136 47560 1336 47632
rect 1136 47508 1148 47560
rect 1200 47508 1272 47560
rect 1324 47508 1336 47560
rect 1136 47445 1336 47508
rect 1136 47389 1146 47445
rect 1202 47389 1270 47445
rect 1326 47389 1336 47445
rect 1136 47384 1148 47389
rect 1200 47384 1272 47389
rect 1324 47384 1336 47389
rect 1136 47321 1336 47384
rect 1136 47265 1146 47321
rect 1202 47265 1270 47321
rect 1326 47265 1336 47321
rect 1136 47260 1148 47265
rect 1200 47260 1272 47265
rect 1324 47260 1336 47265
rect 1136 47197 1336 47260
rect 1136 47141 1146 47197
rect 1202 47141 1270 47197
rect 1326 47141 1336 47197
rect 1136 47136 1148 47141
rect 1200 47136 1272 47141
rect 1324 47136 1336 47141
rect 1136 47073 1336 47136
rect 1136 47017 1146 47073
rect 1202 47017 1270 47073
rect 1326 47017 1336 47073
rect 1136 47012 1148 47017
rect 1200 47012 1272 47017
rect 1324 47012 1336 47017
rect 1136 46949 1336 47012
rect 1136 46893 1146 46949
rect 1202 46893 1270 46949
rect 1326 46893 1336 46949
rect 1136 46888 1148 46893
rect 1200 46888 1272 46893
rect 1324 46888 1336 46893
rect 1136 46825 1336 46888
rect 1136 46769 1146 46825
rect 1202 46769 1270 46825
rect 1326 46769 1336 46825
rect 1136 46764 1148 46769
rect 1200 46764 1272 46769
rect 1324 46764 1336 46769
rect 1136 46701 1336 46764
rect 1136 46645 1146 46701
rect 1202 46645 1270 46701
rect 1326 46645 1336 46701
rect 1136 46640 1148 46645
rect 1200 46640 1272 46645
rect 1324 46640 1336 46645
rect 1136 46577 1336 46640
rect 1136 46521 1146 46577
rect 1202 46521 1270 46577
rect 1326 46521 1336 46577
rect 1136 46516 1148 46521
rect 1200 46516 1272 46521
rect 1324 46516 1336 46521
rect 1136 46453 1336 46516
rect 1136 46397 1146 46453
rect 1202 46397 1270 46453
rect 1326 46397 1336 46453
rect 1136 46392 1148 46397
rect 1200 46392 1272 46397
rect 1324 46392 1336 46397
rect 1136 46329 1336 46392
rect 1136 46273 1146 46329
rect 1202 46273 1270 46329
rect 1326 46273 1336 46329
rect 1136 46268 1148 46273
rect 1200 46268 1272 46273
rect 1324 46268 1336 46273
rect 1136 46205 1336 46268
rect 1136 46149 1146 46205
rect 1202 46149 1270 46205
rect 1326 46149 1336 46205
rect 1136 46144 1148 46149
rect 1200 46144 1272 46149
rect 1324 46144 1336 46149
rect 1136 46072 1336 46144
rect 1136 46020 1148 46072
rect 1200 46020 1272 46072
rect 1324 46020 1336 46072
rect 1136 45948 1336 46020
rect 1136 45896 1148 45948
rect 1200 45896 1272 45948
rect 1324 45896 1336 45948
rect 1136 45824 1336 45896
rect 1136 45772 1148 45824
rect 1200 45772 1272 45824
rect 1324 45772 1336 45824
rect 1136 45700 1336 45772
rect 1136 45648 1148 45700
rect 1200 45648 1272 45700
rect 1324 45648 1336 45700
rect 1136 45576 1336 45648
rect 1136 45524 1148 45576
rect 1200 45524 1272 45576
rect 1324 45524 1336 45576
rect 1136 45452 1336 45524
rect 1136 45400 1148 45452
rect 1200 45400 1272 45452
rect 1324 45400 1336 45452
rect 1136 45328 1336 45400
rect 1136 45276 1148 45328
rect 1200 45276 1272 45328
rect 1324 45276 1336 45328
rect 1136 44480 1336 45276
rect 1136 44428 1148 44480
rect 1200 44428 1272 44480
rect 1324 44428 1336 44480
rect 1136 44356 1336 44428
rect 1136 44304 1148 44356
rect 1200 44304 1272 44356
rect 1324 44304 1336 44356
rect 1136 44245 1336 44304
rect 1136 44189 1146 44245
rect 1202 44189 1270 44245
rect 1326 44189 1336 44245
rect 1136 44180 1148 44189
rect 1200 44180 1272 44189
rect 1324 44180 1336 44189
rect 1136 44121 1336 44180
rect 1136 44065 1146 44121
rect 1202 44065 1270 44121
rect 1326 44065 1336 44121
rect 1136 44056 1148 44065
rect 1200 44056 1272 44065
rect 1324 44056 1336 44065
rect 1136 43997 1336 44056
rect 1136 43941 1146 43997
rect 1202 43941 1270 43997
rect 1326 43941 1336 43997
rect 1136 43932 1148 43941
rect 1200 43932 1272 43941
rect 1324 43932 1336 43941
rect 1136 43873 1336 43932
rect 1136 43817 1146 43873
rect 1202 43817 1270 43873
rect 1326 43817 1336 43873
rect 1136 43808 1148 43817
rect 1200 43808 1272 43817
rect 1324 43808 1336 43817
rect 1136 43749 1336 43808
rect 1136 43693 1146 43749
rect 1202 43693 1270 43749
rect 1326 43693 1336 43749
rect 1136 43684 1148 43693
rect 1200 43684 1272 43693
rect 1324 43684 1336 43693
rect 1136 43625 1336 43684
rect 1136 43569 1146 43625
rect 1202 43569 1270 43625
rect 1326 43569 1336 43625
rect 1136 43560 1148 43569
rect 1200 43560 1272 43569
rect 1324 43560 1336 43569
rect 1136 43501 1336 43560
rect 1136 43445 1146 43501
rect 1202 43445 1270 43501
rect 1326 43445 1336 43501
rect 1136 43436 1148 43445
rect 1200 43436 1272 43445
rect 1324 43436 1336 43445
rect 1136 43377 1336 43436
rect 1136 43321 1146 43377
rect 1202 43321 1270 43377
rect 1326 43321 1336 43377
rect 1136 43312 1148 43321
rect 1200 43312 1272 43321
rect 1324 43312 1336 43321
rect 1136 43253 1336 43312
rect 1136 43197 1146 43253
rect 1202 43197 1270 43253
rect 1326 43197 1336 43253
rect 1136 43188 1148 43197
rect 1200 43188 1272 43197
rect 1324 43188 1336 43197
rect 1136 43129 1336 43188
rect 1136 43073 1146 43129
rect 1202 43073 1270 43129
rect 1326 43073 1336 43129
rect 1136 43064 1148 43073
rect 1200 43064 1272 43073
rect 1324 43064 1336 43073
rect 1136 43005 1336 43064
rect 1136 42949 1146 43005
rect 1202 42949 1270 43005
rect 1326 42949 1336 43005
rect 1136 42940 1148 42949
rect 1200 42940 1272 42949
rect 1324 42940 1336 42949
rect 1136 42868 1336 42940
rect 1136 42816 1148 42868
rect 1200 42816 1272 42868
rect 1324 42816 1336 42868
rect 1136 42744 1336 42816
rect 1136 42692 1148 42744
rect 1200 42692 1272 42744
rect 1324 42692 1336 42744
rect 1136 42645 1336 42692
rect 1136 42589 1146 42645
rect 1202 42589 1270 42645
rect 1326 42589 1336 42645
rect 1136 42568 1148 42589
rect 1200 42568 1272 42589
rect 1324 42568 1336 42589
rect 1136 42521 1336 42568
rect 1136 42465 1146 42521
rect 1202 42465 1270 42521
rect 1326 42465 1336 42521
rect 1136 42444 1148 42465
rect 1200 42444 1272 42465
rect 1324 42444 1336 42465
rect 1136 42397 1336 42444
rect 1136 42341 1146 42397
rect 1202 42341 1270 42397
rect 1326 42341 1336 42397
rect 1136 42320 1148 42341
rect 1200 42320 1272 42341
rect 1324 42320 1336 42341
rect 1136 42273 1336 42320
rect 1136 42217 1146 42273
rect 1202 42217 1270 42273
rect 1326 42217 1336 42273
rect 1136 42196 1148 42217
rect 1200 42196 1272 42217
rect 1324 42196 1336 42217
rect 1136 42149 1336 42196
rect 1136 42093 1146 42149
rect 1202 42093 1270 42149
rect 1326 42093 1336 42149
rect 1136 42072 1148 42093
rect 1200 42072 1272 42093
rect 1324 42072 1336 42093
rect 1136 42025 1336 42072
rect 1136 41969 1146 42025
rect 1202 41969 1270 42025
rect 1326 41969 1336 42025
rect 1136 41948 1148 41969
rect 1200 41948 1272 41969
rect 1324 41948 1336 41969
rect 1136 41901 1336 41948
rect 1136 41845 1146 41901
rect 1202 41845 1270 41901
rect 1326 41845 1336 41901
rect 1136 41824 1148 41845
rect 1200 41824 1272 41845
rect 1324 41824 1336 41845
rect 1136 41777 1336 41824
rect 1136 41721 1146 41777
rect 1202 41721 1270 41777
rect 1326 41721 1336 41777
rect 1136 41700 1148 41721
rect 1200 41700 1272 41721
rect 1324 41700 1336 41721
rect 1136 41653 1336 41700
rect 1136 41597 1146 41653
rect 1202 41597 1270 41653
rect 1326 41597 1336 41653
rect 1136 41576 1148 41597
rect 1200 41576 1272 41597
rect 1324 41576 1336 41597
rect 1136 41529 1336 41576
rect 1136 41473 1146 41529
rect 1202 41473 1270 41529
rect 1326 41473 1336 41529
rect 1136 41452 1148 41473
rect 1200 41452 1272 41473
rect 1324 41452 1336 41473
rect 1136 41405 1336 41452
rect 1136 41349 1146 41405
rect 1202 41349 1270 41405
rect 1326 41349 1336 41405
rect 1136 41328 1148 41349
rect 1200 41328 1272 41349
rect 1324 41328 1336 41349
rect 1136 41045 1336 41328
rect 1136 40989 1146 41045
rect 1202 40989 1270 41045
rect 1326 40989 1336 41045
rect 1136 40921 1336 40989
rect 1136 40865 1146 40921
rect 1202 40865 1270 40921
rect 1326 40865 1336 40921
rect 1136 40797 1336 40865
rect 1136 40741 1146 40797
rect 1202 40741 1270 40797
rect 1326 40741 1336 40797
rect 1136 40673 1336 40741
rect 1136 40617 1146 40673
rect 1202 40617 1270 40673
rect 1326 40617 1336 40673
rect 1136 40549 1336 40617
rect 1136 40493 1146 40549
rect 1202 40493 1270 40549
rect 1326 40493 1336 40549
rect 1136 40480 1148 40493
rect 1200 40480 1272 40493
rect 1324 40480 1336 40493
rect 1136 40425 1336 40480
rect 1136 40369 1146 40425
rect 1202 40369 1270 40425
rect 1326 40369 1336 40425
rect 1136 40356 1148 40369
rect 1200 40356 1272 40369
rect 1324 40356 1336 40369
rect 1136 40301 1336 40356
rect 1136 40245 1146 40301
rect 1202 40245 1270 40301
rect 1326 40245 1336 40301
rect 1136 40232 1148 40245
rect 1200 40232 1272 40245
rect 1324 40232 1336 40245
rect 1136 40177 1336 40232
rect 1136 40121 1146 40177
rect 1202 40121 1270 40177
rect 1326 40121 1336 40177
rect 1136 40108 1148 40121
rect 1200 40108 1272 40121
rect 1324 40108 1336 40121
rect 1136 40053 1336 40108
rect 1136 39997 1146 40053
rect 1202 39997 1270 40053
rect 1326 39997 1336 40053
rect 1136 39984 1148 39997
rect 1200 39984 1272 39997
rect 1324 39984 1336 39997
rect 1136 39929 1336 39984
rect 1136 39873 1146 39929
rect 1202 39873 1270 39929
rect 1326 39873 1336 39929
rect 1136 39860 1148 39873
rect 1200 39860 1272 39873
rect 1324 39860 1336 39873
rect 1136 39805 1336 39860
rect 1136 39749 1146 39805
rect 1202 39749 1270 39805
rect 1326 39749 1336 39805
rect 1136 39736 1148 39749
rect 1200 39736 1272 39749
rect 1324 39736 1336 39749
rect 1136 39664 1336 39736
rect 1136 39612 1148 39664
rect 1200 39612 1272 39664
rect 1324 39612 1336 39664
rect 1136 39540 1336 39612
rect 1136 39488 1148 39540
rect 1200 39488 1272 39540
rect 1324 39488 1336 39540
rect 1136 39416 1336 39488
rect 1136 39364 1148 39416
rect 1200 39364 1272 39416
rect 1324 39364 1336 39416
rect 1136 39292 1336 39364
rect 1136 39240 1148 39292
rect 1200 39240 1272 39292
rect 1324 39240 1336 39292
rect 1136 39168 1336 39240
rect 1136 39116 1148 39168
rect 1200 39116 1272 39168
rect 1324 39116 1336 39168
rect 1136 39044 1336 39116
rect 1136 38992 1148 39044
rect 1200 38992 1272 39044
rect 1324 38992 1336 39044
rect 1136 38920 1336 38992
rect 1136 38868 1148 38920
rect 1200 38868 1272 38920
rect 1324 38868 1336 38920
rect 1136 38796 1336 38868
rect 1136 38744 1148 38796
rect 1200 38744 1272 38796
rect 1324 38744 1336 38796
rect 1136 38672 1336 38744
rect 1136 38620 1148 38672
rect 1200 38620 1272 38672
rect 1324 38620 1336 38672
rect 1136 38548 1336 38620
rect 1136 38496 1148 38548
rect 1200 38496 1272 38548
rect 1324 38496 1336 38548
rect 1136 38424 1336 38496
rect 1136 38372 1148 38424
rect 1200 38372 1272 38424
rect 1324 38372 1336 38424
rect 1136 38300 1336 38372
rect 1136 38248 1148 38300
rect 1200 38248 1272 38300
rect 1324 38248 1336 38300
rect 1136 38176 1336 38248
rect 1136 38124 1148 38176
rect 1200 38124 1272 38176
rect 1324 38124 1336 38176
rect 260 37172 444 37224
rect 496 37172 552 37224
rect 604 37172 660 37224
rect 712 37172 768 37224
rect 260 37116 768 37172
rect 260 37064 444 37116
rect 496 37064 552 37116
rect 604 37064 660 37116
rect 712 37064 768 37116
rect 260 37008 768 37064
rect 260 36956 444 37008
rect 496 36956 552 37008
rect 604 36956 660 37008
rect 712 36956 768 37008
rect 260 36900 768 36956
rect 260 36848 444 36900
rect 496 36848 552 36900
rect 604 36848 660 36900
rect 712 36848 768 36900
rect 260 36792 768 36848
rect 260 36740 444 36792
rect 496 36740 552 36792
rect 604 36740 660 36792
rect 712 36740 768 36792
rect 260 36251 768 36740
rect 1136 38052 1336 38124
rect 1136 38000 1148 38052
rect 1200 38000 1272 38052
rect 1324 38000 1336 38052
rect 1136 37928 1336 38000
rect 1136 37876 1148 37928
rect 1200 37876 1272 37928
rect 1324 37876 1336 37928
rect 1136 37804 1336 37876
rect 1136 37752 1148 37804
rect 1200 37752 1272 37804
rect 1324 37752 1336 37804
rect 1136 37680 1336 37752
rect 1136 37628 1148 37680
rect 1200 37628 1272 37680
rect 1324 37628 1336 37680
rect 1136 37556 1336 37628
rect 1136 37504 1148 37556
rect 1200 37504 1272 37556
rect 1324 37504 1336 37556
rect 1136 37432 1336 37504
rect 1136 37380 1148 37432
rect 1200 37380 1272 37432
rect 1324 37380 1336 37432
rect 1136 36596 1336 37380
rect 260 36195 300 36251
rect 356 36195 424 36251
rect 480 36195 548 36251
rect 604 36195 672 36251
rect 728 36195 768 36251
rect 260 36127 768 36195
rect 260 36071 300 36127
rect 356 36071 424 36127
rect 480 36071 548 36127
rect 604 36071 672 36127
rect 728 36071 768 36127
rect 260 36003 768 36071
rect 260 35947 300 36003
rect 356 35947 424 36003
rect 480 35947 548 36003
rect 604 35947 672 36003
rect 728 35947 768 36003
rect 260 35879 768 35947
rect 260 35823 300 35879
rect 356 35823 424 35879
rect 480 35823 548 35879
rect 604 35823 672 35879
rect 728 35823 768 35879
rect 260 35755 768 35823
rect 260 35699 300 35755
rect 356 35699 424 35755
rect 480 35699 548 35755
rect 604 35699 672 35755
rect 728 35699 768 35755
rect 260 35631 768 35699
rect 260 35575 300 35631
rect 356 35575 424 35631
rect 480 35575 548 35631
rect 604 35575 672 35631
rect 728 35575 768 35631
rect 260 35507 768 35575
rect 260 35451 300 35507
rect 356 35451 424 35507
rect 480 35451 548 35507
rect 604 35451 672 35507
rect 728 35451 768 35507
rect 260 35383 768 35451
rect 260 35327 300 35383
rect 356 35327 424 35383
rect 480 35327 548 35383
rect 604 35327 672 35383
rect 728 35327 768 35383
rect 260 35259 768 35327
rect 260 35203 300 35259
rect 356 35203 424 35259
rect 480 35203 548 35259
rect 604 35203 672 35259
rect 728 35203 768 35259
rect 260 35135 768 35203
rect 260 35079 300 35135
rect 356 35079 424 35135
rect 480 35079 548 35135
rect 604 35079 672 35135
rect 728 35079 768 35135
rect 260 35011 768 35079
rect 260 34955 300 35011
rect 356 34955 424 35011
rect 480 34955 548 35011
rect 604 34955 672 35011
rect 728 34955 768 35011
rect 260 34887 768 34955
rect 260 34831 300 34887
rect 356 34831 424 34887
rect 480 34831 548 34887
rect 604 34831 672 34887
rect 728 34831 768 34887
rect 260 34763 768 34831
rect 260 34707 300 34763
rect 356 34707 424 34763
rect 480 34707 548 34763
rect 604 34707 672 34763
rect 728 34707 768 34763
rect 260 34639 768 34707
rect 260 34583 300 34639
rect 356 34583 424 34639
rect 480 34583 548 34639
rect 604 34583 672 34639
rect 728 34583 768 34639
rect 260 34515 768 34583
rect 260 34459 300 34515
rect 356 34459 424 34515
rect 480 34459 548 34515
rect 604 34459 672 34515
rect 728 34459 768 34515
rect 260 34391 768 34459
rect 260 34335 300 34391
rect 356 34335 424 34391
rect 480 34335 548 34391
rect 604 34335 672 34391
rect 728 34335 768 34391
rect 260 34267 768 34335
rect 260 34211 300 34267
rect 356 34211 424 34267
rect 480 34211 548 34267
rect 604 34211 672 34267
rect 728 34211 768 34267
rect 260 34143 768 34211
rect 260 34087 300 34143
rect 356 34087 424 34143
rect 480 34087 548 34143
rect 604 34087 672 34143
rect 728 34087 768 34143
rect 260 34019 768 34087
rect 260 33963 300 34019
rect 356 33963 424 34019
rect 480 33963 548 34019
rect 604 33963 672 34019
rect 728 33963 768 34019
rect 260 33895 768 33963
rect 260 33839 300 33895
rect 356 33839 424 33895
rect 480 33839 548 33895
rect 604 33839 672 33895
rect 728 33839 768 33895
rect 260 33771 768 33839
rect 260 33715 300 33771
rect 356 33715 424 33771
rect 480 33715 548 33771
rect 604 33715 672 33771
rect 728 33715 768 33771
rect 260 33647 768 33715
rect 260 33591 300 33647
rect 356 33591 424 33647
rect 480 33591 548 33647
rect 604 33591 672 33647
rect 728 33591 768 33647
rect 260 33523 768 33591
rect 260 33467 300 33523
rect 356 33467 424 33523
rect 480 33467 548 33523
rect 604 33467 672 33523
rect 728 33467 768 33523
rect 260 33399 768 33467
rect 966 36584 1336 36596
rect 966 36532 978 36584
rect 1030 36532 1102 36584
rect 1154 36532 1226 36584
rect 1278 36532 1336 36584
rect 966 36460 1336 36532
rect 966 36408 978 36460
rect 1030 36408 1102 36460
rect 1154 36408 1226 36460
rect 1278 36408 1336 36460
rect 966 36336 1336 36408
rect 966 36284 978 36336
rect 1030 36284 1102 36336
rect 1154 36284 1226 36336
rect 1278 36284 1336 36336
rect 966 36212 1336 36284
rect 966 36160 978 36212
rect 1030 36160 1102 36212
rect 1154 36160 1226 36212
rect 1278 36160 1336 36212
rect 966 36088 1336 36160
rect 966 36036 978 36088
rect 1030 36036 1102 36088
rect 1154 36036 1226 36088
rect 1278 36036 1336 36088
rect 966 35964 1336 36036
rect 966 35912 978 35964
rect 1030 35912 1102 35964
rect 1154 35912 1226 35964
rect 1278 35912 1336 35964
rect 966 35840 1336 35912
rect 966 35788 978 35840
rect 1030 35788 1102 35840
rect 1154 35788 1226 35840
rect 1278 35788 1336 35840
rect 966 35716 1336 35788
rect 966 35664 978 35716
rect 1030 35664 1102 35716
rect 1154 35664 1226 35716
rect 1278 35664 1336 35716
rect 966 35592 1336 35664
rect 966 35540 978 35592
rect 1030 35540 1102 35592
rect 1154 35540 1226 35592
rect 1278 35540 1336 35592
rect 966 35468 1336 35540
rect 966 35416 978 35468
rect 1030 35416 1102 35468
rect 1154 35416 1226 35468
rect 1278 35416 1336 35468
rect 966 35344 1336 35416
rect 966 35292 978 35344
rect 1030 35292 1102 35344
rect 1154 35292 1226 35344
rect 1278 35292 1336 35344
rect 966 35220 1336 35292
rect 966 35168 978 35220
rect 1030 35168 1102 35220
rect 1154 35168 1226 35220
rect 1278 35168 1336 35220
rect 966 35096 1336 35168
rect 966 35044 978 35096
rect 1030 35044 1102 35096
rect 1154 35044 1226 35096
rect 1278 35044 1336 35096
rect 966 34972 1336 35044
rect 966 34920 978 34972
rect 1030 34920 1102 34972
rect 1154 34920 1226 34972
rect 1278 34920 1336 34972
rect 966 34848 1336 34920
rect 966 34796 978 34848
rect 1030 34796 1102 34848
rect 1154 34796 1226 34848
rect 1278 34796 1336 34848
rect 966 34724 1336 34796
rect 966 34672 978 34724
rect 1030 34672 1102 34724
rect 1154 34672 1226 34724
rect 1278 34672 1336 34724
rect 966 34600 1336 34672
rect 966 34548 978 34600
rect 1030 34548 1102 34600
rect 1154 34548 1226 34600
rect 1278 34548 1336 34600
rect 966 34476 1336 34548
rect 966 34424 978 34476
rect 1030 34424 1102 34476
rect 1154 34424 1226 34476
rect 1278 34424 1336 34476
rect 966 34352 1336 34424
rect 966 34300 978 34352
rect 1030 34300 1102 34352
rect 1154 34300 1226 34352
rect 1278 34300 1336 34352
rect 966 34228 1336 34300
rect 966 34176 978 34228
rect 1030 34176 1102 34228
rect 1154 34176 1226 34228
rect 1278 34176 1336 34228
rect 966 34104 1336 34176
rect 966 34052 978 34104
rect 1030 34052 1102 34104
rect 1154 34052 1226 34104
rect 1278 34052 1336 34104
rect 966 33980 1336 34052
rect 966 33928 978 33980
rect 1030 33928 1102 33980
rect 1154 33928 1226 33980
rect 1278 33928 1336 33980
rect 966 33856 1336 33928
rect 966 33804 978 33856
rect 1030 33804 1102 33856
rect 1154 33804 1226 33856
rect 1278 33804 1336 33856
rect 966 33732 1336 33804
rect 966 33680 978 33732
rect 1030 33680 1102 33732
rect 1154 33680 1226 33732
rect 1278 33680 1336 33732
rect 966 33608 1336 33680
rect 966 33556 978 33608
rect 1030 33556 1102 33608
rect 1154 33556 1226 33608
rect 1278 33556 1336 33608
rect 966 33484 1336 33556
rect 966 33432 978 33484
rect 1030 33432 1102 33484
rect 1154 33432 1226 33484
rect 1278 33432 1336 33484
rect 966 33420 1336 33432
rect 260 33343 300 33399
rect 356 33343 424 33399
rect 480 33343 548 33399
rect 604 33343 672 33399
rect 728 33343 768 33399
rect 260 33276 768 33343
rect 260 33224 444 33276
rect 496 33224 552 33276
rect 604 33224 660 33276
rect 712 33224 768 33276
rect 260 33168 768 33224
rect 260 33116 444 33168
rect 496 33116 552 33168
rect 604 33116 660 33168
rect 712 33116 768 33168
rect 260 33060 768 33116
rect 1136 33061 1336 33420
rect 260 33008 444 33060
rect 496 33008 552 33060
rect 604 33008 660 33060
rect 712 33008 768 33060
rect 260 32952 768 33008
rect 260 32900 444 32952
rect 496 32900 552 32952
rect 604 32900 660 32952
rect 712 32900 768 32952
rect 260 32844 768 32900
rect 260 32792 444 32844
rect 496 32792 552 32844
rect 604 32792 660 32844
rect 712 32792 768 32844
rect 260 29328 768 32792
rect 858 33051 1336 33061
rect 858 32995 868 33051
rect 924 32995 992 33051
rect 1048 32995 1116 33051
rect 1172 32995 1240 33051
rect 1296 32995 1336 33051
rect 858 32927 1336 32995
rect 858 32871 868 32927
rect 924 32871 992 32927
rect 1048 32871 1116 32927
rect 1172 32871 1240 32927
rect 1296 32871 1336 32927
rect 858 32803 1336 32871
rect 858 32747 868 32803
rect 924 32747 992 32803
rect 1048 32747 1116 32803
rect 1172 32747 1240 32803
rect 1296 32747 1336 32803
rect 858 32679 1336 32747
rect 858 32623 868 32679
rect 924 32636 992 32679
rect 1048 32636 1116 32679
rect 1172 32636 1240 32679
rect 924 32623 978 32636
rect 1048 32623 1102 32636
rect 1172 32623 1226 32636
rect 1296 32623 1336 32679
rect 858 32584 978 32623
rect 1030 32584 1102 32623
rect 1154 32584 1226 32623
rect 1278 32584 1336 32623
rect 858 32555 1336 32584
rect 858 32499 868 32555
rect 924 32512 992 32555
rect 1048 32512 1116 32555
rect 1172 32512 1240 32555
rect 924 32499 978 32512
rect 1048 32499 1102 32512
rect 1172 32499 1226 32512
rect 1296 32499 1336 32555
rect 858 32460 978 32499
rect 1030 32460 1102 32499
rect 1154 32460 1226 32499
rect 1278 32460 1336 32499
rect 858 32431 1336 32460
rect 858 32375 868 32431
rect 924 32388 992 32431
rect 1048 32388 1116 32431
rect 1172 32388 1240 32431
rect 924 32375 978 32388
rect 1048 32375 1102 32388
rect 1172 32375 1226 32388
rect 1296 32375 1336 32431
rect 858 32336 978 32375
rect 1030 32336 1102 32375
rect 1154 32336 1226 32375
rect 1278 32336 1336 32375
rect 858 32307 1336 32336
rect 858 32251 868 32307
rect 924 32264 992 32307
rect 1048 32264 1116 32307
rect 1172 32264 1240 32307
rect 924 32251 978 32264
rect 1048 32251 1102 32264
rect 1172 32251 1226 32264
rect 1296 32251 1336 32307
rect 858 32212 978 32251
rect 1030 32212 1102 32251
rect 1154 32212 1226 32251
rect 1278 32212 1336 32251
rect 858 32183 1336 32212
rect 858 32127 868 32183
rect 924 32140 992 32183
rect 1048 32140 1116 32183
rect 1172 32140 1240 32183
rect 924 32127 978 32140
rect 1048 32127 1102 32140
rect 1172 32127 1226 32140
rect 1296 32127 1336 32183
rect 858 32088 978 32127
rect 1030 32088 1102 32127
rect 1154 32088 1226 32127
rect 1278 32088 1336 32127
rect 858 32059 1336 32088
rect 858 32003 868 32059
rect 924 32016 992 32059
rect 1048 32016 1116 32059
rect 1172 32016 1240 32059
rect 924 32003 978 32016
rect 1048 32003 1102 32016
rect 1172 32003 1226 32016
rect 1296 32003 1336 32059
rect 858 31964 978 32003
rect 1030 31964 1102 32003
rect 1154 31964 1226 32003
rect 1278 31964 1336 32003
rect 858 31935 1336 31964
rect 858 31879 868 31935
rect 924 31892 992 31935
rect 1048 31892 1116 31935
rect 1172 31892 1240 31935
rect 924 31879 978 31892
rect 1048 31879 1102 31892
rect 1172 31879 1226 31892
rect 1296 31879 1336 31935
rect 858 31840 978 31879
rect 1030 31840 1102 31879
rect 1154 31840 1226 31879
rect 1278 31840 1336 31879
rect 858 31811 1336 31840
rect 858 31755 868 31811
rect 924 31768 992 31811
rect 1048 31768 1116 31811
rect 1172 31768 1240 31811
rect 924 31755 978 31768
rect 1048 31755 1102 31768
rect 1172 31755 1226 31768
rect 1296 31755 1336 31811
rect 858 31716 978 31755
rect 1030 31716 1102 31755
rect 1154 31716 1226 31755
rect 1278 31716 1336 31755
rect 858 31687 1336 31716
rect 858 31631 868 31687
rect 924 31644 992 31687
rect 1048 31644 1116 31687
rect 1172 31644 1240 31687
rect 924 31631 978 31644
rect 1048 31631 1102 31644
rect 1172 31631 1226 31644
rect 1296 31631 1336 31687
rect 858 31592 978 31631
rect 1030 31592 1102 31631
rect 1154 31592 1226 31631
rect 1278 31592 1336 31631
rect 858 31563 1336 31592
rect 858 31507 868 31563
rect 924 31520 992 31563
rect 1048 31520 1116 31563
rect 1172 31520 1240 31563
rect 924 31507 978 31520
rect 1048 31507 1102 31520
rect 1172 31507 1226 31520
rect 1296 31507 1336 31563
rect 858 31468 978 31507
rect 1030 31468 1102 31507
rect 1154 31468 1226 31507
rect 1278 31468 1336 31507
rect 858 31439 1336 31468
rect 858 31383 868 31439
rect 924 31396 992 31439
rect 1048 31396 1116 31439
rect 1172 31396 1240 31439
rect 924 31383 978 31396
rect 1048 31383 1102 31396
rect 1172 31383 1226 31396
rect 1296 31383 1336 31439
rect 858 31344 978 31383
rect 1030 31344 1102 31383
rect 1154 31344 1226 31383
rect 1278 31344 1336 31383
rect 858 31315 1336 31344
rect 858 31259 868 31315
rect 924 31272 992 31315
rect 1048 31272 1116 31315
rect 1172 31272 1240 31315
rect 924 31259 978 31272
rect 1048 31259 1102 31272
rect 1172 31259 1226 31272
rect 1296 31259 1336 31315
rect 858 31220 978 31259
rect 1030 31220 1102 31259
rect 1154 31220 1226 31259
rect 1278 31220 1336 31259
rect 858 31191 1336 31220
rect 858 31135 868 31191
rect 924 31148 992 31191
rect 1048 31148 1116 31191
rect 1172 31148 1240 31191
rect 924 31135 978 31148
rect 1048 31135 1102 31148
rect 1172 31135 1226 31148
rect 1296 31135 1336 31191
rect 858 31096 978 31135
rect 1030 31096 1102 31135
rect 1154 31096 1226 31135
rect 1278 31096 1336 31135
rect 858 31067 1336 31096
rect 858 31011 868 31067
rect 924 31024 992 31067
rect 1048 31024 1116 31067
rect 1172 31024 1240 31067
rect 924 31011 978 31024
rect 1048 31011 1102 31024
rect 1172 31011 1226 31024
rect 1296 31011 1336 31067
rect 858 30972 978 31011
rect 1030 30972 1102 31011
rect 1154 30972 1226 31011
rect 1278 30972 1336 31011
rect 858 30943 1336 30972
rect 858 30887 868 30943
rect 924 30900 992 30943
rect 1048 30900 1116 30943
rect 1172 30900 1240 30943
rect 924 30887 978 30900
rect 1048 30887 1102 30900
rect 1172 30887 1226 30900
rect 1296 30887 1336 30943
rect 858 30848 978 30887
rect 1030 30848 1102 30887
rect 1154 30848 1226 30887
rect 1278 30848 1336 30887
rect 858 30819 1336 30848
rect 858 30763 868 30819
rect 924 30776 992 30819
rect 1048 30776 1116 30819
rect 1172 30776 1240 30819
rect 924 30763 978 30776
rect 1048 30763 1102 30776
rect 1172 30763 1226 30776
rect 1296 30763 1336 30819
rect 858 30724 978 30763
rect 1030 30724 1102 30763
rect 1154 30724 1226 30763
rect 1278 30724 1336 30763
rect 858 30695 1336 30724
rect 858 30639 868 30695
rect 924 30652 992 30695
rect 1048 30652 1116 30695
rect 1172 30652 1240 30695
rect 924 30639 978 30652
rect 1048 30639 1102 30652
rect 1172 30639 1226 30652
rect 1296 30639 1336 30695
rect 858 30600 978 30639
rect 1030 30600 1102 30639
rect 1154 30600 1226 30639
rect 1278 30600 1336 30639
rect 858 30571 1336 30600
rect 858 30515 868 30571
rect 924 30528 992 30571
rect 1048 30528 1116 30571
rect 1172 30528 1240 30571
rect 924 30515 978 30528
rect 1048 30515 1102 30528
rect 1172 30515 1226 30528
rect 1296 30515 1336 30571
rect 858 30476 978 30515
rect 1030 30476 1102 30515
rect 1154 30476 1226 30515
rect 1278 30476 1336 30515
rect 858 30447 1336 30476
rect 858 30391 868 30447
rect 924 30404 992 30447
rect 1048 30404 1116 30447
rect 1172 30404 1240 30447
rect 924 30391 978 30404
rect 1048 30391 1102 30404
rect 1172 30391 1226 30404
rect 1296 30391 1336 30447
rect 858 30352 978 30391
rect 1030 30352 1102 30391
rect 1154 30352 1226 30391
rect 1278 30352 1336 30391
rect 858 30323 1336 30352
rect 858 30267 868 30323
rect 924 30280 992 30323
rect 1048 30280 1116 30323
rect 1172 30280 1240 30323
rect 924 30267 978 30280
rect 1048 30267 1102 30280
rect 1172 30267 1226 30280
rect 1296 30267 1336 30323
rect 858 30228 978 30267
rect 1030 30228 1102 30267
rect 1154 30228 1226 30267
rect 1278 30228 1336 30267
rect 858 30199 1336 30228
rect 858 30143 868 30199
rect 924 30156 992 30199
rect 1048 30156 1116 30199
rect 1172 30156 1240 30199
rect 924 30143 978 30156
rect 1048 30143 1102 30156
rect 1172 30143 1226 30156
rect 1296 30143 1336 30199
rect 858 30133 978 30143
rect 966 30104 978 30133
rect 1030 30104 1102 30143
rect 1154 30104 1226 30143
rect 1278 30104 1336 30143
rect 966 30032 1336 30104
rect 966 29980 978 30032
rect 1030 29980 1102 30032
rect 1154 29980 1226 30032
rect 1278 29980 1336 30032
rect 966 29908 1336 29980
rect 966 29856 978 29908
rect 1030 29856 1102 29908
rect 1154 29856 1226 29908
rect 1278 29856 1336 29908
rect 966 29855 1336 29856
rect 260 29276 444 29328
rect 496 29276 552 29328
rect 604 29276 660 29328
rect 712 29276 768 29328
rect 260 29220 768 29276
rect 260 29168 444 29220
rect 496 29168 552 29220
rect 604 29168 660 29220
rect 712 29168 768 29220
rect 260 29112 768 29168
rect 260 29060 444 29112
rect 496 29060 552 29112
rect 604 29060 660 29112
rect 712 29060 768 29112
rect 260 29004 768 29060
rect 260 28952 444 29004
rect 496 28952 552 29004
rect 604 28952 660 29004
rect 712 28952 768 29004
rect 260 28896 768 28952
rect 260 28844 444 28896
rect 496 28844 552 28896
rect 604 28844 660 28896
rect 712 28844 768 28896
rect 260 28245 768 28844
rect 858 29845 1336 29855
rect 858 29789 868 29845
rect 924 29789 992 29845
rect 1048 29789 1116 29845
rect 1172 29789 1240 29845
rect 1296 29789 1336 29845
rect 858 29784 1336 29789
rect 858 29732 978 29784
rect 1030 29732 1102 29784
rect 1154 29732 1226 29784
rect 1278 29732 1336 29784
rect 858 29721 1336 29732
rect 858 29665 868 29721
rect 924 29665 992 29721
rect 1048 29665 1116 29721
rect 1172 29665 1240 29721
rect 1296 29665 1336 29721
rect 858 29660 1336 29665
rect 858 29608 978 29660
rect 1030 29608 1102 29660
rect 1154 29608 1226 29660
rect 1278 29608 1336 29660
rect 858 29597 1336 29608
rect 858 29541 868 29597
rect 924 29541 992 29597
rect 1048 29541 1116 29597
rect 1172 29541 1240 29597
rect 1296 29541 1336 29597
rect 858 29536 1336 29541
rect 858 29484 978 29536
rect 1030 29484 1102 29536
rect 1154 29484 1226 29536
rect 1278 29484 1336 29536
rect 858 29473 1336 29484
rect 858 29417 868 29473
rect 924 29417 992 29473
rect 1048 29417 1116 29473
rect 1172 29417 1240 29473
rect 1296 29417 1336 29473
rect 858 29349 1336 29417
rect 858 29293 868 29349
rect 924 29293 992 29349
rect 1048 29293 1116 29349
rect 1172 29293 1240 29349
rect 1296 29293 1336 29349
rect 858 29225 1336 29293
rect 858 29169 868 29225
rect 924 29169 992 29225
rect 1048 29169 1116 29225
rect 1172 29169 1240 29225
rect 1296 29169 1336 29225
rect 858 29101 1336 29169
rect 858 29045 868 29101
rect 924 29045 992 29101
rect 1048 29045 1116 29101
rect 1172 29045 1240 29101
rect 1296 29045 1336 29101
rect 858 28977 1336 29045
rect 858 28921 868 28977
rect 924 28921 992 28977
rect 1048 28921 1116 28977
rect 1172 28921 1240 28977
rect 1296 28921 1336 28977
rect 858 28853 1336 28921
rect 858 28797 868 28853
rect 924 28797 992 28853
rect 1048 28797 1116 28853
rect 1172 28797 1240 28853
rect 1296 28797 1336 28853
rect 858 28729 1336 28797
rect 858 28673 868 28729
rect 924 28688 992 28729
rect 1048 28688 1116 28729
rect 1172 28688 1240 28729
rect 924 28673 978 28688
rect 1048 28673 1102 28688
rect 1172 28673 1226 28688
rect 1296 28673 1336 28729
rect 858 28636 978 28673
rect 1030 28636 1102 28673
rect 1154 28636 1226 28673
rect 1278 28636 1336 28673
rect 858 28605 1336 28636
rect 858 28549 868 28605
rect 924 28564 992 28605
rect 1048 28564 1116 28605
rect 1172 28564 1240 28605
rect 924 28549 978 28564
rect 1048 28549 1102 28564
rect 1172 28549 1226 28564
rect 1296 28549 1336 28605
rect 858 28539 978 28549
rect 260 28189 300 28245
rect 356 28189 424 28245
rect 480 28189 548 28245
rect 604 28189 672 28245
rect 728 28189 768 28245
rect 260 28121 768 28189
rect 260 28065 300 28121
rect 356 28065 424 28121
rect 480 28065 548 28121
rect 604 28065 672 28121
rect 728 28065 768 28121
rect 260 27997 768 28065
rect 260 27941 300 27997
rect 356 27941 424 27997
rect 480 27941 548 27997
rect 604 27941 672 27997
rect 728 27941 768 27997
rect 260 27873 768 27941
rect 260 27817 300 27873
rect 356 27817 424 27873
rect 480 27817 548 27873
rect 604 27817 672 27873
rect 728 27817 768 27873
rect 260 27749 768 27817
rect 260 27693 300 27749
rect 356 27693 424 27749
rect 480 27693 548 27749
rect 604 27693 672 27749
rect 728 27693 768 27749
rect 260 27625 768 27693
rect 260 27569 300 27625
rect 356 27569 424 27625
rect 480 27569 548 27625
rect 604 27569 672 27625
rect 728 27569 768 27625
rect 260 27501 768 27569
rect 260 27445 300 27501
rect 356 27445 424 27501
rect 480 27445 548 27501
rect 604 27445 672 27501
rect 728 27445 768 27501
rect 260 27377 768 27445
rect 260 27321 300 27377
rect 356 27321 424 27377
rect 480 27321 548 27377
rect 604 27321 672 27377
rect 728 27321 768 27377
rect 260 27253 768 27321
rect 260 27197 300 27253
rect 356 27197 424 27253
rect 480 27197 548 27253
rect 604 27197 672 27253
rect 728 27197 768 27253
rect 260 27129 768 27197
rect 260 27073 300 27129
rect 356 27073 424 27129
rect 480 27073 548 27129
rect 604 27073 672 27129
rect 728 27073 768 27129
rect 260 27005 768 27073
rect 260 26949 300 27005
rect 356 26949 424 27005
rect 480 26949 548 27005
rect 604 26949 672 27005
rect 728 26949 768 27005
rect 260 25380 768 26949
rect 966 28512 978 28539
rect 1030 28512 1102 28549
rect 1154 28512 1226 28549
rect 1278 28512 1336 28549
rect 966 28440 1336 28512
rect 966 28388 978 28440
rect 1030 28388 1102 28440
rect 1154 28388 1226 28440
rect 1278 28388 1336 28440
rect 966 28316 1336 28388
rect 966 28264 978 28316
rect 1030 28264 1102 28316
rect 1154 28264 1226 28316
rect 1278 28264 1336 28316
rect 966 28192 1336 28264
rect 966 28140 978 28192
rect 1030 28140 1102 28192
rect 1154 28140 1226 28192
rect 1278 28140 1336 28192
rect 966 28068 1336 28140
rect 966 28016 978 28068
rect 1030 28016 1102 28068
rect 1154 28016 1226 28068
rect 1278 28016 1336 28068
rect 966 27944 1336 28016
rect 966 27892 978 27944
rect 1030 27892 1102 27944
rect 1154 27892 1226 27944
rect 1278 27892 1336 27944
rect 966 27820 1336 27892
rect 966 27768 978 27820
rect 1030 27768 1102 27820
rect 1154 27768 1226 27820
rect 1278 27768 1336 27820
rect 966 27696 1336 27768
rect 966 27644 978 27696
rect 1030 27644 1102 27696
rect 1154 27644 1226 27696
rect 1278 27644 1336 27696
rect 966 27572 1336 27644
rect 966 27520 978 27572
rect 1030 27520 1102 27572
rect 1154 27520 1226 27572
rect 1278 27520 1336 27572
rect 966 27448 1336 27520
rect 966 27396 978 27448
rect 1030 27396 1102 27448
rect 1154 27396 1226 27448
rect 1278 27396 1336 27448
rect 966 27324 1336 27396
rect 966 27272 978 27324
rect 1030 27272 1102 27324
rect 1154 27272 1226 27324
rect 1278 27272 1336 27324
rect 966 27200 1336 27272
rect 966 27148 978 27200
rect 1030 27148 1102 27200
rect 1154 27148 1226 27200
rect 1278 27148 1336 27200
rect 966 27076 1336 27148
rect 966 27024 978 27076
rect 1030 27024 1102 27076
rect 1154 27024 1226 27076
rect 1278 27024 1336 27076
rect 966 26952 1336 27024
rect 966 26900 978 26952
rect 1030 26900 1102 26952
rect 1154 26900 1226 26952
rect 1278 26900 1336 26952
rect 966 26828 1336 26900
rect 966 26776 978 26828
rect 1030 26776 1102 26828
rect 1154 26776 1226 26828
rect 1278 26776 1336 26828
rect 966 26704 1336 26776
rect 966 26661 978 26704
rect 260 25328 444 25380
rect 496 25328 552 25380
rect 604 25328 660 25380
rect 712 25328 768 25380
rect 260 25272 768 25328
rect 260 25220 444 25272
rect 496 25220 552 25272
rect 604 25220 660 25272
rect 712 25220 768 25272
rect 260 25164 768 25220
rect 260 25112 444 25164
rect 496 25112 552 25164
rect 604 25112 660 25164
rect 712 25112 768 25164
rect 260 25056 768 25112
rect 260 25004 444 25056
rect 496 25004 552 25056
rect 604 25004 660 25056
rect 712 25004 768 25056
rect 260 24948 768 25004
rect 260 24896 444 24948
rect 496 24896 552 24948
rect 604 24896 660 24948
rect 712 24896 768 24948
rect 260 21469 768 24896
rect 858 26652 978 26661
rect 1030 26652 1102 26704
rect 1154 26652 1226 26704
rect 1278 26652 1336 26704
rect 858 26651 1336 26652
rect 858 26595 868 26651
rect 924 26595 992 26651
rect 1048 26595 1116 26651
rect 1172 26595 1240 26651
rect 1296 26595 1336 26651
rect 858 26580 1336 26595
rect 858 26528 978 26580
rect 1030 26528 1102 26580
rect 1154 26528 1226 26580
rect 1278 26528 1336 26580
rect 858 26527 1336 26528
rect 858 26471 868 26527
rect 924 26471 992 26527
rect 1048 26471 1116 26527
rect 1172 26471 1240 26527
rect 1296 26471 1336 26527
rect 858 26456 1336 26471
rect 858 26404 978 26456
rect 1030 26404 1102 26456
rect 1154 26404 1226 26456
rect 1278 26404 1336 26456
rect 858 26403 1336 26404
rect 858 26347 868 26403
rect 924 26347 992 26403
rect 1048 26347 1116 26403
rect 1172 26347 1240 26403
rect 1296 26347 1336 26403
rect 858 26332 1336 26347
rect 858 26280 978 26332
rect 1030 26280 1102 26332
rect 1154 26280 1226 26332
rect 1278 26280 1336 26332
rect 858 26279 1336 26280
rect 858 26223 868 26279
rect 924 26223 992 26279
rect 1048 26223 1116 26279
rect 1172 26223 1240 26279
rect 1296 26223 1336 26279
rect 858 26208 1336 26223
rect 858 26156 978 26208
rect 1030 26156 1102 26208
rect 1154 26156 1226 26208
rect 1278 26156 1336 26208
rect 858 26155 1336 26156
rect 858 26099 868 26155
rect 924 26099 992 26155
rect 1048 26099 1116 26155
rect 1172 26099 1240 26155
rect 1296 26099 1336 26155
rect 858 26084 1336 26099
rect 858 26032 978 26084
rect 1030 26032 1102 26084
rect 1154 26032 1226 26084
rect 1278 26032 1336 26084
rect 858 26031 1336 26032
rect 858 25975 868 26031
rect 924 25975 992 26031
rect 1048 25975 1116 26031
rect 1172 25975 1240 26031
rect 1296 25975 1336 26031
rect 858 25960 1336 25975
rect 858 25908 978 25960
rect 1030 25908 1102 25960
rect 1154 25908 1226 25960
rect 1278 25908 1336 25960
rect 858 25907 1336 25908
rect 858 25851 868 25907
rect 924 25851 992 25907
rect 1048 25851 1116 25907
rect 1172 25851 1240 25907
rect 1296 25851 1336 25907
rect 858 25836 1336 25851
rect 858 25784 978 25836
rect 1030 25784 1102 25836
rect 1154 25784 1226 25836
rect 1278 25784 1336 25836
rect 858 25783 1336 25784
rect 858 25727 868 25783
rect 924 25727 992 25783
rect 1048 25727 1116 25783
rect 1172 25727 1240 25783
rect 1296 25727 1336 25783
rect 858 25712 1336 25727
rect 858 25660 978 25712
rect 1030 25660 1102 25712
rect 1154 25660 1226 25712
rect 1278 25660 1336 25712
rect 858 25659 1336 25660
rect 858 25603 868 25659
rect 924 25603 992 25659
rect 1048 25603 1116 25659
rect 1172 25603 1240 25659
rect 1296 25603 1336 25659
rect 858 25588 1336 25603
rect 858 25536 978 25588
rect 1030 25536 1102 25588
rect 1154 25536 1226 25588
rect 1278 25536 1336 25588
rect 858 25535 1336 25536
rect 858 25479 868 25535
rect 924 25479 992 25535
rect 1048 25479 1116 25535
rect 1172 25479 1240 25535
rect 1296 25479 1336 25535
rect 858 25411 1336 25479
rect 858 25355 868 25411
rect 924 25355 992 25411
rect 1048 25355 1116 25411
rect 1172 25355 1240 25411
rect 1296 25355 1336 25411
rect 858 25287 1336 25355
rect 858 25231 868 25287
rect 924 25231 992 25287
rect 1048 25231 1116 25287
rect 1172 25231 1240 25287
rect 1296 25231 1336 25287
rect 858 25163 1336 25231
rect 858 25107 868 25163
rect 924 25107 992 25163
rect 1048 25107 1116 25163
rect 1172 25107 1240 25163
rect 1296 25107 1336 25163
rect 858 25039 1336 25107
rect 858 24983 868 25039
rect 924 24983 992 25039
rect 1048 24983 1116 25039
rect 1172 24983 1240 25039
rect 1296 24983 1336 25039
rect 858 24915 1336 24983
rect 858 24859 868 24915
rect 924 24859 992 24915
rect 1048 24859 1116 24915
rect 1172 24859 1240 24915
rect 1296 24859 1336 24915
rect 858 24791 1336 24859
rect 858 24735 868 24791
rect 924 24740 992 24791
rect 1048 24740 1116 24791
rect 1172 24740 1240 24791
rect 924 24735 978 24740
rect 1048 24735 1102 24740
rect 1172 24735 1226 24740
rect 1296 24735 1336 24791
rect 858 24688 978 24735
rect 1030 24688 1102 24735
rect 1154 24688 1226 24735
rect 1278 24688 1336 24735
rect 858 24667 1336 24688
rect 858 24611 868 24667
rect 924 24616 992 24667
rect 1048 24616 1116 24667
rect 1172 24616 1240 24667
rect 924 24611 978 24616
rect 1048 24611 1102 24616
rect 1172 24611 1226 24616
rect 1296 24611 1336 24667
rect 858 24564 978 24611
rect 1030 24564 1102 24611
rect 1154 24564 1226 24611
rect 1278 24564 1336 24611
rect 858 24543 1336 24564
rect 858 24487 868 24543
rect 924 24492 992 24543
rect 1048 24492 1116 24543
rect 1172 24492 1240 24543
rect 924 24487 978 24492
rect 1048 24487 1102 24492
rect 1172 24487 1226 24492
rect 1296 24487 1336 24543
rect 858 24440 978 24487
rect 1030 24440 1102 24487
rect 1154 24440 1226 24487
rect 1278 24440 1336 24487
rect 858 24419 1336 24440
rect 858 24363 868 24419
rect 924 24368 992 24419
rect 1048 24368 1116 24419
rect 1172 24368 1240 24419
rect 924 24363 978 24368
rect 1048 24363 1102 24368
rect 1172 24363 1226 24368
rect 1296 24363 1336 24419
rect 858 24316 978 24363
rect 1030 24316 1102 24363
rect 1154 24316 1226 24363
rect 1278 24316 1336 24363
rect 858 24295 1336 24316
rect 858 24239 868 24295
rect 924 24244 992 24295
rect 1048 24244 1116 24295
rect 1172 24244 1240 24295
rect 924 24239 978 24244
rect 1048 24239 1102 24244
rect 1172 24239 1226 24244
rect 1296 24239 1336 24295
rect 858 24192 978 24239
rect 1030 24192 1102 24239
rect 1154 24192 1226 24239
rect 1278 24192 1336 24239
rect 858 24171 1336 24192
rect 858 24115 868 24171
rect 924 24120 992 24171
rect 1048 24120 1116 24171
rect 1172 24120 1240 24171
rect 924 24115 978 24120
rect 1048 24115 1102 24120
rect 1172 24115 1226 24120
rect 1296 24115 1336 24171
rect 858 24068 978 24115
rect 1030 24068 1102 24115
rect 1154 24068 1226 24115
rect 1278 24068 1336 24115
rect 858 24047 1336 24068
rect 858 23991 868 24047
rect 924 23996 992 24047
rect 1048 23996 1116 24047
rect 1172 23996 1240 24047
rect 924 23991 978 23996
rect 1048 23991 1102 23996
rect 1172 23991 1226 23996
rect 1296 23991 1336 24047
rect 858 23944 978 23991
rect 1030 23944 1102 23991
rect 1154 23944 1226 23991
rect 1278 23944 1336 23991
rect 858 23923 1336 23944
rect 858 23867 868 23923
rect 924 23872 992 23923
rect 1048 23872 1116 23923
rect 1172 23872 1240 23923
rect 924 23867 978 23872
rect 1048 23867 1102 23872
rect 1172 23867 1226 23872
rect 1296 23867 1336 23923
rect 858 23820 978 23867
rect 1030 23820 1102 23867
rect 1154 23820 1226 23867
rect 1278 23820 1336 23867
rect 858 23799 1336 23820
rect 858 23743 868 23799
rect 924 23748 992 23799
rect 1048 23748 1116 23799
rect 1172 23748 1240 23799
rect 924 23743 978 23748
rect 1048 23743 1102 23748
rect 1172 23743 1226 23748
rect 1296 23743 1336 23799
rect 858 23733 978 23743
rect 966 23696 978 23733
rect 1030 23696 1102 23743
rect 1154 23696 1226 23743
rect 1278 23696 1336 23743
rect 966 23624 1336 23696
rect 966 23572 978 23624
rect 1030 23572 1102 23624
rect 1154 23572 1226 23624
rect 1278 23572 1336 23624
rect 966 23500 1336 23572
rect 966 23461 978 23500
rect 260 21417 444 21469
rect 496 21417 552 21469
rect 604 21417 660 21469
rect 712 21417 768 21469
rect 260 21361 768 21417
rect 260 21309 444 21361
rect 496 21309 552 21361
rect 604 21309 660 21361
rect 712 21309 768 21361
rect 260 21253 768 21309
rect 260 21201 444 21253
rect 496 21201 552 21253
rect 604 21201 660 21253
rect 712 21201 768 21253
rect 260 13845 768 21201
rect 858 23451 978 23461
rect 1030 23451 1102 23500
rect 1154 23451 1226 23500
rect 1278 23451 1336 23500
rect 858 23395 868 23451
rect 924 23448 978 23451
rect 1048 23448 1102 23451
rect 1172 23448 1226 23451
rect 924 23395 992 23448
rect 1048 23395 1116 23448
rect 1172 23395 1240 23448
rect 1296 23395 1336 23451
rect 858 23376 1336 23395
rect 858 23327 978 23376
rect 1030 23327 1102 23376
rect 1154 23327 1226 23376
rect 1278 23327 1336 23376
rect 858 23271 868 23327
rect 924 23324 978 23327
rect 1048 23324 1102 23327
rect 1172 23324 1226 23327
rect 924 23271 992 23324
rect 1048 23271 1116 23324
rect 1172 23271 1240 23324
rect 1296 23271 1336 23327
rect 858 23252 1336 23271
rect 858 23203 978 23252
rect 1030 23203 1102 23252
rect 1154 23203 1226 23252
rect 1278 23203 1336 23252
rect 858 23147 868 23203
rect 924 23200 978 23203
rect 1048 23200 1102 23203
rect 1172 23200 1226 23203
rect 924 23147 992 23200
rect 1048 23147 1116 23200
rect 1172 23147 1240 23200
rect 1296 23147 1336 23203
rect 858 23128 1336 23147
rect 858 23079 978 23128
rect 1030 23079 1102 23128
rect 1154 23079 1226 23128
rect 1278 23079 1336 23128
rect 858 23023 868 23079
rect 924 23076 978 23079
rect 1048 23076 1102 23079
rect 1172 23076 1226 23079
rect 924 23023 992 23076
rect 1048 23023 1116 23076
rect 1172 23023 1240 23076
rect 1296 23023 1336 23079
rect 858 23004 1336 23023
rect 858 22955 978 23004
rect 1030 22955 1102 23004
rect 1154 22955 1226 23004
rect 1278 22955 1336 23004
rect 858 22899 868 22955
rect 924 22952 978 22955
rect 1048 22952 1102 22955
rect 1172 22952 1226 22955
rect 924 22899 992 22952
rect 1048 22899 1116 22952
rect 1172 22899 1240 22952
rect 1296 22899 1336 22955
rect 858 22880 1336 22899
rect 858 22831 978 22880
rect 1030 22831 1102 22880
rect 1154 22831 1226 22880
rect 1278 22831 1336 22880
rect 858 22775 868 22831
rect 924 22828 978 22831
rect 1048 22828 1102 22831
rect 1172 22828 1226 22831
rect 924 22775 992 22828
rect 1048 22775 1116 22828
rect 1172 22775 1240 22828
rect 1296 22775 1336 22831
rect 858 22756 1336 22775
rect 858 22707 978 22756
rect 1030 22707 1102 22756
rect 1154 22707 1226 22756
rect 1278 22707 1336 22756
rect 858 22651 868 22707
rect 924 22704 978 22707
rect 1048 22704 1102 22707
rect 1172 22704 1226 22707
rect 924 22651 992 22704
rect 1048 22651 1116 22704
rect 1172 22651 1240 22704
rect 1296 22651 1336 22707
rect 858 22632 1336 22651
rect 858 22583 978 22632
rect 1030 22583 1102 22632
rect 1154 22583 1226 22632
rect 1278 22583 1336 22632
rect 858 22527 868 22583
rect 924 22580 978 22583
rect 1048 22580 1102 22583
rect 1172 22580 1226 22583
rect 924 22527 992 22580
rect 1048 22527 1116 22580
rect 1172 22527 1240 22580
rect 1296 22527 1336 22583
rect 858 22508 1336 22527
rect 858 22459 978 22508
rect 1030 22459 1102 22508
rect 1154 22459 1226 22508
rect 1278 22459 1336 22508
rect 858 22403 868 22459
rect 924 22456 978 22459
rect 1048 22456 1102 22459
rect 1172 22456 1226 22459
rect 924 22403 992 22456
rect 1048 22403 1116 22456
rect 1172 22403 1240 22456
rect 1296 22403 1336 22459
rect 858 22384 1336 22403
rect 858 22335 978 22384
rect 1030 22335 1102 22384
rect 1154 22335 1226 22384
rect 1278 22335 1336 22384
rect 858 22279 868 22335
rect 924 22332 978 22335
rect 1048 22332 1102 22335
rect 1172 22332 1226 22335
rect 924 22279 992 22332
rect 1048 22279 1116 22332
rect 1172 22279 1240 22332
rect 1296 22279 1336 22335
rect 858 22260 1336 22279
rect 858 22211 978 22260
rect 1030 22211 1102 22260
rect 1154 22211 1226 22260
rect 1278 22211 1336 22260
rect 858 22155 868 22211
rect 924 22208 978 22211
rect 1048 22208 1102 22211
rect 1172 22208 1226 22211
rect 924 22155 992 22208
rect 1048 22155 1116 22208
rect 1172 22155 1240 22208
rect 1296 22155 1336 22211
rect 858 22136 1336 22155
rect 858 22087 978 22136
rect 1030 22087 1102 22136
rect 1154 22087 1226 22136
rect 1278 22087 1336 22136
rect 858 22031 868 22087
rect 924 22084 978 22087
rect 1048 22084 1102 22087
rect 1172 22084 1226 22087
rect 924 22031 992 22084
rect 1048 22031 1116 22084
rect 1172 22031 1240 22084
rect 1296 22031 1336 22087
rect 858 22012 1336 22031
rect 858 21963 978 22012
rect 1030 21963 1102 22012
rect 1154 21963 1226 22012
rect 1278 21963 1336 22012
rect 858 21907 868 21963
rect 924 21960 978 21963
rect 1048 21960 1102 21963
rect 1172 21960 1226 21963
rect 924 21907 992 21960
rect 1048 21907 1116 21960
rect 1172 21907 1240 21960
rect 1296 21907 1336 21963
rect 858 21888 1336 21907
rect 858 21839 978 21888
rect 1030 21839 1102 21888
rect 1154 21839 1226 21888
rect 1278 21839 1336 21888
rect 858 21783 868 21839
rect 924 21836 978 21839
rect 1048 21836 1102 21839
rect 1172 21836 1226 21839
rect 924 21783 992 21836
rect 1048 21783 1116 21836
rect 1172 21783 1240 21836
rect 1296 21783 1336 21839
rect 858 21764 1336 21783
rect 858 21715 978 21764
rect 1030 21715 1102 21764
rect 1154 21715 1226 21764
rect 1278 21715 1336 21764
rect 858 21659 868 21715
rect 924 21712 978 21715
rect 1048 21712 1102 21715
rect 1172 21712 1226 21715
rect 924 21659 992 21712
rect 1048 21659 1116 21712
rect 1172 21659 1240 21712
rect 1296 21659 1336 21715
rect 858 21640 1336 21659
rect 858 21591 978 21640
rect 1030 21591 1102 21640
rect 1154 21591 1226 21640
rect 1278 21591 1336 21640
rect 858 21535 868 21591
rect 924 21588 978 21591
rect 1048 21588 1102 21591
rect 1172 21588 1226 21591
rect 924 21535 992 21588
rect 1048 21535 1116 21588
rect 1172 21535 1240 21588
rect 1296 21535 1336 21591
rect 858 21467 1336 21535
rect 858 21411 868 21467
rect 924 21411 992 21467
rect 1048 21411 1116 21467
rect 1172 21411 1240 21467
rect 1296 21411 1336 21467
rect 858 21343 1336 21411
rect 858 21287 868 21343
rect 924 21287 992 21343
rect 1048 21287 1116 21343
rect 1172 21287 1240 21343
rect 1296 21287 1336 21343
rect 858 21219 1336 21287
rect 858 21163 868 21219
rect 924 21163 992 21219
rect 1048 21163 1116 21219
rect 1172 21163 1240 21219
rect 1296 21163 1336 21219
rect 858 21095 1336 21163
rect 858 21039 868 21095
rect 924 21039 992 21095
rect 1048 21039 1116 21095
rect 1172 21039 1240 21095
rect 1296 21039 1336 21095
rect 858 20971 1336 21039
rect 858 20915 868 20971
rect 924 20915 992 20971
rect 1048 20915 1116 20971
rect 1172 20915 1240 20971
rect 1296 20915 1336 20971
rect 858 20847 1336 20915
rect 858 20791 868 20847
rect 924 20791 992 20847
rect 1048 20791 1116 20847
rect 1172 20791 1240 20847
rect 1296 20791 1336 20847
rect 858 20723 1336 20791
rect 858 20667 868 20723
rect 924 20667 992 20723
rect 1048 20667 1116 20723
rect 1172 20667 1240 20723
rect 1296 20667 1336 20723
rect 858 20599 1336 20667
rect 858 20543 868 20599
rect 924 20543 992 20599
rect 1048 20543 1116 20599
rect 1172 20543 1240 20599
rect 1296 20543 1336 20599
rect 858 20533 1336 20543
rect 1136 20261 1336 20533
rect 858 20251 1336 20261
rect 858 20195 868 20251
rect 924 20195 992 20251
rect 1048 20195 1116 20251
rect 1172 20195 1240 20251
rect 1296 20195 1336 20251
rect 858 20127 1336 20195
rect 858 20071 868 20127
rect 924 20071 992 20127
rect 1048 20071 1116 20127
rect 1172 20071 1240 20127
rect 1296 20071 1336 20127
rect 858 20003 1336 20071
rect 858 19947 868 20003
rect 924 19947 992 20003
rect 1048 19947 1116 20003
rect 1172 19947 1240 20003
rect 1296 19947 1336 20003
rect 858 19879 1336 19947
rect 858 19823 868 19879
rect 924 19823 992 19879
rect 1048 19823 1116 19879
rect 1172 19823 1240 19879
rect 1296 19823 1336 19879
rect 858 19755 1336 19823
rect 858 19699 868 19755
rect 924 19699 992 19755
rect 1048 19699 1116 19755
rect 1172 19699 1240 19755
rect 1296 19699 1336 19755
rect 858 19631 1336 19699
rect 858 19575 868 19631
rect 924 19575 992 19631
rect 1048 19575 1116 19631
rect 1172 19575 1240 19631
rect 1296 19575 1336 19631
rect 858 19507 1336 19575
rect 858 19451 868 19507
rect 924 19451 992 19507
rect 1048 19451 1116 19507
rect 1172 19451 1240 19507
rect 1296 19451 1336 19507
rect 858 19383 1336 19451
rect 858 19327 868 19383
rect 924 19327 992 19383
rect 1048 19327 1116 19383
rect 1172 19327 1240 19383
rect 1296 19327 1336 19383
rect 858 19259 1336 19327
rect 858 19203 868 19259
rect 924 19203 992 19259
rect 1048 19203 1116 19259
rect 1172 19203 1240 19259
rect 1296 19203 1336 19259
rect 858 19135 1336 19203
rect 858 19079 868 19135
rect 924 19079 992 19135
rect 1048 19079 1116 19135
rect 1172 19079 1240 19135
rect 1296 19079 1336 19135
rect 858 19011 1336 19079
rect 858 18955 868 19011
rect 924 18955 992 19011
rect 1048 18955 1116 19011
rect 1172 18955 1240 19011
rect 1296 18955 1336 19011
rect 858 18887 1336 18955
rect 858 18831 868 18887
rect 924 18831 992 18887
rect 1048 18831 1116 18887
rect 1172 18831 1240 18887
rect 1296 18831 1336 18887
rect 858 18763 1336 18831
rect 858 18707 868 18763
rect 924 18707 992 18763
rect 1048 18707 1116 18763
rect 1172 18707 1240 18763
rect 1296 18707 1336 18763
rect 858 18639 1336 18707
rect 858 18583 868 18639
rect 924 18583 992 18639
rect 1048 18583 1116 18639
rect 1172 18583 1240 18639
rect 1296 18583 1336 18639
rect 858 18515 1336 18583
rect 858 18459 868 18515
rect 924 18459 992 18515
rect 1048 18459 1116 18515
rect 1172 18459 1240 18515
rect 1296 18459 1336 18515
rect 858 18391 1336 18459
rect 858 18335 868 18391
rect 924 18335 992 18391
rect 1048 18335 1116 18391
rect 1172 18335 1240 18391
rect 1296 18335 1336 18391
rect 858 18267 1336 18335
rect 858 18211 868 18267
rect 924 18211 992 18267
rect 1048 18211 1116 18267
rect 1172 18211 1240 18267
rect 1296 18211 1336 18267
rect 858 18143 1336 18211
rect 858 18087 868 18143
rect 924 18087 992 18143
rect 1048 18087 1116 18143
rect 1172 18087 1240 18143
rect 1296 18087 1336 18143
rect 858 18019 1336 18087
rect 858 17963 868 18019
rect 924 17963 992 18019
rect 1048 17963 1116 18019
rect 1172 17963 1240 18019
rect 1296 17963 1336 18019
rect 858 17895 1336 17963
rect 858 17839 868 17895
rect 924 17839 992 17895
rect 1048 17839 1116 17895
rect 1172 17839 1240 17895
rect 1296 17839 1336 17895
rect 858 17771 1336 17839
rect 858 17715 868 17771
rect 924 17715 992 17771
rect 1048 17715 1116 17771
rect 1172 17715 1240 17771
rect 1296 17715 1336 17771
rect 858 17647 1336 17715
rect 858 17591 868 17647
rect 924 17591 992 17647
rect 1048 17591 1116 17647
rect 1172 17591 1240 17647
rect 1296 17591 1336 17647
rect 858 17523 1336 17591
rect 858 17467 868 17523
rect 924 17467 992 17523
rect 1048 17467 1116 17523
rect 1172 17467 1240 17523
rect 1296 17467 1336 17523
rect 858 17399 1336 17467
rect 858 17343 868 17399
rect 924 17343 992 17399
rect 1048 17343 1116 17399
rect 1172 17343 1240 17399
rect 1296 17343 1336 17399
rect 858 17333 1336 17343
rect 1136 17061 1336 17333
rect 858 17051 1336 17061
rect 858 16995 868 17051
rect 924 16995 992 17051
rect 1048 16995 1116 17051
rect 1172 16995 1240 17051
rect 1296 16995 1336 17051
rect 858 16927 1336 16995
rect 858 16871 868 16927
rect 924 16871 992 16927
rect 1048 16871 1116 16927
rect 1172 16871 1240 16927
rect 1296 16871 1336 16927
rect 858 16803 1336 16871
rect 858 16747 868 16803
rect 924 16747 992 16803
rect 1048 16747 1116 16803
rect 1172 16747 1240 16803
rect 1296 16747 1336 16803
rect 858 16679 1336 16747
rect 858 16623 868 16679
rect 924 16623 992 16679
rect 1048 16623 1116 16679
rect 1172 16623 1240 16679
rect 1296 16623 1336 16679
rect 858 16555 1336 16623
rect 858 16499 868 16555
rect 924 16499 992 16555
rect 1048 16499 1116 16555
rect 1172 16499 1240 16555
rect 1296 16499 1336 16555
rect 858 16431 1336 16499
rect 858 16375 868 16431
rect 924 16375 992 16431
rect 1048 16375 1116 16431
rect 1172 16375 1240 16431
rect 1296 16375 1336 16431
rect 858 16307 1336 16375
rect 858 16251 868 16307
rect 924 16251 992 16307
rect 1048 16251 1116 16307
rect 1172 16251 1240 16307
rect 1296 16251 1336 16307
rect 858 16183 1336 16251
rect 858 16127 868 16183
rect 924 16127 992 16183
rect 1048 16127 1116 16183
rect 1172 16127 1240 16183
rect 1296 16127 1336 16183
rect 858 16059 1336 16127
rect 858 16003 868 16059
rect 924 16003 992 16059
rect 1048 16003 1116 16059
rect 1172 16003 1240 16059
rect 1296 16003 1336 16059
rect 858 15935 1336 16003
rect 858 15879 868 15935
rect 924 15879 992 15935
rect 1048 15879 1116 15935
rect 1172 15879 1240 15935
rect 1296 15879 1336 15935
rect 858 15811 1336 15879
rect 858 15755 868 15811
rect 924 15755 992 15811
rect 1048 15755 1116 15811
rect 1172 15755 1240 15811
rect 1296 15755 1336 15811
rect 1396 53101 1904 53169
rect 1396 53045 1436 53101
rect 1492 53045 1560 53101
rect 1616 53045 1684 53101
rect 1740 53045 1808 53101
rect 1864 53045 1904 53101
rect 1396 52996 1438 53045
rect 1490 52996 1562 53045
rect 1614 52996 1686 53045
rect 1738 52996 1810 53045
rect 1862 52996 1904 53045
rect 1396 52977 1904 52996
rect 1396 52921 1436 52977
rect 1492 52921 1560 52977
rect 1616 52921 1684 52977
rect 1740 52921 1808 52977
rect 1864 52921 1904 52977
rect 1396 52872 1438 52921
rect 1490 52872 1562 52921
rect 1614 52872 1686 52921
rect 1738 52872 1810 52921
rect 1862 52872 1904 52921
rect 1396 52853 1904 52872
rect 1396 52797 1436 52853
rect 1492 52797 1560 52853
rect 1616 52797 1684 52853
rect 1740 52797 1808 52853
rect 1864 52797 1904 52853
rect 1396 52748 1438 52797
rect 1490 52748 1562 52797
rect 1614 52748 1686 52797
rect 1738 52748 1810 52797
rect 1862 52748 1904 52797
rect 1396 52729 1904 52748
rect 1396 52673 1436 52729
rect 1492 52673 1560 52729
rect 1616 52673 1684 52729
rect 1740 52673 1808 52729
rect 1864 52673 1904 52729
rect 1396 52624 1438 52673
rect 1490 52624 1562 52673
rect 1614 52624 1686 52673
rect 1738 52624 1810 52673
rect 1862 52624 1904 52673
rect 1396 52605 1904 52624
rect 1396 52549 1436 52605
rect 1492 52549 1560 52605
rect 1616 52549 1684 52605
rect 1740 52549 1808 52605
rect 1864 52549 1904 52605
rect 1396 52500 1438 52549
rect 1490 52500 1562 52549
rect 1614 52500 1686 52549
rect 1738 52500 1810 52549
rect 1862 52500 1904 52549
rect 1396 49100 1904 52500
rect 1396 49048 1438 49100
rect 1490 49048 1562 49100
rect 1614 49048 1686 49100
rect 1738 49048 1810 49100
rect 1862 49048 1904 49100
rect 1396 49045 1904 49048
rect 1396 48989 1436 49045
rect 1492 48989 1560 49045
rect 1616 48989 1684 49045
rect 1740 48989 1808 49045
rect 1864 48989 1904 49045
rect 1396 48976 1904 48989
rect 1396 48924 1438 48976
rect 1490 48924 1562 48976
rect 1614 48924 1686 48976
rect 1738 48924 1810 48976
rect 1862 48924 1904 48976
rect 1396 48921 1904 48924
rect 1396 48865 1436 48921
rect 1492 48865 1560 48921
rect 1616 48865 1684 48921
rect 1740 48865 1808 48921
rect 1864 48865 1904 48921
rect 1396 48852 1904 48865
rect 1396 48800 1438 48852
rect 1490 48800 1562 48852
rect 1614 48800 1686 48852
rect 1738 48800 1810 48852
rect 1862 48800 1904 48852
rect 1396 48797 1904 48800
rect 1396 48741 1436 48797
rect 1492 48741 1560 48797
rect 1616 48741 1684 48797
rect 1740 48741 1808 48797
rect 1864 48741 1904 48797
rect 1396 48728 1904 48741
rect 1396 48676 1438 48728
rect 1490 48676 1562 48728
rect 1614 48676 1686 48728
rect 1738 48676 1810 48728
rect 1862 48676 1904 48728
rect 1396 48673 1904 48676
rect 1396 48617 1436 48673
rect 1492 48617 1560 48673
rect 1616 48617 1684 48673
rect 1740 48617 1808 48673
rect 1864 48617 1904 48673
rect 1396 48604 1904 48617
rect 1396 48552 1438 48604
rect 1490 48552 1562 48604
rect 1614 48552 1686 48604
rect 1738 48552 1810 48604
rect 1862 48552 1904 48604
rect 1396 48549 1904 48552
rect 1396 48493 1436 48549
rect 1492 48493 1560 48549
rect 1616 48493 1684 48549
rect 1740 48493 1808 48549
rect 1864 48493 1904 48549
rect 1396 48425 1904 48493
rect 1396 48369 1436 48425
rect 1492 48369 1560 48425
rect 1616 48369 1684 48425
rect 1740 48369 1808 48425
rect 1864 48369 1904 48425
rect 1396 48301 1904 48369
rect 1396 48245 1436 48301
rect 1492 48245 1560 48301
rect 1616 48245 1684 48301
rect 1740 48245 1808 48301
rect 1864 48245 1904 48301
rect 1396 48177 1904 48245
rect 1396 48121 1436 48177
rect 1492 48121 1560 48177
rect 1616 48121 1684 48177
rect 1740 48121 1808 48177
rect 1864 48121 1904 48177
rect 1396 48053 1904 48121
rect 1396 47997 1436 48053
rect 1492 47997 1560 48053
rect 1616 47997 1684 48053
rect 1740 47997 1808 48053
rect 1864 47997 1904 48053
rect 1396 47929 1904 47997
rect 1396 47873 1436 47929
rect 1492 47873 1560 47929
rect 1616 47873 1684 47929
rect 1740 47873 1808 47929
rect 1864 47873 1904 47929
rect 1396 47805 1904 47873
rect 1396 47749 1436 47805
rect 1492 47749 1560 47805
rect 1616 47749 1684 47805
rect 1740 47749 1808 47805
rect 1864 47749 1904 47805
rect 1396 45845 1904 47749
rect 1396 45789 1436 45845
rect 1492 45789 1560 45845
rect 1616 45789 1684 45845
rect 1740 45789 1808 45845
rect 1864 45789 1904 45845
rect 1396 45721 1904 45789
rect 1396 45665 1436 45721
rect 1492 45665 1560 45721
rect 1616 45665 1684 45721
rect 1740 45665 1808 45721
rect 1864 45665 1904 45721
rect 1396 45597 1904 45665
rect 1396 45541 1436 45597
rect 1492 45541 1560 45597
rect 1616 45541 1684 45597
rect 1740 45541 1808 45597
rect 1864 45541 1904 45597
rect 1396 45473 1904 45541
rect 1396 45417 1436 45473
rect 1492 45417 1560 45473
rect 1616 45417 1684 45473
rect 1740 45417 1808 45473
rect 1864 45417 1904 45473
rect 1396 45349 1904 45417
rect 1396 45293 1436 45349
rect 1492 45293 1560 45349
rect 1616 45293 1684 45349
rect 1740 45293 1808 45349
rect 1864 45293 1904 45349
rect 1396 45225 1904 45293
rect 1396 45169 1436 45225
rect 1492 45169 1560 45225
rect 1616 45169 1684 45225
rect 1740 45169 1808 45225
rect 1864 45169 1904 45225
rect 1396 45152 1904 45169
rect 1396 45101 1438 45152
rect 1490 45101 1562 45152
rect 1614 45101 1686 45152
rect 1738 45101 1810 45152
rect 1862 45101 1904 45152
rect 1396 45045 1436 45101
rect 1492 45045 1560 45101
rect 1616 45045 1684 45101
rect 1740 45045 1808 45101
rect 1864 45045 1904 45101
rect 1396 45028 1904 45045
rect 1396 44977 1438 45028
rect 1490 44977 1562 45028
rect 1614 44977 1686 45028
rect 1738 44977 1810 45028
rect 1862 44977 1904 45028
rect 1396 44921 1436 44977
rect 1492 44921 1560 44977
rect 1616 44921 1684 44977
rect 1740 44921 1808 44977
rect 1864 44921 1904 44977
rect 1396 44904 1904 44921
rect 1396 44853 1438 44904
rect 1490 44853 1562 44904
rect 1614 44853 1686 44904
rect 1738 44853 1810 44904
rect 1862 44853 1904 44904
rect 1396 44797 1436 44853
rect 1492 44797 1560 44853
rect 1616 44797 1684 44853
rect 1740 44797 1808 44853
rect 1864 44797 1904 44853
rect 1396 44780 1904 44797
rect 1396 44729 1438 44780
rect 1490 44729 1562 44780
rect 1614 44729 1686 44780
rect 1738 44729 1810 44780
rect 1862 44729 1904 44780
rect 1396 44673 1436 44729
rect 1492 44673 1560 44729
rect 1616 44673 1684 44729
rect 1740 44673 1808 44729
rect 1864 44673 1904 44729
rect 1396 44656 1904 44673
rect 1396 44605 1438 44656
rect 1490 44605 1562 44656
rect 1614 44605 1686 44656
rect 1738 44605 1810 44656
rect 1862 44605 1904 44656
rect 1396 44549 1436 44605
rect 1492 44549 1560 44605
rect 1616 44549 1684 44605
rect 1740 44549 1808 44605
rect 1864 44549 1904 44605
rect 1396 41204 1904 44549
rect 1396 41152 1438 41204
rect 1490 41152 1562 41204
rect 1614 41152 1686 41204
rect 1738 41152 1810 41204
rect 1862 41152 1904 41204
rect 1396 41080 1904 41152
rect 1396 41028 1438 41080
rect 1490 41028 1562 41080
rect 1614 41028 1686 41080
rect 1738 41028 1810 41080
rect 1862 41028 1904 41080
rect 1396 40956 1904 41028
rect 1396 40904 1438 40956
rect 1490 40904 1562 40956
rect 1614 40904 1686 40956
rect 1738 40904 1810 40956
rect 1862 40904 1904 40956
rect 1396 40832 1904 40904
rect 1396 40780 1438 40832
rect 1490 40780 1562 40832
rect 1614 40780 1686 40832
rect 1738 40780 1810 40832
rect 1862 40780 1904 40832
rect 1396 40708 1904 40780
rect 1396 40656 1438 40708
rect 1490 40656 1562 40708
rect 1614 40656 1686 40708
rect 1738 40656 1810 40708
rect 1862 40656 1904 40708
rect 1396 37256 1904 40656
rect 1396 37204 1438 37256
rect 1490 37204 1562 37256
rect 1614 37204 1686 37256
rect 1738 37204 1810 37256
rect 1862 37204 1904 37256
rect 1396 37132 1904 37204
rect 1396 37080 1438 37132
rect 1490 37080 1562 37132
rect 1614 37080 1686 37132
rect 1738 37080 1810 37132
rect 1862 37080 1904 37132
rect 1396 37008 1904 37080
rect 1396 36956 1438 37008
rect 1490 36956 1562 37008
rect 1614 36956 1686 37008
rect 1738 36956 1810 37008
rect 1862 36956 1904 37008
rect 1396 36884 1904 36956
rect 1396 36832 1438 36884
rect 1490 36832 1562 36884
rect 1614 36832 1686 36884
rect 1738 36832 1810 36884
rect 1862 36832 1904 36884
rect 1396 36760 1904 36832
rect 1396 36708 1438 36760
rect 1490 36708 1562 36760
rect 1614 36708 1686 36760
rect 1738 36708 1810 36760
rect 1862 36708 1904 36760
rect 1396 36251 1904 36708
rect 1396 36195 1436 36251
rect 1492 36195 1560 36251
rect 1616 36195 1684 36251
rect 1740 36195 1808 36251
rect 1864 36195 1904 36251
rect 1396 36127 1904 36195
rect 1396 36071 1436 36127
rect 1492 36071 1560 36127
rect 1616 36071 1684 36127
rect 1740 36071 1808 36127
rect 1864 36071 1904 36127
rect 1396 36003 1904 36071
rect 1396 35947 1436 36003
rect 1492 35947 1560 36003
rect 1616 35947 1684 36003
rect 1740 35947 1808 36003
rect 1864 35947 1904 36003
rect 1396 35879 1904 35947
rect 1396 35823 1436 35879
rect 1492 35823 1560 35879
rect 1616 35823 1684 35879
rect 1740 35823 1808 35879
rect 1864 35823 1904 35879
rect 1396 35755 1904 35823
rect 1396 35699 1436 35755
rect 1492 35699 1560 35755
rect 1616 35699 1684 35755
rect 1740 35699 1808 35755
rect 1864 35699 1904 35755
rect 1396 35631 1904 35699
rect 1396 35575 1436 35631
rect 1492 35575 1560 35631
rect 1616 35575 1684 35631
rect 1740 35575 1808 35631
rect 1864 35575 1904 35631
rect 1396 35507 1904 35575
rect 1396 35451 1436 35507
rect 1492 35451 1560 35507
rect 1616 35451 1684 35507
rect 1740 35451 1808 35507
rect 1864 35451 1904 35507
rect 1396 35383 1904 35451
rect 1396 35327 1436 35383
rect 1492 35327 1560 35383
rect 1616 35327 1684 35383
rect 1740 35327 1808 35383
rect 1864 35327 1904 35383
rect 1396 35259 1904 35327
rect 1396 35203 1436 35259
rect 1492 35203 1560 35259
rect 1616 35203 1684 35259
rect 1740 35203 1808 35259
rect 1864 35203 1904 35259
rect 1396 35135 1904 35203
rect 1396 35079 1436 35135
rect 1492 35079 1560 35135
rect 1616 35079 1684 35135
rect 1740 35079 1808 35135
rect 1864 35079 1904 35135
rect 1396 35011 1904 35079
rect 1396 34955 1436 35011
rect 1492 34955 1560 35011
rect 1616 34955 1684 35011
rect 1740 34955 1808 35011
rect 1864 34955 1904 35011
rect 1396 34887 1904 34955
rect 1396 34831 1436 34887
rect 1492 34831 1560 34887
rect 1616 34831 1684 34887
rect 1740 34831 1808 34887
rect 1864 34831 1904 34887
rect 1396 34763 1904 34831
rect 1396 34707 1436 34763
rect 1492 34707 1560 34763
rect 1616 34707 1684 34763
rect 1740 34707 1808 34763
rect 1864 34707 1904 34763
rect 1396 34639 1904 34707
rect 1396 34583 1436 34639
rect 1492 34583 1560 34639
rect 1616 34583 1684 34639
rect 1740 34583 1808 34639
rect 1864 34583 1904 34639
rect 1396 34515 1904 34583
rect 1396 34459 1436 34515
rect 1492 34459 1560 34515
rect 1616 34459 1684 34515
rect 1740 34459 1808 34515
rect 1864 34459 1904 34515
rect 1396 34391 1904 34459
rect 1396 34335 1436 34391
rect 1492 34335 1560 34391
rect 1616 34335 1684 34391
rect 1740 34335 1808 34391
rect 1864 34335 1904 34391
rect 1396 34267 1904 34335
rect 1396 34211 1436 34267
rect 1492 34211 1560 34267
rect 1616 34211 1684 34267
rect 1740 34211 1808 34267
rect 1864 34211 1904 34267
rect 1396 34143 1904 34211
rect 1396 34087 1436 34143
rect 1492 34087 1560 34143
rect 1616 34087 1684 34143
rect 1740 34087 1808 34143
rect 1864 34087 1904 34143
rect 1396 34019 1904 34087
rect 1396 33963 1436 34019
rect 1492 33963 1560 34019
rect 1616 33963 1684 34019
rect 1740 33963 1808 34019
rect 1864 33963 1904 34019
rect 1396 33895 1904 33963
rect 1396 33839 1436 33895
rect 1492 33839 1560 33895
rect 1616 33839 1684 33895
rect 1740 33839 1808 33895
rect 1864 33839 1904 33895
rect 1396 33771 1904 33839
rect 1396 33715 1436 33771
rect 1492 33715 1560 33771
rect 1616 33715 1684 33771
rect 1740 33715 1808 33771
rect 1864 33715 1904 33771
rect 1396 33647 1904 33715
rect 1396 33591 1436 33647
rect 1492 33591 1560 33647
rect 1616 33591 1684 33647
rect 1740 33591 1808 33647
rect 1864 33591 1904 33647
rect 1396 33523 1904 33591
rect 1396 33467 1436 33523
rect 1492 33467 1560 33523
rect 1616 33467 1684 33523
rect 1740 33467 1808 33523
rect 1864 33467 1904 33523
rect 1396 33399 1904 33467
rect 1396 33343 1436 33399
rect 1492 33343 1560 33399
rect 1616 33343 1684 33399
rect 1740 33343 1808 33399
rect 1864 33343 1904 33399
rect 1396 33308 1904 33343
rect 1396 33256 1438 33308
rect 1490 33256 1562 33308
rect 1614 33256 1686 33308
rect 1738 33256 1810 33308
rect 1862 33256 1904 33308
rect 1396 33184 1904 33256
rect 1396 33132 1438 33184
rect 1490 33132 1562 33184
rect 1614 33132 1686 33184
rect 1738 33132 1810 33184
rect 1862 33132 1904 33184
rect 1396 33060 1904 33132
rect 1396 33008 1438 33060
rect 1490 33008 1562 33060
rect 1614 33008 1686 33060
rect 1738 33008 1810 33060
rect 1862 33008 1904 33060
rect 1396 32936 1904 33008
rect 1396 32884 1438 32936
rect 1490 32884 1562 32936
rect 1614 32884 1686 32936
rect 1738 32884 1810 32936
rect 1862 32884 1904 32936
rect 1396 32812 1904 32884
rect 1396 32760 1438 32812
rect 1490 32760 1562 32812
rect 1614 32760 1686 32812
rect 1738 32760 1810 32812
rect 1862 32760 1904 32812
rect 1396 29360 1904 32760
rect 1396 29308 1438 29360
rect 1490 29308 1562 29360
rect 1614 29308 1686 29360
rect 1738 29308 1810 29360
rect 1862 29308 1904 29360
rect 1396 29236 1904 29308
rect 1396 29184 1438 29236
rect 1490 29184 1562 29236
rect 1614 29184 1686 29236
rect 1738 29184 1810 29236
rect 1862 29184 1904 29236
rect 1396 29112 1904 29184
rect 1396 29060 1438 29112
rect 1490 29060 1562 29112
rect 1614 29060 1686 29112
rect 1738 29060 1810 29112
rect 1862 29060 1904 29112
rect 1396 28988 1904 29060
rect 1396 28936 1438 28988
rect 1490 28936 1562 28988
rect 1614 28936 1686 28988
rect 1738 28936 1810 28988
rect 1862 28936 1904 28988
rect 1396 28864 1904 28936
rect 1396 28812 1438 28864
rect 1490 28812 1562 28864
rect 1614 28812 1686 28864
rect 1738 28812 1810 28864
rect 1862 28812 1904 28864
rect 1396 28245 1904 28812
rect 1396 28189 1436 28245
rect 1492 28189 1560 28245
rect 1616 28189 1684 28245
rect 1740 28189 1808 28245
rect 1864 28189 1904 28245
rect 1396 28121 1904 28189
rect 1396 28065 1436 28121
rect 1492 28065 1560 28121
rect 1616 28065 1684 28121
rect 1740 28065 1808 28121
rect 1864 28065 1904 28121
rect 1396 27997 1904 28065
rect 1396 27941 1436 27997
rect 1492 27941 1560 27997
rect 1616 27941 1684 27997
rect 1740 27941 1808 27997
rect 1864 27941 1904 27997
rect 1396 27873 1904 27941
rect 1396 27817 1436 27873
rect 1492 27817 1560 27873
rect 1616 27817 1684 27873
rect 1740 27817 1808 27873
rect 1864 27817 1904 27873
rect 1396 27749 1904 27817
rect 1396 27693 1436 27749
rect 1492 27693 1560 27749
rect 1616 27693 1684 27749
rect 1740 27693 1808 27749
rect 1864 27693 1904 27749
rect 1396 27625 1904 27693
rect 1396 27569 1436 27625
rect 1492 27569 1560 27625
rect 1616 27569 1684 27625
rect 1740 27569 1808 27625
rect 1864 27569 1904 27625
rect 1396 27501 1904 27569
rect 1396 27445 1436 27501
rect 1492 27445 1560 27501
rect 1616 27445 1684 27501
rect 1740 27445 1808 27501
rect 1864 27445 1904 27501
rect 1396 27377 1904 27445
rect 1396 27321 1436 27377
rect 1492 27321 1560 27377
rect 1616 27321 1684 27377
rect 1740 27321 1808 27377
rect 1864 27321 1904 27377
rect 1396 27253 1904 27321
rect 1396 27197 1436 27253
rect 1492 27197 1560 27253
rect 1616 27197 1684 27253
rect 1740 27197 1808 27253
rect 1864 27197 1904 27253
rect 1396 27129 1904 27197
rect 1396 27073 1436 27129
rect 1492 27073 1560 27129
rect 1616 27073 1684 27129
rect 1740 27073 1808 27129
rect 1864 27073 1904 27129
rect 1396 27005 1904 27073
rect 1396 26949 1436 27005
rect 1492 26949 1560 27005
rect 1616 26949 1684 27005
rect 1740 26949 1808 27005
rect 1864 26949 1904 27005
rect 1396 25412 1904 26949
rect 1396 25360 1438 25412
rect 1490 25360 1562 25412
rect 1614 25360 1686 25412
rect 1738 25360 1810 25412
rect 1862 25360 1904 25412
rect 1396 25288 1904 25360
rect 1396 25236 1438 25288
rect 1490 25236 1562 25288
rect 1614 25236 1686 25288
rect 1738 25236 1810 25288
rect 1862 25236 1904 25288
rect 1396 25164 1904 25236
rect 1396 25112 1438 25164
rect 1490 25112 1562 25164
rect 1614 25112 1686 25164
rect 1738 25112 1810 25164
rect 1862 25112 1904 25164
rect 1396 25040 1904 25112
rect 1396 24988 1438 25040
rect 1490 24988 1562 25040
rect 1614 24988 1686 25040
rect 1738 24988 1810 25040
rect 1862 24988 1904 25040
rect 1396 24916 1904 24988
rect 1396 24864 1438 24916
rect 1490 24864 1562 24916
rect 1614 24864 1686 24916
rect 1738 24864 1810 24916
rect 1862 24864 1904 24916
rect 1396 21469 1904 24864
rect 1396 21417 1408 21469
rect 1460 21417 1516 21469
rect 1568 21417 1624 21469
rect 1676 21417 1732 21469
rect 1784 21417 1840 21469
rect 1892 21417 1904 21469
rect 1396 21361 1904 21417
rect 1396 21309 1408 21361
rect 1460 21309 1516 21361
rect 1568 21309 1624 21361
rect 1676 21309 1732 21361
rect 1784 21309 1840 21361
rect 1892 21309 1904 21361
rect 1396 21253 1904 21309
rect 1396 21201 1408 21253
rect 1460 21201 1516 21253
rect 1568 21201 1624 21253
rect 1676 21201 1732 21253
rect 1784 21201 1840 21253
rect 1892 21201 1904 21253
rect 1396 15762 1904 21201
rect 1964 55445 2472 56975
rect 1964 55389 2004 55445
rect 2060 55389 2128 55445
rect 2184 55389 2252 55445
rect 2308 55389 2376 55445
rect 2432 55389 2472 55445
rect 1964 55321 2472 55389
rect 1964 55265 2004 55321
rect 2060 55265 2128 55321
rect 2184 55265 2252 55321
rect 2308 55265 2376 55321
rect 2432 55265 2472 55321
rect 1964 55197 2472 55265
rect 1964 55141 2004 55197
rect 2060 55141 2128 55197
rect 2184 55141 2252 55197
rect 2308 55141 2376 55197
rect 2432 55141 2472 55197
rect 1964 55073 2472 55141
rect 1964 55017 2004 55073
rect 2060 55017 2128 55073
rect 2184 55017 2252 55073
rect 2308 55017 2376 55073
rect 2432 55017 2472 55073
rect 1964 54949 2472 55017
rect 1964 54893 2004 54949
rect 2060 54893 2128 54949
rect 2184 54893 2252 54949
rect 2308 54893 2376 54949
rect 2432 54893 2472 54949
rect 1964 54825 2472 54893
rect 1964 54769 2004 54825
rect 2060 54769 2128 54825
rect 2184 54769 2252 54825
rect 2308 54769 2376 54825
rect 2432 54769 2472 54825
rect 1964 54701 2472 54769
rect 1964 54645 2004 54701
rect 2060 54645 2128 54701
rect 2184 54645 2252 54701
rect 2308 54645 2376 54701
rect 2432 54645 2472 54701
rect 1964 54577 2472 54645
rect 1964 54521 2004 54577
rect 2060 54521 2128 54577
rect 2184 54521 2252 54577
rect 2308 54521 2376 54577
rect 2432 54521 2472 54577
rect 1964 54453 2472 54521
rect 1964 54397 2004 54453
rect 2060 54397 2128 54453
rect 2184 54397 2252 54453
rect 2308 54397 2376 54453
rect 2432 54397 2472 54453
rect 1964 54329 2472 54397
rect 1964 54273 2004 54329
rect 2060 54273 2128 54329
rect 2184 54273 2252 54329
rect 2308 54273 2376 54329
rect 2432 54273 2472 54329
rect 1964 54205 2472 54273
rect 1964 54149 2004 54205
rect 2060 54149 2128 54205
rect 2184 54149 2252 54205
rect 2308 54149 2376 54205
rect 2432 54149 2472 54205
rect 1964 47445 2472 54149
rect 1964 47389 2004 47445
rect 2060 47389 2128 47445
rect 2184 47389 2252 47445
rect 2308 47389 2376 47445
rect 2432 47389 2472 47445
rect 1964 47321 2472 47389
rect 1964 47265 2004 47321
rect 2060 47265 2128 47321
rect 2184 47265 2252 47321
rect 2308 47265 2376 47321
rect 2432 47265 2472 47321
rect 1964 47197 2472 47265
rect 1964 47141 2004 47197
rect 2060 47141 2128 47197
rect 2184 47141 2252 47197
rect 2308 47141 2376 47197
rect 2432 47141 2472 47197
rect 1964 47073 2472 47141
rect 1964 47017 2004 47073
rect 2060 47017 2128 47073
rect 2184 47017 2252 47073
rect 2308 47017 2376 47073
rect 2432 47017 2472 47073
rect 1964 46949 2472 47017
rect 1964 46893 2004 46949
rect 2060 46893 2128 46949
rect 2184 46893 2252 46949
rect 2308 46893 2376 46949
rect 2432 46893 2472 46949
rect 1964 46825 2472 46893
rect 1964 46769 2004 46825
rect 2060 46769 2128 46825
rect 2184 46769 2252 46825
rect 2308 46769 2376 46825
rect 2432 46769 2472 46825
rect 1964 46701 2472 46769
rect 1964 46645 2004 46701
rect 2060 46645 2128 46701
rect 2184 46645 2252 46701
rect 2308 46645 2376 46701
rect 2432 46645 2472 46701
rect 1964 46577 2472 46645
rect 1964 46521 2004 46577
rect 2060 46521 2128 46577
rect 2184 46521 2252 46577
rect 2308 46521 2376 46577
rect 2432 46521 2472 46577
rect 1964 46453 2472 46521
rect 1964 46397 2004 46453
rect 2060 46397 2128 46453
rect 2184 46397 2252 46453
rect 2308 46397 2376 46453
rect 2432 46397 2472 46453
rect 1964 46329 2472 46397
rect 1964 46273 2004 46329
rect 2060 46273 2128 46329
rect 2184 46273 2252 46329
rect 2308 46273 2376 46329
rect 2432 46273 2472 46329
rect 1964 46205 2472 46273
rect 1964 46149 2004 46205
rect 2060 46149 2128 46205
rect 2184 46149 2252 46205
rect 2308 46149 2376 46205
rect 2432 46149 2472 46205
rect 1964 44245 2472 46149
rect 1964 44189 2004 44245
rect 2060 44189 2128 44245
rect 2184 44189 2252 44245
rect 2308 44189 2376 44245
rect 2432 44189 2472 44245
rect 1964 44121 2472 44189
rect 1964 44065 2004 44121
rect 2060 44065 2128 44121
rect 2184 44065 2252 44121
rect 2308 44065 2376 44121
rect 2432 44065 2472 44121
rect 1964 43997 2472 44065
rect 1964 43941 2004 43997
rect 2060 43941 2128 43997
rect 2184 43941 2252 43997
rect 2308 43941 2376 43997
rect 2432 43941 2472 43997
rect 1964 43873 2472 43941
rect 1964 43817 2004 43873
rect 2060 43817 2128 43873
rect 2184 43817 2252 43873
rect 2308 43817 2376 43873
rect 2432 43817 2472 43873
rect 1964 43749 2472 43817
rect 1964 43693 2004 43749
rect 2060 43693 2128 43749
rect 2184 43693 2252 43749
rect 2308 43693 2376 43749
rect 2432 43693 2472 43749
rect 1964 43625 2472 43693
rect 1964 43569 2004 43625
rect 2060 43569 2128 43625
rect 2184 43569 2252 43625
rect 2308 43569 2376 43625
rect 2432 43569 2472 43625
rect 1964 43501 2472 43569
rect 1964 43445 2004 43501
rect 2060 43445 2128 43501
rect 2184 43445 2252 43501
rect 2308 43445 2376 43501
rect 2432 43445 2472 43501
rect 1964 43377 2472 43445
rect 1964 43321 2004 43377
rect 2060 43321 2128 43377
rect 2184 43321 2252 43377
rect 2308 43321 2376 43377
rect 2432 43321 2472 43377
rect 1964 43253 2472 43321
rect 1964 43197 2004 43253
rect 2060 43197 2128 43253
rect 2184 43197 2252 43253
rect 2308 43197 2376 43253
rect 2432 43197 2472 43253
rect 1964 43129 2472 43197
rect 1964 43073 2004 43129
rect 2060 43073 2128 43129
rect 2184 43073 2252 43129
rect 2308 43073 2376 43129
rect 2432 43073 2472 43129
rect 1964 43005 2472 43073
rect 1964 42949 2004 43005
rect 2060 42949 2128 43005
rect 2184 42949 2252 43005
rect 2308 42949 2376 43005
rect 2432 42949 2472 43005
rect 1964 42645 2472 42949
rect 1964 42589 2004 42645
rect 2060 42589 2128 42645
rect 2184 42589 2252 42645
rect 2308 42589 2376 42645
rect 2432 42589 2472 42645
rect 1964 42521 2472 42589
rect 1964 42465 2004 42521
rect 2060 42465 2128 42521
rect 2184 42465 2252 42521
rect 2308 42465 2376 42521
rect 2432 42465 2472 42521
rect 1964 42397 2472 42465
rect 1964 42341 2004 42397
rect 2060 42341 2128 42397
rect 2184 42341 2252 42397
rect 2308 42341 2376 42397
rect 2432 42341 2472 42397
rect 1964 42273 2472 42341
rect 1964 42217 2004 42273
rect 2060 42217 2128 42273
rect 2184 42217 2252 42273
rect 2308 42217 2376 42273
rect 2432 42217 2472 42273
rect 1964 42149 2472 42217
rect 1964 42093 2004 42149
rect 2060 42093 2128 42149
rect 2184 42093 2252 42149
rect 2308 42093 2376 42149
rect 2432 42093 2472 42149
rect 1964 42025 2472 42093
rect 1964 41969 2004 42025
rect 2060 41969 2128 42025
rect 2184 41969 2252 42025
rect 2308 41969 2376 42025
rect 2432 41969 2472 42025
rect 1964 41901 2472 41969
rect 1964 41845 2004 41901
rect 2060 41845 2128 41901
rect 2184 41845 2252 41901
rect 2308 41845 2376 41901
rect 2432 41845 2472 41901
rect 1964 41777 2472 41845
rect 1964 41721 2004 41777
rect 2060 41721 2128 41777
rect 2184 41721 2252 41777
rect 2308 41721 2376 41777
rect 2432 41721 2472 41777
rect 1964 41653 2472 41721
rect 1964 41597 2004 41653
rect 2060 41597 2128 41653
rect 2184 41597 2252 41653
rect 2308 41597 2376 41653
rect 2432 41597 2472 41653
rect 1964 41529 2472 41597
rect 1964 41473 2004 41529
rect 2060 41473 2128 41529
rect 2184 41473 2252 41529
rect 2308 41473 2376 41529
rect 2432 41473 2472 41529
rect 1964 41405 2472 41473
rect 1964 41349 2004 41405
rect 2060 41349 2128 41405
rect 2184 41349 2252 41405
rect 2308 41349 2376 41405
rect 2432 41349 2472 41405
rect 1964 41045 2472 41349
rect 1964 40989 2004 41045
rect 2060 40989 2128 41045
rect 2184 40989 2252 41045
rect 2308 40989 2376 41045
rect 2432 40989 2472 41045
rect 1964 40921 2472 40989
rect 1964 40865 2004 40921
rect 2060 40865 2128 40921
rect 2184 40865 2252 40921
rect 2308 40865 2376 40921
rect 2432 40865 2472 40921
rect 1964 40797 2472 40865
rect 1964 40741 2004 40797
rect 2060 40741 2128 40797
rect 2184 40741 2252 40797
rect 2308 40741 2376 40797
rect 2432 40741 2472 40797
rect 1964 40673 2472 40741
rect 1964 40617 2004 40673
rect 2060 40617 2128 40673
rect 2184 40617 2252 40673
rect 2308 40617 2376 40673
rect 2432 40617 2472 40673
rect 1964 40549 2472 40617
rect 1964 40493 2004 40549
rect 2060 40493 2128 40549
rect 2184 40493 2252 40549
rect 2308 40493 2376 40549
rect 2432 40493 2472 40549
rect 1964 40425 2472 40493
rect 1964 40369 2004 40425
rect 2060 40369 2128 40425
rect 2184 40369 2252 40425
rect 2308 40369 2376 40425
rect 2432 40369 2472 40425
rect 1964 40301 2472 40369
rect 1964 40245 2004 40301
rect 2060 40245 2128 40301
rect 2184 40245 2252 40301
rect 2308 40245 2376 40301
rect 2432 40245 2472 40301
rect 1964 40177 2472 40245
rect 1964 40121 2004 40177
rect 2060 40121 2128 40177
rect 2184 40121 2252 40177
rect 2308 40121 2376 40177
rect 2432 40121 2472 40177
rect 1964 40053 2472 40121
rect 1964 39997 2004 40053
rect 2060 39997 2128 40053
rect 2184 39997 2252 40053
rect 2308 39997 2376 40053
rect 2432 39997 2472 40053
rect 1964 39929 2472 39997
rect 1964 39873 2004 39929
rect 2060 39873 2128 39929
rect 2184 39873 2252 39929
rect 2308 39873 2376 39929
rect 2432 39873 2472 39929
rect 1964 39805 2472 39873
rect 1964 39749 2004 39805
rect 2060 39749 2128 39805
rect 2184 39749 2252 39805
rect 2308 39749 2376 39805
rect 2432 39749 2472 39805
rect 1964 33051 2472 39749
rect 1964 32995 2004 33051
rect 2060 32995 2128 33051
rect 2184 32995 2252 33051
rect 2308 32995 2376 33051
rect 2432 32995 2472 33051
rect 1964 32927 2472 32995
rect 1964 32871 2004 32927
rect 2060 32871 2128 32927
rect 2184 32871 2252 32927
rect 2308 32871 2376 32927
rect 2432 32871 2472 32927
rect 1964 32803 2472 32871
rect 1964 32747 2004 32803
rect 2060 32747 2128 32803
rect 2184 32747 2252 32803
rect 2308 32747 2376 32803
rect 2432 32747 2472 32803
rect 1964 32679 2472 32747
rect 1964 32623 2004 32679
rect 2060 32623 2128 32679
rect 2184 32623 2252 32679
rect 2308 32623 2376 32679
rect 2432 32623 2472 32679
rect 1964 32555 2472 32623
rect 1964 32499 2004 32555
rect 2060 32499 2128 32555
rect 2184 32499 2252 32555
rect 2308 32499 2376 32555
rect 2432 32499 2472 32555
rect 1964 32431 2472 32499
rect 1964 32375 2004 32431
rect 2060 32375 2128 32431
rect 2184 32375 2252 32431
rect 2308 32375 2376 32431
rect 2432 32375 2472 32431
rect 1964 32307 2472 32375
rect 1964 32251 2004 32307
rect 2060 32251 2128 32307
rect 2184 32251 2252 32307
rect 2308 32251 2376 32307
rect 2432 32251 2472 32307
rect 1964 32183 2472 32251
rect 1964 32127 2004 32183
rect 2060 32127 2128 32183
rect 2184 32127 2252 32183
rect 2308 32127 2376 32183
rect 2432 32127 2472 32183
rect 1964 32059 2472 32127
rect 1964 32003 2004 32059
rect 2060 32003 2128 32059
rect 2184 32003 2252 32059
rect 2308 32003 2376 32059
rect 2432 32003 2472 32059
rect 1964 31935 2472 32003
rect 1964 31879 2004 31935
rect 2060 31879 2128 31935
rect 2184 31879 2252 31935
rect 2308 31879 2376 31935
rect 2432 31879 2472 31935
rect 1964 31811 2472 31879
rect 1964 31755 2004 31811
rect 2060 31755 2128 31811
rect 2184 31755 2252 31811
rect 2308 31755 2376 31811
rect 2432 31755 2472 31811
rect 1964 31687 2472 31755
rect 1964 31631 2004 31687
rect 2060 31631 2128 31687
rect 2184 31631 2252 31687
rect 2308 31631 2376 31687
rect 2432 31631 2472 31687
rect 1964 31563 2472 31631
rect 1964 31507 2004 31563
rect 2060 31507 2128 31563
rect 2184 31507 2252 31563
rect 2308 31507 2376 31563
rect 2432 31507 2472 31563
rect 1964 31439 2472 31507
rect 1964 31383 2004 31439
rect 2060 31383 2128 31439
rect 2184 31383 2252 31439
rect 2308 31383 2376 31439
rect 2432 31383 2472 31439
rect 1964 31315 2472 31383
rect 1964 31259 2004 31315
rect 2060 31259 2128 31315
rect 2184 31259 2252 31315
rect 2308 31259 2376 31315
rect 2432 31259 2472 31315
rect 1964 31191 2472 31259
rect 1964 31135 2004 31191
rect 2060 31135 2128 31191
rect 2184 31135 2252 31191
rect 2308 31135 2376 31191
rect 2432 31135 2472 31191
rect 1964 31067 2472 31135
rect 1964 31011 2004 31067
rect 2060 31011 2128 31067
rect 2184 31011 2252 31067
rect 2308 31011 2376 31067
rect 2432 31011 2472 31067
rect 1964 30943 2472 31011
rect 1964 30887 2004 30943
rect 2060 30887 2128 30943
rect 2184 30887 2252 30943
rect 2308 30887 2376 30943
rect 2432 30887 2472 30943
rect 1964 30819 2472 30887
rect 1964 30763 2004 30819
rect 2060 30763 2128 30819
rect 2184 30763 2252 30819
rect 2308 30763 2376 30819
rect 2432 30763 2472 30819
rect 1964 30695 2472 30763
rect 1964 30639 2004 30695
rect 2060 30639 2128 30695
rect 2184 30639 2252 30695
rect 2308 30639 2376 30695
rect 2432 30639 2472 30695
rect 1964 30571 2472 30639
rect 1964 30515 2004 30571
rect 2060 30515 2128 30571
rect 2184 30515 2252 30571
rect 2308 30515 2376 30571
rect 2432 30515 2472 30571
rect 1964 30447 2472 30515
rect 1964 30391 2004 30447
rect 2060 30391 2128 30447
rect 2184 30391 2252 30447
rect 2308 30391 2376 30447
rect 2432 30391 2472 30447
rect 1964 30323 2472 30391
rect 1964 30267 2004 30323
rect 2060 30267 2128 30323
rect 2184 30267 2252 30323
rect 2308 30267 2376 30323
rect 2432 30267 2472 30323
rect 1964 30199 2472 30267
rect 1964 30143 2004 30199
rect 2060 30143 2128 30199
rect 2184 30143 2252 30199
rect 2308 30143 2376 30199
rect 2432 30143 2472 30199
rect 1964 29845 2472 30143
rect 1964 29789 2004 29845
rect 2060 29789 2128 29845
rect 2184 29789 2252 29845
rect 2308 29789 2376 29845
rect 2432 29789 2472 29845
rect 1964 29721 2472 29789
rect 1964 29665 2004 29721
rect 2060 29665 2128 29721
rect 2184 29665 2252 29721
rect 2308 29665 2376 29721
rect 2432 29665 2472 29721
rect 1964 29597 2472 29665
rect 1964 29541 2004 29597
rect 2060 29541 2128 29597
rect 2184 29541 2252 29597
rect 2308 29541 2376 29597
rect 2432 29541 2472 29597
rect 1964 29473 2472 29541
rect 1964 29417 2004 29473
rect 2060 29417 2128 29473
rect 2184 29417 2252 29473
rect 2308 29417 2376 29473
rect 2432 29417 2472 29473
rect 1964 29349 2472 29417
rect 1964 29293 2004 29349
rect 2060 29293 2128 29349
rect 2184 29293 2252 29349
rect 2308 29293 2376 29349
rect 2432 29293 2472 29349
rect 1964 29225 2472 29293
rect 1964 29169 2004 29225
rect 2060 29169 2128 29225
rect 2184 29169 2252 29225
rect 2308 29169 2376 29225
rect 2432 29169 2472 29225
rect 1964 29101 2472 29169
rect 1964 29045 2004 29101
rect 2060 29045 2128 29101
rect 2184 29045 2252 29101
rect 2308 29045 2376 29101
rect 2432 29045 2472 29101
rect 1964 28977 2472 29045
rect 1964 28921 2004 28977
rect 2060 28921 2128 28977
rect 2184 28921 2252 28977
rect 2308 28921 2376 28977
rect 2432 28921 2472 28977
rect 1964 28853 2472 28921
rect 1964 28797 2004 28853
rect 2060 28797 2128 28853
rect 2184 28797 2252 28853
rect 2308 28797 2376 28853
rect 2432 28797 2472 28853
rect 1964 28729 2472 28797
rect 1964 28673 2004 28729
rect 2060 28673 2128 28729
rect 2184 28673 2252 28729
rect 2308 28673 2376 28729
rect 2432 28673 2472 28729
rect 1964 28605 2472 28673
rect 1964 28549 2004 28605
rect 2060 28549 2128 28605
rect 2184 28549 2252 28605
rect 2308 28549 2376 28605
rect 2432 28549 2472 28605
rect 1964 26651 2472 28549
rect 1964 26595 2004 26651
rect 2060 26595 2128 26651
rect 2184 26595 2252 26651
rect 2308 26595 2376 26651
rect 2432 26595 2472 26651
rect 1964 26527 2472 26595
rect 1964 26471 2004 26527
rect 2060 26471 2128 26527
rect 2184 26471 2252 26527
rect 2308 26471 2376 26527
rect 2432 26471 2472 26527
rect 1964 26403 2472 26471
rect 1964 26347 2004 26403
rect 2060 26347 2128 26403
rect 2184 26347 2252 26403
rect 2308 26347 2376 26403
rect 2432 26347 2472 26403
rect 1964 26279 2472 26347
rect 1964 26223 2004 26279
rect 2060 26223 2128 26279
rect 2184 26223 2252 26279
rect 2308 26223 2376 26279
rect 2432 26223 2472 26279
rect 1964 26155 2472 26223
rect 1964 26099 2004 26155
rect 2060 26099 2128 26155
rect 2184 26099 2252 26155
rect 2308 26099 2376 26155
rect 2432 26099 2472 26155
rect 1964 26031 2472 26099
rect 1964 25975 2004 26031
rect 2060 25975 2128 26031
rect 2184 25975 2252 26031
rect 2308 25975 2376 26031
rect 2432 25975 2472 26031
rect 1964 25907 2472 25975
rect 1964 25851 2004 25907
rect 2060 25851 2128 25907
rect 2184 25851 2252 25907
rect 2308 25851 2376 25907
rect 2432 25851 2472 25907
rect 1964 25783 2472 25851
rect 1964 25727 2004 25783
rect 2060 25727 2128 25783
rect 2184 25727 2252 25783
rect 2308 25727 2376 25783
rect 2432 25727 2472 25783
rect 1964 25659 2472 25727
rect 1964 25603 2004 25659
rect 2060 25603 2128 25659
rect 2184 25603 2252 25659
rect 2308 25603 2376 25659
rect 2432 25603 2472 25659
rect 1964 25535 2472 25603
rect 1964 25479 2004 25535
rect 2060 25479 2128 25535
rect 2184 25479 2252 25535
rect 2308 25479 2376 25535
rect 2432 25479 2472 25535
rect 1964 25411 2472 25479
rect 1964 25355 2004 25411
rect 2060 25355 2128 25411
rect 2184 25355 2252 25411
rect 2308 25355 2376 25411
rect 2432 25355 2472 25411
rect 1964 25287 2472 25355
rect 1964 25231 2004 25287
rect 2060 25231 2128 25287
rect 2184 25231 2252 25287
rect 2308 25231 2376 25287
rect 2432 25231 2472 25287
rect 1964 25163 2472 25231
rect 1964 25107 2004 25163
rect 2060 25107 2128 25163
rect 2184 25107 2252 25163
rect 2308 25107 2376 25163
rect 2432 25107 2472 25163
rect 1964 25039 2472 25107
rect 1964 24983 2004 25039
rect 2060 24983 2128 25039
rect 2184 24983 2252 25039
rect 2308 24983 2376 25039
rect 2432 24983 2472 25039
rect 1964 24915 2472 24983
rect 1964 24859 2004 24915
rect 2060 24859 2128 24915
rect 2184 24859 2252 24915
rect 2308 24859 2376 24915
rect 2432 24859 2472 24915
rect 1964 24791 2472 24859
rect 1964 24735 2004 24791
rect 2060 24735 2128 24791
rect 2184 24735 2252 24791
rect 2308 24735 2376 24791
rect 2432 24735 2472 24791
rect 1964 24667 2472 24735
rect 1964 24611 2004 24667
rect 2060 24611 2128 24667
rect 2184 24611 2252 24667
rect 2308 24611 2376 24667
rect 2432 24611 2472 24667
rect 1964 24543 2472 24611
rect 1964 24487 2004 24543
rect 2060 24487 2128 24543
rect 2184 24487 2252 24543
rect 2308 24487 2376 24543
rect 2432 24487 2472 24543
rect 1964 24419 2472 24487
rect 1964 24363 2004 24419
rect 2060 24363 2128 24419
rect 2184 24363 2252 24419
rect 2308 24363 2376 24419
rect 2432 24363 2472 24419
rect 1964 24295 2472 24363
rect 1964 24239 2004 24295
rect 2060 24239 2128 24295
rect 2184 24239 2252 24295
rect 2308 24239 2376 24295
rect 2432 24239 2472 24295
rect 1964 24171 2472 24239
rect 1964 24115 2004 24171
rect 2060 24115 2128 24171
rect 2184 24115 2252 24171
rect 2308 24115 2376 24171
rect 2432 24115 2472 24171
rect 1964 24047 2472 24115
rect 1964 23991 2004 24047
rect 2060 23991 2128 24047
rect 2184 23991 2252 24047
rect 2308 23991 2376 24047
rect 2432 23991 2472 24047
rect 1964 23923 2472 23991
rect 1964 23867 2004 23923
rect 2060 23867 2128 23923
rect 2184 23867 2252 23923
rect 2308 23867 2376 23923
rect 2432 23867 2472 23923
rect 1964 23799 2472 23867
rect 1964 23743 2004 23799
rect 2060 23743 2128 23799
rect 2184 23743 2252 23799
rect 2308 23743 2376 23799
rect 2432 23743 2472 23799
rect 1964 23451 2472 23743
rect 1964 23395 2004 23451
rect 2060 23395 2128 23451
rect 2184 23395 2252 23451
rect 2308 23395 2376 23451
rect 2432 23395 2472 23451
rect 1964 23327 2472 23395
rect 1964 23271 2004 23327
rect 2060 23271 2128 23327
rect 2184 23271 2252 23327
rect 2308 23271 2376 23327
rect 2432 23271 2472 23327
rect 1964 23203 2472 23271
rect 1964 23147 2004 23203
rect 2060 23147 2128 23203
rect 2184 23147 2252 23203
rect 2308 23147 2376 23203
rect 2432 23147 2472 23203
rect 1964 23079 2472 23147
rect 1964 23023 2004 23079
rect 2060 23023 2128 23079
rect 2184 23023 2252 23079
rect 2308 23023 2376 23079
rect 2432 23023 2472 23079
rect 1964 22955 2472 23023
rect 1964 22899 2004 22955
rect 2060 22899 2128 22955
rect 2184 22899 2252 22955
rect 2308 22899 2376 22955
rect 2432 22899 2472 22955
rect 1964 22831 2472 22899
rect 1964 22775 2004 22831
rect 2060 22775 2128 22831
rect 2184 22775 2252 22831
rect 2308 22775 2376 22831
rect 2432 22775 2472 22831
rect 1964 22707 2472 22775
rect 1964 22651 2004 22707
rect 2060 22651 2128 22707
rect 2184 22651 2252 22707
rect 2308 22651 2376 22707
rect 2432 22651 2472 22707
rect 1964 22583 2472 22651
rect 1964 22527 2004 22583
rect 2060 22527 2128 22583
rect 2184 22527 2252 22583
rect 2308 22527 2376 22583
rect 2432 22527 2472 22583
rect 1964 22459 2472 22527
rect 1964 22403 2004 22459
rect 2060 22403 2128 22459
rect 2184 22403 2252 22459
rect 2308 22403 2376 22459
rect 2432 22403 2472 22459
rect 1964 22335 2472 22403
rect 1964 22279 2004 22335
rect 2060 22279 2128 22335
rect 2184 22279 2252 22335
rect 2308 22279 2376 22335
rect 2432 22279 2472 22335
rect 1964 22211 2472 22279
rect 1964 22155 2004 22211
rect 2060 22155 2128 22211
rect 2184 22155 2252 22211
rect 2308 22155 2376 22211
rect 2432 22155 2472 22211
rect 1964 22087 2472 22155
rect 1964 22031 2004 22087
rect 2060 22031 2128 22087
rect 2184 22031 2252 22087
rect 2308 22031 2376 22087
rect 2432 22031 2472 22087
rect 1964 21963 2472 22031
rect 1964 21907 2004 21963
rect 2060 21907 2128 21963
rect 2184 21907 2252 21963
rect 2308 21907 2376 21963
rect 2432 21907 2472 21963
rect 1964 21839 2472 21907
rect 1964 21783 2004 21839
rect 2060 21783 2128 21839
rect 2184 21783 2252 21839
rect 2308 21783 2376 21839
rect 2432 21783 2472 21839
rect 1964 21715 2472 21783
rect 1964 21659 2004 21715
rect 2060 21659 2128 21715
rect 2184 21659 2252 21715
rect 2308 21659 2376 21715
rect 2432 21659 2472 21715
rect 1964 21591 2472 21659
rect 1964 21535 2004 21591
rect 2060 21535 2128 21591
rect 2184 21535 2252 21591
rect 2308 21535 2376 21591
rect 2432 21535 2472 21591
rect 1964 21467 2472 21535
rect 1964 21411 2004 21467
rect 2060 21411 2128 21467
rect 2184 21411 2252 21467
rect 2308 21411 2376 21467
rect 2432 21411 2472 21467
rect 1964 21343 2472 21411
rect 1964 21287 2004 21343
rect 2060 21287 2128 21343
rect 2184 21287 2252 21343
rect 2308 21287 2376 21343
rect 2432 21287 2472 21343
rect 1964 21219 2472 21287
rect 1964 21163 2004 21219
rect 2060 21163 2128 21219
rect 2184 21163 2252 21219
rect 2308 21163 2376 21219
rect 2432 21163 2472 21219
rect 1964 21095 2472 21163
rect 1964 21039 2004 21095
rect 2060 21039 2128 21095
rect 2184 21039 2252 21095
rect 2308 21039 2376 21095
rect 2432 21039 2472 21095
rect 1964 20971 2472 21039
rect 1964 20915 2004 20971
rect 2060 20915 2128 20971
rect 2184 20915 2252 20971
rect 2308 20915 2376 20971
rect 2432 20915 2472 20971
rect 1964 20847 2472 20915
rect 1964 20791 2004 20847
rect 2060 20791 2128 20847
rect 2184 20791 2252 20847
rect 2308 20791 2376 20847
rect 2432 20791 2472 20847
rect 1964 20723 2472 20791
rect 1964 20667 2004 20723
rect 2060 20667 2128 20723
rect 2184 20667 2252 20723
rect 2308 20667 2376 20723
rect 2432 20667 2472 20723
rect 1964 20599 2472 20667
rect 1964 20543 2004 20599
rect 2060 20543 2128 20599
rect 2184 20543 2252 20599
rect 2308 20543 2376 20599
rect 2432 20543 2472 20599
rect 1964 20251 2472 20543
rect 1964 20195 2004 20251
rect 2060 20195 2128 20251
rect 2184 20195 2252 20251
rect 2308 20195 2376 20251
rect 2432 20195 2472 20251
rect 1964 20127 2472 20195
rect 1964 20071 2004 20127
rect 2060 20071 2128 20127
rect 2184 20071 2252 20127
rect 2308 20071 2376 20127
rect 2432 20071 2472 20127
rect 1964 20003 2472 20071
rect 1964 19947 2004 20003
rect 2060 19947 2128 20003
rect 2184 19947 2252 20003
rect 2308 19947 2376 20003
rect 2432 19947 2472 20003
rect 1964 19879 2472 19947
rect 1964 19823 2004 19879
rect 2060 19823 2128 19879
rect 2184 19823 2252 19879
rect 2308 19823 2376 19879
rect 2432 19823 2472 19879
rect 1964 19755 2472 19823
rect 1964 19699 2004 19755
rect 2060 19699 2128 19755
rect 2184 19699 2252 19755
rect 2308 19699 2376 19755
rect 2432 19699 2472 19755
rect 1964 19631 2472 19699
rect 1964 19575 2004 19631
rect 2060 19575 2128 19631
rect 2184 19575 2252 19631
rect 2308 19575 2376 19631
rect 2432 19575 2472 19631
rect 1964 19507 2472 19575
rect 1964 19451 2004 19507
rect 2060 19451 2128 19507
rect 2184 19451 2252 19507
rect 2308 19451 2376 19507
rect 2432 19451 2472 19507
rect 1964 19383 2472 19451
rect 1964 19327 2004 19383
rect 2060 19327 2128 19383
rect 2184 19327 2252 19383
rect 2308 19327 2376 19383
rect 2432 19327 2472 19383
rect 1964 19259 2472 19327
rect 1964 19203 2004 19259
rect 2060 19203 2128 19259
rect 2184 19203 2252 19259
rect 2308 19203 2376 19259
rect 2432 19203 2472 19259
rect 1964 19135 2472 19203
rect 1964 19079 2004 19135
rect 2060 19079 2128 19135
rect 2184 19079 2252 19135
rect 2308 19079 2376 19135
rect 2432 19079 2472 19135
rect 1964 19011 2472 19079
rect 1964 18955 2004 19011
rect 2060 18955 2128 19011
rect 2184 18955 2252 19011
rect 2308 18955 2376 19011
rect 2432 18955 2472 19011
rect 1964 18887 2472 18955
rect 1964 18831 2004 18887
rect 2060 18831 2128 18887
rect 2184 18831 2252 18887
rect 2308 18831 2376 18887
rect 2432 18831 2472 18887
rect 1964 18763 2472 18831
rect 1964 18707 2004 18763
rect 2060 18707 2128 18763
rect 2184 18707 2252 18763
rect 2308 18707 2376 18763
rect 2432 18707 2472 18763
rect 1964 18639 2472 18707
rect 1964 18583 2004 18639
rect 2060 18583 2128 18639
rect 2184 18583 2252 18639
rect 2308 18583 2376 18639
rect 2432 18583 2472 18639
rect 1964 18515 2472 18583
rect 1964 18459 2004 18515
rect 2060 18459 2128 18515
rect 2184 18459 2252 18515
rect 2308 18459 2376 18515
rect 2432 18459 2472 18515
rect 1964 18391 2472 18459
rect 1964 18335 2004 18391
rect 2060 18335 2128 18391
rect 2184 18335 2252 18391
rect 2308 18335 2376 18391
rect 2432 18335 2472 18391
rect 1964 18267 2472 18335
rect 1964 18211 2004 18267
rect 2060 18211 2128 18267
rect 2184 18211 2252 18267
rect 2308 18211 2376 18267
rect 2432 18211 2472 18267
rect 1964 18143 2472 18211
rect 1964 18087 2004 18143
rect 2060 18087 2128 18143
rect 2184 18087 2252 18143
rect 2308 18087 2376 18143
rect 2432 18087 2472 18143
rect 1964 18019 2472 18087
rect 1964 17963 2004 18019
rect 2060 17963 2128 18019
rect 2184 17963 2252 18019
rect 2308 17963 2376 18019
rect 2432 17963 2472 18019
rect 1964 17895 2472 17963
rect 1964 17839 2004 17895
rect 2060 17839 2128 17895
rect 2184 17839 2252 17895
rect 2308 17839 2376 17895
rect 2432 17839 2472 17895
rect 1964 17771 2472 17839
rect 1964 17715 2004 17771
rect 2060 17715 2128 17771
rect 2184 17715 2252 17771
rect 2308 17715 2376 17771
rect 2432 17715 2472 17771
rect 1964 17647 2472 17715
rect 1964 17591 2004 17647
rect 2060 17591 2128 17647
rect 2184 17591 2252 17647
rect 2308 17591 2376 17647
rect 2432 17591 2472 17647
rect 1964 17523 2472 17591
rect 1964 17467 2004 17523
rect 2060 17467 2128 17523
rect 2184 17467 2252 17523
rect 2308 17467 2376 17523
rect 2432 17467 2472 17523
rect 1964 17399 2472 17467
rect 1964 17343 2004 17399
rect 2060 17343 2128 17399
rect 2184 17343 2252 17399
rect 2308 17343 2376 17399
rect 2432 17343 2472 17399
rect 1964 17051 2472 17343
rect 1964 16995 2004 17051
rect 2060 16995 2128 17051
rect 2184 16995 2252 17051
rect 2308 16995 2376 17051
rect 2432 16995 2472 17051
rect 1964 16927 2472 16995
rect 1964 16871 2004 16927
rect 2060 16871 2128 16927
rect 2184 16871 2252 16927
rect 2308 16871 2376 16927
rect 2432 16871 2472 16927
rect 1964 16803 2472 16871
rect 1964 16747 2004 16803
rect 2060 16747 2128 16803
rect 2184 16747 2252 16803
rect 2308 16747 2376 16803
rect 2432 16747 2472 16803
rect 1964 16679 2472 16747
rect 1964 16623 2004 16679
rect 2060 16623 2128 16679
rect 2184 16623 2252 16679
rect 2308 16623 2376 16679
rect 2432 16623 2472 16679
rect 1964 16555 2472 16623
rect 1964 16499 2004 16555
rect 2060 16499 2128 16555
rect 2184 16499 2252 16555
rect 2308 16499 2376 16555
rect 2432 16499 2472 16555
rect 1964 16431 2472 16499
rect 1964 16375 2004 16431
rect 2060 16375 2128 16431
rect 2184 16375 2252 16431
rect 2308 16375 2376 16431
rect 2432 16375 2472 16431
rect 1964 16307 2472 16375
rect 1964 16251 2004 16307
rect 2060 16251 2128 16307
rect 2184 16251 2252 16307
rect 2308 16251 2376 16307
rect 2432 16251 2472 16307
rect 1964 16183 2472 16251
rect 1964 16127 2004 16183
rect 2060 16127 2128 16183
rect 2184 16127 2252 16183
rect 2308 16127 2376 16183
rect 2432 16127 2472 16183
rect 1964 16059 2472 16127
rect 1964 16003 2004 16059
rect 2060 16003 2128 16059
rect 2184 16003 2252 16059
rect 2308 16003 2376 16059
rect 2432 16003 2472 16059
rect 1964 15935 2472 16003
rect 1964 15879 2004 15935
rect 2060 15879 2128 15935
rect 2184 15879 2252 15935
rect 2308 15879 2376 15935
rect 2432 15879 2472 15935
rect 1964 15811 2472 15879
rect 1964 15762 2004 15811
rect 858 15687 1336 15755
rect 858 15631 868 15687
rect 924 15631 992 15687
rect 1048 15631 1116 15687
rect 1172 15631 1240 15687
rect 1296 15631 1336 15687
rect 858 15563 1336 15631
rect 858 15507 868 15563
rect 924 15507 992 15563
rect 1048 15507 1116 15563
rect 1172 15507 1240 15563
rect 1296 15507 1336 15563
rect 858 15439 1336 15507
rect 858 15383 868 15439
rect 924 15383 992 15439
rect 1048 15383 1116 15439
rect 1172 15383 1240 15439
rect 1296 15383 1336 15439
rect 858 15315 1336 15383
rect 858 15259 868 15315
rect 924 15259 992 15315
rect 1048 15259 1116 15315
rect 1172 15259 1240 15315
rect 1296 15259 1336 15315
rect 858 15191 1336 15259
rect 858 15135 868 15191
rect 924 15135 992 15191
rect 1048 15135 1116 15191
rect 1172 15135 1240 15191
rect 1296 15135 1336 15191
rect 858 15067 1336 15135
rect 858 15011 868 15067
rect 924 15011 992 15067
rect 1048 15011 1116 15067
rect 1172 15011 1240 15067
rect 1296 15011 1336 15067
rect 858 14943 1336 15011
rect 858 14887 868 14943
rect 924 14887 992 14943
rect 1048 14887 1116 14943
rect 1172 14887 1240 14943
rect 1296 14887 1336 14943
rect 858 14819 1336 14887
rect 858 14763 868 14819
rect 924 14763 992 14819
rect 1048 14763 1116 14819
rect 1172 14763 1240 14819
rect 1296 14763 1336 14819
rect 858 14695 1336 14763
rect 858 14639 868 14695
rect 924 14639 992 14695
rect 1048 14639 1116 14695
rect 1172 14639 1240 14695
rect 1296 14639 1336 14695
rect 858 14571 1336 14639
rect 858 14515 868 14571
rect 924 14515 992 14571
rect 1048 14515 1116 14571
rect 1172 14515 1240 14571
rect 1296 14515 1336 14571
rect 858 14447 1336 14515
rect 858 14391 868 14447
rect 924 14391 992 14447
rect 1048 14391 1116 14447
rect 1172 14391 1240 14447
rect 1296 14391 1336 14447
rect 858 14323 1336 14391
rect 858 14267 868 14323
rect 924 14267 992 14323
rect 1048 14267 1116 14323
rect 1172 14267 1240 14323
rect 1296 14267 1336 14323
rect 858 14199 1336 14267
rect 858 14143 868 14199
rect 924 14143 992 14199
rect 1048 14143 1116 14199
rect 1172 14143 1240 14199
rect 1296 14143 1336 14199
rect 858 14133 1336 14143
rect 1994 15755 2004 15762
rect 2060 15755 2128 15811
rect 2184 15755 2252 15811
rect 2308 15755 2376 15811
rect 2432 15762 2472 15811
rect 2532 56922 3040 56975
rect 2532 56866 2572 56922
rect 2628 56866 2696 56922
rect 2752 56866 2820 56922
rect 2876 56866 2944 56922
rect 3000 56866 3040 56922
rect 2532 56798 3040 56866
rect 2532 56742 2572 56798
rect 2628 56742 2696 56798
rect 2752 56742 2820 56798
rect 2876 56742 2944 56798
rect 3000 56742 3040 56798
rect 2532 56711 3040 56742
rect 2532 56659 2544 56711
rect 2596 56674 2652 56711
rect 2704 56674 2760 56711
rect 2628 56659 2652 56674
rect 2752 56659 2760 56674
rect 2812 56674 2868 56711
rect 2920 56674 2976 56711
rect 2812 56659 2820 56674
rect 2920 56659 2944 56674
rect 3028 56659 3040 56711
rect 2532 56618 2572 56659
rect 2628 56618 2696 56659
rect 2752 56618 2820 56659
rect 2876 56618 2944 56659
rect 3000 56618 3040 56659
rect 2532 56603 3040 56618
rect 2532 56551 2544 56603
rect 2596 56551 2652 56603
rect 2704 56551 2760 56603
rect 2812 56551 2868 56603
rect 2920 56551 2976 56603
rect 3028 56551 3040 56603
rect 2532 56550 3040 56551
rect 2532 56495 2572 56550
rect 2628 56495 2696 56550
rect 2752 56495 2820 56550
rect 2876 56495 2944 56550
rect 3000 56495 3040 56550
rect 2532 56443 2544 56495
rect 2628 56494 2652 56495
rect 2752 56494 2760 56495
rect 2596 56443 2652 56494
rect 2704 56443 2760 56494
rect 2812 56494 2820 56495
rect 2920 56494 2944 56495
rect 2812 56443 2868 56494
rect 2920 56443 2976 56494
rect 3028 56443 3040 56495
rect 2532 56426 3040 56443
rect 2532 56370 2572 56426
rect 2628 56370 2696 56426
rect 2752 56370 2820 56426
rect 2876 56370 2944 56426
rect 3000 56370 3040 56426
rect 2532 56302 3040 56370
rect 2532 56246 2572 56302
rect 2628 56246 2696 56302
rect 2752 56246 2820 56302
rect 2876 56246 2944 56302
rect 3000 56246 3040 56302
rect 2532 56178 3040 56246
rect 2532 56122 2572 56178
rect 2628 56122 2696 56178
rect 2752 56122 2820 56178
rect 2876 56122 2944 56178
rect 3000 56122 3040 56178
rect 2532 56054 3040 56122
rect 2532 55998 2572 56054
rect 2628 55998 2696 56054
rect 2752 55998 2820 56054
rect 2876 55998 2944 56054
rect 3000 55998 3040 56054
rect 2532 55930 3040 55998
rect 2532 55874 2572 55930
rect 2628 55874 2696 55930
rect 2752 55874 2820 55930
rect 2876 55874 2944 55930
rect 3000 55874 3040 55930
rect 2532 55806 3040 55874
rect 2532 55750 2572 55806
rect 2628 55750 2696 55806
rect 2752 55750 2820 55806
rect 2876 55750 2944 55806
rect 3000 55750 3040 55806
rect 2532 53845 3040 55750
rect 2532 53789 2572 53845
rect 2628 53789 2696 53845
rect 2752 53789 2820 53845
rect 2876 53789 2944 53845
rect 3000 53789 3040 53845
rect 2532 53721 3040 53789
rect 2532 53665 2572 53721
rect 2628 53665 2696 53721
rect 2752 53665 2820 53721
rect 2876 53665 2944 53721
rect 3000 53665 3040 53721
rect 2532 53597 3040 53665
rect 2532 53541 2572 53597
rect 2628 53541 2696 53597
rect 2752 53541 2820 53597
rect 2876 53541 2944 53597
rect 3000 53541 3040 53597
rect 2532 53473 3040 53541
rect 2532 53417 2572 53473
rect 2628 53417 2696 53473
rect 2752 53417 2820 53473
rect 2876 53417 2944 53473
rect 3000 53417 3040 53473
rect 2532 53349 3040 53417
rect 2532 53293 2572 53349
rect 2628 53293 2696 53349
rect 2752 53293 2820 53349
rect 2876 53293 2944 53349
rect 3000 53293 3040 53349
rect 2532 53225 3040 53293
rect 2532 53169 2572 53225
rect 2628 53169 2696 53225
rect 2752 53169 2820 53225
rect 2876 53169 2944 53225
rect 3000 53169 3040 53225
rect 2532 53101 3040 53169
rect 2532 53045 2572 53101
rect 2628 53045 2696 53101
rect 2752 53045 2820 53101
rect 2876 53045 2944 53101
rect 3000 53045 3040 53101
rect 2532 52996 2574 53045
rect 2626 52996 2698 53045
rect 2750 52996 2822 53045
rect 2874 52996 2946 53045
rect 2998 52996 3040 53045
rect 2532 52977 3040 52996
rect 2532 52921 2572 52977
rect 2628 52921 2696 52977
rect 2752 52921 2820 52977
rect 2876 52921 2944 52977
rect 3000 52921 3040 52977
rect 2532 52872 2574 52921
rect 2626 52872 2698 52921
rect 2750 52872 2822 52921
rect 2874 52872 2946 52921
rect 2998 52872 3040 52921
rect 2532 52853 3040 52872
rect 2532 52797 2572 52853
rect 2628 52797 2696 52853
rect 2752 52797 2820 52853
rect 2876 52797 2944 52853
rect 3000 52797 3040 52853
rect 2532 52748 2574 52797
rect 2626 52748 2698 52797
rect 2750 52748 2822 52797
rect 2874 52748 2946 52797
rect 2998 52748 3040 52797
rect 2532 52729 3040 52748
rect 2532 52673 2572 52729
rect 2628 52673 2696 52729
rect 2752 52673 2820 52729
rect 2876 52673 2944 52729
rect 3000 52673 3040 52729
rect 2532 52624 2574 52673
rect 2626 52624 2698 52673
rect 2750 52624 2822 52673
rect 2874 52624 2946 52673
rect 2998 52624 3040 52673
rect 2532 52605 3040 52624
rect 2532 52549 2572 52605
rect 2628 52549 2696 52605
rect 2752 52549 2820 52605
rect 2876 52549 2944 52605
rect 3000 52549 3040 52605
rect 2532 52500 2574 52549
rect 2626 52500 2698 52549
rect 2750 52500 2822 52549
rect 2874 52500 2946 52549
rect 2998 52500 3040 52549
rect 2532 49100 3040 52500
rect 2532 49048 2574 49100
rect 2626 49048 2698 49100
rect 2750 49048 2822 49100
rect 2874 49048 2946 49100
rect 2998 49048 3040 49100
rect 2532 49045 3040 49048
rect 2532 48989 2572 49045
rect 2628 48989 2696 49045
rect 2752 48989 2820 49045
rect 2876 48989 2944 49045
rect 3000 48989 3040 49045
rect 2532 48976 3040 48989
rect 2532 48924 2574 48976
rect 2626 48924 2698 48976
rect 2750 48924 2822 48976
rect 2874 48924 2946 48976
rect 2998 48924 3040 48976
rect 2532 48921 3040 48924
rect 2532 48865 2572 48921
rect 2628 48865 2696 48921
rect 2752 48865 2820 48921
rect 2876 48865 2944 48921
rect 3000 48865 3040 48921
rect 2532 48852 3040 48865
rect 2532 48800 2574 48852
rect 2626 48800 2698 48852
rect 2750 48800 2822 48852
rect 2874 48800 2946 48852
rect 2998 48800 3040 48852
rect 2532 48797 3040 48800
rect 2532 48741 2572 48797
rect 2628 48741 2696 48797
rect 2752 48741 2820 48797
rect 2876 48741 2944 48797
rect 3000 48741 3040 48797
rect 2532 48728 3040 48741
rect 2532 48676 2574 48728
rect 2626 48676 2698 48728
rect 2750 48676 2822 48728
rect 2874 48676 2946 48728
rect 2998 48676 3040 48728
rect 2532 48673 3040 48676
rect 2532 48617 2572 48673
rect 2628 48617 2696 48673
rect 2752 48617 2820 48673
rect 2876 48617 2944 48673
rect 3000 48617 3040 48673
rect 2532 48604 3040 48617
rect 2532 48552 2574 48604
rect 2626 48552 2698 48604
rect 2750 48552 2822 48604
rect 2874 48552 2946 48604
rect 2998 48552 3040 48604
rect 2532 48549 3040 48552
rect 2532 48493 2572 48549
rect 2628 48493 2696 48549
rect 2752 48493 2820 48549
rect 2876 48493 2944 48549
rect 3000 48493 3040 48549
rect 2532 48425 3040 48493
rect 2532 48369 2572 48425
rect 2628 48369 2696 48425
rect 2752 48369 2820 48425
rect 2876 48369 2944 48425
rect 3000 48369 3040 48425
rect 2532 48301 3040 48369
rect 2532 48245 2572 48301
rect 2628 48245 2696 48301
rect 2752 48245 2820 48301
rect 2876 48245 2944 48301
rect 3000 48245 3040 48301
rect 2532 48177 3040 48245
rect 2532 48121 2572 48177
rect 2628 48121 2696 48177
rect 2752 48121 2820 48177
rect 2876 48121 2944 48177
rect 3000 48121 3040 48177
rect 2532 48053 3040 48121
rect 2532 47997 2572 48053
rect 2628 47997 2696 48053
rect 2752 47997 2820 48053
rect 2876 47997 2944 48053
rect 3000 47997 3040 48053
rect 2532 47929 3040 47997
rect 2532 47873 2572 47929
rect 2628 47873 2696 47929
rect 2752 47873 2820 47929
rect 2876 47873 2944 47929
rect 3000 47873 3040 47929
rect 2532 47805 3040 47873
rect 2532 47749 2572 47805
rect 2628 47749 2696 47805
rect 2752 47749 2820 47805
rect 2876 47749 2944 47805
rect 3000 47749 3040 47805
rect 2532 45845 3040 47749
rect 2532 45789 2572 45845
rect 2628 45789 2696 45845
rect 2752 45789 2820 45845
rect 2876 45789 2944 45845
rect 3000 45789 3040 45845
rect 2532 45721 3040 45789
rect 2532 45665 2572 45721
rect 2628 45665 2696 45721
rect 2752 45665 2820 45721
rect 2876 45665 2944 45721
rect 3000 45665 3040 45721
rect 2532 45597 3040 45665
rect 2532 45541 2572 45597
rect 2628 45541 2696 45597
rect 2752 45541 2820 45597
rect 2876 45541 2944 45597
rect 3000 45541 3040 45597
rect 2532 45473 3040 45541
rect 2532 45417 2572 45473
rect 2628 45417 2696 45473
rect 2752 45417 2820 45473
rect 2876 45417 2944 45473
rect 3000 45417 3040 45473
rect 2532 45349 3040 45417
rect 2532 45293 2572 45349
rect 2628 45293 2696 45349
rect 2752 45293 2820 45349
rect 2876 45293 2944 45349
rect 3000 45293 3040 45349
rect 2532 45225 3040 45293
rect 2532 45169 2572 45225
rect 2628 45169 2696 45225
rect 2752 45169 2820 45225
rect 2876 45169 2944 45225
rect 3000 45169 3040 45225
rect 2532 45152 3040 45169
rect 2532 45101 2574 45152
rect 2626 45101 2698 45152
rect 2750 45101 2822 45152
rect 2874 45101 2946 45152
rect 2998 45101 3040 45152
rect 2532 45045 2572 45101
rect 2628 45045 2696 45101
rect 2752 45045 2820 45101
rect 2876 45045 2944 45101
rect 3000 45045 3040 45101
rect 2532 45028 3040 45045
rect 2532 44977 2574 45028
rect 2626 44977 2698 45028
rect 2750 44977 2822 45028
rect 2874 44977 2946 45028
rect 2998 44977 3040 45028
rect 2532 44921 2572 44977
rect 2628 44921 2696 44977
rect 2752 44921 2820 44977
rect 2876 44921 2944 44977
rect 3000 44921 3040 44977
rect 2532 44904 3040 44921
rect 2532 44853 2574 44904
rect 2626 44853 2698 44904
rect 2750 44853 2822 44904
rect 2874 44853 2946 44904
rect 2998 44853 3040 44904
rect 2532 44797 2572 44853
rect 2628 44797 2696 44853
rect 2752 44797 2820 44853
rect 2876 44797 2944 44853
rect 3000 44797 3040 44853
rect 2532 44780 3040 44797
rect 2532 44729 2574 44780
rect 2626 44729 2698 44780
rect 2750 44729 2822 44780
rect 2874 44729 2946 44780
rect 2998 44729 3040 44780
rect 2532 44673 2572 44729
rect 2628 44673 2696 44729
rect 2752 44673 2820 44729
rect 2876 44673 2944 44729
rect 3000 44673 3040 44729
rect 2532 44656 3040 44673
rect 2532 44605 2574 44656
rect 2626 44605 2698 44656
rect 2750 44605 2822 44656
rect 2874 44605 2946 44656
rect 2998 44605 3040 44656
rect 2532 44549 2572 44605
rect 2628 44549 2696 44605
rect 2752 44549 2820 44605
rect 2876 44549 2944 44605
rect 3000 44549 3040 44605
rect 2532 41204 3040 44549
rect 2532 41152 2574 41204
rect 2626 41152 2698 41204
rect 2750 41152 2822 41204
rect 2874 41152 2946 41204
rect 2998 41152 3040 41204
rect 2532 41080 3040 41152
rect 2532 41028 2574 41080
rect 2626 41028 2698 41080
rect 2750 41028 2822 41080
rect 2874 41028 2946 41080
rect 2998 41028 3040 41080
rect 2532 40956 3040 41028
rect 2532 40904 2574 40956
rect 2626 40904 2698 40956
rect 2750 40904 2822 40956
rect 2874 40904 2946 40956
rect 2998 40904 3040 40956
rect 2532 40832 3040 40904
rect 2532 40780 2574 40832
rect 2626 40780 2698 40832
rect 2750 40780 2822 40832
rect 2874 40780 2946 40832
rect 2998 40780 3040 40832
rect 2532 40708 3040 40780
rect 2532 40656 2574 40708
rect 2626 40656 2698 40708
rect 2750 40656 2822 40708
rect 2874 40656 2946 40708
rect 2998 40656 3040 40708
rect 2532 37256 3040 40656
rect 2532 37204 2574 37256
rect 2626 37204 2698 37256
rect 2750 37204 2822 37256
rect 2874 37204 2946 37256
rect 2998 37204 3040 37256
rect 2532 37132 3040 37204
rect 2532 37080 2574 37132
rect 2626 37080 2698 37132
rect 2750 37080 2822 37132
rect 2874 37080 2946 37132
rect 2998 37080 3040 37132
rect 2532 37008 3040 37080
rect 2532 36956 2574 37008
rect 2626 36956 2698 37008
rect 2750 36956 2822 37008
rect 2874 36956 2946 37008
rect 2998 36956 3040 37008
rect 2532 36884 3040 36956
rect 2532 36832 2574 36884
rect 2626 36832 2698 36884
rect 2750 36832 2822 36884
rect 2874 36832 2946 36884
rect 2998 36832 3040 36884
rect 2532 36760 3040 36832
rect 2532 36708 2574 36760
rect 2626 36708 2698 36760
rect 2750 36708 2822 36760
rect 2874 36708 2946 36760
rect 2998 36708 3040 36760
rect 2532 36251 3040 36708
rect 2532 36195 2572 36251
rect 2628 36195 2696 36251
rect 2752 36195 2820 36251
rect 2876 36195 2944 36251
rect 3000 36195 3040 36251
rect 2532 36127 3040 36195
rect 2532 36071 2572 36127
rect 2628 36071 2696 36127
rect 2752 36071 2820 36127
rect 2876 36071 2944 36127
rect 3000 36071 3040 36127
rect 2532 36003 3040 36071
rect 2532 35947 2572 36003
rect 2628 35947 2696 36003
rect 2752 35947 2820 36003
rect 2876 35947 2944 36003
rect 3000 35947 3040 36003
rect 2532 35879 3040 35947
rect 2532 35823 2572 35879
rect 2628 35823 2696 35879
rect 2752 35823 2820 35879
rect 2876 35823 2944 35879
rect 3000 35823 3040 35879
rect 2532 35755 3040 35823
rect 2532 35699 2572 35755
rect 2628 35699 2696 35755
rect 2752 35699 2820 35755
rect 2876 35699 2944 35755
rect 3000 35699 3040 35755
rect 2532 35631 3040 35699
rect 2532 35575 2572 35631
rect 2628 35575 2696 35631
rect 2752 35575 2820 35631
rect 2876 35575 2944 35631
rect 3000 35575 3040 35631
rect 2532 35507 3040 35575
rect 2532 35451 2572 35507
rect 2628 35451 2696 35507
rect 2752 35451 2820 35507
rect 2876 35451 2944 35507
rect 3000 35451 3040 35507
rect 2532 35383 3040 35451
rect 2532 35327 2572 35383
rect 2628 35327 2696 35383
rect 2752 35327 2820 35383
rect 2876 35327 2944 35383
rect 3000 35327 3040 35383
rect 2532 35259 3040 35327
rect 2532 35203 2572 35259
rect 2628 35203 2696 35259
rect 2752 35203 2820 35259
rect 2876 35203 2944 35259
rect 3000 35203 3040 35259
rect 2532 35135 3040 35203
rect 2532 35079 2572 35135
rect 2628 35079 2696 35135
rect 2752 35079 2820 35135
rect 2876 35079 2944 35135
rect 3000 35079 3040 35135
rect 2532 35011 3040 35079
rect 2532 34955 2572 35011
rect 2628 34955 2696 35011
rect 2752 34955 2820 35011
rect 2876 34955 2944 35011
rect 3000 34955 3040 35011
rect 2532 34887 3040 34955
rect 2532 34831 2572 34887
rect 2628 34831 2696 34887
rect 2752 34831 2820 34887
rect 2876 34831 2944 34887
rect 3000 34831 3040 34887
rect 2532 34763 3040 34831
rect 2532 34707 2572 34763
rect 2628 34707 2696 34763
rect 2752 34707 2820 34763
rect 2876 34707 2944 34763
rect 3000 34707 3040 34763
rect 2532 34639 3040 34707
rect 2532 34583 2572 34639
rect 2628 34583 2696 34639
rect 2752 34583 2820 34639
rect 2876 34583 2944 34639
rect 3000 34583 3040 34639
rect 2532 34515 3040 34583
rect 2532 34459 2572 34515
rect 2628 34459 2696 34515
rect 2752 34459 2820 34515
rect 2876 34459 2944 34515
rect 3000 34459 3040 34515
rect 2532 34391 3040 34459
rect 2532 34335 2572 34391
rect 2628 34335 2696 34391
rect 2752 34335 2820 34391
rect 2876 34335 2944 34391
rect 3000 34335 3040 34391
rect 2532 34267 3040 34335
rect 2532 34211 2572 34267
rect 2628 34211 2696 34267
rect 2752 34211 2820 34267
rect 2876 34211 2944 34267
rect 3000 34211 3040 34267
rect 2532 34143 3040 34211
rect 2532 34087 2572 34143
rect 2628 34087 2696 34143
rect 2752 34087 2820 34143
rect 2876 34087 2944 34143
rect 3000 34087 3040 34143
rect 2532 34019 3040 34087
rect 2532 33963 2572 34019
rect 2628 33963 2696 34019
rect 2752 33963 2820 34019
rect 2876 33963 2944 34019
rect 3000 33963 3040 34019
rect 2532 33895 3040 33963
rect 2532 33839 2572 33895
rect 2628 33839 2696 33895
rect 2752 33839 2820 33895
rect 2876 33839 2944 33895
rect 3000 33839 3040 33895
rect 2532 33771 3040 33839
rect 2532 33715 2572 33771
rect 2628 33715 2696 33771
rect 2752 33715 2820 33771
rect 2876 33715 2944 33771
rect 3000 33715 3040 33771
rect 2532 33647 3040 33715
rect 2532 33591 2572 33647
rect 2628 33591 2696 33647
rect 2752 33591 2820 33647
rect 2876 33591 2944 33647
rect 3000 33591 3040 33647
rect 2532 33523 3040 33591
rect 2532 33467 2572 33523
rect 2628 33467 2696 33523
rect 2752 33467 2820 33523
rect 2876 33467 2944 33523
rect 3000 33467 3040 33523
rect 2532 33399 3040 33467
rect 2532 33343 2572 33399
rect 2628 33343 2696 33399
rect 2752 33343 2820 33399
rect 2876 33343 2944 33399
rect 3000 33343 3040 33399
rect 2532 33308 3040 33343
rect 2532 33256 2574 33308
rect 2626 33256 2698 33308
rect 2750 33256 2822 33308
rect 2874 33256 2946 33308
rect 2998 33256 3040 33308
rect 2532 33184 3040 33256
rect 2532 33132 2574 33184
rect 2626 33132 2698 33184
rect 2750 33132 2822 33184
rect 2874 33132 2946 33184
rect 2998 33132 3040 33184
rect 2532 33060 3040 33132
rect 2532 33008 2574 33060
rect 2626 33008 2698 33060
rect 2750 33008 2822 33060
rect 2874 33008 2946 33060
rect 2998 33008 3040 33060
rect 2532 32936 3040 33008
rect 2532 32884 2574 32936
rect 2626 32884 2698 32936
rect 2750 32884 2822 32936
rect 2874 32884 2946 32936
rect 2998 32884 3040 32936
rect 2532 32812 3040 32884
rect 2532 32760 2574 32812
rect 2626 32760 2698 32812
rect 2750 32760 2822 32812
rect 2874 32760 2946 32812
rect 2998 32760 3040 32812
rect 2532 29360 3040 32760
rect 2532 29308 2574 29360
rect 2626 29308 2698 29360
rect 2750 29308 2822 29360
rect 2874 29308 2946 29360
rect 2998 29308 3040 29360
rect 2532 29236 3040 29308
rect 2532 29184 2574 29236
rect 2626 29184 2698 29236
rect 2750 29184 2822 29236
rect 2874 29184 2946 29236
rect 2998 29184 3040 29236
rect 2532 29112 3040 29184
rect 2532 29060 2574 29112
rect 2626 29060 2698 29112
rect 2750 29060 2822 29112
rect 2874 29060 2946 29112
rect 2998 29060 3040 29112
rect 2532 28988 3040 29060
rect 2532 28936 2574 28988
rect 2626 28936 2698 28988
rect 2750 28936 2822 28988
rect 2874 28936 2946 28988
rect 2998 28936 3040 28988
rect 2532 28864 3040 28936
rect 2532 28812 2574 28864
rect 2626 28812 2698 28864
rect 2750 28812 2822 28864
rect 2874 28812 2946 28864
rect 2998 28812 3040 28864
rect 2532 28245 3040 28812
rect 2532 28189 2572 28245
rect 2628 28189 2696 28245
rect 2752 28189 2820 28245
rect 2876 28189 2944 28245
rect 3000 28189 3040 28245
rect 2532 28121 3040 28189
rect 2532 28065 2572 28121
rect 2628 28065 2696 28121
rect 2752 28065 2820 28121
rect 2876 28065 2944 28121
rect 3000 28065 3040 28121
rect 2532 27997 3040 28065
rect 2532 27941 2572 27997
rect 2628 27941 2696 27997
rect 2752 27941 2820 27997
rect 2876 27941 2944 27997
rect 3000 27941 3040 27997
rect 2532 27873 3040 27941
rect 2532 27817 2572 27873
rect 2628 27817 2696 27873
rect 2752 27817 2820 27873
rect 2876 27817 2944 27873
rect 3000 27817 3040 27873
rect 2532 27749 3040 27817
rect 2532 27693 2572 27749
rect 2628 27693 2696 27749
rect 2752 27693 2820 27749
rect 2876 27693 2944 27749
rect 3000 27693 3040 27749
rect 2532 27625 3040 27693
rect 2532 27569 2572 27625
rect 2628 27569 2696 27625
rect 2752 27569 2820 27625
rect 2876 27569 2944 27625
rect 3000 27569 3040 27625
rect 2532 27501 3040 27569
rect 2532 27445 2572 27501
rect 2628 27445 2696 27501
rect 2752 27445 2820 27501
rect 2876 27445 2944 27501
rect 3000 27445 3040 27501
rect 2532 27377 3040 27445
rect 2532 27321 2572 27377
rect 2628 27321 2696 27377
rect 2752 27321 2820 27377
rect 2876 27321 2944 27377
rect 3000 27321 3040 27377
rect 2532 27253 3040 27321
rect 2532 27197 2572 27253
rect 2628 27197 2696 27253
rect 2752 27197 2820 27253
rect 2876 27197 2944 27253
rect 3000 27197 3040 27253
rect 2532 27129 3040 27197
rect 2532 27073 2572 27129
rect 2628 27073 2696 27129
rect 2752 27073 2820 27129
rect 2876 27073 2944 27129
rect 3000 27073 3040 27129
rect 2532 27005 3040 27073
rect 2532 26949 2572 27005
rect 2628 26949 2696 27005
rect 2752 26949 2820 27005
rect 2876 26949 2944 27005
rect 3000 26949 3040 27005
rect 2532 25412 3040 26949
rect 2532 25360 2574 25412
rect 2626 25360 2698 25412
rect 2750 25360 2822 25412
rect 2874 25360 2946 25412
rect 2998 25360 3040 25412
rect 2532 25288 3040 25360
rect 2532 25236 2574 25288
rect 2626 25236 2698 25288
rect 2750 25236 2822 25288
rect 2874 25236 2946 25288
rect 2998 25236 3040 25288
rect 2532 25164 3040 25236
rect 2532 25112 2574 25164
rect 2626 25112 2698 25164
rect 2750 25112 2822 25164
rect 2874 25112 2946 25164
rect 2998 25112 3040 25164
rect 2532 25040 3040 25112
rect 2532 24988 2574 25040
rect 2626 24988 2698 25040
rect 2750 24988 2822 25040
rect 2874 24988 2946 25040
rect 2998 24988 3040 25040
rect 2532 24916 3040 24988
rect 2532 24864 2574 24916
rect 2626 24864 2698 24916
rect 2750 24864 2822 24916
rect 2874 24864 2946 24916
rect 2998 24864 3040 24916
rect 2532 21469 3040 24864
rect 2532 21417 2544 21469
rect 2596 21417 2652 21469
rect 2704 21417 2760 21469
rect 2812 21417 2868 21469
rect 2920 21417 2976 21469
rect 3028 21417 3040 21469
rect 2532 21361 3040 21417
rect 2532 21309 2544 21361
rect 2596 21309 2652 21361
rect 2704 21309 2760 21361
rect 2812 21309 2868 21361
rect 2920 21309 2976 21361
rect 3028 21309 3040 21361
rect 2532 21253 3040 21309
rect 2532 21201 2544 21253
rect 2596 21201 2652 21253
rect 2704 21201 2760 21253
rect 2812 21201 2868 21253
rect 2920 21201 2976 21253
rect 3028 21201 3040 21253
rect 2532 15762 3040 21201
rect 3668 56286 4176 56975
rect 3668 56234 3729 56286
rect 3781 56234 4176 56286
rect 3668 56178 4176 56234
rect 3668 56126 3729 56178
rect 3781 56126 4176 56178
rect 3668 56070 4176 56126
rect 3668 56018 3729 56070
rect 3781 56018 4176 56070
rect 3668 55962 4176 56018
rect 3668 55910 3729 55962
rect 3781 55910 4176 55962
rect 3668 55854 4176 55910
rect 3668 55802 3729 55854
rect 3781 55802 4176 55854
rect 3668 55746 4176 55802
rect 3668 55694 3729 55746
rect 3781 55694 4176 55746
rect 3668 55638 4176 55694
rect 3668 55586 3729 55638
rect 3781 55586 4176 55638
rect 3668 55530 4176 55586
rect 3668 55478 3729 55530
rect 3781 55478 4176 55530
rect 3668 55445 4176 55478
rect 3668 55389 3708 55445
rect 3764 55422 3832 55445
rect 3781 55389 3832 55422
rect 3888 55389 3956 55445
rect 4012 55389 4080 55445
rect 4136 55389 4176 55445
rect 3668 55370 3729 55389
rect 3781 55370 4176 55389
rect 3668 55321 4176 55370
rect 3668 55265 3708 55321
rect 3764 55314 3832 55321
rect 3781 55265 3832 55314
rect 3888 55265 3956 55321
rect 4012 55265 4080 55321
rect 4136 55265 4176 55321
rect 3668 55262 3729 55265
rect 3781 55262 4176 55265
rect 3668 55206 4176 55262
rect 3668 55197 3729 55206
rect 3781 55197 4176 55206
rect 3668 55141 3708 55197
rect 3781 55154 3832 55197
rect 3764 55141 3832 55154
rect 3888 55141 3956 55197
rect 4012 55141 4080 55197
rect 4136 55141 4176 55197
rect 3668 55098 4176 55141
rect 3668 55073 3729 55098
rect 3781 55073 4176 55098
rect 3668 55017 3708 55073
rect 3781 55046 3832 55073
rect 3764 55017 3832 55046
rect 3888 55017 3956 55073
rect 4012 55017 4080 55073
rect 4136 55017 4176 55073
rect 3668 54990 4176 55017
rect 3668 54949 3729 54990
rect 3781 54949 4176 54990
rect 3668 54893 3708 54949
rect 3781 54938 3832 54949
rect 3764 54893 3832 54938
rect 3888 54893 3956 54949
rect 4012 54893 4080 54949
rect 4136 54893 4176 54949
rect 3668 54882 4176 54893
rect 3668 54830 3729 54882
rect 3781 54830 4176 54882
rect 3668 54825 4176 54830
rect 3668 54769 3708 54825
rect 3764 54774 3832 54825
rect 3781 54769 3832 54774
rect 3888 54769 3956 54825
rect 4012 54769 4080 54825
rect 4136 54769 4176 54825
rect 3668 54722 3729 54769
rect 3781 54722 4176 54769
rect 3668 54701 4176 54722
rect 3668 54645 3708 54701
rect 3764 54666 3832 54701
rect 3781 54645 3832 54666
rect 3888 54645 3956 54701
rect 4012 54645 4080 54701
rect 4136 54645 4176 54701
rect 3668 54614 3729 54645
rect 3781 54614 4176 54645
rect 3668 54577 4176 54614
rect 3668 54521 3708 54577
rect 3764 54558 3832 54577
rect 3781 54521 3832 54558
rect 3888 54521 3956 54577
rect 4012 54521 4080 54577
rect 4136 54521 4176 54577
rect 3668 54506 3729 54521
rect 3781 54506 4176 54521
rect 3668 54453 4176 54506
rect 3668 54397 3708 54453
rect 3764 54450 3832 54453
rect 3781 54398 3832 54450
rect 3764 54397 3832 54398
rect 3888 54397 3956 54453
rect 4012 54397 4080 54453
rect 4136 54397 4176 54453
rect 3668 54342 4176 54397
rect 3668 54329 3729 54342
rect 3781 54329 4176 54342
rect 3668 54273 3708 54329
rect 3781 54290 3832 54329
rect 3764 54273 3832 54290
rect 3888 54273 3956 54329
rect 4012 54273 4080 54329
rect 4136 54273 4176 54329
rect 3668 54234 4176 54273
rect 3668 54205 3729 54234
rect 3781 54205 4176 54234
rect 3668 54149 3708 54205
rect 3781 54182 3832 54205
rect 3764 54149 3832 54182
rect 3888 54149 3956 54205
rect 4012 54149 4080 54205
rect 4136 54149 4176 54205
rect 3668 54126 4176 54149
rect 3668 54074 3729 54126
rect 3781 54074 4176 54126
rect 3668 54018 4176 54074
rect 3668 53966 3729 54018
rect 3781 53966 4176 54018
rect 3668 53910 4176 53966
rect 3668 53858 3729 53910
rect 3781 53858 4176 53910
rect 3668 53802 4176 53858
rect 3668 53750 3729 53802
rect 3781 53750 4176 53802
rect 3668 53694 4176 53750
rect 3668 53642 3729 53694
rect 3781 53642 4176 53694
rect 3668 53586 4176 53642
rect 3668 53534 3729 53586
rect 3781 53534 4176 53586
rect 3668 53478 4176 53534
rect 3668 53426 3729 53478
rect 3781 53426 4176 53478
rect 3668 53370 4176 53426
rect 3668 53318 3729 53370
rect 3781 53318 4176 53370
rect 3668 53262 4176 53318
rect 3668 53210 3729 53262
rect 3781 53210 4176 53262
rect 3668 52338 4176 53210
rect 3668 52286 3729 52338
rect 3781 52286 4176 52338
rect 3668 52230 4176 52286
rect 3668 52178 3729 52230
rect 3781 52178 4176 52230
rect 3668 52122 4176 52178
rect 3668 52070 3729 52122
rect 3781 52070 4176 52122
rect 3668 52014 4176 52070
rect 3668 51962 3729 52014
rect 3781 51962 4176 52014
rect 3668 51906 4176 51962
rect 3668 51854 3729 51906
rect 3781 51854 4176 51906
rect 3668 51798 4176 51854
rect 3668 51746 3729 51798
rect 3781 51746 4176 51798
rect 3668 51690 4176 51746
rect 3668 51638 3729 51690
rect 3781 51638 4176 51690
rect 3668 51582 4176 51638
rect 3668 51530 3729 51582
rect 3781 51530 4176 51582
rect 3668 51474 4176 51530
rect 3668 51422 3729 51474
rect 3781 51422 4176 51474
rect 3668 51366 4176 51422
rect 3668 51314 3729 51366
rect 3781 51314 4176 51366
rect 3668 51258 4176 51314
rect 3668 51206 3729 51258
rect 3781 51206 4176 51258
rect 3668 51150 4176 51206
rect 3668 51098 3729 51150
rect 3781 51098 4176 51150
rect 3668 51042 4176 51098
rect 3668 50990 3729 51042
rect 3781 50990 4176 51042
rect 3668 50934 4176 50990
rect 3668 50882 3729 50934
rect 3781 50882 4176 50934
rect 3668 50826 4176 50882
rect 3668 50774 3729 50826
rect 3781 50774 4176 50826
rect 3668 50718 4176 50774
rect 3668 50666 3729 50718
rect 3781 50666 4176 50718
rect 3668 50610 4176 50666
rect 3668 50558 3729 50610
rect 3781 50558 4176 50610
rect 3668 50502 4176 50558
rect 3668 50450 3729 50502
rect 3781 50450 4176 50502
rect 3668 50394 4176 50450
rect 3668 50342 3729 50394
rect 3781 50342 4176 50394
rect 3668 50286 4176 50342
rect 3668 50234 3729 50286
rect 3781 50234 4176 50286
rect 3668 50178 4176 50234
rect 3668 50126 3729 50178
rect 3781 50126 4176 50178
rect 3668 50070 4176 50126
rect 3668 50018 3729 50070
rect 3781 50018 4176 50070
rect 3668 49962 4176 50018
rect 3668 49910 3729 49962
rect 3781 49910 4176 49962
rect 3668 49854 4176 49910
rect 3668 49802 3729 49854
rect 3781 49802 4176 49854
rect 3668 49746 4176 49802
rect 3668 49694 3729 49746
rect 3781 49694 4176 49746
rect 3668 49638 4176 49694
rect 3668 49586 3729 49638
rect 3781 49586 4176 49638
rect 3668 49530 4176 49586
rect 3668 49478 3729 49530
rect 3781 49478 4176 49530
rect 3668 49422 4176 49478
rect 3668 49370 3729 49422
rect 3781 49370 4176 49422
rect 3668 49314 4176 49370
rect 3668 49262 3729 49314
rect 3781 49262 4176 49314
rect 3668 48390 4176 49262
rect 3668 48338 3729 48390
rect 3781 48338 4176 48390
rect 3668 48282 4176 48338
rect 3668 48230 3729 48282
rect 3781 48230 4176 48282
rect 3668 48174 4176 48230
rect 3668 48122 3729 48174
rect 3781 48122 4176 48174
rect 3668 48066 4176 48122
rect 3668 48014 3729 48066
rect 3781 48014 4176 48066
rect 3668 47958 4176 48014
rect 3668 47906 3729 47958
rect 3781 47906 4176 47958
rect 3668 47850 4176 47906
rect 3668 47798 3729 47850
rect 3781 47798 4176 47850
rect 3668 47742 4176 47798
rect 3668 47690 3729 47742
rect 3781 47690 4176 47742
rect 3668 47634 4176 47690
rect 3668 47582 3729 47634
rect 3781 47582 4176 47634
rect 3668 47526 4176 47582
rect 3668 47474 3729 47526
rect 3781 47474 4176 47526
rect 3668 47445 4176 47474
rect 3668 47389 3708 47445
rect 3764 47418 3832 47445
rect 3781 47389 3832 47418
rect 3888 47389 3956 47445
rect 4012 47389 4080 47445
rect 4136 47389 4176 47445
rect 3668 47366 3729 47389
rect 3781 47366 4176 47389
rect 3668 47321 4176 47366
rect 3668 47265 3708 47321
rect 3764 47310 3832 47321
rect 3781 47265 3832 47310
rect 3888 47265 3956 47321
rect 4012 47265 4080 47321
rect 4136 47265 4176 47321
rect 3668 47258 3729 47265
rect 3781 47258 4176 47265
rect 3668 47202 4176 47258
rect 3668 47197 3729 47202
rect 3781 47197 4176 47202
rect 3668 47141 3708 47197
rect 3781 47150 3832 47197
rect 3764 47141 3832 47150
rect 3888 47141 3956 47197
rect 4012 47141 4080 47197
rect 4136 47141 4176 47197
rect 3668 47094 4176 47141
rect 3668 47073 3729 47094
rect 3781 47073 4176 47094
rect 3668 47017 3708 47073
rect 3781 47042 3832 47073
rect 3764 47017 3832 47042
rect 3888 47017 3956 47073
rect 4012 47017 4080 47073
rect 4136 47017 4176 47073
rect 3668 46986 4176 47017
rect 3668 46949 3729 46986
rect 3781 46949 4176 46986
rect 3668 46893 3708 46949
rect 3781 46934 3832 46949
rect 3764 46893 3832 46934
rect 3888 46893 3956 46949
rect 4012 46893 4080 46949
rect 4136 46893 4176 46949
rect 3668 46878 4176 46893
rect 3668 46826 3729 46878
rect 3781 46826 4176 46878
rect 3668 46825 4176 46826
rect 3668 46769 3708 46825
rect 3764 46770 3832 46825
rect 3781 46769 3832 46770
rect 3888 46769 3956 46825
rect 4012 46769 4080 46825
rect 4136 46769 4176 46825
rect 3668 46718 3729 46769
rect 3781 46718 4176 46769
rect 3668 46701 4176 46718
rect 3668 46645 3708 46701
rect 3764 46662 3832 46701
rect 3781 46645 3832 46662
rect 3888 46645 3956 46701
rect 4012 46645 4080 46701
rect 4136 46645 4176 46701
rect 3668 46610 3729 46645
rect 3781 46610 4176 46645
rect 3668 46577 4176 46610
rect 3668 46521 3708 46577
rect 3764 46554 3832 46577
rect 3781 46521 3832 46554
rect 3888 46521 3956 46577
rect 4012 46521 4080 46577
rect 4136 46521 4176 46577
rect 3668 46502 3729 46521
rect 3781 46502 4176 46521
rect 3668 46453 4176 46502
rect 3668 46397 3708 46453
rect 3764 46446 3832 46453
rect 3781 46397 3832 46446
rect 3888 46397 3956 46453
rect 4012 46397 4080 46453
rect 4136 46397 4176 46453
rect 3668 46394 3729 46397
rect 3781 46394 4176 46397
rect 3668 46338 4176 46394
rect 3668 46329 3729 46338
rect 3781 46329 4176 46338
rect 3668 46273 3708 46329
rect 3781 46286 3832 46329
rect 3764 46273 3832 46286
rect 3888 46273 3956 46329
rect 4012 46273 4080 46329
rect 4136 46273 4176 46329
rect 3668 46230 4176 46273
rect 3668 46205 3729 46230
rect 3781 46205 4176 46230
rect 3668 46149 3708 46205
rect 3781 46178 3832 46205
rect 3764 46149 3832 46178
rect 3888 46149 3956 46205
rect 4012 46149 4080 46205
rect 4136 46149 4176 46205
rect 3668 46122 4176 46149
rect 3668 46070 3729 46122
rect 3781 46070 4176 46122
rect 3668 46014 4176 46070
rect 3668 45962 3729 46014
rect 3781 45962 4176 46014
rect 3668 45906 4176 45962
rect 3668 45854 3729 45906
rect 3781 45854 4176 45906
rect 3668 45798 4176 45854
rect 3668 45746 3729 45798
rect 3781 45746 4176 45798
rect 3668 45690 4176 45746
rect 3668 45638 3729 45690
rect 3781 45638 4176 45690
rect 3668 45582 4176 45638
rect 3668 45530 3729 45582
rect 3781 45530 4176 45582
rect 3668 45474 4176 45530
rect 3668 45422 3729 45474
rect 3781 45422 4176 45474
rect 3668 45366 4176 45422
rect 3668 45314 3729 45366
rect 3781 45314 4176 45366
rect 3668 44442 4176 45314
rect 3668 44390 3729 44442
rect 3781 44390 4176 44442
rect 3668 44334 4176 44390
rect 3668 44282 3729 44334
rect 3781 44282 4176 44334
rect 3668 44245 4176 44282
rect 3668 44189 3708 44245
rect 3764 44226 3832 44245
rect 3781 44189 3832 44226
rect 3888 44189 3956 44245
rect 4012 44189 4080 44245
rect 4136 44189 4176 44245
rect 3668 44174 3729 44189
rect 3781 44174 4176 44189
rect 3668 44121 4176 44174
rect 3668 44065 3708 44121
rect 3764 44118 3832 44121
rect 3781 44066 3832 44118
rect 3764 44065 3832 44066
rect 3888 44065 3956 44121
rect 4012 44065 4080 44121
rect 4136 44065 4176 44121
rect 3668 44010 4176 44065
rect 3668 43997 3729 44010
rect 3781 43997 4176 44010
rect 3668 43941 3708 43997
rect 3781 43958 3832 43997
rect 3764 43941 3832 43958
rect 3888 43941 3956 43997
rect 4012 43941 4080 43997
rect 4136 43941 4176 43997
rect 3668 43902 4176 43941
rect 3668 43873 3729 43902
rect 3781 43873 4176 43902
rect 3668 43817 3708 43873
rect 3781 43850 3832 43873
rect 3764 43817 3832 43850
rect 3888 43817 3956 43873
rect 4012 43817 4080 43873
rect 4136 43817 4176 43873
rect 3668 43794 4176 43817
rect 3668 43749 3729 43794
rect 3781 43749 4176 43794
rect 3668 43693 3708 43749
rect 3781 43742 3832 43749
rect 3764 43693 3832 43742
rect 3888 43693 3956 43749
rect 4012 43693 4080 43749
rect 4136 43693 4176 43749
rect 3668 43686 4176 43693
rect 3668 43634 3729 43686
rect 3781 43634 4176 43686
rect 3668 43625 4176 43634
rect 3668 43569 3708 43625
rect 3764 43578 3832 43625
rect 3781 43569 3832 43578
rect 3888 43569 3956 43625
rect 4012 43569 4080 43625
rect 4136 43569 4176 43625
rect 3668 43526 3729 43569
rect 3781 43526 4176 43569
rect 3668 43501 4176 43526
rect 3668 43445 3708 43501
rect 3764 43470 3832 43501
rect 3781 43445 3832 43470
rect 3888 43445 3956 43501
rect 4012 43445 4080 43501
rect 4136 43445 4176 43501
rect 3668 43418 3729 43445
rect 3781 43418 4176 43445
rect 3668 43377 4176 43418
rect 3668 43321 3708 43377
rect 3764 43362 3832 43377
rect 3781 43321 3832 43362
rect 3888 43321 3956 43377
rect 4012 43321 4080 43377
rect 4136 43321 4176 43377
rect 3668 43310 3729 43321
rect 3781 43310 4176 43321
rect 3668 43254 4176 43310
rect 3668 43253 3729 43254
rect 3781 43253 4176 43254
rect 3668 43197 3708 43253
rect 3781 43202 3832 43253
rect 3764 43197 3832 43202
rect 3888 43197 3956 43253
rect 4012 43197 4080 43253
rect 4136 43197 4176 43253
rect 3668 43146 4176 43197
rect 3668 43129 3729 43146
rect 3781 43129 4176 43146
rect 3668 43073 3708 43129
rect 3781 43094 3832 43129
rect 3764 43073 3832 43094
rect 3888 43073 3956 43129
rect 4012 43073 4080 43129
rect 4136 43073 4176 43129
rect 3668 43038 4176 43073
rect 3668 43005 3729 43038
rect 3781 43005 4176 43038
rect 3668 42949 3708 43005
rect 3781 42986 3832 43005
rect 3764 42949 3832 42986
rect 3888 42949 3956 43005
rect 4012 42949 4080 43005
rect 4136 42949 4176 43005
rect 3668 42930 4176 42949
rect 3668 42878 3729 42930
rect 3781 42878 4176 42930
rect 3668 42822 4176 42878
rect 3668 42770 3729 42822
rect 3781 42770 4176 42822
rect 3668 42714 4176 42770
rect 3668 42662 3729 42714
rect 3781 42662 4176 42714
rect 3668 42645 4176 42662
rect 3668 42589 3708 42645
rect 3764 42606 3832 42645
rect 3781 42589 3832 42606
rect 3888 42589 3956 42645
rect 4012 42589 4080 42645
rect 4136 42589 4176 42645
rect 3668 42554 3729 42589
rect 3781 42554 4176 42589
rect 3668 42521 4176 42554
rect 3668 42465 3708 42521
rect 3764 42498 3832 42521
rect 3781 42465 3832 42498
rect 3888 42465 3956 42521
rect 4012 42465 4080 42521
rect 4136 42465 4176 42521
rect 3668 42446 3729 42465
rect 3781 42446 4176 42465
rect 3668 42397 4176 42446
rect 3668 42341 3708 42397
rect 3764 42390 3832 42397
rect 3781 42341 3832 42390
rect 3888 42341 3956 42397
rect 4012 42341 4080 42397
rect 4136 42341 4176 42397
rect 3668 42338 3729 42341
rect 3781 42338 4176 42341
rect 3668 42282 4176 42338
rect 3668 42273 3729 42282
rect 3781 42273 4176 42282
rect 3668 42217 3708 42273
rect 3781 42230 3832 42273
rect 3764 42217 3832 42230
rect 3888 42217 3956 42273
rect 4012 42217 4080 42273
rect 4136 42217 4176 42273
rect 3668 42174 4176 42217
rect 3668 42149 3729 42174
rect 3781 42149 4176 42174
rect 3668 42093 3708 42149
rect 3781 42122 3832 42149
rect 3764 42093 3832 42122
rect 3888 42093 3956 42149
rect 4012 42093 4080 42149
rect 4136 42093 4176 42149
rect 3668 42066 4176 42093
rect 3668 42025 3729 42066
rect 3781 42025 4176 42066
rect 3668 41969 3708 42025
rect 3781 42014 3832 42025
rect 3764 41969 3832 42014
rect 3888 41969 3956 42025
rect 4012 41969 4080 42025
rect 4136 41969 4176 42025
rect 3668 41958 4176 41969
rect 3668 41906 3729 41958
rect 3781 41906 4176 41958
rect 3668 41901 4176 41906
rect 3668 41845 3708 41901
rect 3764 41850 3832 41901
rect 3781 41845 3832 41850
rect 3888 41845 3956 41901
rect 4012 41845 4080 41901
rect 4136 41845 4176 41901
rect 3668 41798 3729 41845
rect 3781 41798 4176 41845
rect 3668 41777 4176 41798
rect 3668 41721 3708 41777
rect 3764 41742 3832 41777
rect 3781 41721 3832 41742
rect 3888 41721 3956 41777
rect 4012 41721 4080 41777
rect 4136 41721 4176 41777
rect 3668 41690 3729 41721
rect 3781 41690 4176 41721
rect 3668 41653 4176 41690
rect 3668 41597 3708 41653
rect 3764 41634 3832 41653
rect 3781 41597 3832 41634
rect 3888 41597 3956 41653
rect 4012 41597 4080 41653
rect 4136 41597 4176 41653
rect 3668 41582 3729 41597
rect 3781 41582 4176 41597
rect 3668 41529 4176 41582
rect 3668 41473 3708 41529
rect 3764 41526 3832 41529
rect 3781 41474 3832 41526
rect 3764 41473 3832 41474
rect 3888 41473 3956 41529
rect 4012 41473 4080 41529
rect 4136 41473 4176 41529
rect 3668 41418 4176 41473
rect 3668 41405 3729 41418
rect 3781 41405 4176 41418
rect 3668 41349 3708 41405
rect 3781 41366 3832 41405
rect 3764 41349 3832 41366
rect 3888 41349 3956 41405
rect 4012 41349 4080 41405
rect 4136 41349 4176 41405
rect 3668 41045 4176 41349
rect 3668 40989 3708 41045
rect 3764 40989 3832 41045
rect 3888 40989 3956 41045
rect 4012 40989 4080 41045
rect 4136 40989 4176 41045
rect 3668 40921 4176 40989
rect 3668 40865 3708 40921
rect 3764 40865 3832 40921
rect 3888 40865 3956 40921
rect 4012 40865 4080 40921
rect 4136 40865 4176 40921
rect 3668 40797 4176 40865
rect 3668 40741 3708 40797
rect 3764 40741 3832 40797
rect 3888 40741 3956 40797
rect 4012 40741 4080 40797
rect 4136 40741 4176 40797
rect 3668 40673 4176 40741
rect 3668 40617 3708 40673
rect 3764 40617 3832 40673
rect 3888 40617 3956 40673
rect 4012 40617 4080 40673
rect 4136 40617 4176 40673
rect 3668 40549 4176 40617
rect 3668 40493 3708 40549
rect 3764 40494 3832 40549
rect 3781 40493 3832 40494
rect 3888 40493 3956 40549
rect 4012 40493 4080 40549
rect 4136 40493 4176 40549
rect 3668 40442 3729 40493
rect 3781 40442 4176 40493
rect 3668 40425 4176 40442
rect 3668 40369 3708 40425
rect 3764 40386 3832 40425
rect 3781 40369 3832 40386
rect 3888 40369 3956 40425
rect 4012 40369 4080 40425
rect 4136 40369 4176 40425
rect 3668 40334 3729 40369
rect 3781 40334 4176 40369
rect 3668 40301 4176 40334
rect 3668 40245 3708 40301
rect 3764 40278 3832 40301
rect 3781 40245 3832 40278
rect 3888 40245 3956 40301
rect 4012 40245 4080 40301
rect 4136 40245 4176 40301
rect 3668 40226 3729 40245
rect 3781 40226 4176 40245
rect 3668 40177 4176 40226
rect 3668 40121 3708 40177
rect 3764 40170 3832 40177
rect 3781 40121 3832 40170
rect 3888 40121 3956 40177
rect 4012 40121 4080 40177
rect 4136 40121 4176 40177
rect 3668 40118 3729 40121
rect 3781 40118 4176 40121
rect 3668 40062 4176 40118
rect 3668 40053 3729 40062
rect 3781 40053 4176 40062
rect 3668 39997 3708 40053
rect 3781 40010 3832 40053
rect 3764 39997 3832 40010
rect 3888 39997 3956 40053
rect 4012 39997 4080 40053
rect 4136 39997 4176 40053
rect 3668 39954 4176 39997
rect 3668 39929 3729 39954
rect 3781 39929 4176 39954
rect 3668 39873 3708 39929
rect 3781 39902 3832 39929
rect 3764 39873 3832 39902
rect 3888 39873 3956 39929
rect 4012 39873 4080 39929
rect 4136 39873 4176 39929
rect 3668 39846 4176 39873
rect 3668 39805 3729 39846
rect 3781 39805 4176 39846
rect 3668 39749 3708 39805
rect 3781 39794 3832 39805
rect 3764 39749 3832 39794
rect 3888 39749 3956 39805
rect 4012 39749 4080 39805
rect 4136 39749 4176 39805
rect 3668 39738 4176 39749
rect 3668 39686 3729 39738
rect 3781 39686 4176 39738
rect 3668 39630 4176 39686
rect 3668 39578 3729 39630
rect 3781 39578 4176 39630
rect 3668 39522 4176 39578
rect 3668 39470 3729 39522
rect 3781 39470 4176 39522
rect 3668 39414 4176 39470
rect 3668 39362 3729 39414
rect 3781 39362 4176 39414
rect 3668 39306 4176 39362
rect 3668 39254 3729 39306
rect 3781 39254 4176 39306
rect 3668 39198 4176 39254
rect 3668 39146 3729 39198
rect 3781 39146 4176 39198
rect 3668 39090 4176 39146
rect 3668 39038 3729 39090
rect 3781 39038 4176 39090
rect 3668 38982 4176 39038
rect 3668 38930 3729 38982
rect 3781 38930 4176 38982
rect 3668 38874 4176 38930
rect 3668 38822 3729 38874
rect 3781 38822 4176 38874
rect 3668 38766 4176 38822
rect 3668 38714 3729 38766
rect 3781 38714 4176 38766
rect 3668 38658 4176 38714
rect 3668 38606 3729 38658
rect 3781 38606 4176 38658
rect 3668 38550 4176 38606
rect 3668 38498 3729 38550
rect 3781 38498 4176 38550
rect 3668 38442 4176 38498
rect 3668 38390 3729 38442
rect 3781 38390 4176 38442
rect 3668 38334 4176 38390
rect 3668 38282 3729 38334
rect 3781 38282 4176 38334
rect 3668 38226 4176 38282
rect 3668 38174 3729 38226
rect 3781 38174 4176 38226
rect 3668 38118 4176 38174
rect 3668 38066 3729 38118
rect 3781 38066 4176 38118
rect 3668 38010 4176 38066
rect 3668 37958 3729 38010
rect 3781 37958 4176 38010
rect 3668 37902 4176 37958
rect 3668 37850 3729 37902
rect 3781 37850 4176 37902
rect 3668 37794 4176 37850
rect 3668 37742 3729 37794
rect 3781 37742 4176 37794
rect 3668 37686 4176 37742
rect 3668 37634 3729 37686
rect 3781 37634 4176 37686
rect 3668 37578 4176 37634
rect 3668 37526 3729 37578
rect 3781 37526 4176 37578
rect 3668 37470 4176 37526
rect 3668 37418 3729 37470
rect 3781 37418 4176 37470
rect 3668 36546 4176 37418
rect 3668 36494 3729 36546
rect 3781 36494 4176 36546
rect 3668 36438 4176 36494
rect 3668 36386 3729 36438
rect 3781 36386 4176 36438
rect 3668 36330 4176 36386
rect 3668 36278 3729 36330
rect 3781 36278 4176 36330
rect 3668 36222 4176 36278
rect 3668 36170 3729 36222
rect 3781 36170 4176 36222
rect 3668 36114 4176 36170
rect 3668 36062 3729 36114
rect 3781 36062 4176 36114
rect 3668 36006 4176 36062
rect 3668 35954 3729 36006
rect 3781 35954 4176 36006
rect 3668 35898 4176 35954
rect 3668 35846 3729 35898
rect 3781 35846 4176 35898
rect 3668 35790 4176 35846
rect 3668 35738 3729 35790
rect 3781 35738 4176 35790
rect 3668 35682 4176 35738
rect 3668 35630 3729 35682
rect 3781 35630 4176 35682
rect 3668 35574 4176 35630
rect 3668 35522 3729 35574
rect 3781 35522 4176 35574
rect 3668 35466 4176 35522
rect 3668 35414 3729 35466
rect 3781 35414 4176 35466
rect 3668 35358 4176 35414
rect 3668 35306 3729 35358
rect 3781 35306 4176 35358
rect 3668 35250 4176 35306
rect 3668 35198 3729 35250
rect 3781 35198 4176 35250
rect 3668 35142 4176 35198
rect 3668 35090 3729 35142
rect 3781 35090 4176 35142
rect 3668 35034 4176 35090
rect 3668 34982 3729 35034
rect 3781 34982 4176 35034
rect 3668 34926 4176 34982
rect 3668 34874 3729 34926
rect 3781 34874 4176 34926
rect 3668 34818 4176 34874
rect 3668 34766 3729 34818
rect 3781 34766 4176 34818
rect 3668 34710 4176 34766
rect 3668 34658 3729 34710
rect 3781 34658 4176 34710
rect 3668 34602 4176 34658
rect 3668 34550 3729 34602
rect 3781 34550 4176 34602
rect 3668 34494 4176 34550
rect 3668 34442 3729 34494
rect 3781 34442 4176 34494
rect 3668 34386 4176 34442
rect 3668 34334 3729 34386
rect 3781 34334 4176 34386
rect 3668 34278 4176 34334
rect 3668 34226 3729 34278
rect 3781 34226 4176 34278
rect 3668 34170 4176 34226
rect 3668 34118 3729 34170
rect 3781 34118 4176 34170
rect 3668 34062 4176 34118
rect 3668 34010 3729 34062
rect 3781 34010 4176 34062
rect 3668 33954 4176 34010
rect 3668 33902 3729 33954
rect 3781 33902 4176 33954
rect 3668 33846 4176 33902
rect 3668 33794 3729 33846
rect 3781 33794 4176 33846
rect 3668 33738 4176 33794
rect 3668 33686 3729 33738
rect 3781 33686 4176 33738
rect 3668 33630 4176 33686
rect 3668 33578 3729 33630
rect 3781 33578 4176 33630
rect 3668 33522 4176 33578
rect 3668 33470 3729 33522
rect 3781 33470 4176 33522
rect 3668 33051 4176 33470
rect 3668 32995 3708 33051
rect 3764 32995 3832 33051
rect 3888 32995 3956 33051
rect 4012 32995 4080 33051
rect 4136 32995 4176 33051
rect 3668 32927 4176 32995
rect 3668 32871 3708 32927
rect 3764 32871 3832 32927
rect 3888 32871 3956 32927
rect 4012 32871 4080 32927
rect 4136 32871 4176 32927
rect 3668 32803 4176 32871
rect 3668 32747 3708 32803
rect 3764 32747 3832 32803
rect 3888 32747 3956 32803
rect 4012 32747 4080 32803
rect 4136 32747 4176 32803
rect 3668 32679 4176 32747
rect 3668 32623 3708 32679
rect 3764 32623 3832 32679
rect 3888 32623 3956 32679
rect 4012 32623 4080 32679
rect 4136 32623 4176 32679
rect 3668 32598 4176 32623
rect 3668 32555 3729 32598
rect 3781 32555 4176 32598
rect 3668 32499 3708 32555
rect 3781 32546 3832 32555
rect 3764 32499 3832 32546
rect 3888 32499 3956 32555
rect 4012 32499 4080 32555
rect 4136 32499 4176 32555
rect 3668 32490 4176 32499
rect 3668 32438 3729 32490
rect 3781 32438 4176 32490
rect 3668 32431 4176 32438
rect 3668 32375 3708 32431
rect 3764 32382 3832 32431
rect 3781 32375 3832 32382
rect 3888 32375 3956 32431
rect 4012 32375 4080 32431
rect 4136 32375 4176 32431
rect 3668 32330 3729 32375
rect 3781 32330 4176 32375
rect 3668 32307 4176 32330
rect 3668 32251 3708 32307
rect 3764 32274 3832 32307
rect 3781 32251 3832 32274
rect 3888 32251 3956 32307
rect 4012 32251 4080 32307
rect 4136 32251 4176 32307
rect 3668 32222 3729 32251
rect 3781 32222 4176 32251
rect 3668 32183 4176 32222
rect 3668 32127 3708 32183
rect 3764 32166 3832 32183
rect 3781 32127 3832 32166
rect 3888 32127 3956 32183
rect 4012 32127 4080 32183
rect 4136 32127 4176 32183
rect 3668 32114 3729 32127
rect 3781 32114 4176 32127
rect 3668 32059 4176 32114
rect 3668 32003 3708 32059
rect 3764 32058 3832 32059
rect 3781 32006 3832 32058
rect 3764 32003 3832 32006
rect 3888 32003 3956 32059
rect 4012 32003 4080 32059
rect 4136 32003 4176 32059
rect 3668 31950 4176 32003
rect 3668 31935 3729 31950
rect 3781 31935 4176 31950
rect 3668 31879 3708 31935
rect 3781 31898 3832 31935
rect 3764 31879 3832 31898
rect 3888 31879 3956 31935
rect 4012 31879 4080 31935
rect 4136 31879 4176 31935
rect 3668 31842 4176 31879
rect 3668 31811 3729 31842
rect 3781 31811 4176 31842
rect 3668 31755 3708 31811
rect 3781 31790 3832 31811
rect 3764 31755 3832 31790
rect 3888 31755 3956 31811
rect 4012 31755 4080 31811
rect 4136 31755 4176 31811
rect 3668 31734 4176 31755
rect 3668 31687 3729 31734
rect 3781 31687 4176 31734
rect 3668 31631 3708 31687
rect 3781 31682 3832 31687
rect 3764 31631 3832 31682
rect 3888 31631 3956 31687
rect 4012 31631 4080 31687
rect 4136 31631 4176 31687
rect 3668 31626 4176 31631
rect 3668 31574 3729 31626
rect 3781 31574 4176 31626
rect 3668 31563 4176 31574
rect 3668 31507 3708 31563
rect 3764 31518 3832 31563
rect 3781 31507 3832 31518
rect 3888 31507 3956 31563
rect 4012 31507 4080 31563
rect 4136 31507 4176 31563
rect 3668 31466 3729 31507
rect 3781 31466 4176 31507
rect 3668 31439 4176 31466
rect 3668 31383 3708 31439
rect 3764 31410 3832 31439
rect 3781 31383 3832 31410
rect 3888 31383 3956 31439
rect 4012 31383 4080 31439
rect 4136 31383 4176 31439
rect 3668 31358 3729 31383
rect 3781 31358 4176 31383
rect 3668 31315 4176 31358
rect 3668 31259 3708 31315
rect 3764 31302 3832 31315
rect 3781 31259 3832 31302
rect 3888 31259 3956 31315
rect 4012 31259 4080 31315
rect 4136 31259 4176 31315
rect 3668 31250 3729 31259
rect 3781 31250 4176 31259
rect 3668 31194 4176 31250
rect 3668 31191 3729 31194
rect 3781 31191 4176 31194
rect 3668 31135 3708 31191
rect 3781 31142 3832 31191
rect 3764 31135 3832 31142
rect 3888 31135 3956 31191
rect 4012 31135 4080 31191
rect 4136 31135 4176 31191
rect 3668 31086 4176 31135
rect 3668 31067 3729 31086
rect 3781 31067 4176 31086
rect 3668 31011 3708 31067
rect 3781 31034 3832 31067
rect 3764 31011 3832 31034
rect 3888 31011 3956 31067
rect 4012 31011 4080 31067
rect 4136 31011 4176 31067
rect 3668 30978 4176 31011
rect 3668 30943 3729 30978
rect 3781 30943 4176 30978
rect 3668 30887 3708 30943
rect 3781 30926 3832 30943
rect 3764 30887 3832 30926
rect 3888 30887 3956 30943
rect 4012 30887 4080 30943
rect 4136 30887 4176 30943
rect 3668 30870 4176 30887
rect 3668 30819 3729 30870
rect 3781 30819 4176 30870
rect 3668 30763 3708 30819
rect 3781 30818 3832 30819
rect 3764 30763 3832 30818
rect 3888 30763 3956 30819
rect 4012 30763 4080 30819
rect 4136 30763 4176 30819
rect 3668 30762 4176 30763
rect 3668 30710 3729 30762
rect 3781 30710 4176 30762
rect 3668 30695 4176 30710
rect 3668 30639 3708 30695
rect 3764 30654 3832 30695
rect 3781 30639 3832 30654
rect 3888 30639 3956 30695
rect 4012 30639 4080 30695
rect 4136 30639 4176 30695
rect 3668 30602 3729 30639
rect 3781 30602 4176 30639
rect 3668 30571 4176 30602
rect 3668 30515 3708 30571
rect 3764 30546 3832 30571
rect 3781 30515 3832 30546
rect 3888 30515 3956 30571
rect 4012 30515 4080 30571
rect 4136 30515 4176 30571
rect 3668 30494 3729 30515
rect 3781 30494 4176 30515
rect 3668 30447 4176 30494
rect 3668 30391 3708 30447
rect 3764 30438 3832 30447
rect 3781 30391 3832 30438
rect 3888 30391 3956 30447
rect 4012 30391 4080 30447
rect 4136 30391 4176 30447
rect 3668 30386 3729 30391
rect 3781 30386 4176 30391
rect 3668 30330 4176 30386
rect 3668 30323 3729 30330
rect 3781 30323 4176 30330
rect 3668 30267 3708 30323
rect 3781 30278 3832 30323
rect 3764 30267 3832 30278
rect 3888 30267 3956 30323
rect 4012 30267 4080 30323
rect 4136 30267 4176 30323
rect 3668 30222 4176 30267
rect 3668 30199 3729 30222
rect 3781 30199 4176 30222
rect 3668 30143 3708 30199
rect 3781 30170 3832 30199
rect 3764 30143 3832 30170
rect 3888 30143 3956 30199
rect 4012 30143 4080 30199
rect 4136 30143 4176 30199
rect 3668 30114 4176 30143
rect 3668 30062 3729 30114
rect 3781 30062 4176 30114
rect 3668 30006 4176 30062
rect 3668 29954 3729 30006
rect 3781 29954 4176 30006
rect 3668 29898 4176 29954
rect 3668 29846 3729 29898
rect 3781 29846 4176 29898
rect 3668 29845 4176 29846
rect 3668 29789 3708 29845
rect 3764 29790 3832 29845
rect 3781 29789 3832 29790
rect 3888 29789 3956 29845
rect 4012 29789 4080 29845
rect 4136 29789 4176 29845
rect 3668 29738 3729 29789
rect 3781 29738 4176 29789
rect 3668 29721 4176 29738
rect 3668 29665 3708 29721
rect 3764 29682 3832 29721
rect 3781 29665 3832 29682
rect 3888 29665 3956 29721
rect 4012 29665 4080 29721
rect 4136 29665 4176 29721
rect 3668 29630 3729 29665
rect 3781 29630 4176 29665
rect 3668 29597 4176 29630
rect 3668 29541 3708 29597
rect 3764 29574 3832 29597
rect 3781 29541 3832 29574
rect 3888 29541 3956 29597
rect 4012 29541 4080 29597
rect 4136 29541 4176 29597
rect 3668 29522 3729 29541
rect 3781 29522 4176 29541
rect 3668 29473 4176 29522
rect 3668 29417 3708 29473
rect 3764 29417 3832 29473
rect 3888 29417 3956 29473
rect 4012 29417 4080 29473
rect 4136 29417 4176 29473
rect 3668 29349 4176 29417
rect 3668 29293 3708 29349
rect 3764 29293 3832 29349
rect 3888 29293 3956 29349
rect 4012 29293 4080 29349
rect 4136 29293 4176 29349
rect 3668 29225 4176 29293
rect 3668 29169 3708 29225
rect 3764 29169 3832 29225
rect 3888 29169 3956 29225
rect 4012 29169 4080 29225
rect 4136 29169 4176 29225
rect 3668 29101 4176 29169
rect 3668 29045 3708 29101
rect 3764 29045 3832 29101
rect 3888 29045 3956 29101
rect 4012 29045 4080 29101
rect 4136 29045 4176 29101
rect 3668 28977 4176 29045
rect 3668 28921 3708 28977
rect 3764 28921 3832 28977
rect 3888 28921 3956 28977
rect 4012 28921 4080 28977
rect 4136 28921 4176 28977
rect 3668 28853 4176 28921
rect 3668 28797 3708 28853
rect 3764 28797 3832 28853
rect 3888 28797 3956 28853
rect 4012 28797 4080 28853
rect 4136 28797 4176 28853
rect 3668 28729 4176 28797
rect 3668 28673 3708 28729
rect 3764 28673 3832 28729
rect 3888 28673 3956 28729
rect 4012 28673 4080 28729
rect 4136 28673 4176 28729
rect 3668 28650 4176 28673
rect 3668 28605 3729 28650
rect 3781 28605 4176 28650
rect 3668 28549 3708 28605
rect 3781 28598 3832 28605
rect 3764 28549 3832 28598
rect 3888 28549 3956 28605
rect 4012 28549 4080 28605
rect 4136 28549 4176 28605
rect 3668 28542 4176 28549
rect 3668 28490 3729 28542
rect 3781 28490 4176 28542
rect 3668 28434 4176 28490
rect 3668 28382 3729 28434
rect 3781 28382 4176 28434
rect 3668 28326 4176 28382
rect 3668 28274 3729 28326
rect 3781 28274 4176 28326
rect 3668 28218 4176 28274
rect 3668 28166 3729 28218
rect 3781 28166 4176 28218
rect 3668 28110 4176 28166
rect 3668 28058 3729 28110
rect 3781 28058 4176 28110
rect 3668 28002 4176 28058
rect 3668 27950 3729 28002
rect 3781 27950 4176 28002
rect 3668 27894 4176 27950
rect 3668 27842 3729 27894
rect 3781 27842 4176 27894
rect 3668 27786 4176 27842
rect 3668 27734 3729 27786
rect 3781 27734 4176 27786
rect 3668 27678 4176 27734
rect 3668 27626 3729 27678
rect 3781 27626 4176 27678
rect 3668 27570 4176 27626
rect 3668 27518 3729 27570
rect 3781 27518 4176 27570
rect 3668 27462 4176 27518
rect 3668 27410 3729 27462
rect 3781 27410 4176 27462
rect 3668 27354 4176 27410
rect 3668 27302 3729 27354
rect 3781 27302 4176 27354
rect 3668 27246 4176 27302
rect 3668 27194 3729 27246
rect 3781 27194 4176 27246
rect 3668 27138 4176 27194
rect 3668 27086 3729 27138
rect 3781 27086 4176 27138
rect 3668 27030 4176 27086
rect 3668 26978 3729 27030
rect 3781 26978 4176 27030
rect 3668 26922 4176 26978
rect 3668 26870 3729 26922
rect 3781 26870 4176 26922
rect 3668 26814 4176 26870
rect 3668 26762 3729 26814
rect 3781 26762 4176 26814
rect 3668 26706 4176 26762
rect 3668 26654 3729 26706
rect 3781 26654 4176 26706
rect 3668 26651 4176 26654
rect 3668 26595 3708 26651
rect 3764 26598 3832 26651
rect 3781 26595 3832 26598
rect 3888 26595 3956 26651
rect 4012 26595 4080 26651
rect 4136 26595 4176 26651
rect 3668 26546 3729 26595
rect 3781 26546 4176 26595
rect 3668 26527 4176 26546
rect 3668 26471 3708 26527
rect 3764 26490 3832 26527
rect 3781 26471 3832 26490
rect 3888 26471 3956 26527
rect 4012 26471 4080 26527
rect 4136 26471 4176 26527
rect 3668 26438 3729 26471
rect 3781 26438 4176 26471
rect 3668 26403 4176 26438
rect 3668 26347 3708 26403
rect 3764 26382 3832 26403
rect 3781 26347 3832 26382
rect 3888 26347 3956 26403
rect 4012 26347 4080 26403
rect 4136 26347 4176 26403
rect 3668 26330 3729 26347
rect 3781 26330 4176 26347
rect 3668 26279 4176 26330
rect 3668 26223 3708 26279
rect 3764 26274 3832 26279
rect 3781 26223 3832 26274
rect 3888 26223 3956 26279
rect 4012 26223 4080 26279
rect 4136 26223 4176 26279
rect 3668 26222 3729 26223
rect 3781 26222 4176 26223
rect 3668 26166 4176 26222
rect 3668 26155 3729 26166
rect 3781 26155 4176 26166
rect 3668 26099 3708 26155
rect 3781 26114 3832 26155
rect 3764 26099 3832 26114
rect 3888 26099 3956 26155
rect 4012 26099 4080 26155
rect 4136 26099 4176 26155
rect 3668 26058 4176 26099
rect 3668 26031 3729 26058
rect 3781 26031 4176 26058
rect 3668 25975 3708 26031
rect 3781 26006 3832 26031
rect 3764 25975 3832 26006
rect 3888 25975 3956 26031
rect 4012 25975 4080 26031
rect 4136 25975 4176 26031
rect 3668 25950 4176 25975
rect 3668 25907 3729 25950
rect 3781 25907 4176 25950
rect 3668 25851 3708 25907
rect 3781 25898 3832 25907
rect 3764 25851 3832 25898
rect 3888 25851 3956 25907
rect 4012 25851 4080 25907
rect 4136 25851 4176 25907
rect 3668 25842 4176 25851
rect 3668 25790 3729 25842
rect 3781 25790 4176 25842
rect 3668 25783 4176 25790
rect 3668 25727 3708 25783
rect 3764 25734 3832 25783
rect 3781 25727 3832 25734
rect 3888 25727 3956 25783
rect 4012 25727 4080 25783
rect 4136 25727 4176 25783
rect 3668 25682 3729 25727
rect 3781 25682 4176 25727
rect 3668 25659 4176 25682
rect 3668 25603 3708 25659
rect 3764 25626 3832 25659
rect 3781 25603 3832 25626
rect 3888 25603 3956 25659
rect 4012 25603 4080 25659
rect 4136 25603 4176 25659
rect 3668 25574 3729 25603
rect 3781 25574 4176 25603
rect 3668 25535 4176 25574
rect 3668 25479 3708 25535
rect 3764 25479 3832 25535
rect 3888 25479 3956 25535
rect 4012 25479 4080 25535
rect 4136 25479 4176 25535
rect 3668 25411 4176 25479
rect 3668 25355 3708 25411
rect 3764 25355 3832 25411
rect 3888 25355 3956 25411
rect 4012 25355 4080 25411
rect 4136 25355 4176 25411
rect 3668 25287 4176 25355
rect 3668 25231 3708 25287
rect 3764 25231 3832 25287
rect 3888 25231 3956 25287
rect 4012 25231 4080 25287
rect 4136 25231 4176 25287
rect 3668 25163 4176 25231
rect 3668 25107 3708 25163
rect 3764 25107 3832 25163
rect 3888 25107 3956 25163
rect 4012 25107 4080 25163
rect 4136 25107 4176 25163
rect 3668 25039 4176 25107
rect 3668 24983 3708 25039
rect 3764 24983 3832 25039
rect 3888 24983 3956 25039
rect 4012 24983 4080 25039
rect 4136 24983 4176 25039
rect 3668 24915 4176 24983
rect 3668 24859 3708 24915
rect 3764 24859 3832 24915
rect 3888 24859 3956 24915
rect 4012 24859 4080 24915
rect 4136 24859 4176 24915
rect 3668 24791 4176 24859
rect 3668 24735 3708 24791
rect 3764 24735 3832 24791
rect 3888 24735 3956 24791
rect 4012 24735 4080 24791
rect 4136 24735 4176 24791
rect 3668 24702 4176 24735
rect 3668 24667 3729 24702
rect 3781 24667 4176 24702
rect 3668 24611 3708 24667
rect 3781 24650 3832 24667
rect 3764 24611 3832 24650
rect 3888 24611 3956 24667
rect 4012 24611 4080 24667
rect 4136 24611 4176 24667
rect 3668 24594 4176 24611
rect 3668 24543 3729 24594
rect 3781 24543 4176 24594
rect 3668 24487 3708 24543
rect 3781 24542 3832 24543
rect 3764 24487 3832 24542
rect 3888 24487 3956 24543
rect 4012 24487 4080 24543
rect 4136 24487 4176 24543
rect 3668 24486 4176 24487
rect 3668 24434 3729 24486
rect 3781 24434 4176 24486
rect 3668 24419 4176 24434
rect 3668 24363 3708 24419
rect 3764 24378 3832 24419
rect 3781 24363 3832 24378
rect 3888 24363 3956 24419
rect 4012 24363 4080 24419
rect 4136 24363 4176 24419
rect 3668 24326 3729 24363
rect 3781 24326 4176 24363
rect 3668 24295 4176 24326
rect 3668 24239 3708 24295
rect 3764 24270 3832 24295
rect 3781 24239 3832 24270
rect 3888 24239 3956 24295
rect 4012 24239 4080 24295
rect 4136 24239 4176 24295
rect 3668 24218 3729 24239
rect 3781 24218 4176 24239
rect 3668 24171 4176 24218
rect 3668 24115 3708 24171
rect 3764 24162 3832 24171
rect 3781 24115 3832 24162
rect 3888 24115 3956 24171
rect 4012 24115 4080 24171
rect 4136 24115 4176 24171
rect 3668 24110 3729 24115
rect 3781 24110 4176 24115
rect 3668 24054 4176 24110
rect 3668 24047 3729 24054
rect 3781 24047 4176 24054
rect 3668 23991 3708 24047
rect 3781 24002 3832 24047
rect 3764 23991 3832 24002
rect 3888 23991 3956 24047
rect 4012 23991 4080 24047
rect 4136 23991 4176 24047
rect 3668 23946 4176 23991
rect 3668 23923 3729 23946
rect 3781 23923 4176 23946
rect 3668 23867 3708 23923
rect 3781 23894 3832 23923
rect 3764 23867 3832 23894
rect 3888 23867 3956 23923
rect 4012 23867 4080 23923
rect 4136 23867 4176 23923
rect 3668 23838 4176 23867
rect 3668 23799 3729 23838
rect 3781 23799 4176 23838
rect 3668 23743 3708 23799
rect 3781 23786 3832 23799
rect 3764 23743 3832 23786
rect 3888 23743 3956 23799
rect 4012 23743 4080 23799
rect 4136 23743 4176 23799
rect 3668 23730 4176 23743
rect 3668 23678 3729 23730
rect 3781 23678 4176 23730
rect 3668 23622 4176 23678
rect 3668 23570 3729 23622
rect 3781 23570 4176 23622
rect 3668 23514 4176 23570
rect 3668 23462 3729 23514
rect 3781 23462 4176 23514
rect 3668 23451 4176 23462
rect 3668 23395 3708 23451
rect 3764 23406 3832 23451
rect 3781 23395 3832 23406
rect 3888 23395 3956 23451
rect 4012 23395 4080 23451
rect 4136 23395 4176 23451
rect 3668 23354 3729 23395
rect 3781 23354 4176 23395
rect 3668 23327 4176 23354
rect 3668 23271 3708 23327
rect 3764 23298 3832 23327
rect 3781 23271 3832 23298
rect 3888 23271 3956 23327
rect 4012 23271 4080 23327
rect 4136 23271 4176 23327
rect 3668 23246 3729 23271
rect 3781 23246 4176 23271
rect 3668 23203 4176 23246
rect 3668 23147 3708 23203
rect 3764 23190 3832 23203
rect 3781 23147 3832 23190
rect 3888 23147 3956 23203
rect 4012 23147 4080 23203
rect 4136 23147 4176 23203
rect 3668 23138 3729 23147
rect 3781 23138 4176 23147
rect 3668 23082 4176 23138
rect 3668 23079 3729 23082
rect 3781 23079 4176 23082
rect 3668 23023 3708 23079
rect 3781 23030 3832 23079
rect 3764 23023 3832 23030
rect 3888 23023 3956 23079
rect 4012 23023 4080 23079
rect 4136 23023 4176 23079
rect 3668 22974 4176 23023
rect 3668 22955 3729 22974
rect 3781 22955 4176 22974
rect 3668 22899 3708 22955
rect 3781 22922 3832 22955
rect 3764 22899 3832 22922
rect 3888 22899 3956 22955
rect 4012 22899 4080 22955
rect 4136 22899 4176 22955
rect 3668 22866 4176 22899
rect 3668 22831 3729 22866
rect 3781 22831 4176 22866
rect 3668 22775 3708 22831
rect 3781 22814 3832 22831
rect 3764 22775 3832 22814
rect 3888 22775 3956 22831
rect 4012 22775 4080 22831
rect 4136 22775 4176 22831
rect 3668 22758 4176 22775
rect 3668 22707 3729 22758
rect 3781 22707 4176 22758
rect 3668 22651 3708 22707
rect 3781 22706 3832 22707
rect 3764 22651 3832 22706
rect 3888 22651 3956 22707
rect 4012 22651 4080 22707
rect 4136 22651 4176 22707
rect 3668 22650 4176 22651
rect 3668 22598 3729 22650
rect 3781 22598 4176 22650
rect 3668 22583 4176 22598
rect 3668 22527 3708 22583
rect 3764 22542 3832 22583
rect 3781 22527 3832 22542
rect 3888 22527 3956 22583
rect 4012 22527 4080 22583
rect 4136 22527 4176 22583
rect 3668 22490 3729 22527
rect 3781 22490 4176 22527
rect 3668 22459 4176 22490
rect 3668 22403 3708 22459
rect 3764 22434 3832 22459
rect 3781 22403 3832 22434
rect 3888 22403 3956 22459
rect 4012 22403 4080 22459
rect 4136 22403 4176 22459
rect 3668 22382 3729 22403
rect 3781 22382 4176 22403
rect 3668 22335 4176 22382
rect 3668 22279 3708 22335
rect 3764 22326 3832 22335
rect 3781 22279 3832 22326
rect 3888 22279 3956 22335
rect 4012 22279 4080 22335
rect 4136 22279 4176 22335
rect 3668 22274 3729 22279
rect 3781 22274 4176 22279
rect 3668 22218 4176 22274
rect 3668 22211 3729 22218
rect 3781 22211 4176 22218
rect 3668 22155 3708 22211
rect 3781 22166 3832 22211
rect 3764 22155 3832 22166
rect 3888 22155 3956 22211
rect 4012 22155 4080 22211
rect 4136 22155 4176 22211
rect 3668 22110 4176 22155
rect 3668 22087 3729 22110
rect 3781 22087 4176 22110
rect 3668 22031 3708 22087
rect 3781 22058 3832 22087
rect 3764 22031 3832 22058
rect 3888 22031 3956 22087
rect 4012 22031 4080 22087
rect 4136 22031 4176 22087
rect 3668 22002 4176 22031
rect 3668 21963 3729 22002
rect 3781 21963 4176 22002
rect 3668 21907 3708 21963
rect 3781 21950 3832 21963
rect 3764 21907 3832 21950
rect 3888 21907 3956 21963
rect 4012 21907 4080 21963
rect 4136 21907 4176 21963
rect 3668 21894 4176 21907
rect 3668 21842 3729 21894
rect 3781 21842 4176 21894
rect 3668 21839 4176 21842
rect 3668 21783 3708 21839
rect 3764 21786 3832 21839
rect 3781 21783 3832 21786
rect 3888 21783 3956 21839
rect 4012 21783 4080 21839
rect 4136 21783 4176 21839
rect 3668 21734 3729 21783
rect 3781 21734 4176 21783
rect 3668 21715 4176 21734
rect 3668 21659 3708 21715
rect 3764 21678 3832 21715
rect 3781 21659 3832 21678
rect 3888 21659 3956 21715
rect 4012 21659 4080 21715
rect 4136 21659 4176 21715
rect 3668 21626 3729 21659
rect 3781 21626 4176 21659
rect 3668 21591 4176 21626
rect 3668 21535 3708 21591
rect 3764 21535 3832 21591
rect 3888 21535 3956 21591
rect 4012 21535 4080 21591
rect 4136 21535 4176 21591
rect 3668 21467 4176 21535
rect 3668 21411 3708 21467
rect 3764 21411 3832 21467
rect 3888 21411 3956 21467
rect 4012 21411 4080 21467
rect 4136 21411 4176 21467
rect 3668 21343 4176 21411
rect 3668 21287 3708 21343
rect 3764 21287 3832 21343
rect 3888 21287 3956 21343
rect 4012 21287 4080 21343
rect 4136 21287 4176 21343
rect 3668 21219 4176 21287
rect 3668 21163 3708 21219
rect 3764 21163 3832 21219
rect 3888 21163 3956 21219
rect 4012 21163 4080 21219
rect 4136 21163 4176 21219
rect 3668 21095 4176 21163
rect 3668 21039 3708 21095
rect 3764 21039 3832 21095
rect 3888 21039 3956 21095
rect 4012 21039 4080 21095
rect 4136 21039 4176 21095
rect 3668 20971 4176 21039
rect 3668 20915 3708 20971
rect 3764 20915 3832 20971
rect 3888 20915 3956 20971
rect 4012 20915 4080 20971
rect 4136 20915 4176 20971
rect 3668 20847 4176 20915
rect 3668 20791 3708 20847
rect 3764 20791 3832 20847
rect 3888 20791 3956 20847
rect 4012 20791 4080 20847
rect 4136 20791 4176 20847
rect 3668 20723 4176 20791
rect 3668 20667 3708 20723
rect 3764 20667 3832 20723
rect 3888 20667 3956 20723
rect 4012 20667 4080 20723
rect 4136 20667 4176 20723
rect 3668 20599 4176 20667
rect 3668 20577 3708 20599
rect 3764 20577 3832 20599
rect 3888 20577 3956 20599
rect 4012 20577 4080 20599
rect 4136 20577 4176 20599
rect 3668 20525 3680 20577
rect 3764 20543 3788 20577
rect 3888 20543 3896 20577
rect 3732 20525 3788 20543
rect 3840 20525 3896 20543
rect 3948 20543 3956 20577
rect 4056 20543 4080 20577
rect 3948 20525 4004 20543
rect 4056 20525 4112 20543
rect 4164 20525 4176 20577
rect 3668 20469 4176 20525
rect 3668 20417 3680 20469
rect 3732 20417 3788 20469
rect 3840 20417 3896 20469
rect 3948 20417 4004 20469
rect 4056 20417 4112 20469
rect 4164 20417 4176 20469
rect 3668 20361 4176 20417
rect 3668 20309 3680 20361
rect 3732 20309 3788 20361
rect 3840 20309 3896 20361
rect 3948 20309 4004 20361
rect 4056 20309 4112 20361
rect 4164 20309 4176 20361
rect 3668 20251 4176 20309
rect 3668 20195 3708 20251
rect 3764 20195 3832 20251
rect 3888 20195 3956 20251
rect 4012 20195 4080 20251
rect 4136 20195 4176 20251
rect 3668 20127 4176 20195
rect 3668 20071 3708 20127
rect 3764 20071 3832 20127
rect 3888 20071 3956 20127
rect 4012 20071 4080 20127
rect 4136 20071 4176 20127
rect 3668 20003 4176 20071
rect 3668 19947 3708 20003
rect 3764 19947 3832 20003
rect 3888 19947 3956 20003
rect 4012 19947 4080 20003
rect 4136 19947 4176 20003
rect 3668 19879 4176 19947
rect 3668 19823 3708 19879
rect 3764 19823 3832 19879
rect 3888 19823 3956 19879
rect 4012 19823 4080 19879
rect 4136 19823 4176 19879
rect 3668 19755 4176 19823
rect 3668 19699 3708 19755
rect 3764 19699 3832 19755
rect 3888 19699 3956 19755
rect 4012 19699 4080 19755
rect 4136 19699 4176 19755
rect 3668 19631 4176 19699
rect 3668 19584 3708 19631
rect 3764 19584 3832 19631
rect 3888 19584 3956 19631
rect 4012 19584 4080 19631
rect 4136 19584 4176 19631
rect 3668 19532 3680 19584
rect 3764 19575 3788 19584
rect 3888 19575 3896 19584
rect 3732 19532 3788 19575
rect 3840 19532 3896 19575
rect 3948 19575 3956 19584
rect 4056 19575 4080 19584
rect 3948 19532 4004 19575
rect 4056 19532 4112 19575
rect 4164 19532 4176 19584
rect 3668 19507 4176 19532
rect 3668 19476 3708 19507
rect 3764 19476 3832 19507
rect 3888 19476 3956 19507
rect 4012 19476 4080 19507
rect 4136 19476 4176 19507
rect 3668 19424 3680 19476
rect 3764 19451 3788 19476
rect 3888 19451 3896 19476
rect 3732 19424 3788 19451
rect 3840 19424 3896 19451
rect 3948 19451 3956 19476
rect 4056 19451 4080 19476
rect 3948 19424 4004 19451
rect 4056 19424 4112 19451
rect 4164 19424 4176 19476
rect 3668 19383 4176 19424
rect 3668 19327 3708 19383
rect 3764 19327 3832 19383
rect 3888 19327 3956 19383
rect 4012 19327 4080 19383
rect 4136 19327 4176 19383
rect 3668 19259 4176 19327
rect 3668 19203 3708 19259
rect 3764 19203 3832 19259
rect 3888 19203 3956 19259
rect 4012 19203 4080 19259
rect 4136 19203 4176 19259
rect 3668 19135 4176 19203
rect 3668 19079 3708 19135
rect 3764 19079 3832 19135
rect 3888 19079 3956 19135
rect 4012 19079 4080 19135
rect 4136 19079 4176 19135
rect 3668 19011 4176 19079
rect 3668 18955 3708 19011
rect 3764 18955 3832 19011
rect 3888 18955 3956 19011
rect 4012 18955 4080 19011
rect 4136 18955 4176 19011
rect 3668 18887 4176 18955
rect 3668 18831 3708 18887
rect 3764 18831 3832 18887
rect 3888 18831 3956 18887
rect 4012 18831 4080 18887
rect 4136 18831 4176 18887
rect 3668 18763 4176 18831
rect 3668 18712 3708 18763
rect 3764 18712 3832 18763
rect 3888 18712 3956 18763
rect 4012 18712 4080 18763
rect 4136 18712 4176 18763
rect 3668 18660 3680 18712
rect 3764 18707 3788 18712
rect 3888 18707 3896 18712
rect 3732 18660 3788 18707
rect 3840 18660 3896 18707
rect 3948 18707 3956 18712
rect 4056 18707 4080 18712
rect 3948 18660 4004 18707
rect 4056 18660 4112 18707
rect 4164 18660 4176 18712
rect 3668 18639 4176 18660
rect 3668 18604 3708 18639
rect 3764 18604 3832 18639
rect 3888 18604 3956 18639
rect 4012 18604 4080 18639
rect 4136 18604 4176 18639
rect 3668 18552 3680 18604
rect 3764 18583 3788 18604
rect 3888 18583 3896 18604
rect 3732 18552 3788 18583
rect 3840 18552 3896 18583
rect 3948 18583 3956 18604
rect 4056 18583 4080 18604
rect 3948 18552 4004 18583
rect 4056 18552 4112 18583
rect 4164 18552 4176 18604
rect 3668 18515 4176 18552
rect 3668 18459 3708 18515
rect 3764 18459 3832 18515
rect 3888 18459 3956 18515
rect 4012 18459 4080 18515
rect 4136 18459 4176 18515
rect 3668 18391 4176 18459
rect 3668 18335 3708 18391
rect 3764 18335 3832 18391
rect 3888 18335 3956 18391
rect 4012 18335 4080 18391
rect 4136 18335 4176 18391
rect 3668 18267 4176 18335
rect 3668 18211 3708 18267
rect 3764 18211 3832 18267
rect 3888 18211 3956 18267
rect 4012 18211 4080 18267
rect 4136 18211 4176 18267
rect 3668 18143 4176 18211
rect 3668 18087 3708 18143
rect 3764 18087 3832 18143
rect 3888 18087 3956 18143
rect 4012 18087 4080 18143
rect 4136 18087 4176 18143
rect 3668 18019 4176 18087
rect 3668 17963 3708 18019
rect 3764 17963 3832 18019
rect 3888 17963 3956 18019
rect 4012 17963 4080 18019
rect 4136 17963 4176 18019
rect 3668 17895 4176 17963
rect 3668 17840 3708 17895
rect 3764 17840 3832 17895
rect 3888 17840 3956 17895
rect 4012 17840 4080 17895
rect 4136 17840 4176 17895
rect 3668 17788 3680 17840
rect 3764 17839 3788 17840
rect 3888 17839 3896 17840
rect 3732 17788 3788 17839
rect 3840 17788 3896 17839
rect 3948 17839 3956 17840
rect 4056 17839 4080 17840
rect 3948 17788 4004 17839
rect 4056 17788 4112 17839
rect 4164 17788 4176 17840
rect 3668 17771 4176 17788
rect 3668 17732 3708 17771
rect 3764 17732 3832 17771
rect 3888 17732 3956 17771
rect 4012 17732 4080 17771
rect 4136 17732 4176 17771
rect 3668 17680 3680 17732
rect 3764 17715 3788 17732
rect 3888 17715 3896 17732
rect 3732 17680 3788 17715
rect 3840 17680 3896 17715
rect 3948 17715 3956 17732
rect 4056 17715 4080 17732
rect 3948 17680 4004 17715
rect 4056 17680 4112 17715
rect 4164 17680 4176 17732
rect 3668 17647 4176 17680
rect 3668 17591 3708 17647
rect 3764 17591 3832 17647
rect 3888 17591 3956 17647
rect 4012 17591 4080 17647
rect 4136 17591 4176 17647
rect 3668 17523 4176 17591
rect 3668 17467 3708 17523
rect 3764 17467 3832 17523
rect 3888 17467 3956 17523
rect 4012 17467 4080 17523
rect 4136 17467 4176 17523
rect 3668 17399 4176 17467
rect 3668 17343 3708 17399
rect 3764 17343 3832 17399
rect 3888 17343 3956 17399
rect 4012 17343 4080 17399
rect 4136 17343 4176 17399
rect 3668 17051 4176 17343
rect 3668 16995 3708 17051
rect 3764 16995 3832 17051
rect 3888 16995 3956 17051
rect 4012 16995 4080 17051
rect 4136 16995 4176 17051
rect 3668 16968 4176 16995
rect 3668 16916 3680 16968
rect 3732 16927 3788 16968
rect 3840 16927 3896 16968
rect 3764 16916 3788 16927
rect 3888 16916 3896 16927
rect 3948 16927 4004 16968
rect 4056 16927 4112 16968
rect 3948 16916 3956 16927
rect 4056 16916 4080 16927
rect 4164 16916 4176 16968
rect 3668 16871 3708 16916
rect 3764 16871 3832 16916
rect 3888 16871 3956 16916
rect 4012 16871 4080 16916
rect 4136 16871 4176 16916
rect 3668 16860 4176 16871
rect 3668 16808 3680 16860
rect 3732 16808 3788 16860
rect 3840 16808 3896 16860
rect 3948 16808 4004 16860
rect 4056 16808 4112 16860
rect 4164 16808 4176 16860
rect 3668 16803 4176 16808
rect 3668 16747 3708 16803
rect 3764 16747 3832 16803
rect 3888 16747 3956 16803
rect 4012 16747 4080 16803
rect 4136 16747 4176 16803
rect 3668 16679 4176 16747
rect 3668 16623 3708 16679
rect 3764 16623 3832 16679
rect 3888 16623 3956 16679
rect 4012 16623 4080 16679
rect 4136 16623 4176 16679
rect 3668 16555 4176 16623
rect 3668 16499 3708 16555
rect 3764 16499 3832 16555
rect 3888 16499 3956 16555
rect 4012 16499 4080 16555
rect 4136 16499 4176 16555
rect 3668 16431 4176 16499
rect 3668 16375 3708 16431
rect 3764 16375 3832 16431
rect 3888 16375 3956 16431
rect 4012 16375 4080 16431
rect 4136 16375 4176 16431
rect 3668 16307 4176 16375
rect 3668 16251 3708 16307
rect 3764 16251 3832 16307
rect 3888 16251 3956 16307
rect 4012 16251 4080 16307
rect 4136 16251 4176 16307
rect 3668 16183 4176 16251
rect 3668 16127 3708 16183
rect 3764 16127 3832 16183
rect 3888 16127 3956 16183
rect 4012 16127 4080 16183
rect 4136 16127 4176 16183
rect 3668 16083 4176 16127
rect 3668 16031 3680 16083
rect 3732 16059 3788 16083
rect 3840 16059 3896 16083
rect 3764 16031 3788 16059
rect 3888 16031 3896 16059
rect 3948 16059 4004 16083
rect 4056 16059 4112 16083
rect 3948 16031 3956 16059
rect 4056 16031 4080 16059
rect 4164 16031 4176 16083
rect 3668 16003 3708 16031
rect 3764 16003 3832 16031
rect 3888 16003 3956 16031
rect 4012 16003 4080 16031
rect 4136 16003 4176 16031
rect 3668 15975 4176 16003
rect 3668 15923 3680 15975
rect 3732 15935 3788 15975
rect 3840 15935 3896 15975
rect 3764 15923 3788 15935
rect 3888 15923 3896 15935
rect 3948 15935 4004 15975
rect 4056 15935 4112 15975
rect 3948 15923 3956 15935
rect 4056 15923 4080 15935
rect 4164 15923 4176 15975
rect 3668 15879 3708 15923
rect 3764 15879 3832 15923
rect 3888 15879 3956 15923
rect 4012 15879 4080 15923
rect 4136 15879 4176 15923
rect 3668 15867 4176 15879
rect 3668 15815 3680 15867
rect 3732 15815 3788 15867
rect 3840 15815 3896 15867
rect 3948 15815 4004 15867
rect 4056 15815 4112 15867
rect 4164 15815 4176 15867
rect 3668 15811 4176 15815
rect 3668 15762 3708 15811
rect 2432 15755 2442 15762
rect 1994 15687 2442 15755
rect 1994 15631 2004 15687
rect 2060 15631 2128 15687
rect 2184 15631 2252 15687
rect 2308 15631 2376 15687
rect 2432 15631 2442 15687
rect 1994 15563 2442 15631
rect 1994 15507 2004 15563
rect 2060 15507 2128 15563
rect 2184 15507 2252 15563
rect 2308 15507 2376 15563
rect 2432 15507 2442 15563
rect 1994 15439 2442 15507
rect 1994 15383 2004 15439
rect 2060 15383 2128 15439
rect 2184 15383 2252 15439
rect 2308 15383 2376 15439
rect 2432 15383 2442 15439
rect 1994 15315 2442 15383
rect 1994 15259 2004 15315
rect 2060 15259 2128 15315
rect 2184 15259 2252 15315
rect 2308 15259 2376 15315
rect 2432 15259 2442 15315
rect 1994 15191 2442 15259
rect 1994 15135 2004 15191
rect 2060 15135 2128 15191
rect 2184 15135 2252 15191
rect 2308 15135 2376 15191
rect 2432 15135 2442 15191
rect 1994 15067 2442 15135
rect 1994 15011 2004 15067
rect 2060 15011 2128 15067
rect 2184 15011 2252 15067
rect 2308 15011 2376 15067
rect 2432 15011 2442 15067
rect 1994 14943 2442 15011
rect 1994 14887 2004 14943
rect 2060 14887 2128 14943
rect 2184 14887 2252 14943
rect 2308 14887 2376 14943
rect 2432 14887 2442 14943
rect 1994 14819 2442 14887
rect 1994 14763 2004 14819
rect 2060 14763 2128 14819
rect 2184 14763 2252 14819
rect 2308 14763 2376 14819
rect 2432 14763 2442 14819
rect 1994 14695 2442 14763
rect 1994 14639 2004 14695
rect 2060 14639 2128 14695
rect 2184 14639 2252 14695
rect 2308 14639 2376 14695
rect 2432 14639 2442 14695
rect 1994 14571 2442 14639
rect 1994 14515 2004 14571
rect 2060 14515 2128 14571
rect 2184 14515 2252 14571
rect 2308 14515 2376 14571
rect 2432 14515 2442 14571
rect 1994 14447 2442 14515
rect 1994 14391 2004 14447
rect 2060 14391 2128 14447
rect 2184 14391 2252 14447
rect 2308 14391 2376 14447
rect 2432 14391 2442 14447
rect 1994 14323 2442 14391
rect 1994 14267 2004 14323
rect 2060 14267 2128 14323
rect 2184 14267 2252 14323
rect 2308 14267 2376 14323
rect 2432 14267 2442 14323
rect 1994 14199 2442 14267
rect 1994 14143 2004 14199
rect 2060 14143 2128 14199
rect 2184 14143 2252 14199
rect 2308 14143 2376 14199
rect 2432 14143 2442 14199
rect 1994 14133 2442 14143
rect 3698 15755 3708 15762
rect 3764 15755 3832 15811
rect 3888 15755 3956 15811
rect 4012 15755 4080 15811
rect 4136 15762 4176 15811
rect 4804 56922 5312 56975
rect 4804 56866 4844 56922
rect 4900 56866 4968 56922
rect 5024 56866 5092 56922
rect 5148 56866 5216 56922
rect 5272 56866 5312 56922
rect 4804 56798 5312 56866
rect 4804 56742 4844 56798
rect 4900 56742 4968 56798
rect 5024 56742 5092 56798
rect 5148 56742 5216 56798
rect 5272 56742 5312 56798
rect 4804 56711 5312 56742
rect 4804 56659 4816 56711
rect 4868 56674 4924 56711
rect 4976 56674 5032 56711
rect 4900 56659 4924 56674
rect 5024 56659 5032 56674
rect 5084 56674 5140 56711
rect 5192 56674 5248 56711
rect 5084 56659 5092 56674
rect 5192 56659 5216 56674
rect 5300 56659 5312 56711
rect 4804 56618 4844 56659
rect 4900 56618 4968 56659
rect 5024 56618 5092 56659
rect 5148 56618 5216 56659
rect 5272 56618 5312 56659
rect 4804 56603 5312 56618
rect 4804 56551 4816 56603
rect 4868 56551 4924 56603
rect 4976 56551 5032 56603
rect 5084 56551 5140 56603
rect 5192 56551 5248 56603
rect 5300 56551 5312 56603
rect 4804 56550 5312 56551
rect 4804 56495 4844 56550
rect 4900 56495 4968 56550
rect 5024 56495 5092 56550
rect 5148 56495 5216 56550
rect 5272 56495 5312 56550
rect 4804 56443 4816 56495
rect 4900 56494 4924 56495
rect 5024 56494 5032 56495
rect 4868 56443 4924 56494
rect 4976 56443 5032 56494
rect 5084 56494 5092 56495
rect 5192 56494 5216 56495
rect 5084 56443 5140 56494
rect 5192 56443 5248 56494
rect 5300 56443 5312 56495
rect 4804 56426 5312 56443
rect 4804 56370 4844 56426
rect 4900 56370 4968 56426
rect 5024 56370 5092 56426
rect 5148 56370 5216 56426
rect 5272 56370 5312 56426
rect 4804 56302 5312 56370
rect 4804 56246 4844 56302
rect 4900 56246 4968 56302
rect 5024 56246 5092 56302
rect 5148 56246 5216 56302
rect 5272 56246 5312 56302
rect 4804 56178 5312 56246
rect 4804 56122 4844 56178
rect 4900 56122 4968 56178
rect 5024 56122 5092 56178
rect 5148 56122 5216 56178
rect 5272 56122 5312 56178
rect 4804 56054 5312 56122
rect 4804 55998 4844 56054
rect 4900 55998 4968 56054
rect 5024 55998 5092 56054
rect 5148 55998 5216 56054
rect 5272 55998 5312 56054
rect 4804 55930 5312 55998
rect 4804 55874 4844 55930
rect 4900 55874 4968 55930
rect 5024 55874 5092 55930
rect 5148 55874 5216 55930
rect 5272 55874 5312 55930
rect 4804 55806 5312 55874
rect 4804 55750 4844 55806
rect 4900 55750 4968 55806
rect 5024 55750 5092 55806
rect 5148 55750 5216 55806
rect 5272 55750 5312 55806
rect 4804 53845 5312 55750
rect 4804 53789 4844 53845
rect 4900 53789 4968 53845
rect 5024 53789 5092 53845
rect 5148 53789 5216 53845
rect 5272 53789 5312 53845
rect 4804 53721 5312 53789
rect 4804 53665 4844 53721
rect 4900 53665 4968 53721
rect 5024 53665 5092 53721
rect 5148 53665 5216 53721
rect 5272 53665 5312 53721
rect 4804 53597 5312 53665
rect 4804 53541 4844 53597
rect 4900 53541 4968 53597
rect 5024 53541 5092 53597
rect 5148 53541 5216 53597
rect 5272 53541 5312 53597
rect 4804 53473 5312 53541
rect 4804 53417 4844 53473
rect 4900 53417 4968 53473
rect 5024 53417 5092 53473
rect 5148 53417 5216 53473
rect 5272 53417 5312 53473
rect 4804 53349 5312 53417
rect 4804 53293 4844 53349
rect 4900 53293 4968 53349
rect 5024 53293 5092 53349
rect 5148 53293 5216 53349
rect 5272 53293 5312 53349
rect 4804 53225 5312 53293
rect 4804 53169 4844 53225
rect 4900 53169 4968 53225
rect 5024 53169 5092 53225
rect 5148 53169 5216 53225
rect 5272 53169 5312 53225
rect 4804 53101 5312 53169
rect 4804 53045 4844 53101
rect 4900 53045 4968 53101
rect 5024 53045 5092 53101
rect 5148 53045 5216 53101
rect 5272 53045 5312 53101
rect 4804 52996 4846 53045
rect 4898 52996 4970 53045
rect 5022 52996 5094 53045
rect 5146 52996 5218 53045
rect 5270 52996 5312 53045
rect 4804 52977 5312 52996
rect 4804 52921 4844 52977
rect 4900 52921 4968 52977
rect 5024 52921 5092 52977
rect 5148 52921 5216 52977
rect 5272 52921 5312 52977
rect 4804 52872 4846 52921
rect 4898 52872 4970 52921
rect 5022 52872 5094 52921
rect 5146 52872 5218 52921
rect 5270 52872 5312 52921
rect 4804 52853 5312 52872
rect 4804 52797 4844 52853
rect 4900 52797 4968 52853
rect 5024 52797 5092 52853
rect 5148 52797 5216 52853
rect 5272 52797 5312 52853
rect 4804 52748 4846 52797
rect 4898 52748 4970 52797
rect 5022 52748 5094 52797
rect 5146 52748 5218 52797
rect 5270 52748 5312 52797
rect 4804 52729 5312 52748
rect 4804 52673 4844 52729
rect 4900 52673 4968 52729
rect 5024 52673 5092 52729
rect 5148 52673 5216 52729
rect 5272 52673 5312 52729
rect 4804 52624 4846 52673
rect 4898 52624 4970 52673
rect 5022 52624 5094 52673
rect 5146 52624 5218 52673
rect 5270 52624 5312 52673
rect 4804 52605 5312 52624
rect 4804 52549 4844 52605
rect 4900 52549 4968 52605
rect 5024 52549 5092 52605
rect 5148 52549 5216 52605
rect 5272 52549 5312 52605
rect 4804 52500 4846 52549
rect 4898 52500 4970 52549
rect 5022 52500 5094 52549
rect 5146 52500 5218 52549
rect 5270 52500 5312 52549
rect 4804 49100 5312 52500
rect 4804 49048 4846 49100
rect 4898 49048 4970 49100
rect 5022 49048 5094 49100
rect 5146 49048 5218 49100
rect 5270 49048 5312 49100
rect 4804 49045 5312 49048
rect 4804 48989 4844 49045
rect 4900 48989 4968 49045
rect 5024 48989 5092 49045
rect 5148 48989 5216 49045
rect 5272 48989 5312 49045
rect 4804 48976 5312 48989
rect 4804 48924 4846 48976
rect 4898 48924 4970 48976
rect 5022 48924 5094 48976
rect 5146 48924 5218 48976
rect 5270 48924 5312 48976
rect 4804 48921 5312 48924
rect 4804 48865 4844 48921
rect 4900 48865 4968 48921
rect 5024 48865 5092 48921
rect 5148 48865 5216 48921
rect 5272 48865 5312 48921
rect 4804 48852 5312 48865
rect 4804 48800 4846 48852
rect 4898 48800 4970 48852
rect 5022 48800 5094 48852
rect 5146 48800 5218 48852
rect 5270 48800 5312 48852
rect 4804 48797 5312 48800
rect 4804 48741 4844 48797
rect 4900 48741 4968 48797
rect 5024 48741 5092 48797
rect 5148 48741 5216 48797
rect 5272 48741 5312 48797
rect 4804 48728 5312 48741
rect 4804 48676 4846 48728
rect 4898 48676 4970 48728
rect 5022 48676 5094 48728
rect 5146 48676 5218 48728
rect 5270 48676 5312 48728
rect 4804 48673 5312 48676
rect 4804 48617 4844 48673
rect 4900 48617 4968 48673
rect 5024 48617 5092 48673
rect 5148 48617 5216 48673
rect 5272 48617 5312 48673
rect 4804 48604 5312 48617
rect 4804 48552 4846 48604
rect 4898 48552 4970 48604
rect 5022 48552 5094 48604
rect 5146 48552 5218 48604
rect 5270 48552 5312 48604
rect 4804 48549 5312 48552
rect 4804 48493 4844 48549
rect 4900 48493 4968 48549
rect 5024 48493 5092 48549
rect 5148 48493 5216 48549
rect 5272 48493 5312 48549
rect 4804 48425 5312 48493
rect 4804 48369 4844 48425
rect 4900 48369 4968 48425
rect 5024 48369 5092 48425
rect 5148 48369 5216 48425
rect 5272 48369 5312 48425
rect 4804 48301 5312 48369
rect 4804 48245 4844 48301
rect 4900 48245 4968 48301
rect 5024 48245 5092 48301
rect 5148 48245 5216 48301
rect 5272 48245 5312 48301
rect 4804 48177 5312 48245
rect 4804 48121 4844 48177
rect 4900 48121 4968 48177
rect 5024 48121 5092 48177
rect 5148 48121 5216 48177
rect 5272 48121 5312 48177
rect 4804 48053 5312 48121
rect 4804 47997 4844 48053
rect 4900 47997 4968 48053
rect 5024 47997 5092 48053
rect 5148 47997 5216 48053
rect 5272 47997 5312 48053
rect 4804 47929 5312 47997
rect 4804 47873 4844 47929
rect 4900 47873 4968 47929
rect 5024 47873 5092 47929
rect 5148 47873 5216 47929
rect 5272 47873 5312 47929
rect 4804 47805 5312 47873
rect 4804 47749 4844 47805
rect 4900 47749 4968 47805
rect 5024 47749 5092 47805
rect 5148 47749 5216 47805
rect 5272 47749 5312 47805
rect 4804 45845 5312 47749
rect 4804 45789 4844 45845
rect 4900 45789 4968 45845
rect 5024 45789 5092 45845
rect 5148 45789 5216 45845
rect 5272 45789 5312 45845
rect 4804 45721 5312 45789
rect 4804 45665 4844 45721
rect 4900 45665 4968 45721
rect 5024 45665 5092 45721
rect 5148 45665 5216 45721
rect 5272 45665 5312 45721
rect 4804 45597 5312 45665
rect 4804 45541 4844 45597
rect 4900 45541 4968 45597
rect 5024 45541 5092 45597
rect 5148 45541 5216 45597
rect 5272 45541 5312 45597
rect 4804 45473 5312 45541
rect 4804 45417 4844 45473
rect 4900 45417 4968 45473
rect 5024 45417 5092 45473
rect 5148 45417 5216 45473
rect 5272 45417 5312 45473
rect 4804 45349 5312 45417
rect 4804 45293 4844 45349
rect 4900 45293 4968 45349
rect 5024 45293 5092 45349
rect 5148 45293 5216 45349
rect 5272 45293 5312 45349
rect 4804 45225 5312 45293
rect 4804 45169 4844 45225
rect 4900 45169 4968 45225
rect 5024 45169 5092 45225
rect 5148 45169 5216 45225
rect 5272 45169 5312 45225
rect 4804 45152 5312 45169
rect 4804 45101 4846 45152
rect 4898 45101 4970 45152
rect 5022 45101 5094 45152
rect 5146 45101 5218 45152
rect 5270 45101 5312 45152
rect 4804 45045 4844 45101
rect 4900 45045 4968 45101
rect 5024 45045 5092 45101
rect 5148 45045 5216 45101
rect 5272 45045 5312 45101
rect 4804 45028 5312 45045
rect 4804 44977 4846 45028
rect 4898 44977 4970 45028
rect 5022 44977 5094 45028
rect 5146 44977 5218 45028
rect 5270 44977 5312 45028
rect 4804 44921 4844 44977
rect 4900 44921 4968 44977
rect 5024 44921 5092 44977
rect 5148 44921 5216 44977
rect 5272 44921 5312 44977
rect 4804 44904 5312 44921
rect 4804 44853 4846 44904
rect 4898 44853 4970 44904
rect 5022 44853 5094 44904
rect 5146 44853 5218 44904
rect 5270 44853 5312 44904
rect 4804 44797 4844 44853
rect 4900 44797 4968 44853
rect 5024 44797 5092 44853
rect 5148 44797 5216 44853
rect 5272 44797 5312 44853
rect 4804 44780 5312 44797
rect 4804 44729 4846 44780
rect 4898 44729 4970 44780
rect 5022 44729 5094 44780
rect 5146 44729 5218 44780
rect 5270 44729 5312 44780
rect 4804 44673 4844 44729
rect 4900 44673 4968 44729
rect 5024 44673 5092 44729
rect 5148 44673 5216 44729
rect 5272 44673 5312 44729
rect 4804 44656 5312 44673
rect 4804 44605 4846 44656
rect 4898 44605 4970 44656
rect 5022 44605 5094 44656
rect 5146 44605 5218 44656
rect 5270 44605 5312 44656
rect 4804 44549 4844 44605
rect 4900 44549 4968 44605
rect 5024 44549 5092 44605
rect 5148 44549 5216 44605
rect 5272 44549 5312 44605
rect 4804 41204 5312 44549
rect 4804 41152 4846 41204
rect 4898 41152 4970 41204
rect 5022 41152 5094 41204
rect 5146 41152 5218 41204
rect 5270 41152 5312 41204
rect 4804 41080 5312 41152
rect 4804 41028 4846 41080
rect 4898 41028 4970 41080
rect 5022 41028 5094 41080
rect 5146 41028 5218 41080
rect 5270 41028 5312 41080
rect 4804 40956 5312 41028
rect 4804 40904 4846 40956
rect 4898 40904 4970 40956
rect 5022 40904 5094 40956
rect 5146 40904 5218 40956
rect 5270 40904 5312 40956
rect 4804 40832 5312 40904
rect 4804 40780 4846 40832
rect 4898 40780 4970 40832
rect 5022 40780 5094 40832
rect 5146 40780 5218 40832
rect 5270 40780 5312 40832
rect 4804 40708 5312 40780
rect 4804 40656 4846 40708
rect 4898 40656 4970 40708
rect 5022 40656 5094 40708
rect 5146 40656 5218 40708
rect 5270 40656 5312 40708
rect 4804 37256 5312 40656
rect 4804 37204 4846 37256
rect 4898 37204 4970 37256
rect 5022 37204 5094 37256
rect 5146 37204 5218 37256
rect 5270 37204 5312 37256
rect 4804 37132 5312 37204
rect 4804 37080 4846 37132
rect 4898 37080 4970 37132
rect 5022 37080 5094 37132
rect 5146 37080 5218 37132
rect 5270 37080 5312 37132
rect 4804 37008 5312 37080
rect 4804 36956 4846 37008
rect 4898 36956 4970 37008
rect 5022 36956 5094 37008
rect 5146 36956 5218 37008
rect 5270 36956 5312 37008
rect 4804 36884 5312 36956
rect 4804 36832 4846 36884
rect 4898 36832 4970 36884
rect 5022 36832 5094 36884
rect 5146 36832 5218 36884
rect 5270 36832 5312 36884
rect 4804 36760 5312 36832
rect 4804 36708 4846 36760
rect 4898 36708 4970 36760
rect 5022 36708 5094 36760
rect 5146 36708 5218 36760
rect 5270 36708 5312 36760
rect 4804 36251 5312 36708
rect 4804 36195 4844 36251
rect 4900 36195 4968 36251
rect 5024 36195 5092 36251
rect 5148 36195 5216 36251
rect 5272 36195 5312 36251
rect 4804 36127 5312 36195
rect 4804 36071 4844 36127
rect 4900 36071 4968 36127
rect 5024 36071 5092 36127
rect 5148 36071 5216 36127
rect 5272 36071 5312 36127
rect 4804 36003 5312 36071
rect 4804 35947 4844 36003
rect 4900 35947 4968 36003
rect 5024 35947 5092 36003
rect 5148 35947 5216 36003
rect 5272 35947 5312 36003
rect 4804 35879 5312 35947
rect 4804 35823 4844 35879
rect 4900 35823 4968 35879
rect 5024 35823 5092 35879
rect 5148 35823 5216 35879
rect 5272 35823 5312 35879
rect 4804 35755 5312 35823
rect 4804 35699 4844 35755
rect 4900 35699 4968 35755
rect 5024 35699 5092 35755
rect 5148 35699 5216 35755
rect 5272 35699 5312 35755
rect 4804 35631 5312 35699
rect 4804 35575 4844 35631
rect 4900 35575 4968 35631
rect 5024 35575 5092 35631
rect 5148 35575 5216 35631
rect 5272 35575 5312 35631
rect 4804 35507 5312 35575
rect 4804 35451 4844 35507
rect 4900 35451 4968 35507
rect 5024 35451 5092 35507
rect 5148 35451 5216 35507
rect 5272 35451 5312 35507
rect 4804 35383 5312 35451
rect 4804 35327 4844 35383
rect 4900 35327 4968 35383
rect 5024 35327 5092 35383
rect 5148 35327 5216 35383
rect 5272 35327 5312 35383
rect 4804 35259 5312 35327
rect 4804 35203 4844 35259
rect 4900 35203 4968 35259
rect 5024 35203 5092 35259
rect 5148 35203 5216 35259
rect 5272 35203 5312 35259
rect 4804 35135 5312 35203
rect 4804 35079 4844 35135
rect 4900 35079 4968 35135
rect 5024 35079 5092 35135
rect 5148 35079 5216 35135
rect 5272 35079 5312 35135
rect 4804 35011 5312 35079
rect 4804 34955 4844 35011
rect 4900 34955 4968 35011
rect 5024 34955 5092 35011
rect 5148 34955 5216 35011
rect 5272 34955 5312 35011
rect 4804 34887 5312 34955
rect 4804 34831 4844 34887
rect 4900 34831 4968 34887
rect 5024 34831 5092 34887
rect 5148 34831 5216 34887
rect 5272 34831 5312 34887
rect 4804 34763 5312 34831
rect 4804 34707 4844 34763
rect 4900 34707 4968 34763
rect 5024 34707 5092 34763
rect 5148 34707 5216 34763
rect 5272 34707 5312 34763
rect 4804 34639 5312 34707
rect 4804 34583 4844 34639
rect 4900 34583 4968 34639
rect 5024 34583 5092 34639
rect 5148 34583 5216 34639
rect 5272 34583 5312 34639
rect 4804 34515 5312 34583
rect 4804 34459 4844 34515
rect 4900 34459 4968 34515
rect 5024 34459 5092 34515
rect 5148 34459 5216 34515
rect 5272 34459 5312 34515
rect 4804 34391 5312 34459
rect 4804 34335 4844 34391
rect 4900 34335 4968 34391
rect 5024 34335 5092 34391
rect 5148 34335 5216 34391
rect 5272 34335 5312 34391
rect 4804 34267 5312 34335
rect 4804 34211 4844 34267
rect 4900 34211 4968 34267
rect 5024 34211 5092 34267
rect 5148 34211 5216 34267
rect 5272 34211 5312 34267
rect 4804 34143 5312 34211
rect 4804 34087 4844 34143
rect 4900 34087 4968 34143
rect 5024 34087 5092 34143
rect 5148 34087 5216 34143
rect 5272 34087 5312 34143
rect 4804 34019 5312 34087
rect 4804 33963 4844 34019
rect 4900 33963 4968 34019
rect 5024 33963 5092 34019
rect 5148 33963 5216 34019
rect 5272 33963 5312 34019
rect 4804 33895 5312 33963
rect 4804 33839 4844 33895
rect 4900 33839 4968 33895
rect 5024 33839 5092 33895
rect 5148 33839 5216 33895
rect 5272 33839 5312 33895
rect 4804 33771 5312 33839
rect 4804 33715 4844 33771
rect 4900 33715 4968 33771
rect 5024 33715 5092 33771
rect 5148 33715 5216 33771
rect 5272 33715 5312 33771
rect 4804 33647 5312 33715
rect 4804 33591 4844 33647
rect 4900 33591 4968 33647
rect 5024 33591 5092 33647
rect 5148 33591 5216 33647
rect 5272 33591 5312 33647
rect 4804 33523 5312 33591
rect 4804 33467 4844 33523
rect 4900 33467 4968 33523
rect 5024 33467 5092 33523
rect 5148 33467 5216 33523
rect 5272 33467 5312 33523
rect 4804 33399 5312 33467
rect 4804 33343 4844 33399
rect 4900 33343 4968 33399
rect 5024 33343 5092 33399
rect 5148 33343 5216 33399
rect 5272 33343 5312 33399
rect 4804 33308 5312 33343
rect 4804 33256 4846 33308
rect 4898 33256 4970 33308
rect 5022 33256 5094 33308
rect 5146 33256 5218 33308
rect 5270 33256 5312 33308
rect 4804 33184 5312 33256
rect 4804 33132 4846 33184
rect 4898 33132 4970 33184
rect 5022 33132 5094 33184
rect 5146 33132 5218 33184
rect 5270 33132 5312 33184
rect 4804 33060 5312 33132
rect 4804 33008 4846 33060
rect 4898 33008 4970 33060
rect 5022 33008 5094 33060
rect 5146 33008 5218 33060
rect 5270 33008 5312 33060
rect 4804 32936 5312 33008
rect 4804 32884 4846 32936
rect 4898 32884 4970 32936
rect 5022 32884 5094 32936
rect 5146 32884 5218 32936
rect 5270 32884 5312 32936
rect 4804 32812 5312 32884
rect 4804 32760 4846 32812
rect 4898 32760 4970 32812
rect 5022 32760 5094 32812
rect 5146 32760 5218 32812
rect 5270 32760 5312 32812
rect 4804 29360 5312 32760
rect 4804 29308 4846 29360
rect 4898 29308 4970 29360
rect 5022 29308 5094 29360
rect 5146 29308 5218 29360
rect 5270 29308 5312 29360
rect 4804 29236 5312 29308
rect 4804 29184 4846 29236
rect 4898 29184 4970 29236
rect 5022 29184 5094 29236
rect 5146 29184 5218 29236
rect 5270 29184 5312 29236
rect 4804 29112 5312 29184
rect 4804 29060 4846 29112
rect 4898 29060 4970 29112
rect 5022 29060 5094 29112
rect 5146 29060 5218 29112
rect 5270 29060 5312 29112
rect 4804 28988 5312 29060
rect 4804 28936 4846 28988
rect 4898 28936 4970 28988
rect 5022 28936 5094 28988
rect 5146 28936 5218 28988
rect 5270 28936 5312 28988
rect 4804 28864 5312 28936
rect 4804 28812 4846 28864
rect 4898 28812 4970 28864
rect 5022 28812 5094 28864
rect 5146 28812 5218 28864
rect 5270 28812 5312 28864
rect 4804 28245 5312 28812
rect 4804 28189 4844 28245
rect 4900 28189 4968 28245
rect 5024 28189 5092 28245
rect 5148 28189 5216 28245
rect 5272 28189 5312 28245
rect 4804 28121 5312 28189
rect 4804 28065 4844 28121
rect 4900 28065 4968 28121
rect 5024 28065 5092 28121
rect 5148 28065 5216 28121
rect 5272 28065 5312 28121
rect 4804 27997 5312 28065
rect 4804 27941 4844 27997
rect 4900 27941 4968 27997
rect 5024 27941 5092 27997
rect 5148 27941 5216 27997
rect 5272 27941 5312 27997
rect 4804 27873 5312 27941
rect 4804 27817 4844 27873
rect 4900 27817 4968 27873
rect 5024 27817 5092 27873
rect 5148 27817 5216 27873
rect 5272 27817 5312 27873
rect 4804 27749 5312 27817
rect 4804 27693 4844 27749
rect 4900 27693 4968 27749
rect 5024 27693 5092 27749
rect 5148 27693 5216 27749
rect 5272 27693 5312 27749
rect 4804 27625 5312 27693
rect 4804 27569 4844 27625
rect 4900 27569 4968 27625
rect 5024 27569 5092 27625
rect 5148 27569 5216 27625
rect 5272 27569 5312 27625
rect 4804 27501 5312 27569
rect 4804 27445 4844 27501
rect 4900 27445 4968 27501
rect 5024 27445 5092 27501
rect 5148 27445 5216 27501
rect 5272 27445 5312 27501
rect 4804 27377 5312 27445
rect 4804 27321 4844 27377
rect 4900 27321 4968 27377
rect 5024 27321 5092 27377
rect 5148 27321 5216 27377
rect 5272 27321 5312 27377
rect 4804 27253 5312 27321
rect 4804 27197 4844 27253
rect 4900 27197 4968 27253
rect 5024 27197 5092 27253
rect 5148 27197 5216 27253
rect 5272 27197 5312 27253
rect 4804 27129 5312 27197
rect 4804 27073 4844 27129
rect 4900 27073 4968 27129
rect 5024 27073 5092 27129
rect 5148 27073 5216 27129
rect 5272 27073 5312 27129
rect 4804 27005 5312 27073
rect 4804 26949 4844 27005
rect 4900 26949 4968 27005
rect 5024 26949 5092 27005
rect 5148 26949 5216 27005
rect 5272 26949 5312 27005
rect 4804 25412 5312 26949
rect 4804 25360 4846 25412
rect 4898 25360 4970 25412
rect 5022 25360 5094 25412
rect 5146 25360 5218 25412
rect 5270 25360 5312 25412
rect 4804 25288 5312 25360
rect 4804 25236 4846 25288
rect 4898 25236 4970 25288
rect 5022 25236 5094 25288
rect 5146 25236 5218 25288
rect 5270 25236 5312 25288
rect 4804 25164 5312 25236
rect 4804 25112 4846 25164
rect 4898 25112 4970 25164
rect 5022 25112 5094 25164
rect 5146 25112 5218 25164
rect 5270 25112 5312 25164
rect 4804 25040 5312 25112
rect 4804 24988 4846 25040
rect 4898 24988 4970 25040
rect 5022 24988 5094 25040
rect 5146 24988 5218 25040
rect 5270 24988 5312 25040
rect 4804 24916 5312 24988
rect 4804 24864 4846 24916
rect 4898 24864 4970 24916
rect 5022 24864 5094 24916
rect 5146 24864 5218 24916
rect 5270 24864 5312 24916
rect 4804 21469 5312 24864
rect 4804 21417 4816 21469
rect 4868 21417 4924 21469
rect 4976 21417 5032 21469
rect 5084 21417 5140 21469
rect 5192 21417 5248 21469
rect 5300 21417 5312 21469
rect 4804 21361 5312 21417
rect 4804 21309 4816 21361
rect 4868 21309 4924 21361
rect 4976 21309 5032 21361
rect 5084 21309 5140 21361
rect 5192 21309 5248 21361
rect 5300 21309 5312 21361
rect 4804 21253 5312 21309
rect 4804 21201 4816 21253
rect 4868 21201 4924 21253
rect 4976 21201 5032 21253
rect 5084 21201 5140 21253
rect 5192 21201 5248 21253
rect 5300 21201 5312 21253
rect 4804 19951 5312 21201
rect 4804 19899 4816 19951
rect 4868 19899 4924 19951
rect 4976 19899 5032 19951
rect 5084 19899 5140 19951
rect 5192 19899 5248 19951
rect 5300 19899 5312 19951
rect 4804 19843 5312 19899
rect 4804 19791 4816 19843
rect 4868 19791 4924 19843
rect 4976 19791 5032 19843
rect 5084 19791 5140 19843
rect 5192 19791 5248 19843
rect 5300 19791 5312 19843
rect 4804 19202 5312 19791
rect 4804 19150 4816 19202
rect 4868 19150 4924 19202
rect 4976 19150 5032 19202
rect 5084 19150 5140 19202
rect 5192 19150 5248 19202
rect 5300 19150 5312 19202
rect 4804 19094 5312 19150
rect 4804 19042 4816 19094
rect 4868 19042 4924 19094
rect 4976 19042 5032 19094
rect 5084 19042 5140 19094
rect 5192 19042 5248 19094
rect 5300 19042 5312 19094
rect 4804 18986 5312 19042
rect 4804 18934 4816 18986
rect 4868 18934 4924 18986
rect 4976 18934 5032 18986
rect 5084 18934 5140 18986
rect 5192 18934 5248 18986
rect 5300 18934 5312 18986
rect 4804 18330 5312 18934
rect 4804 18278 4816 18330
rect 4868 18278 4924 18330
rect 4976 18278 5032 18330
rect 5084 18278 5140 18330
rect 5192 18278 5248 18330
rect 5300 18278 5312 18330
rect 4804 18222 5312 18278
rect 4804 18170 4816 18222
rect 4868 18170 4924 18222
rect 4976 18170 5032 18222
rect 5084 18170 5140 18222
rect 5192 18170 5248 18222
rect 5300 18170 5312 18222
rect 4804 18114 5312 18170
rect 4804 18062 4816 18114
rect 4868 18062 4924 18114
rect 4976 18062 5032 18114
rect 5084 18062 5140 18114
rect 5192 18062 5248 18114
rect 5300 18062 5312 18114
rect 4804 17458 5312 18062
rect 4804 17406 4816 17458
rect 4868 17406 4924 17458
rect 4976 17406 5032 17458
rect 5084 17406 5140 17458
rect 5192 17406 5248 17458
rect 5300 17406 5312 17458
rect 4804 17350 5312 17406
rect 4804 17298 4816 17350
rect 4868 17298 4924 17350
rect 4976 17298 5032 17350
rect 5084 17298 5140 17350
rect 5192 17298 5248 17350
rect 5300 17298 5312 17350
rect 4804 17242 5312 17298
rect 4804 17190 4816 17242
rect 4868 17190 4924 17242
rect 4976 17190 5032 17242
rect 5084 17190 5140 17242
rect 5192 17190 5248 17242
rect 5300 17190 5312 17242
rect 4804 16601 5312 17190
rect 4804 16549 4816 16601
rect 4868 16549 4924 16601
rect 4976 16549 5032 16601
rect 5084 16549 5140 16601
rect 5192 16549 5248 16601
rect 5300 16549 5312 16601
rect 4804 16493 5312 16549
rect 4804 16441 4816 16493
rect 4868 16441 4924 16493
rect 4976 16441 5032 16493
rect 5084 16441 5140 16493
rect 5192 16441 5248 16493
rect 5300 16441 5312 16493
rect 4804 15762 5312 16441
rect 5940 56286 6448 56975
rect 5940 56234 6335 56286
rect 6387 56234 6448 56286
rect 5940 56178 6448 56234
rect 5940 56126 6335 56178
rect 6387 56126 6448 56178
rect 5940 56070 6448 56126
rect 5940 56018 6335 56070
rect 6387 56018 6448 56070
rect 5940 55962 6448 56018
rect 5940 55910 6335 55962
rect 6387 55910 6448 55962
rect 5940 55854 6448 55910
rect 5940 55802 6335 55854
rect 6387 55802 6448 55854
rect 5940 55746 6448 55802
rect 5940 55694 6335 55746
rect 6387 55694 6448 55746
rect 5940 55638 6448 55694
rect 5940 55586 6335 55638
rect 6387 55586 6448 55638
rect 5940 55530 6448 55586
rect 5940 55478 6335 55530
rect 6387 55478 6448 55530
rect 5940 55445 6448 55478
rect 5940 55389 5980 55445
rect 6036 55389 6104 55445
rect 6160 55389 6228 55445
rect 6284 55422 6352 55445
rect 6284 55389 6335 55422
rect 6408 55389 6448 55445
rect 5940 55370 6335 55389
rect 6387 55370 6448 55389
rect 5940 55321 6448 55370
rect 5940 55265 5980 55321
rect 6036 55265 6104 55321
rect 6160 55265 6228 55321
rect 6284 55314 6352 55321
rect 6284 55265 6335 55314
rect 6408 55265 6448 55321
rect 5940 55262 6335 55265
rect 6387 55262 6448 55265
rect 5940 55206 6448 55262
rect 5940 55197 6335 55206
rect 6387 55197 6448 55206
rect 5940 55141 5980 55197
rect 6036 55141 6104 55197
rect 6160 55141 6228 55197
rect 6284 55154 6335 55197
rect 6284 55141 6352 55154
rect 6408 55141 6448 55197
rect 5940 55098 6448 55141
rect 5940 55073 6335 55098
rect 6387 55073 6448 55098
rect 5940 55017 5980 55073
rect 6036 55017 6104 55073
rect 6160 55017 6228 55073
rect 6284 55046 6335 55073
rect 6284 55017 6352 55046
rect 6408 55017 6448 55073
rect 5940 54990 6448 55017
rect 5940 54949 6335 54990
rect 6387 54949 6448 54990
rect 5940 54893 5980 54949
rect 6036 54893 6104 54949
rect 6160 54893 6228 54949
rect 6284 54938 6335 54949
rect 6284 54893 6352 54938
rect 6408 54893 6448 54949
rect 5940 54882 6448 54893
rect 5940 54830 6335 54882
rect 6387 54830 6448 54882
rect 5940 54825 6448 54830
rect 5940 54769 5980 54825
rect 6036 54769 6104 54825
rect 6160 54769 6228 54825
rect 6284 54774 6352 54825
rect 6284 54769 6335 54774
rect 6408 54769 6448 54825
rect 5940 54722 6335 54769
rect 6387 54722 6448 54769
rect 5940 54701 6448 54722
rect 5940 54645 5980 54701
rect 6036 54645 6104 54701
rect 6160 54645 6228 54701
rect 6284 54666 6352 54701
rect 6284 54645 6335 54666
rect 6408 54645 6448 54701
rect 5940 54614 6335 54645
rect 6387 54614 6448 54645
rect 5940 54577 6448 54614
rect 5940 54521 5980 54577
rect 6036 54521 6104 54577
rect 6160 54521 6228 54577
rect 6284 54558 6352 54577
rect 6284 54521 6335 54558
rect 6408 54521 6448 54577
rect 5940 54506 6335 54521
rect 6387 54506 6448 54521
rect 5940 54453 6448 54506
rect 5940 54397 5980 54453
rect 6036 54397 6104 54453
rect 6160 54397 6228 54453
rect 6284 54450 6352 54453
rect 6284 54398 6335 54450
rect 6284 54397 6352 54398
rect 6408 54397 6448 54453
rect 5940 54342 6448 54397
rect 5940 54329 6335 54342
rect 6387 54329 6448 54342
rect 5940 54273 5980 54329
rect 6036 54273 6104 54329
rect 6160 54273 6228 54329
rect 6284 54290 6335 54329
rect 6284 54273 6352 54290
rect 6408 54273 6448 54329
rect 5940 54234 6448 54273
rect 5940 54205 6335 54234
rect 6387 54205 6448 54234
rect 5940 54149 5980 54205
rect 6036 54149 6104 54205
rect 6160 54149 6228 54205
rect 6284 54182 6335 54205
rect 6284 54149 6352 54182
rect 6408 54149 6448 54205
rect 5940 54126 6448 54149
rect 5940 54074 6335 54126
rect 6387 54074 6448 54126
rect 5940 54018 6448 54074
rect 5940 53966 6335 54018
rect 6387 53966 6448 54018
rect 5940 53910 6448 53966
rect 5940 53858 6335 53910
rect 6387 53858 6448 53910
rect 5940 53802 6448 53858
rect 5940 53750 6335 53802
rect 6387 53750 6448 53802
rect 5940 53694 6448 53750
rect 5940 53642 6335 53694
rect 6387 53642 6448 53694
rect 5940 53586 6448 53642
rect 5940 53534 6335 53586
rect 6387 53534 6448 53586
rect 5940 53478 6448 53534
rect 5940 53426 6335 53478
rect 6387 53426 6448 53478
rect 5940 53370 6448 53426
rect 5940 53318 6335 53370
rect 6387 53318 6448 53370
rect 5940 53262 6448 53318
rect 5940 53210 6335 53262
rect 6387 53210 6448 53262
rect 5940 52338 6448 53210
rect 5940 52286 6335 52338
rect 6387 52286 6448 52338
rect 5940 52230 6448 52286
rect 5940 52178 6335 52230
rect 6387 52178 6448 52230
rect 5940 52122 6448 52178
rect 5940 52070 6335 52122
rect 6387 52070 6448 52122
rect 5940 52014 6448 52070
rect 5940 51962 6335 52014
rect 6387 51962 6448 52014
rect 5940 51906 6448 51962
rect 5940 51854 6335 51906
rect 6387 51854 6448 51906
rect 5940 51798 6448 51854
rect 5940 51746 6335 51798
rect 6387 51746 6448 51798
rect 5940 51690 6448 51746
rect 5940 51638 6335 51690
rect 6387 51638 6448 51690
rect 5940 51582 6448 51638
rect 5940 51530 6335 51582
rect 6387 51530 6448 51582
rect 5940 51474 6448 51530
rect 5940 51422 6335 51474
rect 6387 51422 6448 51474
rect 5940 51366 6448 51422
rect 5940 51314 6335 51366
rect 6387 51314 6448 51366
rect 5940 51258 6448 51314
rect 5940 51206 6335 51258
rect 6387 51206 6448 51258
rect 5940 51150 6448 51206
rect 5940 51098 6335 51150
rect 6387 51098 6448 51150
rect 5940 51042 6448 51098
rect 5940 50990 6335 51042
rect 6387 50990 6448 51042
rect 5940 50934 6448 50990
rect 5940 50882 6335 50934
rect 6387 50882 6448 50934
rect 5940 50826 6448 50882
rect 5940 50774 6335 50826
rect 6387 50774 6448 50826
rect 5940 50718 6448 50774
rect 5940 50666 6335 50718
rect 6387 50666 6448 50718
rect 5940 50610 6448 50666
rect 5940 50558 6335 50610
rect 6387 50558 6448 50610
rect 5940 50502 6448 50558
rect 5940 50450 6335 50502
rect 6387 50450 6448 50502
rect 5940 50394 6448 50450
rect 5940 50342 6335 50394
rect 6387 50342 6448 50394
rect 5940 50286 6448 50342
rect 5940 50234 6335 50286
rect 6387 50234 6448 50286
rect 5940 50178 6448 50234
rect 5940 50126 6335 50178
rect 6387 50126 6448 50178
rect 5940 50070 6448 50126
rect 5940 50018 6335 50070
rect 6387 50018 6448 50070
rect 5940 49962 6448 50018
rect 5940 49910 6335 49962
rect 6387 49910 6448 49962
rect 5940 49854 6448 49910
rect 5940 49802 6335 49854
rect 6387 49802 6448 49854
rect 5940 49746 6448 49802
rect 5940 49694 6335 49746
rect 6387 49694 6448 49746
rect 5940 49638 6448 49694
rect 5940 49586 6335 49638
rect 6387 49586 6448 49638
rect 5940 49530 6448 49586
rect 5940 49478 6335 49530
rect 6387 49478 6448 49530
rect 5940 49422 6448 49478
rect 5940 49370 6335 49422
rect 6387 49370 6448 49422
rect 5940 49314 6448 49370
rect 5940 49262 6335 49314
rect 6387 49262 6448 49314
rect 5940 48390 6448 49262
rect 5940 48338 6335 48390
rect 6387 48338 6448 48390
rect 5940 48282 6448 48338
rect 5940 48230 6335 48282
rect 6387 48230 6448 48282
rect 5940 48174 6448 48230
rect 5940 48122 6335 48174
rect 6387 48122 6448 48174
rect 5940 48066 6448 48122
rect 5940 48014 6335 48066
rect 6387 48014 6448 48066
rect 5940 47958 6448 48014
rect 5940 47906 6335 47958
rect 6387 47906 6448 47958
rect 5940 47850 6448 47906
rect 5940 47798 6335 47850
rect 6387 47798 6448 47850
rect 5940 47742 6448 47798
rect 5940 47690 6335 47742
rect 6387 47690 6448 47742
rect 5940 47634 6448 47690
rect 5940 47582 6335 47634
rect 6387 47582 6448 47634
rect 5940 47526 6448 47582
rect 5940 47474 6335 47526
rect 6387 47474 6448 47526
rect 5940 47445 6448 47474
rect 5940 47389 5980 47445
rect 6036 47389 6104 47445
rect 6160 47389 6228 47445
rect 6284 47418 6352 47445
rect 6284 47389 6335 47418
rect 6408 47389 6448 47445
rect 5940 47366 6335 47389
rect 6387 47366 6448 47389
rect 5940 47321 6448 47366
rect 5940 47265 5980 47321
rect 6036 47265 6104 47321
rect 6160 47265 6228 47321
rect 6284 47310 6352 47321
rect 6284 47265 6335 47310
rect 6408 47265 6448 47321
rect 5940 47258 6335 47265
rect 6387 47258 6448 47265
rect 5940 47202 6448 47258
rect 5940 47197 6335 47202
rect 6387 47197 6448 47202
rect 5940 47141 5980 47197
rect 6036 47141 6104 47197
rect 6160 47141 6228 47197
rect 6284 47150 6335 47197
rect 6284 47141 6352 47150
rect 6408 47141 6448 47197
rect 5940 47094 6448 47141
rect 5940 47073 6335 47094
rect 6387 47073 6448 47094
rect 5940 47017 5980 47073
rect 6036 47017 6104 47073
rect 6160 47017 6228 47073
rect 6284 47042 6335 47073
rect 6284 47017 6352 47042
rect 6408 47017 6448 47073
rect 5940 46986 6448 47017
rect 5940 46949 6335 46986
rect 6387 46949 6448 46986
rect 5940 46893 5980 46949
rect 6036 46893 6104 46949
rect 6160 46893 6228 46949
rect 6284 46934 6335 46949
rect 6284 46893 6352 46934
rect 6408 46893 6448 46949
rect 5940 46878 6448 46893
rect 5940 46826 6335 46878
rect 6387 46826 6448 46878
rect 5940 46825 6448 46826
rect 5940 46769 5980 46825
rect 6036 46769 6104 46825
rect 6160 46769 6228 46825
rect 6284 46770 6352 46825
rect 6284 46769 6335 46770
rect 6408 46769 6448 46825
rect 5940 46718 6335 46769
rect 6387 46718 6448 46769
rect 5940 46701 6448 46718
rect 5940 46645 5980 46701
rect 6036 46645 6104 46701
rect 6160 46645 6228 46701
rect 6284 46662 6352 46701
rect 6284 46645 6335 46662
rect 6408 46645 6448 46701
rect 5940 46610 6335 46645
rect 6387 46610 6448 46645
rect 5940 46577 6448 46610
rect 5940 46521 5980 46577
rect 6036 46521 6104 46577
rect 6160 46521 6228 46577
rect 6284 46554 6352 46577
rect 6284 46521 6335 46554
rect 6408 46521 6448 46577
rect 5940 46502 6335 46521
rect 6387 46502 6448 46521
rect 5940 46453 6448 46502
rect 5940 46397 5980 46453
rect 6036 46397 6104 46453
rect 6160 46397 6228 46453
rect 6284 46446 6352 46453
rect 6284 46397 6335 46446
rect 6408 46397 6448 46453
rect 5940 46394 6335 46397
rect 6387 46394 6448 46397
rect 5940 46338 6448 46394
rect 5940 46329 6335 46338
rect 6387 46329 6448 46338
rect 5940 46273 5980 46329
rect 6036 46273 6104 46329
rect 6160 46273 6228 46329
rect 6284 46286 6335 46329
rect 6284 46273 6352 46286
rect 6408 46273 6448 46329
rect 5940 46230 6448 46273
rect 5940 46205 6335 46230
rect 6387 46205 6448 46230
rect 5940 46149 5980 46205
rect 6036 46149 6104 46205
rect 6160 46149 6228 46205
rect 6284 46178 6335 46205
rect 6284 46149 6352 46178
rect 6408 46149 6448 46205
rect 5940 46122 6448 46149
rect 5940 46070 6335 46122
rect 6387 46070 6448 46122
rect 5940 46014 6448 46070
rect 5940 45962 6335 46014
rect 6387 45962 6448 46014
rect 5940 45906 6448 45962
rect 5940 45854 6335 45906
rect 6387 45854 6448 45906
rect 5940 45798 6448 45854
rect 5940 45746 6335 45798
rect 6387 45746 6448 45798
rect 5940 45690 6448 45746
rect 5940 45638 6335 45690
rect 6387 45638 6448 45690
rect 5940 45582 6448 45638
rect 5940 45530 6335 45582
rect 6387 45530 6448 45582
rect 5940 45474 6448 45530
rect 5940 45422 6335 45474
rect 6387 45422 6448 45474
rect 5940 45366 6448 45422
rect 5940 45314 6335 45366
rect 6387 45314 6448 45366
rect 5940 44442 6448 45314
rect 5940 44390 6335 44442
rect 6387 44390 6448 44442
rect 5940 44334 6448 44390
rect 5940 44282 6335 44334
rect 6387 44282 6448 44334
rect 5940 44245 6448 44282
rect 5940 44189 5980 44245
rect 6036 44189 6104 44245
rect 6160 44189 6228 44245
rect 6284 44226 6352 44245
rect 6284 44189 6335 44226
rect 6408 44189 6448 44245
rect 5940 44174 6335 44189
rect 6387 44174 6448 44189
rect 5940 44121 6448 44174
rect 5940 44065 5980 44121
rect 6036 44065 6104 44121
rect 6160 44065 6228 44121
rect 6284 44118 6352 44121
rect 6284 44066 6335 44118
rect 6284 44065 6352 44066
rect 6408 44065 6448 44121
rect 5940 44010 6448 44065
rect 5940 43997 6335 44010
rect 6387 43997 6448 44010
rect 5940 43941 5980 43997
rect 6036 43941 6104 43997
rect 6160 43941 6228 43997
rect 6284 43958 6335 43997
rect 6284 43941 6352 43958
rect 6408 43941 6448 43997
rect 5940 43902 6448 43941
rect 5940 43873 6335 43902
rect 6387 43873 6448 43902
rect 5940 43817 5980 43873
rect 6036 43817 6104 43873
rect 6160 43817 6228 43873
rect 6284 43850 6335 43873
rect 6284 43817 6352 43850
rect 6408 43817 6448 43873
rect 5940 43794 6448 43817
rect 5940 43749 6335 43794
rect 6387 43749 6448 43794
rect 5940 43693 5980 43749
rect 6036 43693 6104 43749
rect 6160 43693 6228 43749
rect 6284 43742 6335 43749
rect 6284 43693 6352 43742
rect 6408 43693 6448 43749
rect 5940 43686 6448 43693
rect 5940 43634 6335 43686
rect 6387 43634 6448 43686
rect 5940 43625 6448 43634
rect 5940 43569 5980 43625
rect 6036 43569 6104 43625
rect 6160 43569 6228 43625
rect 6284 43578 6352 43625
rect 6284 43569 6335 43578
rect 6408 43569 6448 43625
rect 5940 43526 6335 43569
rect 6387 43526 6448 43569
rect 5940 43501 6448 43526
rect 5940 43445 5980 43501
rect 6036 43445 6104 43501
rect 6160 43445 6228 43501
rect 6284 43470 6352 43501
rect 6284 43445 6335 43470
rect 6408 43445 6448 43501
rect 5940 43418 6335 43445
rect 6387 43418 6448 43445
rect 5940 43377 6448 43418
rect 5940 43321 5980 43377
rect 6036 43321 6104 43377
rect 6160 43321 6228 43377
rect 6284 43362 6352 43377
rect 6284 43321 6335 43362
rect 6408 43321 6448 43377
rect 5940 43310 6335 43321
rect 6387 43310 6448 43321
rect 5940 43254 6448 43310
rect 5940 43253 6335 43254
rect 6387 43253 6448 43254
rect 5940 43197 5980 43253
rect 6036 43197 6104 43253
rect 6160 43197 6228 43253
rect 6284 43202 6335 43253
rect 6284 43197 6352 43202
rect 6408 43197 6448 43253
rect 5940 43146 6448 43197
rect 5940 43129 6335 43146
rect 6387 43129 6448 43146
rect 5940 43073 5980 43129
rect 6036 43073 6104 43129
rect 6160 43073 6228 43129
rect 6284 43094 6335 43129
rect 6284 43073 6352 43094
rect 6408 43073 6448 43129
rect 5940 43038 6448 43073
rect 5940 43005 6335 43038
rect 6387 43005 6448 43038
rect 5940 42949 5980 43005
rect 6036 42949 6104 43005
rect 6160 42949 6228 43005
rect 6284 42986 6335 43005
rect 6284 42949 6352 42986
rect 6408 42949 6448 43005
rect 5940 42930 6448 42949
rect 5940 42878 6335 42930
rect 6387 42878 6448 42930
rect 5940 42822 6448 42878
rect 5940 42770 6335 42822
rect 6387 42770 6448 42822
rect 5940 42714 6448 42770
rect 5940 42662 6335 42714
rect 6387 42662 6448 42714
rect 5940 42645 6448 42662
rect 5940 42589 5980 42645
rect 6036 42589 6104 42645
rect 6160 42589 6228 42645
rect 6284 42606 6352 42645
rect 6284 42589 6335 42606
rect 6408 42589 6448 42645
rect 5940 42554 6335 42589
rect 6387 42554 6448 42589
rect 5940 42521 6448 42554
rect 5940 42465 5980 42521
rect 6036 42465 6104 42521
rect 6160 42465 6228 42521
rect 6284 42498 6352 42521
rect 6284 42465 6335 42498
rect 6408 42465 6448 42521
rect 5940 42446 6335 42465
rect 6387 42446 6448 42465
rect 5940 42397 6448 42446
rect 5940 42341 5980 42397
rect 6036 42341 6104 42397
rect 6160 42341 6228 42397
rect 6284 42390 6352 42397
rect 6284 42341 6335 42390
rect 6408 42341 6448 42397
rect 5940 42338 6335 42341
rect 6387 42338 6448 42341
rect 5940 42282 6448 42338
rect 5940 42273 6335 42282
rect 6387 42273 6448 42282
rect 5940 42217 5980 42273
rect 6036 42217 6104 42273
rect 6160 42217 6228 42273
rect 6284 42230 6335 42273
rect 6284 42217 6352 42230
rect 6408 42217 6448 42273
rect 5940 42174 6448 42217
rect 5940 42149 6335 42174
rect 6387 42149 6448 42174
rect 5940 42093 5980 42149
rect 6036 42093 6104 42149
rect 6160 42093 6228 42149
rect 6284 42122 6335 42149
rect 6284 42093 6352 42122
rect 6408 42093 6448 42149
rect 5940 42066 6448 42093
rect 5940 42025 6335 42066
rect 6387 42025 6448 42066
rect 5940 41969 5980 42025
rect 6036 41969 6104 42025
rect 6160 41969 6228 42025
rect 6284 42014 6335 42025
rect 6284 41969 6352 42014
rect 6408 41969 6448 42025
rect 5940 41958 6448 41969
rect 5940 41906 6335 41958
rect 6387 41906 6448 41958
rect 5940 41901 6448 41906
rect 5940 41845 5980 41901
rect 6036 41845 6104 41901
rect 6160 41845 6228 41901
rect 6284 41850 6352 41901
rect 6284 41845 6335 41850
rect 6408 41845 6448 41901
rect 5940 41798 6335 41845
rect 6387 41798 6448 41845
rect 5940 41777 6448 41798
rect 5940 41721 5980 41777
rect 6036 41721 6104 41777
rect 6160 41721 6228 41777
rect 6284 41742 6352 41777
rect 6284 41721 6335 41742
rect 6408 41721 6448 41777
rect 5940 41690 6335 41721
rect 6387 41690 6448 41721
rect 5940 41653 6448 41690
rect 5940 41597 5980 41653
rect 6036 41597 6104 41653
rect 6160 41597 6228 41653
rect 6284 41634 6352 41653
rect 6284 41597 6335 41634
rect 6408 41597 6448 41653
rect 5940 41582 6335 41597
rect 6387 41582 6448 41597
rect 5940 41529 6448 41582
rect 5940 41473 5980 41529
rect 6036 41473 6104 41529
rect 6160 41473 6228 41529
rect 6284 41526 6352 41529
rect 6284 41474 6335 41526
rect 6284 41473 6352 41474
rect 6408 41473 6448 41529
rect 5940 41418 6448 41473
rect 5940 41405 6335 41418
rect 6387 41405 6448 41418
rect 5940 41349 5980 41405
rect 6036 41349 6104 41405
rect 6160 41349 6228 41405
rect 6284 41366 6335 41405
rect 6284 41349 6352 41366
rect 6408 41349 6448 41405
rect 5940 41045 6448 41349
rect 5940 40989 5980 41045
rect 6036 40989 6104 41045
rect 6160 40989 6228 41045
rect 6284 40989 6352 41045
rect 6408 40989 6448 41045
rect 5940 40921 6448 40989
rect 5940 40865 5980 40921
rect 6036 40865 6104 40921
rect 6160 40865 6228 40921
rect 6284 40865 6352 40921
rect 6408 40865 6448 40921
rect 5940 40797 6448 40865
rect 5940 40741 5980 40797
rect 6036 40741 6104 40797
rect 6160 40741 6228 40797
rect 6284 40741 6352 40797
rect 6408 40741 6448 40797
rect 5940 40673 6448 40741
rect 5940 40617 5980 40673
rect 6036 40617 6104 40673
rect 6160 40617 6228 40673
rect 6284 40617 6352 40673
rect 6408 40617 6448 40673
rect 5940 40549 6448 40617
rect 5940 40493 5980 40549
rect 6036 40493 6104 40549
rect 6160 40493 6228 40549
rect 6284 40494 6352 40549
rect 6284 40493 6335 40494
rect 6408 40493 6448 40549
rect 5940 40442 6335 40493
rect 6387 40442 6448 40493
rect 5940 40425 6448 40442
rect 5940 40369 5980 40425
rect 6036 40369 6104 40425
rect 6160 40369 6228 40425
rect 6284 40386 6352 40425
rect 6284 40369 6335 40386
rect 6408 40369 6448 40425
rect 5940 40334 6335 40369
rect 6387 40334 6448 40369
rect 5940 40301 6448 40334
rect 5940 40245 5980 40301
rect 6036 40245 6104 40301
rect 6160 40245 6228 40301
rect 6284 40278 6352 40301
rect 6284 40245 6335 40278
rect 6408 40245 6448 40301
rect 5940 40226 6335 40245
rect 6387 40226 6448 40245
rect 5940 40177 6448 40226
rect 5940 40121 5980 40177
rect 6036 40121 6104 40177
rect 6160 40121 6228 40177
rect 6284 40170 6352 40177
rect 6284 40121 6335 40170
rect 6408 40121 6448 40177
rect 5940 40118 6335 40121
rect 6387 40118 6448 40121
rect 5940 40062 6448 40118
rect 5940 40053 6335 40062
rect 6387 40053 6448 40062
rect 5940 39997 5980 40053
rect 6036 39997 6104 40053
rect 6160 39997 6228 40053
rect 6284 40010 6335 40053
rect 6284 39997 6352 40010
rect 6408 39997 6448 40053
rect 5940 39954 6448 39997
rect 5940 39929 6335 39954
rect 6387 39929 6448 39954
rect 5940 39873 5980 39929
rect 6036 39873 6104 39929
rect 6160 39873 6228 39929
rect 6284 39902 6335 39929
rect 6284 39873 6352 39902
rect 6408 39873 6448 39929
rect 5940 39846 6448 39873
rect 5940 39805 6335 39846
rect 6387 39805 6448 39846
rect 5940 39749 5980 39805
rect 6036 39749 6104 39805
rect 6160 39749 6228 39805
rect 6284 39794 6335 39805
rect 6284 39749 6352 39794
rect 6408 39749 6448 39805
rect 5940 39738 6448 39749
rect 5940 39686 6335 39738
rect 6387 39686 6448 39738
rect 5940 39630 6448 39686
rect 5940 39578 6335 39630
rect 6387 39578 6448 39630
rect 5940 39522 6448 39578
rect 5940 39470 6335 39522
rect 6387 39470 6448 39522
rect 5940 39414 6448 39470
rect 5940 39362 6335 39414
rect 6387 39362 6448 39414
rect 5940 39306 6448 39362
rect 5940 39254 6335 39306
rect 6387 39254 6448 39306
rect 5940 39198 6448 39254
rect 5940 39146 6335 39198
rect 6387 39146 6448 39198
rect 5940 39090 6448 39146
rect 5940 39038 6335 39090
rect 6387 39038 6448 39090
rect 5940 38982 6448 39038
rect 5940 38930 6335 38982
rect 6387 38930 6448 38982
rect 5940 38874 6448 38930
rect 5940 38822 6335 38874
rect 6387 38822 6448 38874
rect 5940 38766 6448 38822
rect 5940 38714 6335 38766
rect 6387 38714 6448 38766
rect 5940 38658 6448 38714
rect 5940 38606 6335 38658
rect 6387 38606 6448 38658
rect 5940 38550 6448 38606
rect 5940 38498 6335 38550
rect 6387 38498 6448 38550
rect 5940 38442 6448 38498
rect 5940 38390 6335 38442
rect 6387 38390 6448 38442
rect 5940 38334 6448 38390
rect 5940 38282 6335 38334
rect 6387 38282 6448 38334
rect 5940 38226 6448 38282
rect 5940 38174 6335 38226
rect 6387 38174 6448 38226
rect 5940 38118 6448 38174
rect 5940 38066 6335 38118
rect 6387 38066 6448 38118
rect 5940 38010 6448 38066
rect 5940 37958 6335 38010
rect 6387 37958 6448 38010
rect 5940 37902 6448 37958
rect 5940 37850 6335 37902
rect 6387 37850 6448 37902
rect 5940 37794 6448 37850
rect 5940 37742 6335 37794
rect 6387 37742 6448 37794
rect 5940 37686 6448 37742
rect 5940 37634 6335 37686
rect 6387 37634 6448 37686
rect 5940 37578 6448 37634
rect 5940 37526 6335 37578
rect 6387 37526 6448 37578
rect 5940 37470 6448 37526
rect 5940 37418 6335 37470
rect 6387 37418 6448 37470
rect 5940 36546 6448 37418
rect 5940 36494 6335 36546
rect 6387 36494 6448 36546
rect 5940 36438 6448 36494
rect 5940 36386 6335 36438
rect 6387 36386 6448 36438
rect 5940 36330 6448 36386
rect 5940 36278 6335 36330
rect 6387 36278 6448 36330
rect 5940 36222 6448 36278
rect 5940 36170 6335 36222
rect 6387 36170 6448 36222
rect 5940 36114 6448 36170
rect 5940 36062 6335 36114
rect 6387 36062 6448 36114
rect 5940 36006 6448 36062
rect 5940 35954 6335 36006
rect 6387 35954 6448 36006
rect 5940 35898 6448 35954
rect 5940 35846 6335 35898
rect 6387 35846 6448 35898
rect 5940 35790 6448 35846
rect 5940 35738 6335 35790
rect 6387 35738 6448 35790
rect 5940 35682 6448 35738
rect 5940 35630 6335 35682
rect 6387 35630 6448 35682
rect 5940 35574 6448 35630
rect 5940 35522 6335 35574
rect 6387 35522 6448 35574
rect 5940 35466 6448 35522
rect 5940 35414 6335 35466
rect 6387 35414 6448 35466
rect 5940 35358 6448 35414
rect 5940 35306 6335 35358
rect 6387 35306 6448 35358
rect 5940 35250 6448 35306
rect 5940 35198 6335 35250
rect 6387 35198 6448 35250
rect 5940 35142 6448 35198
rect 5940 35090 6335 35142
rect 6387 35090 6448 35142
rect 5940 35034 6448 35090
rect 5940 34982 6335 35034
rect 6387 34982 6448 35034
rect 5940 34926 6448 34982
rect 5940 34874 6335 34926
rect 6387 34874 6448 34926
rect 5940 34818 6448 34874
rect 5940 34766 6335 34818
rect 6387 34766 6448 34818
rect 5940 34710 6448 34766
rect 5940 34658 6335 34710
rect 6387 34658 6448 34710
rect 5940 34602 6448 34658
rect 5940 34550 6335 34602
rect 6387 34550 6448 34602
rect 5940 34494 6448 34550
rect 5940 34442 6335 34494
rect 6387 34442 6448 34494
rect 5940 34386 6448 34442
rect 5940 34334 6335 34386
rect 6387 34334 6448 34386
rect 5940 34278 6448 34334
rect 5940 34226 6335 34278
rect 6387 34226 6448 34278
rect 5940 34170 6448 34226
rect 5940 34118 6335 34170
rect 6387 34118 6448 34170
rect 5940 34062 6448 34118
rect 5940 34010 6335 34062
rect 6387 34010 6448 34062
rect 5940 33954 6448 34010
rect 5940 33902 6335 33954
rect 6387 33902 6448 33954
rect 5940 33846 6448 33902
rect 5940 33794 6335 33846
rect 6387 33794 6448 33846
rect 5940 33738 6448 33794
rect 5940 33686 6335 33738
rect 6387 33686 6448 33738
rect 5940 33630 6448 33686
rect 5940 33578 6335 33630
rect 6387 33578 6448 33630
rect 5940 33522 6448 33578
rect 5940 33470 6335 33522
rect 6387 33470 6448 33522
rect 5940 33051 6448 33470
rect 5940 32995 5980 33051
rect 6036 32995 6104 33051
rect 6160 32995 6228 33051
rect 6284 32995 6352 33051
rect 6408 32995 6448 33051
rect 5940 32927 6448 32995
rect 5940 32871 5980 32927
rect 6036 32871 6104 32927
rect 6160 32871 6228 32927
rect 6284 32871 6352 32927
rect 6408 32871 6448 32927
rect 5940 32803 6448 32871
rect 5940 32747 5980 32803
rect 6036 32747 6104 32803
rect 6160 32747 6228 32803
rect 6284 32747 6352 32803
rect 6408 32747 6448 32803
rect 5940 32679 6448 32747
rect 5940 32623 5980 32679
rect 6036 32623 6104 32679
rect 6160 32623 6228 32679
rect 6284 32623 6352 32679
rect 6408 32623 6448 32679
rect 5940 32598 6448 32623
rect 5940 32555 6335 32598
rect 6387 32555 6448 32598
rect 5940 32499 5980 32555
rect 6036 32499 6104 32555
rect 6160 32499 6228 32555
rect 6284 32546 6335 32555
rect 6284 32499 6352 32546
rect 6408 32499 6448 32555
rect 5940 32490 6448 32499
rect 5940 32438 6335 32490
rect 6387 32438 6448 32490
rect 5940 32431 6448 32438
rect 5940 32375 5980 32431
rect 6036 32375 6104 32431
rect 6160 32375 6228 32431
rect 6284 32382 6352 32431
rect 6284 32375 6335 32382
rect 6408 32375 6448 32431
rect 5940 32330 6335 32375
rect 6387 32330 6448 32375
rect 5940 32307 6448 32330
rect 5940 32251 5980 32307
rect 6036 32251 6104 32307
rect 6160 32251 6228 32307
rect 6284 32274 6352 32307
rect 6284 32251 6335 32274
rect 6408 32251 6448 32307
rect 5940 32222 6335 32251
rect 6387 32222 6448 32251
rect 5940 32183 6448 32222
rect 5940 32127 5980 32183
rect 6036 32127 6104 32183
rect 6160 32127 6228 32183
rect 6284 32166 6352 32183
rect 6284 32127 6335 32166
rect 6408 32127 6448 32183
rect 5940 32114 6335 32127
rect 6387 32114 6448 32127
rect 5940 32059 6448 32114
rect 5940 32003 5980 32059
rect 6036 32003 6104 32059
rect 6160 32003 6228 32059
rect 6284 32058 6352 32059
rect 6284 32006 6335 32058
rect 6284 32003 6352 32006
rect 6408 32003 6448 32059
rect 5940 31950 6448 32003
rect 5940 31935 6335 31950
rect 6387 31935 6448 31950
rect 5940 31879 5980 31935
rect 6036 31879 6104 31935
rect 6160 31879 6228 31935
rect 6284 31898 6335 31935
rect 6284 31879 6352 31898
rect 6408 31879 6448 31935
rect 5940 31842 6448 31879
rect 5940 31811 6335 31842
rect 6387 31811 6448 31842
rect 5940 31755 5980 31811
rect 6036 31755 6104 31811
rect 6160 31755 6228 31811
rect 6284 31790 6335 31811
rect 6284 31755 6352 31790
rect 6408 31755 6448 31811
rect 5940 31734 6448 31755
rect 5940 31687 6335 31734
rect 6387 31687 6448 31734
rect 5940 31631 5980 31687
rect 6036 31631 6104 31687
rect 6160 31631 6228 31687
rect 6284 31682 6335 31687
rect 6284 31631 6352 31682
rect 6408 31631 6448 31687
rect 5940 31626 6448 31631
rect 5940 31574 6335 31626
rect 6387 31574 6448 31626
rect 5940 31563 6448 31574
rect 5940 31507 5980 31563
rect 6036 31507 6104 31563
rect 6160 31507 6228 31563
rect 6284 31518 6352 31563
rect 6284 31507 6335 31518
rect 6408 31507 6448 31563
rect 5940 31466 6335 31507
rect 6387 31466 6448 31507
rect 5940 31439 6448 31466
rect 5940 31383 5980 31439
rect 6036 31383 6104 31439
rect 6160 31383 6228 31439
rect 6284 31410 6352 31439
rect 6284 31383 6335 31410
rect 6408 31383 6448 31439
rect 5940 31358 6335 31383
rect 6387 31358 6448 31383
rect 5940 31315 6448 31358
rect 5940 31259 5980 31315
rect 6036 31259 6104 31315
rect 6160 31259 6228 31315
rect 6284 31302 6352 31315
rect 6284 31259 6335 31302
rect 6408 31259 6448 31315
rect 5940 31250 6335 31259
rect 6387 31250 6448 31259
rect 5940 31194 6448 31250
rect 5940 31191 6335 31194
rect 6387 31191 6448 31194
rect 5940 31135 5980 31191
rect 6036 31135 6104 31191
rect 6160 31135 6228 31191
rect 6284 31142 6335 31191
rect 6284 31135 6352 31142
rect 6408 31135 6448 31191
rect 5940 31086 6448 31135
rect 5940 31067 6335 31086
rect 6387 31067 6448 31086
rect 5940 31011 5980 31067
rect 6036 31011 6104 31067
rect 6160 31011 6228 31067
rect 6284 31034 6335 31067
rect 6284 31011 6352 31034
rect 6408 31011 6448 31067
rect 5940 30978 6448 31011
rect 5940 30943 6335 30978
rect 6387 30943 6448 30978
rect 5940 30887 5980 30943
rect 6036 30887 6104 30943
rect 6160 30887 6228 30943
rect 6284 30926 6335 30943
rect 6284 30887 6352 30926
rect 6408 30887 6448 30943
rect 5940 30870 6448 30887
rect 5940 30819 6335 30870
rect 6387 30819 6448 30870
rect 5940 30763 5980 30819
rect 6036 30763 6104 30819
rect 6160 30763 6228 30819
rect 6284 30818 6335 30819
rect 6284 30763 6352 30818
rect 6408 30763 6448 30819
rect 5940 30762 6448 30763
rect 5940 30710 6335 30762
rect 6387 30710 6448 30762
rect 5940 30695 6448 30710
rect 5940 30639 5980 30695
rect 6036 30639 6104 30695
rect 6160 30639 6228 30695
rect 6284 30654 6352 30695
rect 6284 30639 6335 30654
rect 6408 30639 6448 30695
rect 5940 30602 6335 30639
rect 6387 30602 6448 30639
rect 5940 30571 6448 30602
rect 5940 30515 5980 30571
rect 6036 30515 6104 30571
rect 6160 30515 6228 30571
rect 6284 30546 6352 30571
rect 6284 30515 6335 30546
rect 6408 30515 6448 30571
rect 5940 30494 6335 30515
rect 6387 30494 6448 30515
rect 5940 30447 6448 30494
rect 5940 30391 5980 30447
rect 6036 30391 6104 30447
rect 6160 30391 6228 30447
rect 6284 30438 6352 30447
rect 6284 30391 6335 30438
rect 6408 30391 6448 30447
rect 5940 30386 6335 30391
rect 6387 30386 6448 30391
rect 5940 30330 6448 30386
rect 5940 30323 6335 30330
rect 6387 30323 6448 30330
rect 5940 30267 5980 30323
rect 6036 30267 6104 30323
rect 6160 30267 6228 30323
rect 6284 30278 6335 30323
rect 6284 30267 6352 30278
rect 6408 30267 6448 30323
rect 5940 30222 6448 30267
rect 5940 30199 6335 30222
rect 6387 30199 6448 30222
rect 5940 30143 5980 30199
rect 6036 30143 6104 30199
rect 6160 30143 6228 30199
rect 6284 30170 6335 30199
rect 6284 30143 6352 30170
rect 6408 30143 6448 30199
rect 5940 30114 6448 30143
rect 5940 30062 6335 30114
rect 6387 30062 6448 30114
rect 5940 30006 6448 30062
rect 5940 29954 6335 30006
rect 6387 29954 6448 30006
rect 5940 29898 6448 29954
rect 5940 29846 6335 29898
rect 6387 29846 6448 29898
rect 5940 29845 6448 29846
rect 5940 29789 5980 29845
rect 6036 29789 6104 29845
rect 6160 29789 6228 29845
rect 6284 29790 6352 29845
rect 6284 29789 6335 29790
rect 6408 29789 6448 29845
rect 5940 29738 6335 29789
rect 6387 29738 6448 29789
rect 5940 29721 6448 29738
rect 5940 29665 5980 29721
rect 6036 29665 6104 29721
rect 6160 29665 6228 29721
rect 6284 29682 6352 29721
rect 6284 29665 6335 29682
rect 6408 29665 6448 29721
rect 5940 29630 6335 29665
rect 6387 29630 6448 29665
rect 5940 29597 6448 29630
rect 5940 29541 5980 29597
rect 6036 29541 6104 29597
rect 6160 29541 6228 29597
rect 6284 29574 6352 29597
rect 6284 29541 6335 29574
rect 6408 29541 6448 29597
rect 5940 29522 6335 29541
rect 6387 29522 6448 29541
rect 5940 29473 6448 29522
rect 5940 29417 5980 29473
rect 6036 29417 6104 29473
rect 6160 29417 6228 29473
rect 6284 29417 6352 29473
rect 6408 29417 6448 29473
rect 5940 29349 6448 29417
rect 5940 29293 5980 29349
rect 6036 29293 6104 29349
rect 6160 29293 6228 29349
rect 6284 29293 6352 29349
rect 6408 29293 6448 29349
rect 5940 29225 6448 29293
rect 5940 29169 5980 29225
rect 6036 29169 6104 29225
rect 6160 29169 6228 29225
rect 6284 29169 6352 29225
rect 6408 29169 6448 29225
rect 5940 29101 6448 29169
rect 5940 29045 5980 29101
rect 6036 29045 6104 29101
rect 6160 29045 6228 29101
rect 6284 29045 6352 29101
rect 6408 29045 6448 29101
rect 5940 28977 6448 29045
rect 5940 28921 5980 28977
rect 6036 28921 6104 28977
rect 6160 28921 6228 28977
rect 6284 28921 6352 28977
rect 6408 28921 6448 28977
rect 5940 28853 6448 28921
rect 5940 28797 5980 28853
rect 6036 28797 6104 28853
rect 6160 28797 6228 28853
rect 6284 28797 6352 28853
rect 6408 28797 6448 28853
rect 5940 28729 6448 28797
rect 5940 28673 5980 28729
rect 6036 28673 6104 28729
rect 6160 28673 6228 28729
rect 6284 28673 6352 28729
rect 6408 28673 6448 28729
rect 5940 28650 6448 28673
rect 5940 28605 6335 28650
rect 6387 28605 6448 28650
rect 5940 28549 5980 28605
rect 6036 28549 6104 28605
rect 6160 28549 6228 28605
rect 6284 28598 6335 28605
rect 6284 28549 6352 28598
rect 6408 28549 6448 28605
rect 5940 28542 6448 28549
rect 5940 28490 6335 28542
rect 6387 28490 6448 28542
rect 5940 28434 6448 28490
rect 5940 28382 6335 28434
rect 6387 28382 6448 28434
rect 5940 28326 6448 28382
rect 5940 28274 6335 28326
rect 6387 28274 6448 28326
rect 5940 28218 6448 28274
rect 5940 28166 6335 28218
rect 6387 28166 6448 28218
rect 5940 28110 6448 28166
rect 5940 28058 6335 28110
rect 6387 28058 6448 28110
rect 5940 28002 6448 28058
rect 5940 27950 6335 28002
rect 6387 27950 6448 28002
rect 5940 27894 6448 27950
rect 5940 27842 6335 27894
rect 6387 27842 6448 27894
rect 5940 27786 6448 27842
rect 5940 27734 6335 27786
rect 6387 27734 6448 27786
rect 5940 27678 6448 27734
rect 5940 27626 6335 27678
rect 6387 27626 6448 27678
rect 5940 27570 6448 27626
rect 5940 27518 6335 27570
rect 6387 27518 6448 27570
rect 5940 27462 6448 27518
rect 5940 27410 6335 27462
rect 6387 27410 6448 27462
rect 5940 27354 6448 27410
rect 5940 27302 6335 27354
rect 6387 27302 6448 27354
rect 5940 27246 6448 27302
rect 5940 27194 6335 27246
rect 6387 27194 6448 27246
rect 5940 27138 6448 27194
rect 5940 27086 6335 27138
rect 6387 27086 6448 27138
rect 5940 27030 6448 27086
rect 5940 26978 6335 27030
rect 6387 26978 6448 27030
rect 5940 26922 6448 26978
rect 5940 26870 6335 26922
rect 6387 26870 6448 26922
rect 5940 26814 6448 26870
rect 5940 26762 6335 26814
rect 6387 26762 6448 26814
rect 5940 26706 6448 26762
rect 5940 26654 6335 26706
rect 6387 26654 6448 26706
rect 5940 26651 6448 26654
rect 5940 26595 5980 26651
rect 6036 26595 6104 26651
rect 6160 26595 6228 26651
rect 6284 26598 6352 26651
rect 6284 26595 6335 26598
rect 6408 26595 6448 26651
rect 5940 26546 6335 26595
rect 6387 26546 6448 26595
rect 5940 26527 6448 26546
rect 5940 26471 5980 26527
rect 6036 26471 6104 26527
rect 6160 26471 6228 26527
rect 6284 26490 6352 26527
rect 6284 26471 6335 26490
rect 6408 26471 6448 26527
rect 5940 26438 6335 26471
rect 6387 26438 6448 26471
rect 5940 26403 6448 26438
rect 5940 26347 5980 26403
rect 6036 26347 6104 26403
rect 6160 26347 6228 26403
rect 6284 26382 6352 26403
rect 6284 26347 6335 26382
rect 6408 26347 6448 26403
rect 5940 26330 6335 26347
rect 6387 26330 6448 26347
rect 5940 26279 6448 26330
rect 5940 26223 5980 26279
rect 6036 26223 6104 26279
rect 6160 26223 6228 26279
rect 6284 26274 6352 26279
rect 6284 26223 6335 26274
rect 6408 26223 6448 26279
rect 5940 26222 6335 26223
rect 6387 26222 6448 26223
rect 5940 26166 6448 26222
rect 5940 26155 6335 26166
rect 6387 26155 6448 26166
rect 5940 26099 5980 26155
rect 6036 26099 6104 26155
rect 6160 26099 6228 26155
rect 6284 26114 6335 26155
rect 6284 26099 6352 26114
rect 6408 26099 6448 26155
rect 5940 26058 6448 26099
rect 5940 26031 6335 26058
rect 6387 26031 6448 26058
rect 5940 25975 5980 26031
rect 6036 25975 6104 26031
rect 6160 25975 6228 26031
rect 6284 26006 6335 26031
rect 6284 25975 6352 26006
rect 6408 25975 6448 26031
rect 5940 25950 6448 25975
rect 5940 25907 6335 25950
rect 6387 25907 6448 25950
rect 5940 25851 5980 25907
rect 6036 25851 6104 25907
rect 6160 25851 6228 25907
rect 6284 25898 6335 25907
rect 6284 25851 6352 25898
rect 6408 25851 6448 25907
rect 5940 25842 6448 25851
rect 5940 25790 6335 25842
rect 6387 25790 6448 25842
rect 5940 25783 6448 25790
rect 5940 25727 5980 25783
rect 6036 25727 6104 25783
rect 6160 25727 6228 25783
rect 6284 25734 6352 25783
rect 6284 25727 6335 25734
rect 6408 25727 6448 25783
rect 5940 25682 6335 25727
rect 6387 25682 6448 25727
rect 5940 25659 6448 25682
rect 5940 25603 5980 25659
rect 6036 25603 6104 25659
rect 6160 25603 6228 25659
rect 6284 25626 6352 25659
rect 6284 25603 6335 25626
rect 6408 25603 6448 25659
rect 5940 25574 6335 25603
rect 6387 25574 6448 25603
rect 5940 25535 6448 25574
rect 5940 25479 5980 25535
rect 6036 25479 6104 25535
rect 6160 25479 6228 25535
rect 6284 25479 6352 25535
rect 6408 25479 6448 25535
rect 5940 25411 6448 25479
rect 5940 25355 5980 25411
rect 6036 25355 6104 25411
rect 6160 25355 6228 25411
rect 6284 25355 6352 25411
rect 6408 25355 6448 25411
rect 5940 25287 6448 25355
rect 5940 25231 5980 25287
rect 6036 25231 6104 25287
rect 6160 25231 6228 25287
rect 6284 25231 6352 25287
rect 6408 25231 6448 25287
rect 5940 25163 6448 25231
rect 5940 25107 5980 25163
rect 6036 25107 6104 25163
rect 6160 25107 6228 25163
rect 6284 25107 6352 25163
rect 6408 25107 6448 25163
rect 5940 25039 6448 25107
rect 5940 24983 5980 25039
rect 6036 24983 6104 25039
rect 6160 24983 6228 25039
rect 6284 24983 6352 25039
rect 6408 24983 6448 25039
rect 5940 24915 6448 24983
rect 5940 24859 5980 24915
rect 6036 24859 6104 24915
rect 6160 24859 6228 24915
rect 6284 24859 6352 24915
rect 6408 24859 6448 24915
rect 5940 24791 6448 24859
rect 5940 24735 5980 24791
rect 6036 24735 6104 24791
rect 6160 24735 6228 24791
rect 6284 24735 6352 24791
rect 6408 24735 6448 24791
rect 5940 24702 6448 24735
rect 5940 24667 6335 24702
rect 6387 24667 6448 24702
rect 5940 24611 5980 24667
rect 6036 24611 6104 24667
rect 6160 24611 6228 24667
rect 6284 24650 6335 24667
rect 6284 24611 6352 24650
rect 6408 24611 6448 24667
rect 5940 24594 6448 24611
rect 5940 24543 6335 24594
rect 6387 24543 6448 24594
rect 5940 24487 5980 24543
rect 6036 24487 6104 24543
rect 6160 24487 6228 24543
rect 6284 24542 6335 24543
rect 6284 24487 6352 24542
rect 6408 24487 6448 24543
rect 5940 24486 6448 24487
rect 5940 24434 6335 24486
rect 6387 24434 6448 24486
rect 5940 24419 6448 24434
rect 5940 24363 5980 24419
rect 6036 24363 6104 24419
rect 6160 24363 6228 24419
rect 6284 24378 6352 24419
rect 6284 24363 6335 24378
rect 6408 24363 6448 24419
rect 5940 24326 6335 24363
rect 6387 24326 6448 24363
rect 5940 24295 6448 24326
rect 5940 24239 5980 24295
rect 6036 24239 6104 24295
rect 6160 24239 6228 24295
rect 6284 24270 6352 24295
rect 6284 24239 6335 24270
rect 6408 24239 6448 24295
rect 5940 24218 6335 24239
rect 6387 24218 6448 24239
rect 5940 24171 6448 24218
rect 5940 24115 5980 24171
rect 6036 24115 6104 24171
rect 6160 24115 6228 24171
rect 6284 24162 6352 24171
rect 6284 24115 6335 24162
rect 6408 24115 6448 24171
rect 5940 24110 6335 24115
rect 6387 24110 6448 24115
rect 5940 24054 6448 24110
rect 5940 24047 6335 24054
rect 6387 24047 6448 24054
rect 5940 23991 5980 24047
rect 6036 23991 6104 24047
rect 6160 23991 6228 24047
rect 6284 24002 6335 24047
rect 6284 23991 6352 24002
rect 6408 23991 6448 24047
rect 5940 23946 6448 23991
rect 5940 23923 6335 23946
rect 6387 23923 6448 23946
rect 5940 23867 5980 23923
rect 6036 23867 6104 23923
rect 6160 23867 6228 23923
rect 6284 23894 6335 23923
rect 6284 23867 6352 23894
rect 6408 23867 6448 23923
rect 5940 23838 6448 23867
rect 5940 23799 6335 23838
rect 6387 23799 6448 23838
rect 5940 23743 5980 23799
rect 6036 23743 6104 23799
rect 6160 23743 6228 23799
rect 6284 23786 6335 23799
rect 6284 23743 6352 23786
rect 6408 23743 6448 23799
rect 5940 23730 6448 23743
rect 5940 23678 6335 23730
rect 6387 23678 6448 23730
rect 5940 23622 6448 23678
rect 5940 23570 6335 23622
rect 6387 23570 6448 23622
rect 5940 23514 6448 23570
rect 5940 23462 6335 23514
rect 6387 23462 6448 23514
rect 5940 23451 6448 23462
rect 5940 23395 5980 23451
rect 6036 23395 6104 23451
rect 6160 23395 6228 23451
rect 6284 23406 6352 23451
rect 6284 23395 6335 23406
rect 6408 23395 6448 23451
rect 5940 23354 6335 23395
rect 6387 23354 6448 23395
rect 5940 23327 6448 23354
rect 5940 23271 5980 23327
rect 6036 23271 6104 23327
rect 6160 23271 6228 23327
rect 6284 23298 6352 23327
rect 6284 23271 6335 23298
rect 6408 23271 6448 23327
rect 5940 23246 6335 23271
rect 6387 23246 6448 23271
rect 5940 23203 6448 23246
rect 5940 23147 5980 23203
rect 6036 23147 6104 23203
rect 6160 23147 6228 23203
rect 6284 23190 6352 23203
rect 6284 23147 6335 23190
rect 6408 23147 6448 23203
rect 5940 23138 6335 23147
rect 6387 23138 6448 23147
rect 5940 23082 6448 23138
rect 5940 23079 6335 23082
rect 6387 23079 6448 23082
rect 5940 23023 5980 23079
rect 6036 23023 6104 23079
rect 6160 23023 6228 23079
rect 6284 23030 6335 23079
rect 6284 23023 6352 23030
rect 6408 23023 6448 23079
rect 5940 22974 6448 23023
rect 5940 22955 6335 22974
rect 6387 22955 6448 22974
rect 5940 22899 5980 22955
rect 6036 22899 6104 22955
rect 6160 22899 6228 22955
rect 6284 22922 6335 22955
rect 6284 22899 6352 22922
rect 6408 22899 6448 22955
rect 5940 22866 6448 22899
rect 5940 22831 6335 22866
rect 6387 22831 6448 22866
rect 5940 22775 5980 22831
rect 6036 22775 6104 22831
rect 6160 22775 6228 22831
rect 6284 22814 6335 22831
rect 6284 22775 6352 22814
rect 6408 22775 6448 22831
rect 5940 22758 6448 22775
rect 5940 22707 6335 22758
rect 6387 22707 6448 22758
rect 5940 22651 5980 22707
rect 6036 22651 6104 22707
rect 6160 22651 6228 22707
rect 6284 22706 6335 22707
rect 6284 22651 6352 22706
rect 6408 22651 6448 22707
rect 5940 22650 6448 22651
rect 5940 22598 6335 22650
rect 6387 22598 6448 22650
rect 5940 22583 6448 22598
rect 5940 22527 5980 22583
rect 6036 22527 6104 22583
rect 6160 22527 6228 22583
rect 6284 22542 6352 22583
rect 6284 22527 6335 22542
rect 6408 22527 6448 22583
rect 5940 22490 6335 22527
rect 6387 22490 6448 22527
rect 5940 22459 6448 22490
rect 5940 22403 5980 22459
rect 6036 22403 6104 22459
rect 6160 22403 6228 22459
rect 6284 22434 6352 22459
rect 6284 22403 6335 22434
rect 6408 22403 6448 22459
rect 5940 22382 6335 22403
rect 6387 22382 6448 22403
rect 5940 22335 6448 22382
rect 5940 22279 5980 22335
rect 6036 22279 6104 22335
rect 6160 22279 6228 22335
rect 6284 22326 6352 22335
rect 6284 22279 6335 22326
rect 6408 22279 6448 22335
rect 5940 22274 6335 22279
rect 6387 22274 6448 22279
rect 5940 22218 6448 22274
rect 5940 22211 6335 22218
rect 6387 22211 6448 22218
rect 5940 22155 5980 22211
rect 6036 22155 6104 22211
rect 6160 22155 6228 22211
rect 6284 22166 6335 22211
rect 6284 22155 6352 22166
rect 6408 22155 6448 22211
rect 5940 22110 6448 22155
rect 5940 22087 6335 22110
rect 6387 22087 6448 22110
rect 5940 22031 5980 22087
rect 6036 22031 6104 22087
rect 6160 22031 6228 22087
rect 6284 22058 6335 22087
rect 6284 22031 6352 22058
rect 6408 22031 6448 22087
rect 5940 22002 6448 22031
rect 5940 21963 6335 22002
rect 6387 21963 6448 22002
rect 5940 21907 5980 21963
rect 6036 21907 6104 21963
rect 6160 21907 6228 21963
rect 6284 21950 6335 21963
rect 6284 21907 6352 21950
rect 6408 21907 6448 21963
rect 5940 21894 6448 21907
rect 5940 21842 6335 21894
rect 6387 21842 6448 21894
rect 5940 21839 6448 21842
rect 5940 21783 5980 21839
rect 6036 21783 6104 21839
rect 6160 21783 6228 21839
rect 6284 21786 6352 21839
rect 6284 21783 6335 21786
rect 6408 21783 6448 21839
rect 5940 21734 6335 21783
rect 6387 21734 6448 21783
rect 5940 21715 6448 21734
rect 5940 21659 5980 21715
rect 6036 21659 6104 21715
rect 6160 21659 6228 21715
rect 6284 21678 6352 21715
rect 6284 21659 6335 21678
rect 6408 21659 6448 21715
rect 5940 21626 6335 21659
rect 6387 21626 6448 21659
rect 5940 21591 6448 21626
rect 5940 21535 5980 21591
rect 6036 21535 6104 21591
rect 6160 21535 6228 21591
rect 6284 21535 6352 21591
rect 6408 21535 6448 21591
rect 5940 21467 6448 21535
rect 5940 21411 5980 21467
rect 6036 21411 6104 21467
rect 6160 21411 6228 21467
rect 6284 21411 6352 21467
rect 6408 21411 6448 21467
rect 5940 21343 6448 21411
rect 5940 21287 5980 21343
rect 6036 21287 6104 21343
rect 6160 21287 6228 21343
rect 6284 21287 6352 21343
rect 6408 21287 6448 21343
rect 5940 21219 6448 21287
rect 5940 21163 5980 21219
rect 6036 21163 6104 21219
rect 6160 21163 6228 21219
rect 6284 21163 6352 21219
rect 6408 21163 6448 21219
rect 5940 21095 6448 21163
rect 5940 21039 5980 21095
rect 6036 21039 6104 21095
rect 6160 21039 6228 21095
rect 6284 21039 6352 21095
rect 6408 21039 6448 21095
rect 5940 20971 6448 21039
rect 5940 20915 5980 20971
rect 6036 20915 6104 20971
rect 6160 20915 6228 20971
rect 6284 20915 6352 20971
rect 6408 20915 6448 20971
rect 5940 20847 6448 20915
rect 5940 20791 5980 20847
rect 6036 20791 6104 20847
rect 6160 20791 6228 20847
rect 6284 20791 6352 20847
rect 6408 20791 6448 20847
rect 5940 20723 6448 20791
rect 5940 20667 5980 20723
rect 6036 20667 6104 20723
rect 6160 20667 6228 20723
rect 6284 20667 6352 20723
rect 6408 20667 6448 20723
rect 5940 20599 6448 20667
rect 5940 20577 5980 20599
rect 6036 20577 6104 20599
rect 6160 20577 6228 20599
rect 6284 20577 6352 20599
rect 6408 20577 6448 20599
rect 5940 20525 5952 20577
rect 6036 20543 6060 20577
rect 6160 20543 6168 20577
rect 6004 20525 6060 20543
rect 6112 20525 6168 20543
rect 6220 20543 6228 20577
rect 6328 20543 6352 20577
rect 6220 20525 6276 20543
rect 6328 20525 6384 20543
rect 6436 20525 6448 20577
rect 5940 20469 6448 20525
rect 5940 20417 5952 20469
rect 6004 20417 6060 20469
rect 6112 20417 6168 20469
rect 6220 20417 6276 20469
rect 6328 20417 6384 20469
rect 6436 20417 6448 20469
rect 5940 20361 6448 20417
rect 5940 20309 5952 20361
rect 6004 20309 6060 20361
rect 6112 20309 6168 20361
rect 6220 20309 6276 20361
rect 6328 20309 6384 20361
rect 6436 20309 6448 20361
rect 5940 20251 6448 20309
rect 5940 20195 5980 20251
rect 6036 20195 6104 20251
rect 6160 20195 6228 20251
rect 6284 20195 6352 20251
rect 6408 20195 6448 20251
rect 5940 20127 6448 20195
rect 5940 20071 5980 20127
rect 6036 20071 6104 20127
rect 6160 20071 6228 20127
rect 6284 20071 6352 20127
rect 6408 20071 6448 20127
rect 5940 20003 6448 20071
rect 5940 19947 5980 20003
rect 6036 19947 6104 20003
rect 6160 19947 6228 20003
rect 6284 19947 6352 20003
rect 6408 19947 6448 20003
rect 5940 19879 6448 19947
rect 5940 19823 5980 19879
rect 6036 19823 6104 19879
rect 6160 19823 6228 19879
rect 6284 19823 6352 19879
rect 6408 19823 6448 19879
rect 5940 19755 6448 19823
rect 5940 19699 5980 19755
rect 6036 19699 6104 19755
rect 6160 19699 6228 19755
rect 6284 19699 6352 19755
rect 6408 19699 6448 19755
rect 5940 19631 6448 19699
rect 5940 19584 5980 19631
rect 6036 19584 6104 19631
rect 6160 19584 6228 19631
rect 6284 19584 6352 19631
rect 6408 19584 6448 19631
rect 5940 19532 5952 19584
rect 6036 19575 6060 19584
rect 6160 19575 6168 19584
rect 6004 19532 6060 19575
rect 6112 19532 6168 19575
rect 6220 19575 6228 19584
rect 6328 19575 6352 19584
rect 6220 19532 6276 19575
rect 6328 19532 6384 19575
rect 6436 19532 6448 19584
rect 5940 19507 6448 19532
rect 5940 19476 5980 19507
rect 6036 19476 6104 19507
rect 6160 19476 6228 19507
rect 6284 19476 6352 19507
rect 6408 19476 6448 19507
rect 5940 19424 5952 19476
rect 6036 19451 6060 19476
rect 6160 19451 6168 19476
rect 6004 19424 6060 19451
rect 6112 19424 6168 19451
rect 6220 19451 6228 19476
rect 6328 19451 6352 19476
rect 6220 19424 6276 19451
rect 6328 19424 6384 19451
rect 6436 19424 6448 19476
rect 5940 19383 6448 19424
rect 5940 19327 5980 19383
rect 6036 19327 6104 19383
rect 6160 19327 6228 19383
rect 6284 19327 6352 19383
rect 6408 19327 6448 19383
rect 5940 19259 6448 19327
rect 5940 19203 5980 19259
rect 6036 19203 6104 19259
rect 6160 19203 6228 19259
rect 6284 19203 6352 19259
rect 6408 19203 6448 19259
rect 5940 19135 6448 19203
rect 5940 19079 5980 19135
rect 6036 19079 6104 19135
rect 6160 19079 6228 19135
rect 6284 19079 6352 19135
rect 6408 19079 6448 19135
rect 5940 19011 6448 19079
rect 5940 18955 5980 19011
rect 6036 18955 6104 19011
rect 6160 18955 6228 19011
rect 6284 18955 6352 19011
rect 6408 18955 6448 19011
rect 5940 18887 6448 18955
rect 5940 18831 5980 18887
rect 6036 18831 6104 18887
rect 6160 18831 6228 18887
rect 6284 18831 6352 18887
rect 6408 18831 6448 18887
rect 5940 18763 6448 18831
rect 5940 18712 5980 18763
rect 6036 18712 6104 18763
rect 6160 18712 6228 18763
rect 6284 18712 6352 18763
rect 6408 18712 6448 18763
rect 5940 18660 5952 18712
rect 6036 18707 6060 18712
rect 6160 18707 6168 18712
rect 6004 18660 6060 18707
rect 6112 18660 6168 18707
rect 6220 18707 6228 18712
rect 6328 18707 6352 18712
rect 6220 18660 6276 18707
rect 6328 18660 6384 18707
rect 6436 18660 6448 18712
rect 5940 18639 6448 18660
rect 5940 18604 5980 18639
rect 6036 18604 6104 18639
rect 6160 18604 6228 18639
rect 6284 18604 6352 18639
rect 6408 18604 6448 18639
rect 5940 18552 5952 18604
rect 6036 18583 6060 18604
rect 6160 18583 6168 18604
rect 6004 18552 6060 18583
rect 6112 18552 6168 18583
rect 6220 18583 6228 18604
rect 6328 18583 6352 18604
rect 6220 18552 6276 18583
rect 6328 18552 6384 18583
rect 6436 18552 6448 18604
rect 5940 18515 6448 18552
rect 5940 18459 5980 18515
rect 6036 18459 6104 18515
rect 6160 18459 6228 18515
rect 6284 18459 6352 18515
rect 6408 18459 6448 18515
rect 5940 18391 6448 18459
rect 5940 18335 5980 18391
rect 6036 18335 6104 18391
rect 6160 18335 6228 18391
rect 6284 18335 6352 18391
rect 6408 18335 6448 18391
rect 5940 18267 6448 18335
rect 5940 18211 5980 18267
rect 6036 18211 6104 18267
rect 6160 18211 6228 18267
rect 6284 18211 6352 18267
rect 6408 18211 6448 18267
rect 5940 18143 6448 18211
rect 5940 18087 5980 18143
rect 6036 18087 6104 18143
rect 6160 18087 6228 18143
rect 6284 18087 6352 18143
rect 6408 18087 6448 18143
rect 5940 18019 6448 18087
rect 5940 17963 5980 18019
rect 6036 17963 6104 18019
rect 6160 17963 6228 18019
rect 6284 17963 6352 18019
rect 6408 17963 6448 18019
rect 5940 17895 6448 17963
rect 5940 17840 5980 17895
rect 6036 17840 6104 17895
rect 6160 17840 6228 17895
rect 6284 17840 6352 17895
rect 6408 17840 6448 17895
rect 5940 17788 5952 17840
rect 6036 17839 6060 17840
rect 6160 17839 6168 17840
rect 6004 17788 6060 17839
rect 6112 17788 6168 17839
rect 6220 17839 6228 17840
rect 6328 17839 6352 17840
rect 6220 17788 6276 17839
rect 6328 17788 6384 17839
rect 6436 17788 6448 17840
rect 5940 17771 6448 17788
rect 5940 17732 5980 17771
rect 6036 17732 6104 17771
rect 6160 17732 6228 17771
rect 6284 17732 6352 17771
rect 6408 17732 6448 17771
rect 5940 17680 5952 17732
rect 6036 17715 6060 17732
rect 6160 17715 6168 17732
rect 6004 17680 6060 17715
rect 6112 17680 6168 17715
rect 6220 17715 6228 17732
rect 6328 17715 6352 17732
rect 6220 17680 6276 17715
rect 6328 17680 6384 17715
rect 6436 17680 6448 17732
rect 5940 17647 6448 17680
rect 5940 17591 5980 17647
rect 6036 17591 6104 17647
rect 6160 17591 6228 17647
rect 6284 17591 6352 17647
rect 6408 17591 6448 17647
rect 5940 17523 6448 17591
rect 5940 17467 5980 17523
rect 6036 17467 6104 17523
rect 6160 17467 6228 17523
rect 6284 17467 6352 17523
rect 6408 17467 6448 17523
rect 5940 17399 6448 17467
rect 5940 17343 5980 17399
rect 6036 17343 6104 17399
rect 6160 17343 6228 17399
rect 6284 17343 6352 17399
rect 6408 17343 6448 17399
rect 5940 17051 6448 17343
rect 5940 16995 5980 17051
rect 6036 16995 6104 17051
rect 6160 16995 6228 17051
rect 6284 16995 6352 17051
rect 6408 16995 6448 17051
rect 5940 16968 6448 16995
rect 5940 16916 5952 16968
rect 6004 16927 6060 16968
rect 6112 16927 6168 16968
rect 6036 16916 6060 16927
rect 6160 16916 6168 16927
rect 6220 16927 6276 16968
rect 6328 16927 6384 16968
rect 6220 16916 6228 16927
rect 6328 16916 6352 16927
rect 6436 16916 6448 16968
rect 5940 16871 5980 16916
rect 6036 16871 6104 16916
rect 6160 16871 6228 16916
rect 6284 16871 6352 16916
rect 6408 16871 6448 16916
rect 5940 16860 6448 16871
rect 5940 16808 5952 16860
rect 6004 16808 6060 16860
rect 6112 16808 6168 16860
rect 6220 16808 6276 16860
rect 6328 16808 6384 16860
rect 6436 16808 6448 16860
rect 5940 16803 6448 16808
rect 5940 16747 5980 16803
rect 6036 16747 6104 16803
rect 6160 16747 6228 16803
rect 6284 16747 6352 16803
rect 6408 16747 6448 16803
rect 5940 16679 6448 16747
rect 5940 16623 5980 16679
rect 6036 16623 6104 16679
rect 6160 16623 6228 16679
rect 6284 16623 6352 16679
rect 6408 16623 6448 16679
rect 5940 16555 6448 16623
rect 5940 16499 5980 16555
rect 6036 16499 6104 16555
rect 6160 16499 6228 16555
rect 6284 16499 6352 16555
rect 6408 16499 6448 16555
rect 5940 16431 6448 16499
rect 5940 16375 5980 16431
rect 6036 16375 6104 16431
rect 6160 16375 6228 16431
rect 6284 16375 6352 16431
rect 6408 16375 6448 16431
rect 5940 16307 6448 16375
rect 5940 16251 5980 16307
rect 6036 16251 6104 16307
rect 6160 16251 6228 16307
rect 6284 16251 6352 16307
rect 6408 16251 6448 16307
rect 5940 16183 6448 16251
rect 5940 16127 5980 16183
rect 6036 16127 6104 16183
rect 6160 16127 6228 16183
rect 6284 16127 6352 16183
rect 6408 16127 6448 16183
rect 5940 16083 6448 16127
rect 5940 16031 5952 16083
rect 6004 16059 6060 16083
rect 6112 16059 6168 16083
rect 6036 16031 6060 16059
rect 6160 16031 6168 16059
rect 6220 16059 6276 16083
rect 6328 16059 6384 16083
rect 6220 16031 6228 16059
rect 6328 16031 6352 16059
rect 6436 16031 6448 16083
rect 5940 16003 5980 16031
rect 6036 16003 6104 16031
rect 6160 16003 6228 16031
rect 6284 16003 6352 16031
rect 6408 16003 6448 16031
rect 5940 15975 6448 16003
rect 5940 15923 5952 15975
rect 6004 15935 6060 15975
rect 6112 15935 6168 15975
rect 6036 15923 6060 15935
rect 6160 15923 6168 15935
rect 6220 15935 6276 15975
rect 6328 15935 6384 15975
rect 6220 15923 6228 15935
rect 6328 15923 6352 15935
rect 6436 15923 6448 15975
rect 5940 15879 5980 15923
rect 6036 15879 6104 15923
rect 6160 15879 6228 15923
rect 6284 15879 6352 15923
rect 6408 15879 6448 15923
rect 5940 15867 6448 15879
rect 5940 15815 5952 15867
rect 6004 15815 6060 15867
rect 6112 15815 6168 15867
rect 6220 15815 6276 15867
rect 6328 15815 6384 15867
rect 6436 15815 6448 15867
rect 5940 15811 6448 15815
rect 5940 15762 5980 15811
rect 4136 15755 4146 15762
rect 3698 15687 4146 15755
rect 3698 15631 3708 15687
rect 3764 15631 3832 15687
rect 3888 15631 3956 15687
rect 4012 15631 4080 15687
rect 4136 15631 4146 15687
rect 3698 15563 4146 15631
rect 3698 15507 3708 15563
rect 3764 15507 3832 15563
rect 3888 15507 3956 15563
rect 4012 15507 4080 15563
rect 4136 15507 4146 15563
rect 3698 15439 4146 15507
rect 3698 15383 3708 15439
rect 3764 15383 3832 15439
rect 3888 15383 3956 15439
rect 4012 15383 4080 15439
rect 4136 15383 4146 15439
rect 3698 15315 4146 15383
rect 3698 15259 3708 15315
rect 3764 15259 3832 15315
rect 3888 15259 3956 15315
rect 4012 15259 4080 15315
rect 4136 15259 4146 15315
rect 3698 15191 4146 15259
rect 3698 15135 3708 15191
rect 3764 15135 3832 15191
rect 3888 15135 3956 15191
rect 4012 15135 4080 15191
rect 4136 15135 4146 15191
rect 3698 15067 4146 15135
rect 3698 15011 3708 15067
rect 3764 15011 3832 15067
rect 3888 15011 3956 15067
rect 4012 15011 4080 15067
rect 4136 15011 4146 15067
rect 3698 14943 4146 15011
rect 3698 14887 3708 14943
rect 3764 14887 3832 14943
rect 3888 14887 3956 14943
rect 4012 14887 4080 14943
rect 4136 14887 4146 14943
rect 3698 14819 4146 14887
rect 3698 14763 3708 14819
rect 3764 14763 3832 14819
rect 3888 14763 3956 14819
rect 4012 14763 4080 14819
rect 4136 14763 4146 14819
rect 3698 14695 4146 14763
rect 3698 14639 3708 14695
rect 3764 14639 3832 14695
rect 3888 14639 3956 14695
rect 4012 14639 4080 14695
rect 4136 14639 4146 14695
rect 3698 14571 4146 14639
rect 3698 14515 3708 14571
rect 3764 14515 3832 14571
rect 3888 14515 3956 14571
rect 4012 14515 4080 14571
rect 4136 14515 4146 14571
rect 3698 14447 4146 14515
rect 3698 14391 3708 14447
rect 3764 14391 3832 14447
rect 3888 14391 3956 14447
rect 4012 14391 4080 14447
rect 4136 14391 4146 14447
rect 3698 14323 4146 14391
rect 3698 14267 3708 14323
rect 3764 14267 3832 14323
rect 3888 14267 3956 14323
rect 4012 14267 4080 14323
rect 4136 14267 4146 14323
rect 3698 14199 4146 14267
rect 3698 14143 3708 14199
rect 3764 14143 3832 14199
rect 3888 14143 3956 14199
rect 4012 14143 4080 14199
rect 4136 14143 4146 14199
rect 3698 14133 4146 14143
rect 5970 15755 5980 15762
rect 6036 15755 6104 15811
rect 6160 15755 6228 15811
rect 6284 15755 6352 15811
rect 6408 15762 6448 15811
rect 7076 56922 7502 56975
rect 7076 56866 7137 56922
rect 7193 56866 7261 56922
rect 7317 56866 7385 56922
rect 7441 56866 7502 56922
rect 7076 56798 7502 56866
rect 7076 56742 7137 56798
rect 7193 56742 7261 56798
rect 7317 56742 7385 56798
rect 7441 56742 7502 56798
rect 7076 56711 7502 56742
rect 7076 56659 7101 56711
rect 7153 56674 7209 56711
rect 7193 56659 7209 56674
rect 7261 56674 7317 56711
rect 7076 56618 7137 56659
rect 7193 56618 7261 56659
rect 7369 56674 7425 56711
rect 7369 56659 7385 56674
rect 7477 56659 7502 56711
rect 7317 56618 7385 56659
rect 7441 56618 7502 56659
rect 7076 56603 7502 56618
rect 7076 56551 7101 56603
rect 7153 56551 7209 56603
rect 7261 56551 7317 56603
rect 7369 56551 7425 56603
rect 7477 56551 7502 56603
rect 7076 56550 7502 56551
rect 7076 56495 7137 56550
rect 7193 56495 7261 56550
rect 7076 56443 7101 56495
rect 7193 56494 7209 56495
rect 7153 56443 7209 56494
rect 7317 56495 7385 56550
rect 7441 56495 7502 56550
rect 7261 56443 7317 56494
rect 7369 56494 7385 56495
rect 7369 56443 7425 56494
rect 7477 56443 7502 56495
rect 7076 56426 7502 56443
rect 7076 56370 7137 56426
rect 7193 56370 7261 56426
rect 7317 56370 7385 56426
rect 7441 56370 7502 56426
rect 7076 56302 7502 56370
rect 7076 56246 7137 56302
rect 7193 56246 7261 56302
rect 7317 56246 7385 56302
rect 7441 56246 7502 56302
rect 7076 56232 7502 56246
rect 7076 56180 7388 56232
rect 7440 56180 7502 56232
rect 7076 56178 7502 56180
rect 7076 56122 7137 56178
rect 7193 56122 7261 56178
rect 7317 56122 7385 56178
rect 7441 56122 7502 56178
rect 7076 56072 7388 56122
rect 7440 56072 7502 56122
rect 7076 56054 7502 56072
rect 7076 55998 7137 56054
rect 7193 55998 7261 56054
rect 7317 55998 7385 56054
rect 7441 55998 7502 56054
rect 7076 55964 7388 55998
rect 7440 55964 7502 55998
rect 7076 55930 7502 55964
rect 7076 55874 7137 55930
rect 7193 55874 7261 55930
rect 7317 55874 7385 55930
rect 7441 55874 7502 55930
rect 7076 55856 7388 55874
rect 7440 55856 7502 55874
rect 7076 55806 7502 55856
rect 7076 55750 7137 55806
rect 7193 55750 7261 55806
rect 7317 55750 7385 55806
rect 7441 55750 7502 55806
rect 7076 55748 7388 55750
rect 7440 55748 7502 55750
rect 7076 55692 7502 55748
rect 7076 55640 7388 55692
rect 7440 55640 7502 55692
rect 7076 55584 7502 55640
rect 7076 55532 7388 55584
rect 7440 55532 7502 55584
rect 7076 55476 7502 55532
rect 7076 55424 7388 55476
rect 7440 55424 7502 55476
rect 7076 55368 7502 55424
rect 7076 55316 7388 55368
rect 7440 55316 7502 55368
rect 7076 55260 7502 55316
rect 7076 55208 7388 55260
rect 7440 55208 7502 55260
rect 7076 55152 7502 55208
rect 7076 55100 7388 55152
rect 7440 55100 7502 55152
rect 7076 55044 7502 55100
rect 7076 54992 7388 55044
rect 7440 54992 7502 55044
rect 7076 54936 7502 54992
rect 7076 54884 7388 54936
rect 7440 54884 7502 54936
rect 7076 54828 7502 54884
rect 7076 54776 7388 54828
rect 7440 54776 7502 54828
rect 7076 54720 7502 54776
rect 7076 54668 7388 54720
rect 7440 54668 7502 54720
rect 7076 54612 7502 54668
rect 7076 54560 7388 54612
rect 7440 54560 7502 54612
rect 7076 54504 7502 54560
rect 7076 54452 7388 54504
rect 7440 54452 7502 54504
rect 7076 54396 7502 54452
rect 7076 54344 7388 54396
rect 7440 54344 7502 54396
rect 7076 54288 7502 54344
rect 7076 54236 7388 54288
rect 7440 54236 7502 54288
rect 7076 54180 7502 54236
rect 7076 54128 7388 54180
rect 7440 54128 7502 54180
rect 7076 54072 7502 54128
rect 7076 54020 7388 54072
rect 7440 54020 7502 54072
rect 7076 53964 7502 54020
rect 7076 53912 7388 53964
rect 7440 53912 7502 53964
rect 7076 53856 7502 53912
rect 7076 53845 7388 53856
rect 7440 53845 7502 53856
rect 7076 53789 7137 53845
rect 7193 53789 7261 53845
rect 7317 53789 7385 53845
rect 7441 53789 7502 53845
rect 7076 53748 7502 53789
rect 7076 53721 7388 53748
rect 7440 53721 7502 53748
rect 7076 53665 7137 53721
rect 7193 53665 7261 53721
rect 7317 53665 7385 53721
rect 7441 53665 7502 53721
rect 7076 53640 7502 53665
rect 7076 53597 7388 53640
rect 7440 53597 7502 53640
rect 7076 53541 7137 53597
rect 7193 53541 7261 53597
rect 7317 53541 7385 53597
rect 7441 53541 7502 53597
rect 7076 53532 7502 53541
rect 7076 53480 7388 53532
rect 7440 53480 7502 53532
rect 7076 53473 7502 53480
rect 7076 53417 7137 53473
rect 7193 53417 7261 53473
rect 7317 53417 7385 53473
rect 7441 53417 7502 53473
rect 7076 53372 7388 53417
rect 7440 53372 7502 53417
rect 7076 53349 7502 53372
rect 7076 53293 7137 53349
rect 7193 53293 7261 53349
rect 7317 53293 7385 53349
rect 7441 53293 7502 53349
rect 7076 53264 7388 53293
rect 7440 53264 7502 53293
rect 7076 53225 7502 53264
rect 7076 53169 7137 53225
rect 7193 53169 7261 53225
rect 7317 53169 7385 53225
rect 7441 53169 7502 53225
rect 7076 53101 7502 53169
rect 7076 53045 7137 53101
rect 7193 53045 7261 53101
rect 7317 53045 7385 53101
rect 7441 53045 7502 53101
rect 7076 52996 7139 53045
rect 7191 52996 7263 53045
rect 7315 52996 7387 53045
rect 7439 52996 7502 53045
rect 7076 52977 7502 52996
rect 7076 52921 7137 52977
rect 7193 52921 7261 52977
rect 7317 52921 7385 52977
rect 7441 52921 7502 52977
rect 7076 52872 7139 52921
rect 7191 52872 7263 52921
rect 7315 52872 7387 52921
rect 7439 52872 7502 52921
rect 7076 52853 7502 52872
rect 7076 52797 7137 52853
rect 7193 52797 7261 52853
rect 7317 52797 7385 52853
rect 7441 52797 7502 52853
rect 7076 52748 7139 52797
rect 7191 52748 7263 52797
rect 7315 52748 7387 52797
rect 7439 52748 7502 52797
rect 7076 52729 7502 52748
rect 7076 52673 7137 52729
rect 7193 52673 7261 52729
rect 7317 52673 7385 52729
rect 7441 52673 7502 52729
rect 7076 52624 7139 52673
rect 7191 52624 7263 52673
rect 7315 52624 7387 52673
rect 7439 52624 7502 52673
rect 7076 52605 7502 52624
rect 7076 52549 7137 52605
rect 7193 52549 7261 52605
rect 7317 52549 7385 52605
rect 7441 52549 7502 52605
rect 7076 52500 7139 52549
rect 7191 52500 7263 52549
rect 7315 52500 7387 52549
rect 7439 52500 7502 52549
rect 7076 52284 7502 52500
rect 7076 52232 7388 52284
rect 7440 52232 7502 52284
rect 7076 52176 7502 52232
rect 7076 52124 7388 52176
rect 7440 52124 7502 52176
rect 7076 52068 7502 52124
rect 7076 52016 7388 52068
rect 7440 52016 7502 52068
rect 7076 51960 7502 52016
rect 7076 51908 7388 51960
rect 7440 51908 7502 51960
rect 7076 51852 7502 51908
rect 7076 51800 7388 51852
rect 7440 51800 7502 51852
rect 7076 51744 7502 51800
rect 7076 51692 7388 51744
rect 7440 51692 7502 51744
rect 7076 51636 7502 51692
rect 7076 51584 7388 51636
rect 7440 51584 7502 51636
rect 7076 51528 7502 51584
rect 7076 51476 7388 51528
rect 7440 51476 7502 51528
rect 7076 51420 7502 51476
rect 7076 51368 7388 51420
rect 7440 51368 7502 51420
rect 7076 51312 7502 51368
rect 7076 51260 7388 51312
rect 7440 51260 7502 51312
rect 7076 51204 7502 51260
rect 7076 51152 7388 51204
rect 7440 51152 7502 51204
rect 7076 51096 7502 51152
rect 7076 51044 7388 51096
rect 7440 51044 7502 51096
rect 7076 50988 7502 51044
rect 7076 50936 7388 50988
rect 7440 50936 7502 50988
rect 7076 50880 7502 50936
rect 7076 50828 7388 50880
rect 7440 50828 7502 50880
rect 7076 50772 7502 50828
rect 7076 50720 7388 50772
rect 7440 50720 7502 50772
rect 7076 50664 7502 50720
rect 7076 50612 7388 50664
rect 7440 50612 7502 50664
rect 7076 50556 7502 50612
rect 7076 50504 7388 50556
rect 7440 50504 7502 50556
rect 7076 50448 7502 50504
rect 7076 50396 7388 50448
rect 7440 50396 7502 50448
rect 7076 50340 7502 50396
rect 7076 50288 7388 50340
rect 7440 50288 7502 50340
rect 7076 50232 7502 50288
rect 7076 50180 7388 50232
rect 7440 50180 7502 50232
rect 7076 50124 7502 50180
rect 7076 50072 7388 50124
rect 7440 50072 7502 50124
rect 7076 50016 7502 50072
rect 7076 49964 7388 50016
rect 7440 49964 7502 50016
rect 7076 49908 7502 49964
rect 7076 49856 7388 49908
rect 7440 49856 7502 49908
rect 7076 49800 7502 49856
rect 7076 49748 7388 49800
rect 7440 49748 7502 49800
rect 7076 49692 7502 49748
rect 7076 49640 7388 49692
rect 7440 49640 7502 49692
rect 7076 49584 7502 49640
rect 7076 49532 7388 49584
rect 7440 49532 7502 49584
rect 7076 49476 7502 49532
rect 7076 49424 7388 49476
rect 7440 49424 7502 49476
rect 7076 49368 7502 49424
rect 7076 49316 7388 49368
rect 7440 49316 7502 49368
rect 7076 49100 7502 49316
rect 7076 49048 7139 49100
rect 7191 49048 7263 49100
rect 7315 49048 7387 49100
rect 7439 49048 7502 49100
rect 7076 49045 7502 49048
rect 7076 48989 7137 49045
rect 7193 48989 7261 49045
rect 7317 48989 7385 49045
rect 7441 48989 7502 49045
rect 7076 48976 7502 48989
rect 7076 48924 7139 48976
rect 7191 48924 7263 48976
rect 7315 48924 7387 48976
rect 7439 48924 7502 48976
rect 7076 48921 7502 48924
rect 7076 48865 7137 48921
rect 7193 48865 7261 48921
rect 7317 48865 7385 48921
rect 7441 48865 7502 48921
rect 7076 48852 7502 48865
rect 7076 48800 7139 48852
rect 7191 48800 7263 48852
rect 7315 48800 7387 48852
rect 7439 48800 7502 48852
rect 7076 48797 7502 48800
rect 7076 48741 7137 48797
rect 7193 48741 7261 48797
rect 7317 48741 7385 48797
rect 7441 48741 7502 48797
rect 7076 48728 7502 48741
rect 7076 48676 7139 48728
rect 7191 48676 7263 48728
rect 7315 48676 7387 48728
rect 7439 48676 7502 48728
rect 7076 48673 7502 48676
rect 7076 48617 7137 48673
rect 7193 48617 7261 48673
rect 7317 48617 7385 48673
rect 7441 48617 7502 48673
rect 7076 48604 7502 48617
rect 7076 48552 7139 48604
rect 7191 48552 7263 48604
rect 7315 48552 7387 48604
rect 7439 48552 7502 48604
rect 7076 48549 7502 48552
rect 7076 48493 7137 48549
rect 7193 48493 7261 48549
rect 7317 48493 7385 48549
rect 7441 48493 7502 48549
rect 7076 48425 7502 48493
rect 7076 48369 7137 48425
rect 7193 48369 7261 48425
rect 7317 48369 7385 48425
rect 7441 48369 7502 48425
rect 7076 48336 7502 48369
rect 7076 48301 7388 48336
rect 7440 48301 7502 48336
rect 7076 48245 7137 48301
rect 7193 48245 7261 48301
rect 7317 48245 7385 48301
rect 7441 48245 7502 48301
rect 7076 48228 7502 48245
rect 7076 48177 7388 48228
rect 7440 48177 7502 48228
rect 7076 48121 7137 48177
rect 7193 48121 7261 48177
rect 7317 48121 7385 48177
rect 7441 48121 7502 48177
rect 7076 48120 7502 48121
rect 7076 48068 7388 48120
rect 7440 48068 7502 48120
rect 7076 48053 7502 48068
rect 7076 47997 7137 48053
rect 7193 47997 7261 48053
rect 7317 47997 7385 48053
rect 7441 47997 7502 48053
rect 7076 47960 7388 47997
rect 7440 47960 7502 47997
rect 7076 47929 7502 47960
rect 7076 47873 7137 47929
rect 7193 47873 7261 47929
rect 7317 47873 7385 47929
rect 7441 47873 7502 47929
rect 7076 47852 7388 47873
rect 7440 47852 7502 47873
rect 7076 47805 7502 47852
rect 7076 47749 7137 47805
rect 7193 47749 7261 47805
rect 7317 47749 7385 47805
rect 7441 47749 7502 47805
rect 7076 47744 7388 47749
rect 7440 47744 7502 47749
rect 7076 47688 7502 47744
rect 7076 47636 7388 47688
rect 7440 47636 7502 47688
rect 7076 47580 7502 47636
rect 7076 47528 7388 47580
rect 7440 47528 7502 47580
rect 7076 47472 7502 47528
rect 7076 47420 7388 47472
rect 7440 47420 7502 47472
rect 7076 47364 7502 47420
rect 7076 47312 7388 47364
rect 7440 47312 7502 47364
rect 7076 47256 7502 47312
rect 7076 47204 7388 47256
rect 7440 47204 7502 47256
rect 7076 47148 7502 47204
rect 7076 47096 7388 47148
rect 7440 47096 7502 47148
rect 7076 47040 7502 47096
rect 7076 46988 7388 47040
rect 7440 46988 7502 47040
rect 7076 46932 7502 46988
rect 7076 46880 7388 46932
rect 7440 46880 7502 46932
rect 7076 46824 7502 46880
rect 7076 46772 7388 46824
rect 7440 46772 7502 46824
rect 7076 46716 7502 46772
rect 7076 46664 7388 46716
rect 7440 46664 7502 46716
rect 7076 46608 7502 46664
rect 7076 46556 7388 46608
rect 7440 46556 7502 46608
rect 7076 46500 7502 46556
rect 7076 46448 7388 46500
rect 7440 46448 7502 46500
rect 7076 46392 7502 46448
rect 7076 46340 7388 46392
rect 7440 46340 7502 46392
rect 7076 46284 7502 46340
rect 7076 46232 7388 46284
rect 7440 46232 7502 46284
rect 7076 46176 7502 46232
rect 7076 46124 7388 46176
rect 7440 46124 7502 46176
rect 7076 46068 7502 46124
rect 7076 46016 7388 46068
rect 7440 46016 7502 46068
rect 7076 45960 7502 46016
rect 7076 45908 7388 45960
rect 7440 45908 7502 45960
rect 7076 45852 7502 45908
rect 7076 45845 7388 45852
rect 7440 45845 7502 45852
rect 7076 45789 7137 45845
rect 7193 45789 7261 45845
rect 7317 45789 7385 45845
rect 7441 45789 7502 45845
rect 7076 45744 7502 45789
rect 7076 45721 7388 45744
rect 7440 45721 7502 45744
rect 7076 45665 7137 45721
rect 7193 45665 7261 45721
rect 7317 45665 7385 45721
rect 7441 45665 7502 45721
rect 7076 45636 7502 45665
rect 7076 45597 7388 45636
rect 7440 45597 7502 45636
rect 7076 45541 7137 45597
rect 7193 45541 7261 45597
rect 7317 45541 7385 45597
rect 7441 45541 7502 45597
rect 7076 45528 7502 45541
rect 7076 45476 7388 45528
rect 7440 45476 7502 45528
rect 7076 45473 7502 45476
rect 7076 45417 7137 45473
rect 7193 45417 7261 45473
rect 7317 45417 7385 45473
rect 7441 45417 7502 45473
rect 7076 45368 7388 45417
rect 7440 45368 7502 45417
rect 7076 45349 7502 45368
rect 7076 45293 7137 45349
rect 7193 45293 7261 45349
rect 7317 45293 7385 45349
rect 7441 45293 7502 45349
rect 7076 45225 7502 45293
rect 7076 45169 7137 45225
rect 7193 45169 7261 45225
rect 7317 45169 7385 45225
rect 7441 45169 7502 45225
rect 7076 45152 7502 45169
rect 7076 45101 7139 45152
rect 7191 45101 7263 45152
rect 7315 45101 7387 45152
rect 7439 45101 7502 45152
rect 7076 45045 7137 45101
rect 7193 45045 7261 45101
rect 7317 45045 7385 45101
rect 7441 45045 7502 45101
rect 7076 45028 7502 45045
rect 7076 44977 7139 45028
rect 7191 44977 7263 45028
rect 7315 44977 7387 45028
rect 7439 44977 7502 45028
rect 7076 44921 7137 44977
rect 7193 44921 7261 44977
rect 7317 44921 7385 44977
rect 7441 44921 7502 44977
rect 7076 44904 7502 44921
rect 7076 44853 7139 44904
rect 7191 44853 7263 44904
rect 7315 44853 7387 44904
rect 7439 44853 7502 44904
rect 7076 44797 7137 44853
rect 7193 44797 7261 44853
rect 7317 44797 7385 44853
rect 7441 44797 7502 44853
rect 7076 44780 7502 44797
rect 7076 44729 7139 44780
rect 7191 44729 7263 44780
rect 7315 44729 7387 44780
rect 7439 44729 7502 44780
rect 7076 44673 7137 44729
rect 7193 44673 7261 44729
rect 7317 44673 7385 44729
rect 7441 44673 7502 44729
rect 7076 44656 7502 44673
rect 7076 44605 7139 44656
rect 7191 44605 7263 44656
rect 7315 44605 7387 44656
rect 7439 44605 7502 44656
rect 7076 44549 7137 44605
rect 7193 44549 7261 44605
rect 7317 44549 7385 44605
rect 7441 44549 7502 44605
rect 7076 44388 7502 44549
rect 7076 44336 7388 44388
rect 7440 44336 7502 44388
rect 7076 44280 7502 44336
rect 7076 44228 7388 44280
rect 7440 44228 7502 44280
rect 7076 44172 7502 44228
rect 7076 44120 7388 44172
rect 7440 44120 7502 44172
rect 7076 44064 7502 44120
rect 7076 44012 7388 44064
rect 7440 44012 7502 44064
rect 7076 43956 7502 44012
rect 7076 43904 7388 43956
rect 7440 43904 7502 43956
rect 7076 43848 7502 43904
rect 7076 43796 7388 43848
rect 7440 43796 7502 43848
rect 7076 43740 7502 43796
rect 7076 43688 7388 43740
rect 7440 43688 7502 43740
rect 7076 43632 7502 43688
rect 7076 43580 7388 43632
rect 7440 43580 7502 43632
rect 7076 43524 7502 43580
rect 7076 43472 7388 43524
rect 7440 43472 7502 43524
rect 7076 43416 7502 43472
rect 7076 43364 7388 43416
rect 7440 43364 7502 43416
rect 7076 43308 7502 43364
rect 7076 43256 7388 43308
rect 7440 43256 7502 43308
rect 7076 43200 7502 43256
rect 7076 43148 7388 43200
rect 7440 43148 7502 43200
rect 7076 43092 7502 43148
rect 7076 43040 7388 43092
rect 7440 43040 7502 43092
rect 7076 42984 7502 43040
rect 7076 42932 7388 42984
rect 7440 42932 7502 42984
rect 7076 42876 7502 42932
rect 7076 42824 7388 42876
rect 7440 42824 7502 42876
rect 7076 42768 7502 42824
rect 7076 42716 7388 42768
rect 7440 42716 7502 42768
rect 7076 42660 7502 42716
rect 7076 42608 7388 42660
rect 7440 42608 7502 42660
rect 7076 42552 7502 42608
rect 7076 42500 7388 42552
rect 7440 42500 7502 42552
rect 7076 42444 7502 42500
rect 7076 42392 7388 42444
rect 7440 42392 7502 42444
rect 7076 42336 7502 42392
rect 7076 42284 7388 42336
rect 7440 42284 7502 42336
rect 7076 42228 7502 42284
rect 7076 42176 7388 42228
rect 7440 42176 7502 42228
rect 7076 42120 7502 42176
rect 7076 42068 7388 42120
rect 7440 42068 7502 42120
rect 7076 42012 7502 42068
rect 7076 41960 7388 42012
rect 7440 41960 7502 42012
rect 7076 41904 7502 41960
rect 7076 41852 7388 41904
rect 7440 41852 7502 41904
rect 7076 41796 7502 41852
rect 7076 41744 7388 41796
rect 7440 41744 7502 41796
rect 7076 41688 7502 41744
rect 7076 41636 7388 41688
rect 7440 41636 7502 41688
rect 7076 41580 7502 41636
rect 7076 41528 7388 41580
rect 7440 41528 7502 41580
rect 7076 41472 7502 41528
rect 7076 41420 7388 41472
rect 7440 41420 7502 41472
rect 7076 41204 7502 41420
rect 7076 41152 7139 41204
rect 7191 41152 7263 41204
rect 7315 41152 7387 41204
rect 7439 41152 7502 41204
rect 7076 41080 7502 41152
rect 7076 41028 7139 41080
rect 7191 41028 7263 41080
rect 7315 41028 7387 41080
rect 7439 41028 7502 41080
rect 7076 40956 7502 41028
rect 7076 40904 7139 40956
rect 7191 40904 7263 40956
rect 7315 40904 7387 40956
rect 7439 40904 7502 40956
rect 7076 40832 7502 40904
rect 7076 40780 7139 40832
rect 7191 40780 7263 40832
rect 7315 40780 7387 40832
rect 7439 40780 7502 40832
rect 7076 40708 7502 40780
rect 7076 40656 7139 40708
rect 7191 40656 7263 40708
rect 7315 40656 7387 40708
rect 7439 40656 7502 40708
rect 7076 40440 7502 40656
rect 7076 40388 7388 40440
rect 7440 40388 7502 40440
rect 7076 40332 7502 40388
rect 7076 40280 7388 40332
rect 7440 40280 7502 40332
rect 7076 40224 7502 40280
rect 7076 40172 7388 40224
rect 7440 40172 7502 40224
rect 7076 40116 7502 40172
rect 7076 40064 7388 40116
rect 7440 40064 7502 40116
rect 7076 40008 7502 40064
rect 7076 39956 7388 40008
rect 7440 39956 7502 40008
rect 7076 39900 7502 39956
rect 7076 39848 7388 39900
rect 7440 39848 7502 39900
rect 7076 39792 7502 39848
rect 7076 39740 7388 39792
rect 7440 39740 7502 39792
rect 7076 39684 7502 39740
rect 7076 39632 7388 39684
rect 7440 39632 7502 39684
rect 7076 39576 7502 39632
rect 7076 39524 7388 39576
rect 7440 39524 7502 39576
rect 7076 39468 7502 39524
rect 7076 39416 7388 39468
rect 7440 39416 7502 39468
rect 7076 39360 7502 39416
rect 7076 39308 7388 39360
rect 7440 39308 7502 39360
rect 7076 39252 7502 39308
rect 7076 39200 7388 39252
rect 7440 39200 7502 39252
rect 7076 39144 7502 39200
rect 7076 39092 7388 39144
rect 7440 39092 7502 39144
rect 7076 39036 7502 39092
rect 7076 38984 7388 39036
rect 7440 38984 7502 39036
rect 7076 38928 7502 38984
rect 7076 38876 7388 38928
rect 7440 38876 7502 38928
rect 7076 38820 7502 38876
rect 7076 38768 7388 38820
rect 7440 38768 7502 38820
rect 7076 38712 7502 38768
rect 7076 38660 7388 38712
rect 7440 38660 7502 38712
rect 7076 38604 7502 38660
rect 7076 38552 7388 38604
rect 7440 38552 7502 38604
rect 7076 38496 7502 38552
rect 7076 38444 7388 38496
rect 7440 38444 7502 38496
rect 7076 38388 7502 38444
rect 7076 38336 7388 38388
rect 7440 38336 7502 38388
rect 7076 38280 7502 38336
rect 7076 38228 7388 38280
rect 7440 38228 7502 38280
rect 7076 38172 7502 38228
rect 7076 38120 7388 38172
rect 7440 38120 7502 38172
rect 7076 38064 7502 38120
rect 7076 38012 7388 38064
rect 7440 38012 7502 38064
rect 7076 37956 7502 38012
rect 7076 37904 7388 37956
rect 7440 37904 7502 37956
rect 7076 37848 7502 37904
rect 7076 37796 7388 37848
rect 7440 37796 7502 37848
rect 7076 37740 7502 37796
rect 7076 37688 7388 37740
rect 7440 37688 7502 37740
rect 7076 37632 7502 37688
rect 7076 37580 7388 37632
rect 7440 37580 7502 37632
rect 7076 37524 7502 37580
rect 7076 37472 7388 37524
rect 7440 37472 7502 37524
rect 7076 37256 7502 37472
rect 7076 37204 7139 37256
rect 7191 37204 7263 37256
rect 7315 37204 7387 37256
rect 7439 37204 7502 37256
rect 7076 37132 7502 37204
rect 7076 37080 7139 37132
rect 7191 37080 7263 37132
rect 7315 37080 7387 37132
rect 7439 37080 7502 37132
rect 7076 37008 7502 37080
rect 7076 36956 7139 37008
rect 7191 36956 7263 37008
rect 7315 36956 7387 37008
rect 7439 36956 7502 37008
rect 7076 36884 7502 36956
rect 7076 36832 7139 36884
rect 7191 36832 7263 36884
rect 7315 36832 7387 36884
rect 7439 36832 7502 36884
rect 7076 36760 7502 36832
rect 7076 36708 7139 36760
rect 7191 36708 7263 36760
rect 7315 36708 7387 36760
rect 7439 36708 7502 36760
rect 7076 36492 7502 36708
rect 7076 36440 7388 36492
rect 7440 36440 7502 36492
rect 7076 36384 7502 36440
rect 7076 36332 7388 36384
rect 7440 36332 7502 36384
rect 7076 36276 7502 36332
rect 7076 36251 7388 36276
rect 7440 36251 7502 36276
rect 7076 36195 7137 36251
rect 7193 36195 7261 36251
rect 7317 36195 7385 36251
rect 7441 36195 7502 36251
rect 7076 36168 7502 36195
rect 7076 36127 7388 36168
rect 7440 36127 7502 36168
rect 7076 36071 7137 36127
rect 7193 36071 7261 36127
rect 7317 36071 7385 36127
rect 7441 36071 7502 36127
rect 7076 36060 7502 36071
rect 7076 36008 7388 36060
rect 7440 36008 7502 36060
rect 7076 36003 7502 36008
rect 7076 35947 7137 36003
rect 7193 35947 7261 36003
rect 7317 35947 7385 36003
rect 7441 35947 7502 36003
rect 7076 35900 7388 35947
rect 7440 35900 7502 35947
rect 7076 35879 7502 35900
rect 7076 35823 7137 35879
rect 7193 35823 7261 35879
rect 7317 35823 7385 35879
rect 7441 35823 7502 35879
rect 7076 35792 7388 35823
rect 7440 35792 7502 35823
rect 7076 35755 7502 35792
rect 7076 35699 7137 35755
rect 7193 35699 7261 35755
rect 7317 35699 7385 35755
rect 7441 35699 7502 35755
rect 7076 35684 7388 35699
rect 7440 35684 7502 35699
rect 7076 35631 7502 35684
rect 7076 35575 7137 35631
rect 7193 35575 7261 35631
rect 7317 35575 7385 35631
rect 7441 35575 7502 35631
rect 7076 35520 7502 35575
rect 7076 35507 7388 35520
rect 7440 35507 7502 35520
rect 7076 35451 7137 35507
rect 7193 35451 7261 35507
rect 7317 35451 7385 35507
rect 7441 35451 7502 35507
rect 7076 35412 7502 35451
rect 7076 35383 7388 35412
rect 7440 35383 7502 35412
rect 7076 35327 7137 35383
rect 7193 35327 7261 35383
rect 7317 35327 7385 35383
rect 7441 35327 7502 35383
rect 7076 35304 7502 35327
rect 7076 35259 7388 35304
rect 7440 35259 7502 35304
rect 7076 35203 7137 35259
rect 7193 35203 7261 35259
rect 7317 35203 7385 35259
rect 7441 35203 7502 35259
rect 7076 35196 7502 35203
rect 7076 35144 7388 35196
rect 7440 35144 7502 35196
rect 7076 35135 7502 35144
rect 7076 35079 7137 35135
rect 7193 35079 7261 35135
rect 7317 35079 7385 35135
rect 7441 35079 7502 35135
rect 7076 35036 7388 35079
rect 7440 35036 7502 35079
rect 7076 35011 7502 35036
rect 7076 34955 7137 35011
rect 7193 34955 7261 35011
rect 7317 34955 7385 35011
rect 7441 34955 7502 35011
rect 7076 34928 7388 34955
rect 7440 34928 7502 34955
rect 7076 34887 7502 34928
rect 7076 34831 7137 34887
rect 7193 34831 7261 34887
rect 7317 34831 7385 34887
rect 7441 34831 7502 34887
rect 7076 34820 7388 34831
rect 7440 34820 7502 34831
rect 7076 34764 7502 34820
rect 7076 34763 7388 34764
rect 7440 34763 7502 34764
rect 7076 34707 7137 34763
rect 7193 34707 7261 34763
rect 7317 34707 7385 34763
rect 7441 34707 7502 34763
rect 7076 34656 7502 34707
rect 7076 34639 7388 34656
rect 7440 34639 7502 34656
rect 7076 34583 7137 34639
rect 7193 34583 7261 34639
rect 7317 34583 7385 34639
rect 7441 34583 7502 34639
rect 7076 34548 7502 34583
rect 7076 34515 7388 34548
rect 7440 34515 7502 34548
rect 7076 34459 7137 34515
rect 7193 34459 7261 34515
rect 7317 34459 7385 34515
rect 7441 34459 7502 34515
rect 7076 34440 7502 34459
rect 7076 34391 7388 34440
rect 7440 34391 7502 34440
rect 7076 34335 7137 34391
rect 7193 34335 7261 34391
rect 7317 34335 7385 34391
rect 7441 34335 7502 34391
rect 7076 34332 7502 34335
rect 7076 34280 7388 34332
rect 7440 34280 7502 34332
rect 7076 34267 7502 34280
rect 7076 34211 7137 34267
rect 7193 34211 7261 34267
rect 7317 34211 7385 34267
rect 7441 34211 7502 34267
rect 7076 34172 7388 34211
rect 7440 34172 7502 34211
rect 7076 34143 7502 34172
rect 7076 34087 7137 34143
rect 7193 34087 7261 34143
rect 7317 34087 7385 34143
rect 7441 34087 7502 34143
rect 7076 34064 7388 34087
rect 7440 34064 7502 34087
rect 7076 34019 7502 34064
rect 7076 33963 7137 34019
rect 7193 33963 7261 34019
rect 7317 33963 7385 34019
rect 7441 33963 7502 34019
rect 7076 33956 7388 33963
rect 7440 33956 7502 33963
rect 7076 33900 7502 33956
rect 7076 33895 7388 33900
rect 7440 33895 7502 33900
rect 7076 33839 7137 33895
rect 7193 33839 7261 33895
rect 7317 33839 7385 33895
rect 7441 33839 7502 33895
rect 7076 33792 7502 33839
rect 7076 33771 7388 33792
rect 7440 33771 7502 33792
rect 7076 33715 7137 33771
rect 7193 33715 7261 33771
rect 7317 33715 7385 33771
rect 7441 33715 7502 33771
rect 7076 33684 7502 33715
rect 7076 33647 7388 33684
rect 7440 33647 7502 33684
rect 7076 33591 7137 33647
rect 7193 33591 7261 33647
rect 7317 33591 7385 33647
rect 7441 33591 7502 33647
rect 7076 33576 7502 33591
rect 7076 33524 7388 33576
rect 7440 33524 7502 33576
rect 7076 33523 7502 33524
rect 7076 33467 7137 33523
rect 7193 33467 7261 33523
rect 7317 33467 7385 33523
rect 7441 33467 7502 33523
rect 7076 33399 7502 33467
rect 7076 33343 7137 33399
rect 7193 33343 7261 33399
rect 7317 33343 7385 33399
rect 7441 33343 7502 33399
rect 7076 33308 7502 33343
rect 7076 33256 7139 33308
rect 7191 33256 7263 33308
rect 7315 33256 7387 33308
rect 7439 33256 7502 33308
rect 7076 33184 7502 33256
rect 7076 33132 7139 33184
rect 7191 33132 7263 33184
rect 7315 33132 7387 33184
rect 7439 33132 7502 33184
rect 7076 33060 7502 33132
rect 7076 33008 7139 33060
rect 7191 33008 7263 33060
rect 7315 33008 7387 33060
rect 7439 33008 7502 33060
rect 7076 32936 7502 33008
rect 7076 32884 7139 32936
rect 7191 32884 7263 32936
rect 7315 32884 7387 32936
rect 7439 32884 7502 32936
rect 7076 32812 7502 32884
rect 7076 32760 7139 32812
rect 7191 32760 7263 32812
rect 7315 32760 7387 32812
rect 7439 32760 7502 32812
rect 7076 32544 7502 32760
rect 7076 32492 7388 32544
rect 7440 32492 7502 32544
rect 7076 32436 7502 32492
rect 7076 32384 7388 32436
rect 7440 32384 7502 32436
rect 7076 32328 7502 32384
rect 7076 32276 7388 32328
rect 7440 32276 7502 32328
rect 7076 32220 7502 32276
rect 7076 32168 7388 32220
rect 7440 32168 7502 32220
rect 7076 32112 7502 32168
rect 7076 32060 7388 32112
rect 7440 32060 7502 32112
rect 7076 32004 7502 32060
rect 7076 31952 7388 32004
rect 7440 31952 7502 32004
rect 7076 31896 7502 31952
rect 7076 31844 7388 31896
rect 7440 31844 7502 31896
rect 7076 31788 7502 31844
rect 7076 31736 7388 31788
rect 7440 31736 7502 31788
rect 7076 31680 7502 31736
rect 7076 31628 7388 31680
rect 7440 31628 7502 31680
rect 7076 31572 7502 31628
rect 7076 31520 7388 31572
rect 7440 31520 7502 31572
rect 7076 31464 7502 31520
rect 7076 31412 7388 31464
rect 7440 31412 7502 31464
rect 7076 31356 7502 31412
rect 7076 31304 7388 31356
rect 7440 31304 7502 31356
rect 7076 31248 7502 31304
rect 7076 31196 7388 31248
rect 7440 31196 7502 31248
rect 7076 31140 7502 31196
rect 7076 31088 7388 31140
rect 7440 31088 7502 31140
rect 7076 31032 7502 31088
rect 7076 30980 7388 31032
rect 7440 30980 7502 31032
rect 7076 30924 7502 30980
rect 7076 30872 7388 30924
rect 7440 30872 7502 30924
rect 7076 30816 7502 30872
rect 7076 30764 7388 30816
rect 7440 30764 7502 30816
rect 7076 30708 7502 30764
rect 7076 30656 7388 30708
rect 7440 30656 7502 30708
rect 7076 30600 7502 30656
rect 7076 30548 7388 30600
rect 7440 30548 7502 30600
rect 7076 30492 7502 30548
rect 7076 30440 7388 30492
rect 7440 30440 7502 30492
rect 7076 30384 7502 30440
rect 7076 30332 7388 30384
rect 7440 30332 7502 30384
rect 7076 30276 7502 30332
rect 7076 30224 7388 30276
rect 7440 30224 7502 30276
rect 7076 30168 7502 30224
rect 7076 30116 7388 30168
rect 7440 30116 7502 30168
rect 7076 30060 7502 30116
rect 7076 30008 7388 30060
rect 7440 30008 7502 30060
rect 7076 29952 7502 30008
rect 7076 29900 7388 29952
rect 7440 29900 7502 29952
rect 7076 29844 7502 29900
rect 7076 29792 7388 29844
rect 7440 29792 7502 29844
rect 7076 29736 7502 29792
rect 7076 29684 7388 29736
rect 7440 29684 7502 29736
rect 7076 29628 7502 29684
rect 7076 29576 7388 29628
rect 7440 29576 7502 29628
rect 7076 29360 7502 29576
rect 7076 29308 7139 29360
rect 7191 29308 7263 29360
rect 7315 29308 7387 29360
rect 7439 29308 7502 29360
rect 7076 29236 7502 29308
rect 7076 29184 7139 29236
rect 7191 29184 7263 29236
rect 7315 29184 7387 29236
rect 7439 29184 7502 29236
rect 7076 29112 7502 29184
rect 7076 29060 7139 29112
rect 7191 29060 7263 29112
rect 7315 29060 7387 29112
rect 7439 29060 7502 29112
rect 7076 28988 7502 29060
rect 7076 28936 7139 28988
rect 7191 28936 7263 28988
rect 7315 28936 7387 28988
rect 7439 28936 7502 28988
rect 7076 28864 7502 28936
rect 7076 28812 7139 28864
rect 7191 28812 7263 28864
rect 7315 28812 7387 28864
rect 7439 28812 7502 28864
rect 7076 28596 7502 28812
rect 7076 28544 7388 28596
rect 7440 28544 7502 28596
rect 7076 28488 7502 28544
rect 7076 28436 7388 28488
rect 7440 28436 7502 28488
rect 7076 28380 7502 28436
rect 7076 28328 7388 28380
rect 7440 28328 7502 28380
rect 7076 28272 7502 28328
rect 7076 28245 7388 28272
rect 7440 28245 7502 28272
rect 7076 28189 7137 28245
rect 7193 28189 7261 28245
rect 7317 28189 7385 28245
rect 7441 28189 7502 28245
rect 7076 28164 7502 28189
rect 7076 28121 7388 28164
rect 7440 28121 7502 28164
rect 7076 28065 7137 28121
rect 7193 28065 7261 28121
rect 7317 28065 7385 28121
rect 7441 28065 7502 28121
rect 7076 28056 7502 28065
rect 7076 28004 7388 28056
rect 7440 28004 7502 28056
rect 7076 27997 7502 28004
rect 7076 27941 7137 27997
rect 7193 27941 7261 27997
rect 7317 27941 7385 27997
rect 7441 27941 7502 27997
rect 7076 27896 7388 27941
rect 7440 27896 7502 27941
rect 7076 27873 7502 27896
rect 7076 27817 7137 27873
rect 7193 27817 7261 27873
rect 7317 27817 7385 27873
rect 7441 27817 7502 27873
rect 7076 27788 7388 27817
rect 7440 27788 7502 27817
rect 7076 27749 7502 27788
rect 7076 27693 7137 27749
rect 7193 27693 7261 27749
rect 7317 27693 7385 27749
rect 7441 27693 7502 27749
rect 7076 27680 7388 27693
rect 7440 27680 7502 27693
rect 7076 27625 7502 27680
rect 7076 27569 7137 27625
rect 7193 27569 7261 27625
rect 7317 27569 7385 27625
rect 7441 27569 7502 27625
rect 7076 27516 7502 27569
rect 7076 27501 7388 27516
rect 7440 27501 7502 27516
rect 7076 27445 7137 27501
rect 7193 27445 7261 27501
rect 7317 27445 7385 27501
rect 7441 27445 7502 27501
rect 7076 27408 7502 27445
rect 7076 27377 7388 27408
rect 7440 27377 7502 27408
rect 7076 27321 7137 27377
rect 7193 27321 7261 27377
rect 7317 27321 7385 27377
rect 7441 27321 7502 27377
rect 7076 27300 7502 27321
rect 7076 27253 7388 27300
rect 7440 27253 7502 27300
rect 7076 27197 7137 27253
rect 7193 27197 7261 27253
rect 7317 27197 7385 27253
rect 7441 27197 7502 27253
rect 7076 27192 7502 27197
rect 7076 27140 7388 27192
rect 7440 27140 7502 27192
rect 7076 27129 7502 27140
rect 7076 27073 7137 27129
rect 7193 27073 7261 27129
rect 7317 27073 7385 27129
rect 7441 27073 7502 27129
rect 7076 27032 7388 27073
rect 7440 27032 7502 27073
rect 7076 27005 7502 27032
rect 7076 26949 7137 27005
rect 7193 26949 7261 27005
rect 7317 26949 7385 27005
rect 7441 26949 7502 27005
rect 7076 26924 7388 26949
rect 7440 26924 7502 26949
rect 7076 26868 7502 26924
rect 7076 26816 7388 26868
rect 7440 26816 7502 26868
rect 7076 26760 7502 26816
rect 7076 26708 7388 26760
rect 7440 26708 7502 26760
rect 7076 26652 7502 26708
rect 7076 26600 7388 26652
rect 7440 26600 7502 26652
rect 7076 26544 7502 26600
rect 7076 26492 7388 26544
rect 7440 26492 7502 26544
rect 7076 26436 7502 26492
rect 7076 26384 7388 26436
rect 7440 26384 7502 26436
rect 7076 26328 7502 26384
rect 7076 26276 7388 26328
rect 7440 26276 7502 26328
rect 7076 26220 7502 26276
rect 7076 26168 7388 26220
rect 7440 26168 7502 26220
rect 7076 26112 7502 26168
rect 7076 26060 7388 26112
rect 7440 26060 7502 26112
rect 7076 26004 7502 26060
rect 7076 25952 7388 26004
rect 7440 25952 7502 26004
rect 7076 25896 7502 25952
rect 7076 25844 7388 25896
rect 7440 25844 7502 25896
rect 7076 25788 7502 25844
rect 7076 25736 7388 25788
rect 7440 25736 7502 25788
rect 7076 25680 7502 25736
rect 7076 25628 7388 25680
rect 7440 25628 7502 25680
rect 7076 25412 7502 25628
rect 7076 25360 7139 25412
rect 7191 25360 7263 25412
rect 7315 25360 7387 25412
rect 7439 25360 7502 25412
rect 7076 25288 7502 25360
rect 7076 25236 7139 25288
rect 7191 25236 7263 25288
rect 7315 25236 7387 25288
rect 7439 25236 7502 25288
rect 7076 25164 7502 25236
rect 7076 25112 7139 25164
rect 7191 25112 7263 25164
rect 7315 25112 7387 25164
rect 7439 25112 7502 25164
rect 7076 25040 7502 25112
rect 7076 24988 7139 25040
rect 7191 24988 7263 25040
rect 7315 24988 7387 25040
rect 7439 24988 7502 25040
rect 7076 24916 7502 24988
rect 7076 24864 7139 24916
rect 7191 24864 7263 24916
rect 7315 24864 7387 24916
rect 7439 24864 7502 24916
rect 7076 24648 7502 24864
rect 7076 24596 7388 24648
rect 7440 24596 7502 24648
rect 7076 24540 7502 24596
rect 7076 24488 7388 24540
rect 7440 24488 7502 24540
rect 7076 24432 7502 24488
rect 7076 24380 7388 24432
rect 7440 24380 7502 24432
rect 7076 24324 7502 24380
rect 7076 24272 7388 24324
rect 7440 24272 7502 24324
rect 7076 24216 7502 24272
rect 7076 24164 7388 24216
rect 7440 24164 7502 24216
rect 7076 24108 7502 24164
rect 7076 24056 7388 24108
rect 7440 24056 7502 24108
rect 7076 24000 7502 24056
rect 7076 23948 7388 24000
rect 7440 23948 7502 24000
rect 7076 23892 7502 23948
rect 7076 23840 7388 23892
rect 7440 23840 7502 23892
rect 7076 23784 7502 23840
rect 7076 23732 7388 23784
rect 7440 23732 7502 23784
rect 7076 23676 7502 23732
rect 7076 23624 7388 23676
rect 7440 23624 7502 23676
rect 7076 23568 7502 23624
rect 7076 23516 7388 23568
rect 7440 23516 7502 23568
rect 7076 23460 7502 23516
rect 7076 23408 7388 23460
rect 7440 23408 7502 23460
rect 7076 23352 7502 23408
rect 7076 23300 7388 23352
rect 7440 23300 7502 23352
rect 7076 23244 7502 23300
rect 7076 23192 7388 23244
rect 7440 23192 7502 23244
rect 7076 23136 7502 23192
rect 7076 23084 7388 23136
rect 7440 23084 7502 23136
rect 7076 23028 7502 23084
rect 7076 22976 7388 23028
rect 7440 22976 7502 23028
rect 7076 22920 7502 22976
rect 7076 22868 7388 22920
rect 7440 22868 7502 22920
rect 7076 22812 7502 22868
rect 7076 22760 7388 22812
rect 7440 22760 7502 22812
rect 7076 22704 7502 22760
rect 7076 22652 7388 22704
rect 7440 22652 7502 22704
rect 7076 22596 7502 22652
rect 7076 22544 7388 22596
rect 7440 22544 7502 22596
rect 7076 22488 7502 22544
rect 7076 22436 7388 22488
rect 7440 22436 7502 22488
rect 7076 22380 7502 22436
rect 7076 22328 7388 22380
rect 7440 22328 7502 22380
rect 7076 22272 7502 22328
rect 7076 22220 7388 22272
rect 7440 22220 7502 22272
rect 7076 22164 7502 22220
rect 7076 22112 7388 22164
rect 7440 22112 7502 22164
rect 7076 22056 7502 22112
rect 7076 22004 7388 22056
rect 7440 22004 7502 22056
rect 7076 21948 7502 22004
rect 7076 21896 7388 21948
rect 7440 21896 7502 21948
rect 7076 21840 7502 21896
rect 7076 21788 7388 21840
rect 7440 21788 7502 21840
rect 7076 21732 7502 21788
rect 7076 21680 7388 21732
rect 7440 21680 7502 21732
rect 7076 21469 7502 21680
rect 7076 21417 7101 21469
rect 7153 21417 7209 21469
rect 7261 21417 7317 21469
rect 7369 21417 7425 21469
rect 7477 21417 7502 21469
rect 7076 21361 7502 21417
rect 7076 21309 7101 21361
rect 7153 21309 7209 21361
rect 7261 21309 7317 21361
rect 7369 21309 7425 21361
rect 7477 21309 7502 21361
rect 7076 21253 7502 21309
rect 7076 21201 7101 21253
rect 7153 21201 7209 21253
rect 7261 21201 7317 21253
rect 7369 21201 7425 21253
rect 7477 21201 7502 21253
rect 7076 19951 7502 21201
rect 7076 19899 7101 19951
rect 7153 19899 7209 19951
rect 7261 19899 7317 19951
rect 7369 19899 7425 19951
rect 7477 19899 7502 19951
rect 7076 19843 7502 19899
rect 7076 19791 7101 19843
rect 7153 19791 7209 19843
rect 7261 19791 7317 19843
rect 7369 19791 7425 19843
rect 7477 19791 7502 19843
rect 7076 19202 7502 19791
rect 7076 19150 7101 19202
rect 7153 19150 7209 19202
rect 7261 19150 7317 19202
rect 7369 19150 7425 19202
rect 7477 19150 7502 19202
rect 7076 19094 7502 19150
rect 7076 19042 7101 19094
rect 7153 19042 7209 19094
rect 7261 19042 7317 19094
rect 7369 19042 7425 19094
rect 7477 19042 7502 19094
rect 7076 18986 7502 19042
rect 7076 18934 7101 18986
rect 7153 18934 7209 18986
rect 7261 18934 7317 18986
rect 7369 18934 7425 18986
rect 7477 18934 7502 18986
rect 7076 18330 7502 18934
rect 7076 18278 7101 18330
rect 7153 18278 7209 18330
rect 7261 18278 7317 18330
rect 7369 18278 7425 18330
rect 7477 18278 7502 18330
rect 7076 18222 7502 18278
rect 7076 18170 7101 18222
rect 7153 18170 7209 18222
rect 7261 18170 7317 18222
rect 7369 18170 7425 18222
rect 7477 18170 7502 18222
rect 7076 18114 7502 18170
rect 7076 18062 7101 18114
rect 7153 18062 7209 18114
rect 7261 18062 7317 18114
rect 7369 18062 7425 18114
rect 7477 18062 7502 18114
rect 7076 17458 7502 18062
rect 7076 17406 7101 17458
rect 7153 17406 7209 17458
rect 7261 17406 7317 17458
rect 7369 17406 7425 17458
rect 7477 17406 7502 17458
rect 7076 17350 7502 17406
rect 7076 17298 7101 17350
rect 7153 17298 7209 17350
rect 7261 17298 7317 17350
rect 7369 17298 7425 17350
rect 7477 17298 7502 17350
rect 7076 17242 7502 17298
rect 7076 17190 7101 17242
rect 7153 17190 7209 17242
rect 7261 17190 7317 17242
rect 7369 17190 7425 17242
rect 7477 17190 7502 17242
rect 7076 16601 7502 17190
rect 7076 16549 7101 16601
rect 7153 16549 7209 16601
rect 7261 16549 7317 16601
rect 7369 16549 7425 16601
rect 7477 16549 7502 16601
rect 7076 16493 7502 16549
rect 7076 16441 7101 16493
rect 7153 16441 7209 16493
rect 7261 16441 7317 16493
rect 7369 16441 7425 16493
rect 7477 16441 7502 16493
rect 7076 15762 7502 16441
rect 7562 56922 7988 56975
rect 7562 56866 7623 56922
rect 7679 56866 7747 56922
rect 7803 56866 7871 56922
rect 7927 56866 7988 56922
rect 7562 56798 7988 56866
rect 7562 56742 7623 56798
rect 7679 56742 7747 56798
rect 7803 56742 7871 56798
rect 7927 56742 7988 56798
rect 7562 56711 7988 56742
rect 7562 56659 7587 56711
rect 7639 56674 7695 56711
rect 7679 56659 7695 56674
rect 7747 56674 7803 56711
rect 7562 56618 7623 56659
rect 7679 56618 7747 56659
rect 7855 56674 7911 56711
rect 7855 56659 7871 56674
rect 7963 56659 7988 56711
rect 7803 56618 7871 56659
rect 7927 56618 7988 56659
rect 7562 56603 7988 56618
rect 7562 56551 7587 56603
rect 7639 56551 7695 56603
rect 7747 56551 7803 56603
rect 7855 56551 7911 56603
rect 7963 56551 7988 56603
rect 7562 56550 7988 56551
rect 7562 56495 7623 56550
rect 7679 56495 7747 56550
rect 7562 56443 7587 56495
rect 7679 56494 7695 56495
rect 7639 56443 7695 56494
rect 7803 56495 7871 56550
rect 7927 56495 7988 56550
rect 7747 56443 7803 56494
rect 7855 56494 7871 56495
rect 7855 56443 7911 56494
rect 7963 56443 7988 56495
rect 7562 56426 7988 56443
rect 7562 56370 7623 56426
rect 7679 56370 7747 56426
rect 7803 56370 7871 56426
rect 7927 56370 7988 56426
rect 7562 56302 7988 56370
rect 7562 56246 7623 56302
rect 7679 56246 7747 56302
rect 7803 56246 7871 56302
rect 7927 56246 7988 56302
rect 7562 56232 7988 56246
rect 7562 56180 7624 56232
rect 7676 56180 7988 56232
rect 7562 56178 7988 56180
rect 7562 56122 7623 56178
rect 7679 56122 7747 56178
rect 7803 56122 7871 56178
rect 7927 56122 7988 56178
rect 7562 56072 7624 56122
rect 7676 56072 7988 56122
rect 7562 56054 7988 56072
rect 7562 55998 7623 56054
rect 7679 55998 7747 56054
rect 7803 55998 7871 56054
rect 7927 55998 7988 56054
rect 7562 55964 7624 55998
rect 7676 55964 7988 55998
rect 7562 55930 7988 55964
rect 7562 55874 7623 55930
rect 7679 55874 7747 55930
rect 7803 55874 7871 55930
rect 7927 55874 7988 55930
rect 7562 55856 7624 55874
rect 7676 55856 7988 55874
rect 7562 55806 7988 55856
rect 7562 55750 7623 55806
rect 7679 55750 7747 55806
rect 7803 55750 7871 55806
rect 7927 55750 7988 55806
rect 7562 55748 7624 55750
rect 7676 55748 7988 55750
rect 7562 55692 7988 55748
rect 7562 55640 7624 55692
rect 7676 55640 7988 55692
rect 7562 55584 7988 55640
rect 7562 55532 7624 55584
rect 7676 55532 7988 55584
rect 7562 55476 7988 55532
rect 7562 55424 7624 55476
rect 7676 55424 7988 55476
rect 7562 55368 7988 55424
rect 7562 55316 7624 55368
rect 7676 55316 7988 55368
rect 7562 55260 7988 55316
rect 7562 55208 7624 55260
rect 7676 55208 7988 55260
rect 7562 55152 7988 55208
rect 7562 55100 7624 55152
rect 7676 55100 7988 55152
rect 7562 55044 7988 55100
rect 7562 54992 7624 55044
rect 7676 54992 7988 55044
rect 7562 54936 7988 54992
rect 7562 54884 7624 54936
rect 7676 54884 7988 54936
rect 7562 54828 7988 54884
rect 7562 54776 7624 54828
rect 7676 54776 7988 54828
rect 7562 54720 7988 54776
rect 7562 54668 7624 54720
rect 7676 54668 7988 54720
rect 7562 54612 7988 54668
rect 7562 54560 7624 54612
rect 7676 54560 7988 54612
rect 7562 54504 7988 54560
rect 7562 54452 7624 54504
rect 7676 54452 7988 54504
rect 7562 54396 7988 54452
rect 7562 54344 7624 54396
rect 7676 54344 7988 54396
rect 7562 54288 7988 54344
rect 7562 54236 7624 54288
rect 7676 54236 7988 54288
rect 7562 54180 7988 54236
rect 7562 54128 7624 54180
rect 7676 54128 7988 54180
rect 7562 54072 7988 54128
rect 7562 54020 7624 54072
rect 7676 54020 7988 54072
rect 7562 53964 7988 54020
rect 7562 53912 7624 53964
rect 7676 53912 7988 53964
rect 7562 53856 7988 53912
rect 7562 53845 7624 53856
rect 7676 53845 7988 53856
rect 7562 53789 7623 53845
rect 7679 53789 7747 53845
rect 7803 53789 7871 53845
rect 7927 53789 7988 53845
rect 7562 53748 7988 53789
rect 7562 53721 7624 53748
rect 7676 53721 7988 53748
rect 7562 53665 7623 53721
rect 7679 53665 7747 53721
rect 7803 53665 7871 53721
rect 7927 53665 7988 53721
rect 7562 53640 7988 53665
rect 7562 53597 7624 53640
rect 7676 53597 7988 53640
rect 7562 53541 7623 53597
rect 7679 53541 7747 53597
rect 7803 53541 7871 53597
rect 7927 53541 7988 53597
rect 7562 53532 7988 53541
rect 7562 53480 7624 53532
rect 7676 53480 7988 53532
rect 7562 53473 7988 53480
rect 7562 53417 7623 53473
rect 7679 53417 7747 53473
rect 7803 53417 7871 53473
rect 7927 53417 7988 53473
rect 7562 53372 7624 53417
rect 7676 53372 7988 53417
rect 7562 53349 7988 53372
rect 7562 53293 7623 53349
rect 7679 53293 7747 53349
rect 7803 53293 7871 53349
rect 7927 53293 7988 53349
rect 7562 53264 7624 53293
rect 7676 53264 7988 53293
rect 7562 53225 7988 53264
rect 7562 53169 7623 53225
rect 7679 53169 7747 53225
rect 7803 53169 7871 53225
rect 7927 53169 7988 53225
rect 7562 53101 7988 53169
rect 7562 53045 7623 53101
rect 7679 53045 7747 53101
rect 7803 53045 7871 53101
rect 7927 53045 7988 53101
rect 7562 52996 7625 53045
rect 7677 52996 7749 53045
rect 7801 52996 7873 53045
rect 7925 52996 7988 53045
rect 7562 52977 7988 52996
rect 7562 52921 7623 52977
rect 7679 52921 7747 52977
rect 7803 52921 7871 52977
rect 7927 52921 7988 52977
rect 7562 52872 7625 52921
rect 7677 52872 7749 52921
rect 7801 52872 7873 52921
rect 7925 52872 7988 52921
rect 7562 52853 7988 52872
rect 7562 52797 7623 52853
rect 7679 52797 7747 52853
rect 7803 52797 7871 52853
rect 7927 52797 7988 52853
rect 7562 52748 7625 52797
rect 7677 52748 7749 52797
rect 7801 52748 7873 52797
rect 7925 52748 7988 52797
rect 7562 52729 7988 52748
rect 7562 52673 7623 52729
rect 7679 52673 7747 52729
rect 7803 52673 7871 52729
rect 7927 52673 7988 52729
rect 7562 52624 7625 52673
rect 7677 52624 7749 52673
rect 7801 52624 7873 52673
rect 7925 52624 7988 52673
rect 7562 52605 7988 52624
rect 7562 52549 7623 52605
rect 7679 52549 7747 52605
rect 7803 52549 7871 52605
rect 7927 52549 7988 52605
rect 7562 52500 7625 52549
rect 7677 52500 7749 52549
rect 7801 52500 7873 52549
rect 7925 52500 7988 52549
rect 7562 52284 7988 52500
rect 7562 52232 7624 52284
rect 7676 52232 7988 52284
rect 7562 52176 7988 52232
rect 7562 52124 7624 52176
rect 7676 52124 7988 52176
rect 7562 52068 7988 52124
rect 7562 52016 7624 52068
rect 7676 52016 7988 52068
rect 7562 51960 7988 52016
rect 7562 51908 7624 51960
rect 7676 51908 7988 51960
rect 7562 51852 7988 51908
rect 7562 51800 7624 51852
rect 7676 51800 7988 51852
rect 7562 51744 7988 51800
rect 7562 51692 7624 51744
rect 7676 51692 7988 51744
rect 7562 51636 7988 51692
rect 7562 51584 7624 51636
rect 7676 51584 7988 51636
rect 7562 51528 7988 51584
rect 7562 51476 7624 51528
rect 7676 51476 7988 51528
rect 7562 51420 7988 51476
rect 7562 51368 7624 51420
rect 7676 51368 7988 51420
rect 7562 51312 7988 51368
rect 7562 51260 7624 51312
rect 7676 51260 7988 51312
rect 7562 51204 7988 51260
rect 7562 51152 7624 51204
rect 7676 51152 7988 51204
rect 7562 51096 7988 51152
rect 7562 51044 7624 51096
rect 7676 51044 7988 51096
rect 7562 50988 7988 51044
rect 7562 50936 7624 50988
rect 7676 50936 7988 50988
rect 7562 50880 7988 50936
rect 7562 50828 7624 50880
rect 7676 50828 7988 50880
rect 7562 50772 7988 50828
rect 7562 50720 7624 50772
rect 7676 50720 7988 50772
rect 7562 50664 7988 50720
rect 7562 50612 7624 50664
rect 7676 50612 7988 50664
rect 7562 50556 7988 50612
rect 7562 50504 7624 50556
rect 7676 50504 7988 50556
rect 7562 50448 7988 50504
rect 7562 50396 7624 50448
rect 7676 50396 7988 50448
rect 7562 50340 7988 50396
rect 7562 50288 7624 50340
rect 7676 50288 7988 50340
rect 7562 50232 7988 50288
rect 7562 50180 7624 50232
rect 7676 50180 7988 50232
rect 7562 50124 7988 50180
rect 7562 50072 7624 50124
rect 7676 50072 7988 50124
rect 7562 50016 7988 50072
rect 7562 49964 7624 50016
rect 7676 49964 7988 50016
rect 7562 49908 7988 49964
rect 7562 49856 7624 49908
rect 7676 49856 7988 49908
rect 7562 49800 7988 49856
rect 7562 49748 7624 49800
rect 7676 49748 7988 49800
rect 7562 49692 7988 49748
rect 7562 49640 7624 49692
rect 7676 49640 7988 49692
rect 7562 49584 7988 49640
rect 7562 49532 7624 49584
rect 7676 49532 7988 49584
rect 7562 49476 7988 49532
rect 7562 49424 7624 49476
rect 7676 49424 7988 49476
rect 7562 49368 7988 49424
rect 7562 49316 7624 49368
rect 7676 49316 7988 49368
rect 7562 49100 7988 49316
rect 7562 49048 7625 49100
rect 7677 49048 7749 49100
rect 7801 49048 7873 49100
rect 7925 49048 7988 49100
rect 7562 49045 7988 49048
rect 7562 48989 7623 49045
rect 7679 48989 7747 49045
rect 7803 48989 7871 49045
rect 7927 48989 7988 49045
rect 7562 48976 7988 48989
rect 7562 48924 7625 48976
rect 7677 48924 7749 48976
rect 7801 48924 7873 48976
rect 7925 48924 7988 48976
rect 7562 48921 7988 48924
rect 7562 48865 7623 48921
rect 7679 48865 7747 48921
rect 7803 48865 7871 48921
rect 7927 48865 7988 48921
rect 7562 48852 7988 48865
rect 7562 48800 7625 48852
rect 7677 48800 7749 48852
rect 7801 48800 7873 48852
rect 7925 48800 7988 48852
rect 7562 48797 7988 48800
rect 7562 48741 7623 48797
rect 7679 48741 7747 48797
rect 7803 48741 7871 48797
rect 7927 48741 7988 48797
rect 7562 48728 7988 48741
rect 7562 48676 7625 48728
rect 7677 48676 7749 48728
rect 7801 48676 7873 48728
rect 7925 48676 7988 48728
rect 7562 48673 7988 48676
rect 7562 48617 7623 48673
rect 7679 48617 7747 48673
rect 7803 48617 7871 48673
rect 7927 48617 7988 48673
rect 7562 48604 7988 48617
rect 7562 48552 7625 48604
rect 7677 48552 7749 48604
rect 7801 48552 7873 48604
rect 7925 48552 7988 48604
rect 7562 48549 7988 48552
rect 7562 48493 7623 48549
rect 7679 48493 7747 48549
rect 7803 48493 7871 48549
rect 7927 48493 7988 48549
rect 7562 48425 7988 48493
rect 7562 48369 7623 48425
rect 7679 48369 7747 48425
rect 7803 48369 7871 48425
rect 7927 48369 7988 48425
rect 7562 48336 7988 48369
rect 7562 48301 7624 48336
rect 7676 48301 7988 48336
rect 7562 48245 7623 48301
rect 7679 48245 7747 48301
rect 7803 48245 7871 48301
rect 7927 48245 7988 48301
rect 7562 48228 7988 48245
rect 7562 48177 7624 48228
rect 7676 48177 7988 48228
rect 7562 48121 7623 48177
rect 7679 48121 7747 48177
rect 7803 48121 7871 48177
rect 7927 48121 7988 48177
rect 7562 48120 7988 48121
rect 7562 48068 7624 48120
rect 7676 48068 7988 48120
rect 7562 48053 7988 48068
rect 7562 47997 7623 48053
rect 7679 47997 7747 48053
rect 7803 47997 7871 48053
rect 7927 47997 7988 48053
rect 7562 47960 7624 47997
rect 7676 47960 7988 47997
rect 7562 47929 7988 47960
rect 7562 47873 7623 47929
rect 7679 47873 7747 47929
rect 7803 47873 7871 47929
rect 7927 47873 7988 47929
rect 7562 47852 7624 47873
rect 7676 47852 7988 47873
rect 7562 47805 7988 47852
rect 7562 47749 7623 47805
rect 7679 47749 7747 47805
rect 7803 47749 7871 47805
rect 7927 47749 7988 47805
rect 7562 47744 7624 47749
rect 7676 47744 7988 47749
rect 7562 47688 7988 47744
rect 7562 47636 7624 47688
rect 7676 47636 7988 47688
rect 7562 47580 7988 47636
rect 7562 47528 7624 47580
rect 7676 47528 7988 47580
rect 7562 47472 7988 47528
rect 7562 47420 7624 47472
rect 7676 47420 7988 47472
rect 7562 47364 7988 47420
rect 7562 47312 7624 47364
rect 7676 47312 7988 47364
rect 7562 47256 7988 47312
rect 7562 47204 7624 47256
rect 7676 47204 7988 47256
rect 7562 47148 7988 47204
rect 7562 47096 7624 47148
rect 7676 47096 7988 47148
rect 7562 47040 7988 47096
rect 7562 46988 7624 47040
rect 7676 46988 7988 47040
rect 7562 46932 7988 46988
rect 7562 46880 7624 46932
rect 7676 46880 7988 46932
rect 7562 46824 7988 46880
rect 7562 46772 7624 46824
rect 7676 46772 7988 46824
rect 7562 46716 7988 46772
rect 7562 46664 7624 46716
rect 7676 46664 7988 46716
rect 7562 46608 7988 46664
rect 7562 46556 7624 46608
rect 7676 46556 7988 46608
rect 7562 46500 7988 46556
rect 7562 46448 7624 46500
rect 7676 46448 7988 46500
rect 7562 46392 7988 46448
rect 7562 46340 7624 46392
rect 7676 46340 7988 46392
rect 7562 46284 7988 46340
rect 7562 46232 7624 46284
rect 7676 46232 7988 46284
rect 7562 46176 7988 46232
rect 7562 46124 7624 46176
rect 7676 46124 7988 46176
rect 7562 46068 7988 46124
rect 7562 46016 7624 46068
rect 7676 46016 7988 46068
rect 7562 45960 7988 46016
rect 7562 45908 7624 45960
rect 7676 45908 7988 45960
rect 7562 45852 7988 45908
rect 7562 45845 7624 45852
rect 7676 45845 7988 45852
rect 7562 45789 7623 45845
rect 7679 45789 7747 45845
rect 7803 45789 7871 45845
rect 7927 45789 7988 45845
rect 7562 45744 7988 45789
rect 7562 45721 7624 45744
rect 7676 45721 7988 45744
rect 7562 45665 7623 45721
rect 7679 45665 7747 45721
rect 7803 45665 7871 45721
rect 7927 45665 7988 45721
rect 7562 45636 7988 45665
rect 7562 45597 7624 45636
rect 7676 45597 7988 45636
rect 7562 45541 7623 45597
rect 7679 45541 7747 45597
rect 7803 45541 7871 45597
rect 7927 45541 7988 45597
rect 7562 45528 7988 45541
rect 7562 45476 7624 45528
rect 7676 45476 7988 45528
rect 7562 45473 7988 45476
rect 7562 45417 7623 45473
rect 7679 45417 7747 45473
rect 7803 45417 7871 45473
rect 7927 45417 7988 45473
rect 7562 45368 7624 45417
rect 7676 45368 7988 45417
rect 7562 45349 7988 45368
rect 7562 45293 7623 45349
rect 7679 45293 7747 45349
rect 7803 45293 7871 45349
rect 7927 45293 7988 45349
rect 7562 45225 7988 45293
rect 7562 45169 7623 45225
rect 7679 45169 7747 45225
rect 7803 45169 7871 45225
rect 7927 45169 7988 45225
rect 7562 45152 7988 45169
rect 7562 45101 7625 45152
rect 7677 45101 7749 45152
rect 7801 45101 7873 45152
rect 7925 45101 7988 45152
rect 7562 45045 7623 45101
rect 7679 45045 7747 45101
rect 7803 45045 7871 45101
rect 7927 45045 7988 45101
rect 7562 45028 7988 45045
rect 7562 44977 7625 45028
rect 7677 44977 7749 45028
rect 7801 44977 7873 45028
rect 7925 44977 7988 45028
rect 7562 44921 7623 44977
rect 7679 44921 7747 44977
rect 7803 44921 7871 44977
rect 7927 44921 7988 44977
rect 7562 44904 7988 44921
rect 7562 44853 7625 44904
rect 7677 44853 7749 44904
rect 7801 44853 7873 44904
rect 7925 44853 7988 44904
rect 7562 44797 7623 44853
rect 7679 44797 7747 44853
rect 7803 44797 7871 44853
rect 7927 44797 7988 44853
rect 7562 44780 7988 44797
rect 7562 44729 7625 44780
rect 7677 44729 7749 44780
rect 7801 44729 7873 44780
rect 7925 44729 7988 44780
rect 7562 44673 7623 44729
rect 7679 44673 7747 44729
rect 7803 44673 7871 44729
rect 7927 44673 7988 44729
rect 7562 44656 7988 44673
rect 7562 44605 7625 44656
rect 7677 44605 7749 44656
rect 7801 44605 7873 44656
rect 7925 44605 7988 44656
rect 7562 44549 7623 44605
rect 7679 44549 7747 44605
rect 7803 44549 7871 44605
rect 7927 44549 7988 44605
rect 7562 44388 7988 44549
rect 7562 44336 7624 44388
rect 7676 44336 7988 44388
rect 7562 44280 7988 44336
rect 7562 44228 7624 44280
rect 7676 44228 7988 44280
rect 7562 44172 7988 44228
rect 7562 44120 7624 44172
rect 7676 44120 7988 44172
rect 7562 44064 7988 44120
rect 7562 44012 7624 44064
rect 7676 44012 7988 44064
rect 7562 43956 7988 44012
rect 7562 43904 7624 43956
rect 7676 43904 7988 43956
rect 7562 43848 7988 43904
rect 7562 43796 7624 43848
rect 7676 43796 7988 43848
rect 7562 43740 7988 43796
rect 7562 43688 7624 43740
rect 7676 43688 7988 43740
rect 7562 43632 7988 43688
rect 7562 43580 7624 43632
rect 7676 43580 7988 43632
rect 7562 43524 7988 43580
rect 7562 43472 7624 43524
rect 7676 43472 7988 43524
rect 7562 43416 7988 43472
rect 7562 43364 7624 43416
rect 7676 43364 7988 43416
rect 7562 43308 7988 43364
rect 7562 43256 7624 43308
rect 7676 43256 7988 43308
rect 7562 43200 7988 43256
rect 7562 43148 7624 43200
rect 7676 43148 7988 43200
rect 7562 43092 7988 43148
rect 7562 43040 7624 43092
rect 7676 43040 7988 43092
rect 7562 42984 7988 43040
rect 7562 42932 7624 42984
rect 7676 42932 7988 42984
rect 7562 42876 7988 42932
rect 7562 42824 7624 42876
rect 7676 42824 7988 42876
rect 7562 42768 7988 42824
rect 7562 42716 7624 42768
rect 7676 42716 7988 42768
rect 7562 42660 7988 42716
rect 7562 42608 7624 42660
rect 7676 42608 7988 42660
rect 7562 42552 7988 42608
rect 7562 42500 7624 42552
rect 7676 42500 7988 42552
rect 7562 42444 7988 42500
rect 7562 42392 7624 42444
rect 7676 42392 7988 42444
rect 7562 42336 7988 42392
rect 7562 42284 7624 42336
rect 7676 42284 7988 42336
rect 7562 42228 7988 42284
rect 7562 42176 7624 42228
rect 7676 42176 7988 42228
rect 7562 42120 7988 42176
rect 7562 42068 7624 42120
rect 7676 42068 7988 42120
rect 7562 42012 7988 42068
rect 7562 41960 7624 42012
rect 7676 41960 7988 42012
rect 7562 41904 7988 41960
rect 7562 41852 7624 41904
rect 7676 41852 7988 41904
rect 7562 41796 7988 41852
rect 7562 41744 7624 41796
rect 7676 41744 7988 41796
rect 7562 41688 7988 41744
rect 7562 41636 7624 41688
rect 7676 41636 7988 41688
rect 7562 41580 7988 41636
rect 7562 41528 7624 41580
rect 7676 41528 7988 41580
rect 7562 41472 7988 41528
rect 7562 41420 7624 41472
rect 7676 41420 7988 41472
rect 7562 41204 7988 41420
rect 7562 41152 7625 41204
rect 7677 41152 7749 41204
rect 7801 41152 7873 41204
rect 7925 41152 7988 41204
rect 7562 41080 7988 41152
rect 7562 41028 7625 41080
rect 7677 41028 7749 41080
rect 7801 41028 7873 41080
rect 7925 41028 7988 41080
rect 7562 40956 7988 41028
rect 7562 40904 7625 40956
rect 7677 40904 7749 40956
rect 7801 40904 7873 40956
rect 7925 40904 7988 40956
rect 7562 40832 7988 40904
rect 7562 40780 7625 40832
rect 7677 40780 7749 40832
rect 7801 40780 7873 40832
rect 7925 40780 7988 40832
rect 7562 40708 7988 40780
rect 7562 40656 7625 40708
rect 7677 40656 7749 40708
rect 7801 40656 7873 40708
rect 7925 40656 7988 40708
rect 7562 40440 7988 40656
rect 7562 40388 7624 40440
rect 7676 40388 7988 40440
rect 7562 40332 7988 40388
rect 7562 40280 7624 40332
rect 7676 40280 7988 40332
rect 7562 40224 7988 40280
rect 7562 40172 7624 40224
rect 7676 40172 7988 40224
rect 7562 40116 7988 40172
rect 7562 40064 7624 40116
rect 7676 40064 7988 40116
rect 7562 40008 7988 40064
rect 7562 39956 7624 40008
rect 7676 39956 7988 40008
rect 7562 39900 7988 39956
rect 7562 39848 7624 39900
rect 7676 39848 7988 39900
rect 7562 39792 7988 39848
rect 7562 39740 7624 39792
rect 7676 39740 7988 39792
rect 7562 39684 7988 39740
rect 7562 39632 7624 39684
rect 7676 39632 7988 39684
rect 7562 39576 7988 39632
rect 7562 39524 7624 39576
rect 7676 39524 7988 39576
rect 7562 39468 7988 39524
rect 7562 39416 7624 39468
rect 7676 39416 7988 39468
rect 7562 39360 7988 39416
rect 7562 39308 7624 39360
rect 7676 39308 7988 39360
rect 7562 39252 7988 39308
rect 7562 39200 7624 39252
rect 7676 39200 7988 39252
rect 7562 39144 7988 39200
rect 7562 39092 7624 39144
rect 7676 39092 7988 39144
rect 7562 39036 7988 39092
rect 7562 38984 7624 39036
rect 7676 38984 7988 39036
rect 7562 38928 7988 38984
rect 7562 38876 7624 38928
rect 7676 38876 7988 38928
rect 7562 38820 7988 38876
rect 7562 38768 7624 38820
rect 7676 38768 7988 38820
rect 7562 38712 7988 38768
rect 7562 38660 7624 38712
rect 7676 38660 7988 38712
rect 7562 38604 7988 38660
rect 7562 38552 7624 38604
rect 7676 38552 7988 38604
rect 7562 38496 7988 38552
rect 7562 38444 7624 38496
rect 7676 38444 7988 38496
rect 7562 38388 7988 38444
rect 7562 38336 7624 38388
rect 7676 38336 7988 38388
rect 7562 38280 7988 38336
rect 7562 38228 7624 38280
rect 7676 38228 7988 38280
rect 7562 38172 7988 38228
rect 7562 38120 7624 38172
rect 7676 38120 7988 38172
rect 7562 38064 7988 38120
rect 7562 38012 7624 38064
rect 7676 38012 7988 38064
rect 7562 37956 7988 38012
rect 7562 37904 7624 37956
rect 7676 37904 7988 37956
rect 7562 37848 7988 37904
rect 7562 37796 7624 37848
rect 7676 37796 7988 37848
rect 7562 37740 7988 37796
rect 7562 37688 7624 37740
rect 7676 37688 7988 37740
rect 7562 37632 7988 37688
rect 7562 37580 7624 37632
rect 7676 37580 7988 37632
rect 7562 37524 7988 37580
rect 7562 37472 7624 37524
rect 7676 37472 7988 37524
rect 7562 37256 7988 37472
rect 7562 37204 7625 37256
rect 7677 37204 7749 37256
rect 7801 37204 7873 37256
rect 7925 37204 7988 37256
rect 7562 37132 7988 37204
rect 7562 37080 7625 37132
rect 7677 37080 7749 37132
rect 7801 37080 7873 37132
rect 7925 37080 7988 37132
rect 7562 37008 7988 37080
rect 7562 36956 7625 37008
rect 7677 36956 7749 37008
rect 7801 36956 7873 37008
rect 7925 36956 7988 37008
rect 7562 36884 7988 36956
rect 7562 36832 7625 36884
rect 7677 36832 7749 36884
rect 7801 36832 7873 36884
rect 7925 36832 7988 36884
rect 7562 36760 7988 36832
rect 7562 36708 7625 36760
rect 7677 36708 7749 36760
rect 7801 36708 7873 36760
rect 7925 36708 7988 36760
rect 7562 36492 7988 36708
rect 7562 36440 7624 36492
rect 7676 36440 7988 36492
rect 7562 36384 7988 36440
rect 7562 36332 7624 36384
rect 7676 36332 7988 36384
rect 7562 36276 7988 36332
rect 7562 36251 7624 36276
rect 7676 36251 7988 36276
rect 7562 36195 7623 36251
rect 7679 36195 7747 36251
rect 7803 36195 7871 36251
rect 7927 36195 7988 36251
rect 7562 36168 7988 36195
rect 7562 36127 7624 36168
rect 7676 36127 7988 36168
rect 7562 36071 7623 36127
rect 7679 36071 7747 36127
rect 7803 36071 7871 36127
rect 7927 36071 7988 36127
rect 7562 36060 7988 36071
rect 7562 36008 7624 36060
rect 7676 36008 7988 36060
rect 7562 36003 7988 36008
rect 7562 35947 7623 36003
rect 7679 35947 7747 36003
rect 7803 35947 7871 36003
rect 7927 35947 7988 36003
rect 7562 35900 7624 35947
rect 7676 35900 7988 35947
rect 7562 35879 7988 35900
rect 7562 35823 7623 35879
rect 7679 35823 7747 35879
rect 7803 35823 7871 35879
rect 7927 35823 7988 35879
rect 7562 35792 7624 35823
rect 7676 35792 7988 35823
rect 7562 35755 7988 35792
rect 7562 35699 7623 35755
rect 7679 35699 7747 35755
rect 7803 35699 7871 35755
rect 7927 35699 7988 35755
rect 7562 35684 7624 35699
rect 7676 35684 7988 35699
rect 7562 35631 7988 35684
rect 7562 35575 7623 35631
rect 7679 35575 7747 35631
rect 7803 35575 7871 35631
rect 7927 35575 7988 35631
rect 7562 35520 7988 35575
rect 7562 35507 7624 35520
rect 7676 35507 7988 35520
rect 7562 35451 7623 35507
rect 7679 35451 7747 35507
rect 7803 35451 7871 35507
rect 7927 35451 7988 35507
rect 7562 35412 7988 35451
rect 7562 35383 7624 35412
rect 7676 35383 7988 35412
rect 7562 35327 7623 35383
rect 7679 35327 7747 35383
rect 7803 35327 7871 35383
rect 7927 35327 7988 35383
rect 7562 35304 7988 35327
rect 7562 35259 7624 35304
rect 7676 35259 7988 35304
rect 7562 35203 7623 35259
rect 7679 35203 7747 35259
rect 7803 35203 7871 35259
rect 7927 35203 7988 35259
rect 7562 35196 7988 35203
rect 7562 35144 7624 35196
rect 7676 35144 7988 35196
rect 7562 35135 7988 35144
rect 7562 35079 7623 35135
rect 7679 35079 7747 35135
rect 7803 35079 7871 35135
rect 7927 35079 7988 35135
rect 7562 35036 7624 35079
rect 7676 35036 7988 35079
rect 7562 35011 7988 35036
rect 7562 34955 7623 35011
rect 7679 34955 7747 35011
rect 7803 34955 7871 35011
rect 7927 34955 7988 35011
rect 7562 34928 7624 34955
rect 7676 34928 7988 34955
rect 7562 34887 7988 34928
rect 7562 34831 7623 34887
rect 7679 34831 7747 34887
rect 7803 34831 7871 34887
rect 7927 34831 7988 34887
rect 7562 34820 7624 34831
rect 7676 34820 7988 34831
rect 7562 34764 7988 34820
rect 7562 34763 7624 34764
rect 7676 34763 7988 34764
rect 7562 34707 7623 34763
rect 7679 34707 7747 34763
rect 7803 34707 7871 34763
rect 7927 34707 7988 34763
rect 7562 34656 7988 34707
rect 7562 34639 7624 34656
rect 7676 34639 7988 34656
rect 7562 34583 7623 34639
rect 7679 34583 7747 34639
rect 7803 34583 7871 34639
rect 7927 34583 7988 34639
rect 7562 34548 7988 34583
rect 7562 34515 7624 34548
rect 7676 34515 7988 34548
rect 7562 34459 7623 34515
rect 7679 34459 7747 34515
rect 7803 34459 7871 34515
rect 7927 34459 7988 34515
rect 7562 34440 7988 34459
rect 7562 34391 7624 34440
rect 7676 34391 7988 34440
rect 7562 34335 7623 34391
rect 7679 34335 7747 34391
rect 7803 34335 7871 34391
rect 7927 34335 7988 34391
rect 7562 34332 7988 34335
rect 7562 34280 7624 34332
rect 7676 34280 7988 34332
rect 7562 34267 7988 34280
rect 7562 34211 7623 34267
rect 7679 34211 7747 34267
rect 7803 34211 7871 34267
rect 7927 34211 7988 34267
rect 7562 34172 7624 34211
rect 7676 34172 7988 34211
rect 7562 34143 7988 34172
rect 7562 34087 7623 34143
rect 7679 34087 7747 34143
rect 7803 34087 7871 34143
rect 7927 34087 7988 34143
rect 7562 34064 7624 34087
rect 7676 34064 7988 34087
rect 7562 34019 7988 34064
rect 7562 33963 7623 34019
rect 7679 33963 7747 34019
rect 7803 33963 7871 34019
rect 7927 33963 7988 34019
rect 7562 33956 7624 33963
rect 7676 33956 7988 33963
rect 7562 33900 7988 33956
rect 7562 33895 7624 33900
rect 7676 33895 7988 33900
rect 7562 33839 7623 33895
rect 7679 33839 7747 33895
rect 7803 33839 7871 33895
rect 7927 33839 7988 33895
rect 7562 33792 7988 33839
rect 7562 33771 7624 33792
rect 7676 33771 7988 33792
rect 7562 33715 7623 33771
rect 7679 33715 7747 33771
rect 7803 33715 7871 33771
rect 7927 33715 7988 33771
rect 7562 33684 7988 33715
rect 7562 33647 7624 33684
rect 7676 33647 7988 33684
rect 7562 33591 7623 33647
rect 7679 33591 7747 33647
rect 7803 33591 7871 33647
rect 7927 33591 7988 33647
rect 7562 33576 7988 33591
rect 7562 33524 7624 33576
rect 7676 33524 7988 33576
rect 7562 33523 7988 33524
rect 7562 33467 7623 33523
rect 7679 33467 7747 33523
rect 7803 33467 7871 33523
rect 7927 33467 7988 33523
rect 7562 33399 7988 33467
rect 7562 33343 7623 33399
rect 7679 33343 7747 33399
rect 7803 33343 7871 33399
rect 7927 33343 7988 33399
rect 7562 33308 7988 33343
rect 7562 33256 7625 33308
rect 7677 33256 7749 33308
rect 7801 33256 7873 33308
rect 7925 33256 7988 33308
rect 7562 33184 7988 33256
rect 7562 33132 7625 33184
rect 7677 33132 7749 33184
rect 7801 33132 7873 33184
rect 7925 33132 7988 33184
rect 7562 33060 7988 33132
rect 7562 33008 7625 33060
rect 7677 33008 7749 33060
rect 7801 33008 7873 33060
rect 7925 33008 7988 33060
rect 7562 32936 7988 33008
rect 7562 32884 7625 32936
rect 7677 32884 7749 32936
rect 7801 32884 7873 32936
rect 7925 32884 7988 32936
rect 7562 32812 7988 32884
rect 7562 32760 7625 32812
rect 7677 32760 7749 32812
rect 7801 32760 7873 32812
rect 7925 32760 7988 32812
rect 7562 32544 7988 32760
rect 7562 32492 7624 32544
rect 7676 32492 7988 32544
rect 7562 32436 7988 32492
rect 7562 32384 7624 32436
rect 7676 32384 7988 32436
rect 7562 32328 7988 32384
rect 7562 32276 7624 32328
rect 7676 32276 7988 32328
rect 7562 32220 7988 32276
rect 7562 32168 7624 32220
rect 7676 32168 7988 32220
rect 7562 32112 7988 32168
rect 7562 32060 7624 32112
rect 7676 32060 7988 32112
rect 7562 32004 7988 32060
rect 7562 31952 7624 32004
rect 7676 31952 7988 32004
rect 7562 31896 7988 31952
rect 7562 31844 7624 31896
rect 7676 31844 7988 31896
rect 7562 31788 7988 31844
rect 7562 31736 7624 31788
rect 7676 31736 7988 31788
rect 7562 31680 7988 31736
rect 7562 31628 7624 31680
rect 7676 31628 7988 31680
rect 7562 31572 7988 31628
rect 7562 31520 7624 31572
rect 7676 31520 7988 31572
rect 7562 31464 7988 31520
rect 7562 31412 7624 31464
rect 7676 31412 7988 31464
rect 7562 31356 7988 31412
rect 7562 31304 7624 31356
rect 7676 31304 7988 31356
rect 7562 31248 7988 31304
rect 7562 31196 7624 31248
rect 7676 31196 7988 31248
rect 7562 31140 7988 31196
rect 7562 31088 7624 31140
rect 7676 31088 7988 31140
rect 7562 31032 7988 31088
rect 7562 30980 7624 31032
rect 7676 30980 7988 31032
rect 7562 30924 7988 30980
rect 7562 30872 7624 30924
rect 7676 30872 7988 30924
rect 7562 30816 7988 30872
rect 7562 30764 7624 30816
rect 7676 30764 7988 30816
rect 7562 30708 7988 30764
rect 7562 30656 7624 30708
rect 7676 30656 7988 30708
rect 7562 30600 7988 30656
rect 7562 30548 7624 30600
rect 7676 30548 7988 30600
rect 7562 30492 7988 30548
rect 7562 30440 7624 30492
rect 7676 30440 7988 30492
rect 7562 30384 7988 30440
rect 7562 30332 7624 30384
rect 7676 30332 7988 30384
rect 7562 30276 7988 30332
rect 7562 30224 7624 30276
rect 7676 30224 7988 30276
rect 7562 30168 7988 30224
rect 7562 30116 7624 30168
rect 7676 30116 7988 30168
rect 7562 30060 7988 30116
rect 7562 30008 7624 30060
rect 7676 30008 7988 30060
rect 7562 29952 7988 30008
rect 7562 29900 7624 29952
rect 7676 29900 7988 29952
rect 7562 29844 7988 29900
rect 7562 29792 7624 29844
rect 7676 29792 7988 29844
rect 7562 29736 7988 29792
rect 7562 29684 7624 29736
rect 7676 29684 7988 29736
rect 7562 29628 7988 29684
rect 7562 29576 7624 29628
rect 7676 29576 7988 29628
rect 7562 29360 7988 29576
rect 7562 29308 7625 29360
rect 7677 29308 7749 29360
rect 7801 29308 7873 29360
rect 7925 29308 7988 29360
rect 7562 29236 7988 29308
rect 7562 29184 7625 29236
rect 7677 29184 7749 29236
rect 7801 29184 7873 29236
rect 7925 29184 7988 29236
rect 7562 29112 7988 29184
rect 7562 29060 7625 29112
rect 7677 29060 7749 29112
rect 7801 29060 7873 29112
rect 7925 29060 7988 29112
rect 7562 28988 7988 29060
rect 7562 28936 7625 28988
rect 7677 28936 7749 28988
rect 7801 28936 7873 28988
rect 7925 28936 7988 28988
rect 7562 28864 7988 28936
rect 7562 28812 7625 28864
rect 7677 28812 7749 28864
rect 7801 28812 7873 28864
rect 7925 28812 7988 28864
rect 7562 28596 7988 28812
rect 7562 28544 7624 28596
rect 7676 28544 7988 28596
rect 7562 28488 7988 28544
rect 7562 28436 7624 28488
rect 7676 28436 7988 28488
rect 7562 28380 7988 28436
rect 7562 28328 7624 28380
rect 7676 28328 7988 28380
rect 7562 28272 7988 28328
rect 7562 28245 7624 28272
rect 7676 28245 7988 28272
rect 7562 28189 7623 28245
rect 7679 28189 7747 28245
rect 7803 28189 7871 28245
rect 7927 28189 7988 28245
rect 7562 28164 7988 28189
rect 7562 28121 7624 28164
rect 7676 28121 7988 28164
rect 7562 28065 7623 28121
rect 7679 28065 7747 28121
rect 7803 28065 7871 28121
rect 7927 28065 7988 28121
rect 7562 28056 7988 28065
rect 7562 28004 7624 28056
rect 7676 28004 7988 28056
rect 7562 27997 7988 28004
rect 7562 27941 7623 27997
rect 7679 27941 7747 27997
rect 7803 27941 7871 27997
rect 7927 27941 7988 27997
rect 7562 27896 7624 27941
rect 7676 27896 7988 27941
rect 7562 27873 7988 27896
rect 7562 27817 7623 27873
rect 7679 27817 7747 27873
rect 7803 27817 7871 27873
rect 7927 27817 7988 27873
rect 7562 27788 7624 27817
rect 7676 27788 7988 27817
rect 7562 27749 7988 27788
rect 7562 27693 7623 27749
rect 7679 27693 7747 27749
rect 7803 27693 7871 27749
rect 7927 27693 7988 27749
rect 7562 27680 7624 27693
rect 7676 27680 7988 27693
rect 7562 27625 7988 27680
rect 7562 27569 7623 27625
rect 7679 27569 7747 27625
rect 7803 27569 7871 27625
rect 7927 27569 7988 27625
rect 7562 27516 7988 27569
rect 7562 27501 7624 27516
rect 7676 27501 7988 27516
rect 7562 27445 7623 27501
rect 7679 27445 7747 27501
rect 7803 27445 7871 27501
rect 7927 27445 7988 27501
rect 7562 27408 7988 27445
rect 7562 27377 7624 27408
rect 7676 27377 7988 27408
rect 7562 27321 7623 27377
rect 7679 27321 7747 27377
rect 7803 27321 7871 27377
rect 7927 27321 7988 27377
rect 7562 27300 7988 27321
rect 7562 27253 7624 27300
rect 7676 27253 7988 27300
rect 7562 27197 7623 27253
rect 7679 27197 7747 27253
rect 7803 27197 7871 27253
rect 7927 27197 7988 27253
rect 7562 27192 7988 27197
rect 7562 27140 7624 27192
rect 7676 27140 7988 27192
rect 7562 27129 7988 27140
rect 7562 27073 7623 27129
rect 7679 27073 7747 27129
rect 7803 27073 7871 27129
rect 7927 27073 7988 27129
rect 7562 27032 7624 27073
rect 7676 27032 7988 27073
rect 7562 27005 7988 27032
rect 7562 26949 7623 27005
rect 7679 26949 7747 27005
rect 7803 26949 7871 27005
rect 7927 26949 7988 27005
rect 7562 26924 7624 26949
rect 7676 26924 7988 26949
rect 7562 26868 7988 26924
rect 7562 26816 7624 26868
rect 7676 26816 7988 26868
rect 7562 26760 7988 26816
rect 7562 26708 7624 26760
rect 7676 26708 7988 26760
rect 7562 26652 7988 26708
rect 7562 26600 7624 26652
rect 7676 26600 7988 26652
rect 7562 26544 7988 26600
rect 7562 26492 7624 26544
rect 7676 26492 7988 26544
rect 7562 26436 7988 26492
rect 7562 26384 7624 26436
rect 7676 26384 7988 26436
rect 7562 26328 7988 26384
rect 7562 26276 7624 26328
rect 7676 26276 7988 26328
rect 7562 26220 7988 26276
rect 7562 26168 7624 26220
rect 7676 26168 7988 26220
rect 7562 26112 7988 26168
rect 7562 26060 7624 26112
rect 7676 26060 7988 26112
rect 7562 26004 7988 26060
rect 7562 25952 7624 26004
rect 7676 25952 7988 26004
rect 7562 25896 7988 25952
rect 7562 25844 7624 25896
rect 7676 25844 7988 25896
rect 7562 25788 7988 25844
rect 7562 25736 7624 25788
rect 7676 25736 7988 25788
rect 7562 25680 7988 25736
rect 7562 25628 7624 25680
rect 7676 25628 7988 25680
rect 7562 25412 7988 25628
rect 7562 25360 7625 25412
rect 7677 25360 7749 25412
rect 7801 25360 7873 25412
rect 7925 25360 7988 25412
rect 7562 25288 7988 25360
rect 7562 25236 7625 25288
rect 7677 25236 7749 25288
rect 7801 25236 7873 25288
rect 7925 25236 7988 25288
rect 7562 25164 7988 25236
rect 7562 25112 7625 25164
rect 7677 25112 7749 25164
rect 7801 25112 7873 25164
rect 7925 25112 7988 25164
rect 7562 25040 7988 25112
rect 7562 24988 7625 25040
rect 7677 24988 7749 25040
rect 7801 24988 7873 25040
rect 7925 24988 7988 25040
rect 7562 24916 7988 24988
rect 7562 24864 7625 24916
rect 7677 24864 7749 24916
rect 7801 24864 7873 24916
rect 7925 24864 7988 24916
rect 7562 24648 7988 24864
rect 7562 24596 7624 24648
rect 7676 24596 7988 24648
rect 7562 24540 7988 24596
rect 7562 24488 7624 24540
rect 7676 24488 7988 24540
rect 7562 24432 7988 24488
rect 7562 24380 7624 24432
rect 7676 24380 7988 24432
rect 7562 24324 7988 24380
rect 7562 24272 7624 24324
rect 7676 24272 7988 24324
rect 7562 24216 7988 24272
rect 7562 24164 7624 24216
rect 7676 24164 7988 24216
rect 7562 24108 7988 24164
rect 7562 24056 7624 24108
rect 7676 24056 7988 24108
rect 7562 24000 7988 24056
rect 7562 23948 7624 24000
rect 7676 23948 7988 24000
rect 7562 23892 7988 23948
rect 7562 23840 7624 23892
rect 7676 23840 7988 23892
rect 7562 23784 7988 23840
rect 7562 23732 7624 23784
rect 7676 23732 7988 23784
rect 7562 23676 7988 23732
rect 7562 23624 7624 23676
rect 7676 23624 7988 23676
rect 7562 23568 7988 23624
rect 7562 23516 7624 23568
rect 7676 23516 7988 23568
rect 7562 23460 7988 23516
rect 7562 23408 7624 23460
rect 7676 23408 7988 23460
rect 7562 23352 7988 23408
rect 7562 23300 7624 23352
rect 7676 23300 7988 23352
rect 7562 23244 7988 23300
rect 7562 23192 7624 23244
rect 7676 23192 7988 23244
rect 7562 23136 7988 23192
rect 7562 23084 7624 23136
rect 7676 23084 7988 23136
rect 7562 23028 7988 23084
rect 7562 22976 7624 23028
rect 7676 22976 7988 23028
rect 7562 22920 7988 22976
rect 7562 22868 7624 22920
rect 7676 22868 7988 22920
rect 7562 22812 7988 22868
rect 7562 22760 7624 22812
rect 7676 22760 7988 22812
rect 7562 22704 7988 22760
rect 7562 22652 7624 22704
rect 7676 22652 7988 22704
rect 7562 22596 7988 22652
rect 7562 22544 7624 22596
rect 7676 22544 7988 22596
rect 7562 22488 7988 22544
rect 7562 22436 7624 22488
rect 7676 22436 7988 22488
rect 7562 22380 7988 22436
rect 7562 22328 7624 22380
rect 7676 22328 7988 22380
rect 7562 22272 7988 22328
rect 7562 22220 7624 22272
rect 7676 22220 7988 22272
rect 7562 22164 7988 22220
rect 7562 22112 7624 22164
rect 7676 22112 7988 22164
rect 7562 22056 7988 22112
rect 7562 22004 7624 22056
rect 7676 22004 7988 22056
rect 7562 21948 7988 22004
rect 7562 21896 7624 21948
rect 7676 21896 7988 21948
rect 7562 21840 7988 21896
rect 7562 21788 7624 21840
rect 7676 21788 7988 21840
rect 7562 21732 7988 21788
rect 7562 21680 7624 21732
rect 7676 21680 7988 21732
rect 7562 21469 7988 21680
rect 7562 21417 7587 21469
rect 7639 21417 7695 21469
rect 7747 21417 7803 21469
rect 7855 21417 7911 21469
rect 7963 21417 7988 21469
rect 7562 21361 7988 21417
rect 7562 21309 7587 21361
rect 7639 21309 7695 21361
rect 7747 21309 7803 21361
rect 7855 21309 7911 21361
rect 7963 21309 7988 21361
rect 7562 21253 7988 21309
rect 7562 21201 7587 21253
rect 7639 21201 7695 21253
rect 7747 21201 7803 21253
rect 7855 21201 7911 21253
rect 7963 21201 7988 21253
rect 7562 19951 7988 21201
rect 7562 19899 7587 19951
rect 7639 19899 7695 19951
rect 7747 19899 7803 19951
rect 7855 19899 7911 19951
rect 7963 19899 7988 19951
rect 7562 19843 7988 19899
rect 7562 19791 7587 19843
rect 7639 19791 7695 19843
rect 7747 19791 7803 19843
rect 7855 19791 7911 19843
rect 7963 19791 7988 19843
rect 7562 19202 7988 19791
rect 7562 19150 7587 19202
rect 7639 19150 7695 19202
rect 7747 19150 7803 19202
rect 7855 19150 7911 19202
rect 7963 19150 7988 19202
rect 7562 19094 7988 19150
rect 7562 19042 7587 19094
rect 7639 19042 7695 19094
rect 7747 19042 7803 19094
rect 7855 19042 7911 19094
rect 7963 19042 7988 19094
rect 7562 18986 7988 19042
rect 7562 18934 7587 18986
rect 7639 18934 7695 18986
rect 7747 18934 7803 18986
rect 7855 18934 7911 18986
rect 7963 18934 7988 18986
rect 7562 18330 7988 18934
rect 7562 18278 7587 18330
rect 7639 18278 7695 18330
rect 7747 18278 7803 18330
rect 7855 18278 7911 18330
rect 7963 18278 7988 18330
rect 7562 18222 7988 18278
rect 7562 18170 7587 18222
rect 7639 18170 7695 18222
rect 7747 18170 7803 18222
rect 7855 18170 7911 18222
rect 7963 18170 7988 18222
rect 7562 18114 7988 18170
rect 7562 18062 7587 18114
rect 7639 18062 7695 18114
rect 7747 18062 7803 18114
rect 7855 18062 7911 18114
rect 7963 18062 7988 18114
rect 7562 17458 7988 18062
rect 7562 17406 7587 17458
rect 7639 17406 7695 17458
rect 7747 17406 7803 17458
rect 7855 17406 7911 17458
rect 7963 17406 7988 17458
rect 7562 17350 7988 17406
rect 7562 17298 7587 17350
rect 7639 17298 7695 17350
rect 7747 17298 7803 17350
rect 7855 17298 7911 17350
rect 7963 17298 7988 17350
rect 7562 17242 7988 17298
rect 7562 17190 7587 17242
rect 7639 17190 7695 17242
rect 7747 17190 7803 17242
rect 7855 17190 7911 17242
rect 7963 17190 7988 17242
rect 7562 16601 7988 17190
rect 7562 16549 7587 16601
rect 7639 16549 7695 16601
rect 7747 16549 7803 16601
rect 7855 16549 7911 16601
rect 7963 16549 7988 16601
rect 7562 16493 7988 16549
rect 7562 16441 7587 16493
rect 7639 16441 7695 16493
rect 7747 16441 7803 16493
rect 7855 16441 7911 16493
rect 7963 16441 7988 16493
rect 7562 15762 7988 16441
rect 8616 56286 9124 56975
rect 8616 56234 8677 56286
rect 8729 56234 9124 56286
rect 8616 56178 9124 56234
rect 8616 56126 8677 56178
rect 8729 56126 9124 56178
rect 8616 56070 9124 56126
rect 8616 56018 8677 56070
rect 8729 56018 9124 56070
rect 8616 55962 9124 56018
rect 8616 55910 8677 55962
rect 8729 55910 9124 55962
rect 8616 55854 9124 55910
rect 8616 55802 8677 55854
rect 8729 55802 9124 55854
rect 8616 55746 9124 55802
rect 8616 55694 8677 55746
rect 8729 55694 9124 55746
rect 8616 55638 9124 55694
rect 8616 55586 8677 55638
rect 8729 55586 9124 55638
rect 8616 55530 9124 55586
rect 8616 55478 8677 55530
rect 8729 55478 9124 55530
rect 8616 55445 9124 55478
rect 8616 55389 8656 55445
rect 8712 55422 8780 55445
rect 8729 55389 8780 55422
rect 8836 55389 8904 55445
rect 8960 55389 9028 55445
rect 9084 55389 9124 55445
rect 8616 55370 8677 55389
rect 8729 55370 9124 55389
rect 8616 55321 9124 55370
rect 8616 55265 8656 55321
rect 8712 55314 8780 55321
rect 8729 55265 8780 55314
rect 8836 55265 8904 55321
rect 8960 55265 9028 55321
rect 9084 55265 9124 55321
rect 8616 55262 8677 55265
rect 8729 55262 9124 55265
rect 8616 55206 9124 55262
rect 8616 55197 8677 55206
rect 8729 55197 9124 55206
rect 8616 55141 8656 55197
rect 8729 55154 8780 55197
rect 8712 55141 8780 55154
rect 8836 55141 8904 55197
rect 8960 55141 9028 55197
rect 9084 55141 9124 55197
rect 8616 55098 9124 55141
rect 8616 55073 8677 55098
rect 8729 55073 9124 55098
rect 8616 55017 8656 55073
rect 8729 55046 8780 55073
rect 8712 55017 8780 55046
rect 8836 55017 8904 55073
rect 8960 55017 9028 55073
rect 9084 55017 9124 55073
rect 8616 54990 9124 55017
rect 8616 54949 8677 54990
rect 8729 54949 9124 54990
rect 8616 54893 8656 54949
rect 8729 54938 8780 54949
rect 8712 54893 8780 54938
rect 8836 54893 8904 54949
rect 8960 54893 9028 54949
rect 9084 54893 9124 54949
rect 8616 54882 9124 54893
rect 8616 54830 8677 54882
rect 8729 54830 9124 54882
rect 8616 54825 9124 54830
rect 8616 54769 8656 54825
rect 8712 54774 8780 54825
rect 8729 54769 8780 54774
rect 8836 54769 8904 54825
rect 8960 54769 9028 54825
rect 9084 54769 9124 54825
rect 8616 54722 8677 54769
rect 8729 54722 9124 54769
rect 8616 54701 9124 54722
rect 8616 54645 8656 54701
rect 8712 54666 8780 54701
rect 8729 54645 8780 54666
rect 8836 54645 8904 54701
rect 8960 54645 9028 54701
rect 9084 54645 9124 54701
rect 8616 54614 8677 54645
rect 8729 54614 9124 54645
rect 8616 54577 9124 54614
rect 8616 54521 8656 54577
rect 8712 54558 8780 54577
rect 8729 54521 8780 54558
rect 8836 54521 8904 54577
rect 8960 54521 9028 54577
rect 9084 54521 9124 54577
rect 8616 54506 8677 54521
rect 8729 54506 9124 54521
rect 8616 54453 9124 54506
rect 8616 54397 8656 54453
rect 8712 54450 8780 54453
rect 8729 54398 8780 54450
rect 8712 54397 8780 54398
rect 8836 54397 8904 54453
rect 8960 54397 9028 54453
rect 9084 54397 9124 54453
rect 8616 54342 9124 54397
rect 8616 54329 8677 54342
rect 8729 54329 9124 54342
rect 8616 54273 8656 54329
rect 8729 54290 8780 54329
rect 8712 54273 8780 54290
rect 8836 54273 8904 54329
rect 8960 54273 9028 54329
rect 9084 54273 9124 54329
rect 8616 54234 9124 54273
rect 8616 54205 8677 54234
rect 8729 54205 9124 54234
rect 8616 54149 8656 54205
rect 8729 54182 8780 54205
rect 8712 54149 8780 54182
rect 8836 54149 8904 54205
rect 8960 54149 9028 54205
rect 9084 54149 9124 54205
rect 8616 54126 9124 54149
rect 8616 54074 8677 54126
rect 8729 54074 9124 54126
rect 8616 54018 9124 54074
rect 8616 53966 8677 54018
rect 8729 53966 9124 54018
rect 8616 53910 9124 53966
rect 8616 53858 8677 53910
rect 8729 53858 9124 53910
rect 8616 53802 9124 53858
rect 8616 53750 8677 53802
rect 8729 53750 9124 53802
rect 8616 53694 9124 53750
rect 8616 53642 8677 53694
rect 8729 53642 9124 53694
rect 8616 53586 9124 53642
rect 8616 53534 8677 53586
rect 8729 53534 9124 53586
rect 8616 53478 9124 53534
rect 8616 53426 8677 53478
rect 8729 53426 9124 53478
rect 8616 53370 9124 53426
rect 8616 53318 8677 53370
rect 8729 53318 9124 53370
rect 8616 53262 9124 53318
rect 8616 53210 8677 53262
rect 8729 53210 9124 53262
rect 8616 52338 9124 53210
rect 8616 52286 8677 52338
rect 8729 52286 9124 52338
rect 8616 52230 9124 52286
rect 8616 52178 8677 52230
rect 8729 52178 9124 52230
rect 8616 52122 9124 52178
rect 8616 52070 8677 52122
rect 8729 52070 9124 52122
rect 8616 52014 9124 52070
rect 8616 51962 8677 52014
rect 8729 51962 9124 52014
rect 8616 51906 9124 51962
rect 8616 51854 8677 51906
rect 8729 51854 9124 51906
rect 8616 51798 9124 51854
rect 8616 51746 8677 51798
rect 8729 51746 9124 51798
rect 8616 51690 9124 51746
rect 8616 51638 8677 51690
rect 8729 51638 9124 51690
rect 8616 51582 9124 51638
rect 8616 51530 8677 51582
rect 8729 51530 9124 51582
rect 8616 51474 9124 51530
rect 8616 51422 8677 51474
rect 8729 51422 9124 51474
rect 8616 51366 9124 51422
rect 8616 51314 8677 51366
rect 8729 51314 9124 51366
rect 8616 51258 9124 51314
rect 8616 51206 8677 51258
rect 8729 51206 9124 51258
rect 8616 51150 9124 51206
rect 8616 51098 8677 51150
rect 8729 51098 9124 51150
rect 8616 51042 9124 51098
rect 8616 50990 8677 51042
rect 8729 50990 9124 51042
rect 8616 50934 9124 50990
rect 8616 50882 8677 50934
rect 8729 50882 9124 50934
rect 8616 50826 9124 50882
rect 8616 50774 8677 50826
rect 8729 50774 9124 50826
rect 8616 50718 9124 50774
rect 8616 50666 8677 50718
rect 8729 50666 9124 50718
rect 8616 50610 9124 50666
rect 8616 50558 8677 50610
rect 8729 50558 9124 50610
rect 8616 50502 9124 50558
rect 8616 50450 8677 50502
rect 8729 50450 9124 50502
rect 8616 50394 9124 50450
rect 8616 50342 8677 50394
rect 8729 50342 9124 50394
rect 8616 50286 9124 50342
rect 8616 50234 8677 50286
rect 8729 50234 9124 50286
rect 8616 50178 9124 50234
rect 8616 50126 8677 50178
rect 8729 50126 9124 50178
rect 8616 50070 9124 50126
rect 8616 50018 8677 50070
rect 8729 50018 9124 50070
rect 8616 49962 9124 50018
rect 8616 49910 8677 49962
rect 8729 49910 9124 49962
rect 8616 49854 9124 49910
rect 8616 49802 8677 49854
rect 8729 49802 9124 49854
rect 8616 49746 9124 49802
rect 8616 49694 8677 49746
rect 8729 49694 9124 49746
rect 8616 49638 9124 49694
rect 8616 49586 8677 49638
rect 8729 49586 9124 49638
rect 8616 49530 9124 49586
rect 8616 49478 8677 49530
rect 8729 49478 9124 49530
rect 8616 49422 9124 49478
rect 8616 49370 8677 49422
rect 8729 49370 9124 49422
rect 8616 49314 9124 49370
rect 8616 49262 8677 49314
rect 8729 49262 9124 49314
rect 8616 48390 9124 49262
rect 8616 48338 8677 48390
rect 8729 48338 9124 48390
rect 8616 48282 9124 48338
rect 8616 48230 8677 48282
rect 8729 48230 9124 48282
rect 8616 48174 9124 48230
rect 8616 48122 8677 48174
rect 8729 48122 9124 48174
rect 8616 48066 9124 48122
rect 8616 48014 8677 48066
rect 8729 48014 9124 48066
rect 8616 47958 9124 48014
rect 8616 47906 8677 47958
rect 8729 47906 9124 47958
rect 8616 47850 9124 47906
rect 8616 47798 8677 47850
rect 8729 47798 9124 47850
rect 8616 47742 9124 47798
rect 8616 47690 8677 47742
rect 8729 47690 9124 47742
rect 8616 47634 9124 47690
rect 8616 47582 8677 47634
rect 8729 47582 9124 47634
rect 8616 47526 9124 47582
rect 8616 47474 8677 47526
rect 8729 47474 9124 47526
rect 8616 47445 9124 47474
rect 8616 47389 8656 47445
rect 8712 47418 8780 47445
rect 8729 47389 8780 47418
rect 8836 47389 8904 47445
rect 8960 47389 9028 47445
rect 9084 47389 9124 47445
rect 8616 47366 8677 47389
rect 8729 47366 9124 47389
rect 8616 47321 9124 47366
rect 8616 47265 8656 47321
rect 8712 47310 8780 47321
rect 8729 47265 8780 47310
rect 8836 47265 8904 47321
rect 8960 47265 9028 47321
rect 9084 47265 9124 47321
rect 8616 47258 8677 47265
rect 8729 47258 9124 47265
rect 8616 47202 9124 47258
rect 8616 47197 8677 47202
rect 8729 47197 9124 47202
rect 8616 47141 8656 47197
rect 8729 47150 8780 47197
rect 8712 47141 8780 47150
rect 8836 47141 8904 47197
rect 8960 47141 9028 47197
rect 9084 47141 9124 47197
rect 8616 47094 9124 47141
rect 8616 47073 8677 47094
rect 8729 47073 9124 47094
rect 8616 47017 8656 47073
rect 8729 47042 8780 47073
rect 8712 47017 8780 47042
rect 8836 47017 8904 47073
rect 8960 47017 9028 47073
rect 9084 47017 9124 47073
rect 8616 46986 9124 47017
rect 8616 46949 8677 46986
rect 8729 46949 9124 46986
rect 8616 46893 8656 46949
rect 8729 46934 8780 46949
rect 8712 46893 8780 46934
rect 8836 46893 8904 46949
rect 8960 46893 9028 46949
rect 9084 46893 9124 46949
rect 8616 46878 9124 46893
rect 8616 46826 8677 46878
rect 8729 46826 9124 46878
rect 8616 46825 9124 46826
rect 8616 46769 8656 46825
rect 8712 46770 8780 46825
rect 8729 46769 8780 46770
rect 8836 46769 8904 46825
rect 8960 46769 9028 46825
rect 9084 46769 9124 46825
rect 8616 46718 8677 46769
rect 8729 46718 9124 46769
rect 8616 46701 9124 46718
rect 8616 46645 8656 46701
rect 8712 46662 8780 46701
rect 8729 46645 8780 46662
rect 8836 46645 8904 46701
rect 8960 46645 9028 46701
rect 9084 46645 9124 46701
rect 8616 46610 8677 46645
rect 8729 46610 9124 46645
rect 8616 46577 9124 46610
rect 8616 46521 8656 46577
rect 8712 46554 8780 46577
rect 8729 46521 8780 46554
rect 8836 46521 8904 46577
rect 8960 46521 9028 46577
rect 9084 46521 9124 46577
rect 8616 46502 8677 46521
rect 8729 46502 9124 46521
rect 8616 46453 9124 46502
rect 8616 46397 8656 46453
rect 8712 46446 8780 46453
rect 8729 46397 8780 46446
rect 8836 46397 8904 46453
rect 8960 46397 9028 46453
rect 9084 46397 9124 46453
rect 8616 46394 8677 46397
rect 8729 46394 9124 46397
rect 8616 46338 9124 46394
rect 8616 46329 8677 46338
rect 8729 46329 9124 46338
rect 8616 46273 8656 46329
rect 8729 46286 8780 46329
rect 8712 46273 8780 46286
rect 8836 46273 8904 46329
rect 8960 46273 9028 46329
rect 9084 46273 9124 46329
rect 8616 46230 9124 46273
rect 8616 46205 8677 46230
rect 8729 46205 9124 46230
rect 8616 46149 8656 46205
rect 8729 46178 8780 46205
rect 8712 46149 8780 46178
rect 8836 46149 8904 46205
rect 8960 46149 9028 46205
rect 9084 46149 9124 46205
rect 8616 46122 9124 46149
rect 8616 46070 8677 46122
rect 8729 46070 9124 46122
rect 8616 46014 9124 46070
rect 8616 45962 8677 46014
rect 8729 45962 9124 46014
rect 8616 45906 9124 45962
rect 8616 45854 8677 45906
rect 8729 45854 9124 45906
rect 8616 45798 9124 45854
rect 8616 45746 8677 45798
rect 8729 45746 9124 45798
rect 8616 45690 9124 45746
rect 8616 45638 8677 45690
rect 8729 45638 9124 45690
rect 8616 45582 9124 45638
rect 8616 45530 8677 45582
rect 8729 45530 9124 45582
rect 8616 45474 9124 45530
rect 8616 45422 8677 45474
rect 8729 45422 9124 45474
rect 8616 45366 9124 45422
rect 8616 45314 8677 45366
rect 8729 45314 9124 45366
rect 8616 44442 9124 45314
rect 8616 44390 8677 44442
rect 8729 44390 9124 44442
rect 8616 44334 9124 44390
rect 8616 44282 8677 44334
rect 8729 44282 9124 44334
rect 8616 44245 9124 44282
rect 8616 44189 8656 44245
rect 8712 44226 8780 44245
rect 8729 44189 8780 44226
rect 8836 44189 8904 44245
rect 8960 44189 9028 44245
rect 9084 44189 9124 44245
rect 8616 44174 8677 44189
rect 8729 44174 9124 44189
rect 8616 44121 9124 44174
rect 8616 44065 8656 44121
rect 8712 44118 8780 44121
rect 8729 44066 8780 44118
rect 8712 44065 8780 44066
rect 8836 44065 8904 44121
rect 8960 44065 9028 44121
rect 9084 44065 9124 44121
rect 8616 44010 9124 44065
rect 8616 43997 8677 44010
rect 8729 43997 9124 44010
rect 8616 43941 8656 43997
rect 8729 43958 8780 43997
rect 8712 43941 8780 43958
rect 8836 43941 8904 43997
rect 8960 43941 9028 43997
rect 9084 43941 9124 43997
rect 8616 43902 9124 43941
rect 8616 43873 8677 43902
rect 8729 43873 9124 43902
rect 8616 43817 8656 43873
rect 8729 43850 8780 43873
rect 8712 43817 8780 43850
rect 8836 43817 8904 43873
rect 8960 43817 9028 43873
rect 9084 43817 9124 43873
rect 8616 43794 9124 43817
rect 8616 43749 8677 43794
rect 8729 43749 9124 43794
rect 8616 43693 8656 43749
rect 8729 43742 8780 43749
rect 8712 43693 8780 43742
rect 8836 43693 8904 43749
rect 8960 43693 9028 43749
rect 9084 43693 9124 43749
rect 8616 43686 9124 43693
rect 8616 43634 8677 43686
rect 8729 43634 9124 43686
rect 8616 43625 9124 43634
rect 8616 43569 8656 43625
rect 8712 43578 8780 43625
rect 8729 43569 8780 43578
rect 8836 43569 8904 43625
rect 8960 43569 9028 43625
rect 9084 43569 9124 43625
rect 8616 43526 8677 43569
rect 8729 43526 9124 43569
rect 8616 43501 9124 43526
rect 8616 43445 8656 43501
rect 8712 43470 8780 43501
rect 8729 43445 8780 43470
rect 8836 43445 8904 43501
rect 8960 43445 9028 43501
rect 9084 43445 9124 43501
rect 8616 43418 8677 43445
rect 8729 43418 9124 43445
rect 8616 43377 9124 43418
rect 8616 43321 8656 43377
rect 8712 43362 8780 43377
rect 8729 43321 8780 43362
rect 8836 43321 8904 43377
rect 8960 43321 9028 43377
rect 9084 43321 9124 43377
rect 8616 43310 8677 43321
rect 8729 43310 9124 43321
rect 8616 43254 9124 43310
rect 8616 43253 8677 43254
rect 8729 43253 9124 43254
rect 8616 43197 8656 43253
rect 8729 43202 8780 43253
rect 8712 43197 8780 43202
rect 8836 43197 8904 43253
rect 8960 43197 9028 43253
rect 9084 43197 9124 43253
rect 8616 43146 9124 43197
rect 8616 43129 8677 43146
rect 8729 43129 9124 43146
rect 8616 43073 8656 43129
rect 8729 43094 8780 43129
rect 8712 43073 8780 43094
rect 8836 43073 8904 43129
rect 8960 43073 9028 43129
rect 9084 43073 9124 43129
rect 8616 43038 9124 43073
rect 8616 43005 8677 43038
rect 8729 43005 9124 43038
rect 8616 42949 8656 43005
rect 8729 42986 8780 43005
rect 8712 42949 8780 42986
rect 8836 42949 8904 43005
rect 8960 42949 9028 43005
rect 9084 42949 9124 43005
rect 8616 42930 9124 42949
rect 8616 42878 8677 42930
rect 8729 42878 9124 42930
rect 8616 42822 9124 42878
rect 8616 42770 8677 42822
rect 8729 42770 9124 42822
rect 8616 42714 9124 42770
rect 8616 42662 8677 42714
rect 8729 42662 9124 42714
rect 8616 42645 9124 42662
rect 8616 42589 8656 42645
rect 8712 42606 8780 42645
rect 8729 42589 8780 42606
rect 8836 42589 8904 42645
rect 8960 42589 9028 42645
rect 9084 42589 9124 42645
rect 8616 42554 8677 42589
rect 8729 42554 9124 42589
rect 8616 42521 9124 42554
rect 8616 42465 8656 42521
rect 8712 42498 8780 42521
rect 8729 42465 8780 42498
rect 8836 42465 8904 42521
rect 8960 42465 9028 42521
rect 9084 42465 9124 42521
rect 8616 42446 8677 42465
rect 8729 42446 9124 42465
rect 8616 42397 9124 42446
rect 8616 42341 8656 42397
rect 8712 42390 8780 42397
rect 8729 42341 8780 42390
rect 8836 42341 8904 42397
rect 8960 42341 9028 42397
rect 9084 42341 9124 42397
rect 8616 42338 8677 42341
rect 8729 42338 9124 42341
rect 8616 42282 9124 42338
rect 8616 42273 8677 42282
rect 8729 42273 9124 42282
rect 8616 42217 8656 42273
rect 8729 42230 8780 42273
rect 8712 42217 8780 42230
rect 8836 42217 8904 42273
rect 8960 42217 9028 42273
rect 9084 42217 9124 42273
rect 8616 42174 9124 42217
rect 8616 42149 8677 42174
rect 8729 42149 9124 42174
rect 8616 42093 8656 42149
rect 8729 42122 8780 42149
rect 8712 42093 8780 42122
rect 8836 42093 8904 42149
rect 8960 42093 9028 42149
rect 9084 42093 9124 42149
rect 8616 42066 9124 42093
rect 8616 42025 8677 42066
rect 8729 42025 9124 42066
rect 8616 41969 8656 42025
rect 8729 42014 8780 42025
rect 8712 41969 8780 42014
rect 8836 41969 8904 42025
rect 8960 41969 9028 42025
rect 9084 41969 9124 42025
rect 8616 41958 9124 41969
rect 8616 41906 8677 41958
rect 8729 41906 9124 41958
rect 8616 41901 9124 41906
rect 8616 41845 8656 41901
rect 8712 41850 8780 41901
rect 8729 41845 8780 41850
rect 8836 41845 8904 41901
rect 8960 41845 9028 41901
rect 9084 41845 9124 41901
rect 8616 41798 8677 41845
rect 8729 41798 9124 41845
rect 8616 41777 9124 41798
rect 8616 41721 8656 41777
rect 8712 41742 8780 41777
rect 8729 41721 8780 41742
rect 8836 41721 8904 41777
rect 8960 41721 9028 41777
rect 9084 41721 9124 41777
rect 8616 41690 8677 41721
rect 8729 41690 9124 41721
rect 8616 41653 9124 41690
rect 8616 41597 8656 41653
rect 8712 41634 8780 41653
rect 8729 41597 8780 41634
rect 8836 41597 8904 41653
rect 8960 41597 9028 41653
rect 9084 41597 9124 41653
rect 8616 41582 8677 41597
rect 8729 41582 9124 41597
rect 8616 41529 9124 41582
rect 8616 41473 8656 41529
rect 8712 41526 8780 41529
rect 8729 41474 8780 41526
rect 8712 41473 8780 41474
rect 8836 41473 8904 41529
rect 8960 41473 9028 41529
rect 9084 41473 9124 41529
rect 8616 41418 9124 41473
rect 8616 41405 8677 41418
rect 8729 41405 9124 41418
rect 8616 41349 8656 41405
rect 8729 41366 8780 41405
rect 8712 41349 8780 41366
rect 8836 41349 8904 41405
rect 8960 41349 9028 41405
rect 9084 41349 9124 41405
rect 8616 41045 9124 41349
rect 8616 40989 8656 41045
rect 8712 40989 8780 41045
rect 8836 40989 8904 41045
rect 8960 40989 9028 41045
rect 9084 40989 9124 41045
rect 8616 40921 9124 40989
rect 8616 40865 8656 40921
rect 8712 40865 8780 40921
rect 8836 40865 8904 40921
rect 8960 40865 9028 40921
rect 9084 40865 9124 40921
rect 8616 40797 9124 40865
rect 8616 40741 8656 40797
rect 8712 40741 8780 40797
rect 8836 40741 8904 40797
rect 8960 40741 9028 40797
rect 9084 40741 9124 40797
rect 8616 40673 9124 40741
rect 8616 40617 8656 40673
rect 8712 40617 8780 40673
rect 8836 40617 8904 40673
rect 8960 40617 9028 40673
rect 9084 40617 9124 40673
rect 8616 40549 9124 40617
rect 8616 40493 8656 40549
rect 8712 40494 8780 40549
rect 8729 40493 8780 40494
rect 8836 40493 8904 40549
rect 8960 40493 9028 40549
rect 9084 40493 9124 40549
rect 8616 40442 8677 40493
rect 8729 40442 9124 40493
rect 8616 40425 9124 40442
rect 8616 40369 8656 40425
rect 8712 40386 8780 40425
rect 8729 40369 8780 40386
rect 8836 40369 8904 40425
rect 8960 40369 9028 40425
rect 9084 40369 9124 40425
rect 8616 40334 8677 40369
rect 8729 40334 9124 40369
rect 8616 40301 9124 40334
rect 8616 40245 8656 40301
rect 8712 40278 8780 40301
rect 8729 40245 8780 40278
rect 8836 40245 8904 40301
rect 8960 40245 9028 40301
rect 9084 40245 9124 40301
rect 8616 40226 8677 40245
rect 8729 40226 9124 40245
rect 8616 40177 9124 40226
rect 8616 40121 8656 40177
rect 8712 40170 8780 40177
rect 8729 40121 8780 40170
rect 8836 40121 8904 40177
rect 8960 40121 9028 40177
rect 9084 40121 9124 40177
rect 8616 40118 8677 40121
rect 8729 40118 9124 40121
rect 8616 40062 9124 40118
rect 8616 40053 8677 40062
rect 8729 40053 9124 40062
rect 8616 39997 8656 40053
rect 8729 40010 8780 40053
rect 8712 39997 8780 40010
rect 8836 39997 8904 40053
rect 8960 39997 9028 40053
rect 9084 39997 9124 40053
rect 8616 39954 9124 39997
rect 8616 39929 8677 39954
rect 8729 39929 9124 39954
rect 8616 39873 8656 39929
rect 8729 39902 8780 39929
rect 8712 39873 8780 39902
rect 8836 39873 8904 39929
rect 8960 39873 9028 39929
rect 9084 39873 9124 39929
rect 8616 39846 9124 39873
rect 8616 39805 8677 39846
rect 8729 39805 9124 39846
rect 8616 39749 8656 39805
rect 8729 39794 8780 39805
rect 8712 39749 8780 39794
rect 8836 39749 8904 39805
rect 8960 39749 9028 39805
rect 9084 39749 9124 39805
rect 8616 39738 9124 39749
rect 8616 39686 8677 39738
rect 8729 39686 9124 39738
rect 8616 39630 9124 39686
rect 8616 39578 8677 39630
rect 8729 39578 9124 39630
rect 8616 39522 9124 39578
rect 8616 39470 8677 39522
rect 8729 39470 9124 39522
rect 8616 39414 9124 39470
rect 8616 39362 8677 39414
rect 8729 39362 9124 39414
rect 8616 39306 9124 39362
rect 8616 39254 8677 39306
rect 8729 39254 9124 39306
rect 8616 39198 9124 39254
rect 8616 39146 8677 39198
rect 8729 39146 9124 39198
rect 8616 39090 9124 39146
rect 8616 39038 8677 39090
rect 8729 39038 9124 39090
rect 8616 38982 9124 39038
rect 8616 38930 8677 38982
rect 8729 38930 9124 38982
rect 8616 38874 9124 38930
rect 8616 38822 8677 38874
rect 8729 38822 9124 38874
rect 8616 38766 9124 38822
rect 8616 38714 8677 38766
rect 8729 38714 9124 38766
rect 8616 38658 9124 38714
rect 8616 38606 8677 38658
rect 8729 38606 9124 38658
rect 8616 38550 9124 38606
rect 8616 38498 8677 38550
rect 8729 38498 9124 38550
rect 8616 38442 9124 38498
rect 8616 38390 8677 38442
rect 8729 38390 9124 38442
rect 8616 38334 9124 38390
rect 8616 38282 8677 38334
rect 8729 38282 9124 38334
rect 8616 38226 9124 38282
rect 8616 38174 8677 38226
rect 8729 38174 9124 38226
rect 8616 38118 9124 38174
rect 8616 38066 8677 38118
rect 8729 38066 9124 38118
rect 8616 38010 9124 38066
rect 8616 37958 8677 38010
rect 8729 37958 9124 38010
rect 8616 37902 9124 37958
rect 8616 37850 8677 37902
rect 8729 37850 9124 37902
rect 8616 37794 9124 37850
rect 8616 37742 8677 37794
rect 8729 37742 9124 37794
rect 8616 37686 9124 37742
rect 8616 37634 8677 37686
rect 8729 37634 9124 37686
rect 8616 37578 9124 37634
rect 8616 37526 8677 37578
rect 8729 37526 9124 37578
rect 8616 37470 9124 37526
rect 8616 37418 8677 37470
rect 8729 37418 9124 37470
rect 8616 36546 9124 37418
rect 8616 36494 8677 36546
rect 8729 36494 9124 36546
rect 8616 36438 9124 36494
rect 8616 36386 8677 36438
rect 8729 36386 9124 36438
rect 8616 36330 9124 36386
rect 8616 36278 8677 36330
rect 8729 36278 9124 36330
rect 8616 36222 9124 36278
rect 8616 36170 8677 36222
rect 8729 36170 9124 36222
rect 8616 36114 9124 36170
rect 8616 36062 8677 36114
rect 8729 36062 9124 36114
rect 8616 36006 9124 36062
rect 8616 35954 8677 36006
rect 8729 35954 9124 36006
rect 8616 35898 9124 35954
rect 8616 35846 8677 35898
rect 8729 35846 9124 35898
rect 8616 35790 9124 35846
rect 8616 35738 8677 35790
rect 8729 35738 9124 35790
rect 8616 35682 9124 35738
rect 8616 35630 8677 35682
rect 8729 35630 9124 35682
rect 8616 35574 9124 35630
rect 8616 35522 8677 35574
rect 8729 35522 9124 35574
rect 8616 35466 9124 35522
rect 8616 35414 8677 35466
rect 8729 35414 9124 35466
rect 8616 35358 9124 35414
rect 8616 35306 8677 35358
rect 8729 35306 9124 35358
rect 8616 35250 9124 35306
rect 8616 35198 8677 35250
rect 8729 35198 9124 35250
rect 8616 35142 9124 35198
rect 8616 35090 8677 35142
rect 8729 35090 9124 35142
rect 8616 35034 9124 35090
rect 8616 34982 8677 35034
rect 8729 34982 9124 35034
rect 8616 34926 9124 34982
rect 8616 34874 8677 34926
rect 8729 34874 9124 34926
rect 8616 34818 9124 34874
rect 8616 34766 8677 34818
rect 8729 34766 9124 34818
rect 8616 34710 9124 34766
rect 8616 34658 8677 34710
rect 8729 34658 9124 34710
rect 8616 34602 9124 34658
rect 8616 34550 8677 34602
rect 8729 34550 9124 34602
rect 8616 34494 9124 34550
rect 8616 34442 8677 34494
rect 8729 34442 9124 34494
rect 8616 34386 9124 34442
rect 8616 34334 8677 34386
rect 8729 34334 9124 34386
rect 8616 34278 9124 34334
rect 8616 34226 8677 34278
rect 8729 34226 9124 34278
rect 8616 34170 9124 34226
rect 8616 34118 8677 34170
rect 8729 34118 9124 34170
rect 8616 34062 9124 34118
rect 8616 34010 8677 34062
rect 8729 34010 9124 34062
rect 8616 33954 9124 34010
rect 8616 33902 8677 33954
rect 8729 33902 9124 33954
rect 8616 33846 9124 33902
rect 8616 33794 8677 33846
rect 8729 33794 9124 33846
rect 8616 33738 9124 33794
rect 8616 33686 8677 33738
rect 8729 33686 9124 33738
rect 8616 33630 9124 33686
rect 8616 33578 8677 33630
rect 8729 33578 9124 33630
rect 8616 33522 9124 33578
rect 8616 33470 8677 33522
rect 8729 33470 9124 33522
rect 8616 33051 9124 33470
rect 8616 32995 8656 33051
rect 8712 32995 8780 33051
rect 8836 32995 8904 33051
rect 8960 32995 9028 33051
rect 9084 32995 9124 33051
rect 8616 32927 9124 32995
rect 8616 32871 8656 32927
rect 8712 32871 8780 32927
rect 8836 32871 8904 32927
rect 8960 32871 9028 32927
rect 9084 32871 9124 32927
rect 8616 32803 9124 32871
rect 8616 32747 8656 32803
rect 8712 32747 8780 32803
rect 8836 32747 8904 32803
rect 8960 32747 9028 32803
rect 9084 32747 9124 32803
rect 8616 32679 9124 32747
rect 8616 32623 8656 32679
rect 8712 32623 8780 32679
rect 8836 32623 8904 32679
rect 8960 32623 9028 32679
rect 9084 32623 9124 32679
rect 8616 32598 9124 32623
rect 8616 32555 8677 32598
rect 8729 32555 9124 32598
rect 8616 32499 8656 32555
rect 8729 32546 8780 32555
rect 8712 32499 8780 32546
rect 8836 32499 8904 32555
rect 8960 32499 9028 32555
rect 9084 32499 9124 32555
rect 8616 32490 9124 32499
rect 8616 32438 8677 32490
rect 8729 32438 9124 32490
rect 8616 32431 9124 32438
rect 8616 32375 8656 32431
rect 8712 32382 8780 32431
rect 8729 32375 8780 32382
rect 8836 32375 8904 32431
rect 8960 32375 9028 32431
rect 9084 32375 9124 32431
rect 8616 32330 8677 32375
rect 8729 32330 9124 32375
rect 8616 32307 9124 32330
rect 8616 32251 8656 32307
rect 8712 32274 8780 32307
rect 8729 32251 8780 32274
rect 8836 32251 8904 32307
rect 8960 32251 9028 32307
rect 9084 32251 9124 32307
rect 8616 32222 8677 32251
rect 8729 32222 9124 32251
rect 8616 32183 9124 32222
rect 8616 32127 8656 32183
rect 8712 32166 8780 32183
rect 8729 32127 8780 32166
rect 8836 32127 8904 32183
rect 8960 32127 9028 32183
rect 9084 32127 9124 32183
rect 8616 32114 8677 32127
rect 8729 32114 9124 32127
rect 8616 32059 9124 32114
rect 8616 32003 8656 32059
rect 8712 32058 8780 32059
rect 8729 32006 8780 32058
rect 8712 32003 8780 32006
rect 8836 32003 8904 32059
rect 8960 32003 9028 32059
rect 9084 32003 9124 32059
rect 8616 31950 9124 32003
rect 8616 31935 8677 31950
rect 8729 31935 9124 31950
rect 8616 31879 8656 31935
rect 8729 31898 8780 31935
rect 8712 31879 8780 31898
rect 8836 31879 8904 31935
rect 8960 31879 9028 31935
rect 9084 31879 9124 31935
rect 8616 31842 9124 31879
rect 8616 31811 8677 31842
rect 8729 31811 9124 31842
rect 8616 31755 8656 31811
rect 8729 31790 8780 31811
rect 8712 31755 8780 31790
rect 8836 31755 8904 31811
rect 8960 31755 9028 31811
rect 9084 31755 9124 31811
rect 8616 31734 9124 31755
rect 8616 31687 8677 31734
rect 8729 31687 9124 31734
rect 8616 31631 8656 31687
rect 8729 31682 8780 31687
rect 8712 31631 8780 31682
rect 8836 31631 8904 31687
rect 8960 31631 9028 31687
rect 9084 31631 9124 31687
rect 8616 31626 9124 31631
rect 8616 31574 8677 31626
rect 8729 31574 9124 31626
rect 8616 31563 9124 31574
rect 8616 31507 8656 31563
rect 8712 31518 8780 31563
rect 8729 31507 8780 31518
rect 8836 31507 8904 31563
rect 8960 31507 9028 31563
rect 9084 31507 9124 31563
rect 8616 31466 8677 31507
rect 8729 31466 9124 31507
rect 8616 31439 9124 31466
rect 8616 31383 8656 31439
rect 8712 31410 8780 31439
rect 8729 31383 8780 31410
rect 8836 31383 8904 31439
rect 8960 31383 9028 31439
rect 9084 31383 9124 31439
rect 8616 31358 8677 31383
rect 8729 31358 9124 31383
rect 8616 31315 9124 31358
rect 8616 31259 8656 31315
rect 8712 31302 8780 31315
rect 8729 31259 8780 31302
rect 8836 31259 8904 31315
rect 8960 31259 9028 31315
rect 9084 31259 9124 31315
rect 8616 31250 8677 31259
rect 8729 31250 9124 31259
rect 8616 31194 9124 31250
rect 8616 31191 8677 31194
rect 8729 31191 9124 31194
rect 8616 31135 8656 31191
rect 8729 31142 8780 31191
rect 8712 31135 8780 31142
rect 8836 31135 8904 31191
rect 8960 31135 9028 31191
rect 9084 31135 9124 31191
rect 8616 31086 9124 31135
rect 8616 31067 8677 31086
rect 8729 31067 9124 31086
rect 8616 31011 8656 31067
rect 8729 31034 8780 31067
rect 8712 31011 8780 31034
rect 8836 31011 8904 31067
rect 8960 31011 9028 31067
rect 9084 31011 9124 31067
rect 8616 30978 9124 31011
rect 8616 30943 8677 30978
rect 8729 30943 9124 30978
rect 8616 30887 8656 30943
rect 8729 30926 8780 30943
rect 8712 30887 8780 30926
rect 8836 30887 8904 30943
rect 8960 30887 9028 30943
rect 9084 30887 9124 30943
rect 8616 30870 9124 30887
rect 8616 30819 8677 30870
rect 8729 30819 9124 30870
rect 8616 30763 8656 30819
rect 8729 30818 8780 30819
rect 8712 30763 8780 30818
rect 8836 30763 8904 30819
rect 8960 30763 9028 30819
rect 9084 30763 9124 30819
rect 8616 30762 9124 30763
rect 8616 30710 8677 30762
rect 8729 30710 9124 30762
rect 8616 30695 9124 30710
rect 8616 30639 8656 30695
rect 8712 30654 8780 30695
rect 8729 30639 8780 30654
rect 8836 30639 8904 30695
rect 8960 30639 9028 30695
rect 9084 30639 9124 30695
rect 8616 30602 8677 30639
rect 8729 30602 9124 30639
rect 8616 30571 9124 30602
rect 8616 30515 8656 30571
rect 8712 30546 8780 30571
rect 8729 30515 8780 30546
rect 8836 30515 8904 30571
rect 8960 30515 9028 30571
rect 9084 30515 9124 30571
rect 8616 30494 8677 30515
rect 8729 30494 9124 30515
rect 8616 30447 9124 30494
rect 8616 30391 8656 30447
rect 8712 30438 8780 30447
rect 8729 30391 8780 30438
rect 8836 30391 8904 30447
rect 8960 30391 9028 30447
rect 9084 30391 9124 30447
rect 8616 30386 8677 30391
rect 8729 30386 9124 30391
rect 8616 30330 9124 30386
rect 8616 30323 8677 30330
rect 8729 30323 9124 30330
rect 8616 30267 8656 30323
rect 8729 30278 8780 30323
rect 8712 30267 8780 30278
rect 8836 30267 8904 30323
rect 8960 30267 9028 30323
rect 9084 30267 9124 30323
rect 8616 30222 9124 30267
rect 8616 30199 8677 30222
rect 8729 30199 9124 30222
rect 8616 30143 8656 30199
rect 8729 30170 8780 30199
rect 8712 30143 8780 30170
rect 8836 30143 8904 30199
rect 8960 30143 9028 30199
rect 9084 30143 9124 30199
rect 8616 30114 9124 30143
rect 8616 30062 8677 30114
rect 8729 30062 9124 30114
rect 8616 30006 9124 30062
rect 8616 29954 8677 30006
rect 8729 29954 9124 30006
rect 8616 29898 9124 29954
rect 8616 29846 8677 29898
rect 8729 29846 9124 29898
rect 8616 29845 9124 29846
rect 8616 29789 8656 29845
rect 8712 29790 8780 29845
rect 8729 29789 8780 29790
rect 8836 29789 8904 29845
rect 8960 29789 9028 29845
rect 9084 29789 9124 29845
rect 8616 29738 8677 29789
rect 8729 29738 9124 29789
rect 8616 29721 9124 29738
rect 8616 29665 8656 29721
rect 8712 29682 8780 29721
rect 8729 29665 8780 29682
rect 8836 29665 8904 29721
rect 8960 29665 9028 29721
rect 9084 29665 9124 29721
rect 8616 29630 8677 29665
rect 8729 29630 9124 29665
rect 8616 29597 9124 29630
rect 8616 29541 8656 29597
rect 8712 29574 8780 29597
rect 8729 29541 8780 29574
rect 8836 29541 8904 29597
rect 8960 29541 9028 29597
rect 9084 29541 9124 29597
rect 8616 29522 8677 29541
rect 8729 29522 9124 29541
rect 8616 29473 9124 29522
rect 8616 29417 8656 29473
rect 8712 29417 8780 29473
rect 8836 29417 8904 29473
rect 8960 29417 9028 29473
rect 9084 29417 9124 29473
rect 8616 29349 9124 29417
rect 8616 29293 8656 29349
rect 8712 29293 8780 29349
rect 8836 29293 8904 29349
rect 8960 29293 9028 29349
rect 9084 29293 9124 29349
rect 8616 29225 9124 29293
rect 8616 29169 8656 29225
rect 8712 29169 8780 29225
rect 8836 29169 8904 29225
rect 8960 29169 9028 29225
rect 9084 29169 9124 29225
rect 8616 29101 9124 29169
rect 8616 29045 8656 29101
rect 8712 29045 8780 29101
rect 8836 29045 8904 29101
rect 8960 29045 9028 29101
rect 9084 29045 9124 29101
rect 8616 28977 9124 29045
rect 8616 28921 8656 28977
rect 8712 28921 8780 28977
rect 8836 28921 8904 28977
rect 8960 28921 9028 28977
rect 9084 28921 9124 28977
rect 8616 28853 9124 28921
rect 8616 28797 8656 28853
rect 8712 28797 8780 28853
rect 8836 28797 8904 28853
rect 8960 28797 9028 28853
rect 9084 28797 9124 28853
rect 8616 28729 9124 28797
rect 8616 28673 8656 28729
rect 8712 28673 8780 28729
rect 8836 28673 8904 28729
rect 8960 28673 9028 28729
rect 9084 28673 9124 28729
rect 8616 28650 9124 28673
rect 8616 28605 8677 28650
rect 8729 28605 9124 28650
rect 8616 28549 8656 28605
rect 8729 28598 8780 28605
rect 8712 28549 8780 28598
rect 8836 28549 8904 28605
rect 8960 28549 9028 28605
rect 9084 28549 9124 28605
rect 8616 28542 9124 28549
rect 8616 28490 8677 28542
rect 8729 28490 9124 28542
rect 8616 28434 9124 28490
rect 8616 28382 8677 28434
rect 8729 28382 9124 28434
rect 8616 28326 9124 28382
rect 8616 28274 8677 28326
rect 8729 28274 9124 28326
rect 8616 28218 9124 28274
rect 8616 28166 8677 28218
rect 8729 28166 9124 28218
rect 8616 28110 9124 28166
rect 8616 28058 8677 28110
rect 8729 28058 9124 28110
rect 8616 28002 9124 28058
rect 8616 27950 8677 28002
rect 8729 27950 9124 28002
rect 8616 27894 9124 27950
rect 8616 27842 8677 27894
rect 8729 27842 9124 27894
rect 8616 27786 9124 27842
rect 8616 27734 8677 27786
rect 8729 27734 9124 27786
rect 8616 27678 9124 27734
rect 8616 27626 8677 27678
rect 8729 27626 9124 27678
rect 8616 27570 9124 27626
rect 8616 27518 8677 27570
rect 8729 27518 9124 27570
rect 8616 27462 9124 27518
rect 8616 27410 8677 27462
rect 8729 27410 9124 27462
rect 8616 27354 9124 27410
rect 8616 27302 8677 27354
rect 8729 27302 9124 27354
rect 8616 27246 9124 27302
rect 8616 27194 8677 27246
rect 8729 27194 9124 27246
rect 8616 27138 9124 27194
rect 8616 27086 8677 27138
rect 8729 27086 9124 27138
rect 8616 27030 9124 27086
rect 8616 26978 8677 27030
rect 8729 26978 9124 27030
rect 8616 26922 9124 26978
rect 8616 26870 8677 26922
rect 8729 26870 9124 26922
rect 8616 26814 9124 26870
rect 8616 26762 8677 26814
rect 8729 26762 9124 26814
rect 8616 26706 9124 26762
rect 8616 26654 8677 26706
rect 8729 26654 9124 26706
rect 8616 26651 9124 26654
rect 8616 26595 8656 26651
rect 8712 26598 8780 26651
rect 8729 26595 8780 26598
rect 8836 26595 8904 26651
rect 8960 26595 9028 26651
rect 9084 26595 9124 26651
rect 8616 26546 8677 26595
rect 8729 26546 9124 26595
rect 8616 26527 9124 26546
rect 8616 26471 8656 26527
rect 8712 26490 8780 26527
rect 8729 26471 8780 26490
rect 8836 26471 8904 26527
rect 8960 26471 9028 26527
rect 9084 26471 9124 26527
rect 8616 26438 8677 26471
rect 8729 26438 9124 26471
rect 8616 26403 9124 26438
rect 8616 26347 8656 26403
rect 8712 26382 8780 26403
rect 8729 26347 8780 26382
rect 8836 26347 8904 26403
rect 8960 26347 9028 26403
rect 9084 26347 9124 26403
rect 8616 26330 8677 26347
rect 8729 26330 9124 26347
rect 8616 26279 9124 26330
rect 8616 26223 8656 26279
rect 8712 26274 8780 26279
rect 8729 26223 8780 26274
rect 8836 26223 8904 26279
rect 8960 26223 9028 26279
rect 9084 26223 9124 26279
rect 8616 26222 8677 26223
rect 8729 26222 9124 26223
rect 8616 26166 9124 26222
rect 8616 26155 8677 26166
rect 8729 26155 9124 26166
rect 8616 26099 8656 26155
rect 8729 26114 8780 26155
rect 8712 26099 8780 26114
rect 8836 26099 8904 26155
rect 8960 26099 9028 26155
rect 9084 26099 9124 26155
rect 8616 26058 9124 26099
rect 8616 26031 8677 26058
rect 8729 26031 9124 26058
rect 8616 25975 8656 26031
rect 8729 26006 8780 26031
rect 8712 25975 8780 26006
rect 8836 25975 8904 26031
rect 8960 25975 9028 26031
rect 9084 25975 9124 26031
rect 8616 25950 9124 25975
rect 8616 25907 8677 25950
rect 8729 25907 9124 25950
rect 8616 25851 8656 25907
rect 8729 25898 8780 25907
rect 8712 25851 8780 25898
rect 8836 25851 8904 25907
rect 8960 25851 9028 25907
rect 9084 25851 9124 25907
rect 8616 25842 9124 25851
rect 8616 25790 8677 25842
rect 8729 25790 9124 25842
rect 8616 25783 9124 25790
rect 8616 25727 8656 25783
rect 8712 25734 8780 25783
rect 8729 25727 8780 25734
rect 8836 25727 8904 25783
rect 8960 25727 9028 25783
rect 9084 25727 9124 25783
rect 8616 25682 8677 25727
rect 8729 25682 9124 25727
rect 8616 25659 9124 25682
rect 8616 25603 8656 25659
rect 8712 25626 8780 25659
rect 8729 25603 8780 25626
rect 8836 25603 8904 25659
rect 8960 25603 9028 25659
rect 9084 25603 9124 25659
rect 8616 25574 8677 25603
rect 8729 25574 9124 25603
rect 8616 25535 9124 25574
rect 8616 25479 8656 25535
rect 8712 25479 8780 25535
rect 8836 25479 8904 25535
rect 8960 25479 9028 25535
rect 9084 25479 9124 25535
rect 8616 25411 9124 25479
rect 8616 25355 8656 25411
rect 8712 25355 8780 25411
rect 8836 25355 8904 25411
rect 8960 25355 9028 25411
rect 9084 25355 9124 25411
rect 8616 25287 9124 25355
rect 8616 25231 8656 25287
rect 8712 25231 8780 25287
rect 8836 25231 8904 25287
rect 8960 25231 9028 25287
rect 9084 25231 9124 25287
rect 8616 25163 9124 25231
rect 8616 25107 8656 25163
rect 8712 25107 8780 25163
rect 8836 25107 8904 25163
rect 8960 25107 9028 25163
rect 9084 25107 9124 25163
rect 8616 25039 9124 25107
rect 8616 24983 8656 25039
rect 8712 24983 8780 25039
rect 8836 24983 8904 25039
rect 8960 24983 9028 25039
rect 9084 24983 9124 25039
rect 8616 24915 9124 24983
rect 8616 24859 8656 24915
rect 8712 24859 8780 24915
rect 8836 24859 8904 24915
rect 8960 24859 9028 24915
rect 9084 24859 9124 24915
rect 8616 24791 9124 24859
rect 8616 24735 8656 24791
rect 8712 24735 8780 24791
rect 8836 24735 8904 24791
rect 8960 24735 9028 24791
rect 9084 24735 9124 24791
rect 8616 24702 9124 24735
rect 8616 24667 8677 24702
rect 8729 24667 9124 24702
rect 8616 24611 8656 24667
rect 8729 24650 8780 24667
rect 8712 24611 8780 24650
rect 8836 24611 8904 24667
rect 8960 24611 9028 24667
rect 9084 24611 9124 24667
rect 8616 24594 9124 24611
rect 8616 24543 8677 24594
rect 8729 24543 9124 24594
rect 8616 24487 8656 24543
rect 8729 24542 8780 24543
rect 8712 24487 8780 24542
rect 8836 24487 8904 24543
rect 8960 24487 9028 24543
rect 9084 24487 9124 24543
rect 8616 24486 9124 24487
rect 8616 24434 8677 24486
rect 8729 24434 9124 24486
rect 8616 24419 9124 24434
rect 8616 24363 8656 24419
rect 8712 24378 8780 24419
rect 8729 24363 8780 24378
rect 8836 24363 8904 24419
rect 8960 24363 9028 24419
rect 9084 24363 9124 24419
rect 8616 24326 8677 24363
rect 8729 24326 9124 24363
rect 8616 24295 9124 24326
rect 8616 24239 8656 24295
rect 8712 24270 8780 24295
rect 8729 24239 8780 24270
rect 8836 24239 8904 24295
rect 8960 24239 9028 24295
rect 9084 24239 9124 24295
rect 8616 24218 8677 24239
rect 8729 24218 9124 24239
rect 8616 24171 9124 24218
rect 8616 24115 8656 24171
rect 8712 24162 8780 24171
rect 8729 24115 8780 24162
rect 8836 24115 8904 24171
rect 8960 24115 9028 24171
rect 9084 24115 9124 24171
rect 8616 24110 8677 24115
rect 8729 24110 9124 24115
rect 8616 24054 9124 24110
rect 8616 24047 8677 24054
rect 8729 24047 9124 24054
rect 8616 23991 8656 24047
rect 8729 24002 8780 24047
rect 8712 23991 8780 24002
rect 8836 23991 8904 24047
rect 8960 23991 9028 24047
rect 9084 23991 9124 24047
rect 8616 23946 9124 23991
rect 8616 23923 8677 23946
rect 8729 23923 9124 23946
rect 8616 23867 8656 23923
rect 8729 23894 8780 23923
rect 8712 23867 8780 23894
rect 8836 23867 8904 23923
rect 8960 23867 9028 23923
rect 9084 23867 9124 23923
rect 8616 23838 9124 23867
rect 8616 23799 8677 23838
rect 8729 23799 9124 23838
rect 8616 23743 8656 23799
rect 8729 23786 8780 23799
rect 8712 23743 8780 23786
rect 8836 23743 8904 23799
rect 8960 23743 9028 23799
rect 9084 23743 9124 23799
rect 8616 23730 9124 23743
rect 8616 23678 8677 23730
rect 8729 23678 9124 23730
rect 8616 23622 9124 23678
rect 8616 23570 8677 23622
rect 8729 23570 9124 23622
rect 8616 23514 9124 23570
rect 8616 23462 8677 23514
rect 8729 23462 9124 23514
rect 8616 23451 9124 23462
rect 8616 23395 8656 23451
rect 8712 23406 8780 23451
rect 8729 23395 8780 23406
rect 8836 23395 8904 23451
rect 8960 23395 9028 23451
rect 9084 23395 9124 23451
rect 8616 23354 8677 23395
rect 8729 23354 9124 23395
rect 8616 23327 9124 23354
rect 8616 23271 8656 23327
rect 8712 23298 8780 23327
rect 8729 23271 8780 23298
rect 8836 23271 8904 23327
rect 8960 23271 9028 23327
rect 9084 23271 9124 23327
rect 8616 23246 8677 23271
rect 8729 23246 9124 23271
rect 8616 23203 9124 23246
rect 8616 23147 8656 23203
rect 8712 23190 8780 23203
rect 8729 23147 8780 23190
rect 8836 23147 8904 23203
rect 8960 23147 9028 23203
rect 9084 23147 9124 23203
rect 8616 23138 8677 23147
rect 8729 23138 9124 23147
rect 8616 23082 9124 23138
rect 8616 23079 8677 23082
rect 8729 23079 9124 23082
rect 8616 23023 8656 23079
rect 8729 23030 8780 23079
rect 8712 23023 8780 23030
rect 8836 23023 8904 23079
rect 8960 23023 9028 23079
rect 9084 23023 9124 23079
rect 8616 22974 9124 23023
rect 8616 22955 8677 22974
rect 8729 22955 9124 22974
rect 8616 22899 8656 22955
rect 8729 22922 8780 22955
rect 8712 22899 8780 22922
rect 8836 22899 8904 22955
rect 8960 22899 9028 22955
rect 9084 22899 9124 22955
rect 8616 22866 9124 22899
rect 8616 22831 8677 22866
rect 8729 22831 9124 22866
rect 8616 22775 8656 22831
rect 8729 22814 8780 22831
rect 8712 22775 8780 22814
rect 8836 22775 8904 22831
rect 8960 22775 9028 22831
rect 9084 22775 9124 22831
rect 8616 22758 9124 22775
rect 8616 22707 8677 22758
rect 8729 22707 9124 22758
rect 8616 22651 8656 22707
rect 8729 22706 8780 22707
rect 8712 22651 8780 22706
rect 8836 22651 8904 22707
rect 8960 22651 9028 22707
rect 9084 22651 9124 22707
rect 8616 22650 9124 22651
rect 8616 22598 8677 22650
rect 8729 22598 9124 22650
rect 8616 22583 9124 22598
rect 8616 22527 8656 22583
rect 8712 22542 8780 22583
rect 8729 22527 8780 22542
rect 8836 22527 8904 22583
rect 8960 22527 9028 22583
rect 9084 22527 9124 22583
rect 8616 22490 8677 22527
rect 8729 22490 9124 22527
rect 8616 22459 9124 22490
rect 8616 22403 8656 22459
rect 8712 22434 8780 22459
rect 8729 22403 8780 22434
rect 8836 22403 8904 22459
rect 8960 22403 9028 22459
rect 9084 22403 9124 22459
rect 8616 22382 8677 22403
rect 8729 22382 9124 22403
rect 8616 22335 9124 22382
rect 8616 22279 8656 22335
rect 8712 22326 8780 22335
rect 8729 22279 8780 22326
rect 8836 22279 8904 22335
rect 8960 22279 9028 22335
rect 9084 22279 9124 22335
rect 8616 22274 8677 22279
rect 8729 22274 9124 22279
rect 8616 22218 9124 22274
rect 8616 22211 8677 22218
rect 8729 22211 9124 22218
rect 8616 22155 8656 22211
rect 8729 22166 8780 22211
rect 8712 22155 8780 22166
rect 8836 22155 8904 22211
rect 8960 22155 9028 22211
rect 9084 22155 9124 22211
rect 8616 22110 9124 22155
rect 8616 22087 8677 22110
rect 8729 22087 9124 22110
rect 8616 22031 8656 22087
rect 8729 22058 8780 22087
rect 8712 22031 8780 22058
rect 8836 22031 8904 22087
rect 8960 22031 9028 22087
rect 9084 22031 9124 22087
rect 8616 22002 9124 22031
rect 8616 21963 8677 22002
rect 8729 21963 9124 22002
rect 8616 21907 8656 21963
rect 8729 21950 8780 21963
rect 8712 21907 8780 21950
rect 8836 21907 8904 21963
rect 8960 21907 9028 21963
rect 9084 21907 9124 21963
rect 8616 21894 9124 21907
rect 8616 21842 8677 21894
rect 8729 21842 9124 21894
rect 8616 21839 9124 21842
rect 8616 21783 8656 21839
rect 8712 21786 8780 21839
rect 8729 21783 8780 21786
rect 8836 21783 8904 21839
rect 8960 21783 9028 21839
rect 9084 21783 9124 21839
rect 8616 21734 8677 21783
rect 8729 21734 9124 21783
rect 8616 21715 9124 21734
rect 8616 21659 8656 21715
rect 8712 21678 8780 21715
rect 8729 21659 8780 21678
rect 8836 21659 8904 21715
rect 8960 21659 9028 21715
rect 9084 21659 9124 21715
rect 8616 21626 8677 21659
rect 8729 21626 9124 21659
rect 8616 21591 9124 21626
rect 8616 21535 8656 21591
rect 8712 21535 8780 21591
rect 8836 21535 8904 21591
rect 8960 21535 9028 21591
rect 9084 21535 9124 21591
rect 8616 21467 9124 21535
rect 8616 21411 8656 21467
rect 8712 21411 8780 21467
rect 8836 21411 8904 21467
rect 8960 21411 9028 21467
rect 9084 21411 9124 21467
rect 8616 21343 9124 21411
rect 8616 21287 8656 21343
rect 8712 21287 8780 21343
rect 8836 21287 8904 21343
rect 8960 21287 9028 21343
rect 9084 21287 9124 21343
rect 8616 21219 9124 21287
rect 8616 21163 8656 21219
rect 8712 21163 8780 21219
rect 8836 21163 8904 21219
rect 8960 21163 9028 21219
rect 9084 21163 9124 21219
rect 8616 21095 9124 21163
rect 8616 21039 8656 21095
rect 8712 21039 8780 21095
rect 8836 21039 8904 21095
rect 8960 21039 9028 21095
rect 9084 21039 9124 21095
rect 8616 20971 9124 21039
rect 8616 20915 8656 20971
rect 8712 20915 8780 20971
rect 8836 20915 8904 20971
rect 8960 20915 9028 20971
rect 9084 20915 9124 20971
rect 8616 20847 9124 20915
rect 8616 20791 8656 20847
rect 8712 20791 8780 20847
rect 8836 20791 8904 20847
rect 8960 20791 9028 20847
rect 9084 20791 9124 20847
rect 8616 20723 9124 20791
rect 8616 20667 8656 20723
rect 8712 20667 8780 20723
rect 8836 20667 8904 20723
rect 8960 20667 9028 20723
rect 9084 20667 9124 20723
rect 8616 20599 9124 20667
rect 8616 20577 8656 20599
rect 8712 20577 8780 20599
rect 8836 20577 8904 20599
rect 8960 20577 9028 20599
rect 9084 20577 9124 20599
rect 8616 20525 8628 20577
rect 8712 20543 8736 20577
rect 8836 20543 8844 20577
rect 8680 20525 8736 20543
rect 8788 20525 8844 20543
rect 8896 20543 8904 20577
rect 9004 20543 9028 20577
rect 8896 20525 8952 20543
rect 9004 20525 9060 20543
rect 9112 20525 9124 20577
rect 8616 20469 9124 20525
rect 8616 20417 8628 20469
rect 8680 20417 8736 20469
rect 8788 20417 8844 20469
rect 8896 20417 8952 20469
rect 9004 20417 9060 20469
rect 9112 20417 9124 20469
rect 8616 20361 9124 20417
rect 8616 20309 8628 20361
rect 8680 20309 8736 20361
rect 8788 20309 8844 20361
rect 8896 20309 8952 20361
rect 9004 20309 9060 20361
rect 9112 20309 9124 20361
rect 8616 20251 9124 20309
rect 8616 20195 8656 20251
rect 8712 20195 8780 20251
rect 8836 20195 8904 20251
rect 8960 20195 9028 20251
rect 9084 20195 9124 20251
rect 8616 20127 9124 20195
rect 8616 20071 8656 20127
rect 8712 20071 8780 20127
rect 8836 20071 8904 20127
rect 8960 20071 9028 20127
rect 9084 20071 9124 20127
rect 8616 20003 9124 20071
rect 8616 19947 8656 20003
rect 8712 19947 8780 20003
rect 8836 19947 8904 20003
rect 8960 19947 9028 20003
rect 9084 19947 9124 20003
rect 8616 19879 9124 19947
rect 8616 19823 8656 19879
rect 8712 19823 8780 19879
rect 8836 19823 8904 19879
rect 8960 19823 9028 19879
rect 9084 19823 9124 19879
rect 8616 19755 9124 19823
rect 8616 19699 8656 19755
rect 8712 19699 8780 19755
rect 8836 19699 8904 19755
rect 8960 19699 9028 19755
rect 9084 19699 9124 19755
rect 8616 19631 9124 19699
rect 8616 19584 8656 19631
rect 8712 19584 8780 19631
rect 8836 19584 8904 19631
rect 8960 19584 9028 19631
rect 9084 19584 9124 19631
rect 8616 19532 8628 19584
rect 8712 19575 8736 19584
rect 8836 19575 8844 19584
rect 8680 19532 8736 19575
rect 8788 19532 8844 19575
rect 8896 19575 8904 19584
rect 9004 19575 9028 19584
rect 8896 19532 8952 19575
rect 9004 19532 9060 19575
rect 9112 19532 9124 19584
rect 8616 19507 9124 19532
rect 8616 19476 8656 19507
rect 8712 19476 8780 19507
rect 8836 19476 8904 19507
rect 8960 19476 9028 19507
rect 9084 19476 9124 19507
rect 8616 19424 8628 19476
rect 8712 19451 8736 19476
rect 8836 19451 8844 19476
rect 8680 19424 8736 19451
rect 8788 19424 8844 19451
rect 8896 19451 8904 19476
rect 9004 19451 9028 19476
rect 8896 19424 8952 19451
rect 9004 19424 9060 19451
rect 9112 19424 9124 19476
rect 8616 19383 9124 19424
rect 8616 19327 8656 19383
rect 8712 19327 8780 19383
rect 8836 19327 8904 19383
rect 8960 19327 9028 19383
rect 9084 19327 9124 19383
rect 8616 19259 9124 19327
rect 8616 19203 8656 19259
rect 8712 19203 8780 19259
rect 8836 19203 8904 19259
rect 8960 19203 9028 19259
rect 9084 19203 9124 19259
rect 8616 19135 9124 19203
rect 8616 19079 8656 19135
rect 8712 19079 8780 19135
rect 8836 19079 8904 19135
rect 8960 19079 9028 19135
rect 9084 19079 9124 19135
rect 8616 19011 9124 19079
rect 8616 18955 8656 19011
rect 8712 18955 8780 19011
rect 8836 18955 8904 19011
rect 8960 18955 9028 19011
rect 9084 18955 9124 19011
rect 8616 18887 9124 18955
rect 8616 18831 8656 18887
rect 8712 18831 8780 18887
rect 8836 18831 8904 18887
rect 8960 18831 9028 18887
rect 9084 18831 9124 18887
rect 8616 18763 9124 18831
rect 8616 18712 8656 18763
rect 8712 18712 8780 18763
rect 8836 18712 8904 18763
rect 8960 18712 9028 18763
rect 9084 18712 9124 18763
rect 8616 18660 8628 18712
rect 8712 18707 8736 18712
rect 8836 18707 8844 18712
rect 8680 18660 8736 18707
rect 8788 18660 8844 18707
rect 8896 18707 8904 18712
rect 9004 18707 9028 18712
rect 8896 18660 8952 18707
rect 9004 18660 9060 18707
rect 9112 18660 9124 18712
rect 8616 18639 9124 18660
rect 8616 18604 8656 18639
rect 8712 18604 8780 18639
rect 8836 18604 8904 18639
rect 8960 18604 9028 18639
rect 9084 18604 9124 18639
rect 8616 18552 8628 18604
rect 8712 18583 8736 18604
rect 8836 18583 8844 18604
rect 8680 18552 8736 18583
rect 8788 18552 8844 18583
rect 8896 18583 8904 18604
rect 9004 18583 9028 18604
rect 8896 18552 8952 18583
rect 9004 18552 9060 18583
rect 9112 18552 9124 18604
rect 8616 18515 9124 18552
rect 8616 18459 8656 18515
rect 8712 18459 8780 18515
rect 8836 18459 8904 18515
rect 8960 18459 9028 18515
rect 9084 18459 9124 18515
rect 8616 18391 9124 18459
rect 8616 18335 8656 18391
rect 8712 18335 8780 18391
rect 8836 18335 8904 18391
rect 8960 18335 9028 18391
rect 9084 18335 9124 18391
rect 8616 18267 9124 18335
rect 8616 18211 8656 18267
rect 8712 18211 8780 18267
rect 8836 18211 8904 18267
rect 8960 18211 9028 18267
rect 9084 18211 9124 18267
rect 8616 18143 9124 18211
rect 8616 18087 8656 18143
rect 8712 18087 8780 18143
rect 8836 18087 8904 18143
rect 8960 18087 9028 18143
rect 9084 18087 9124 18143
rect 8616 18019 9124 18087
rect 8616 17963 8656 18019
rect 8712 17963 8780 18019
rect 8836 17963 8904 18019
rect 8960 17963 9028 18019
rect 9084 17963 9124 18019
rect 8616 17895 9124 17963
rect 8616 17840 8656 17895
rect 8712 17840 8780 17895
rect 8836 17840 8904 17895
rect 8960 17840 9028 17895
rect 9084 17840 9124 17895
rect 8616 17788 8628 17840
rect 8712 17839 8736 17840
rect 8836 17839 8844 17840
rect 8680 17788 8736 17839
rect 8788 17788 8844 17839
rect 8896 17839 8904 17840
rect 9004 17839 9028 17840
rect 8896 17788 8952 17839
rect 9004 17788 9060 17839
rect 9112 17788 9124 17840
rect 8616 17771 9124 17788
rect 8616 17732 8656 17771
rect 8712 17732 8780 17771
rect 8836 17732 8904 17771
rect 8960 17732 9028 17771
rect 9084 17732 9124 17771
rect 8616 17680 8628 17732
rect 8712 17715 8736 17732
rect 8836 17715 8844 17732
rect 8680 17680 8736 17715
rect 8788 17680 8844 17715
rect 8896 17715 8904 17732
rect 9004 17715 9028 17732
rect 8896 17680 8952 17715
rect 9004 17680 9060 17715
rect 9112 17680 9124 17732
rect 8616 17647 9124 17680
rect 8616 17591 8656 17647
rect 8712 17591 8780 17647
rect 8836 17591 8904 17647
rect 8960 17591 9028 17647
rect 9084 17591 9124 17647
rect 8616 17523 9124 17591
rect 8616 17467 8656 17523
rect 8712 17467 8780 17523
rect 8836 17467 8904 17523
rect 8960 17467 9028 17523
rect 9084 17467 9124 17523
rect 8616 17399 9124 17467
rect 8616 17343 8656 17399
rect 8712 17343 8780 17399
rect 8836 17343 8904 17399
rect 8960 17343 9028 17399
rect 9084 17343 9124 17399
rect 8616 17051 9124 17343
rect 8616 16995 8656 17051
rect 8712 16995 8780 17051
rect 8836 16995 8904 17051
rect 8960 16995 9028 17051
rect 9084 16995 9124 17051
rect 8616 16968 9124 16995
rect 8616 16916 8628 16968
rect 8680 16927 8736 16968
rect 8788 16927 8844 16968
rect 8712 16916 8736 16927
rect 8836 16916 8844 16927
rect 8896 16927 8952 16968
rect 9004 16927 9060 16968
rect 8896 16916 8904 16927
rect 9004 16916 9028 16927
rect 9112 16916 9124 16968
rect 8616 16871 8656 16916
rect 8712 16871 8780 16916
rect 8836 16871 8904 16916
rect 8960 16871 9028 16916
rect 9084 16871 9124 16916
rect 8616 16860 9124 16871
rect 8616 16808 8628 16860
rect 8680 16808 8736 16860
rect 8788 16808 8844 16860
rect 8896 16808 8952 16860
rect 9004 16808 9060 16860
rect 9112 16808 9124 16860
rect 8616 16803 9124 16808
rect 8616 16747 8656 16803
rect 8712 16747 8780 16803
rect 8836 16747 8904 16803
rect 8960 16747 9028 16803
rect 9084 16747 9124 16803
rect 8616 16679 9124 16747
rect 8616 16623 8656 16679
rect 8712 16623 8780 16679
rect 8836 16623 8904 16679
rect 8960 16623 9028 16679
rect 9084 16623 9124 16679
rect 8616 16555 9124 16623
rect 8616 16499 8656 16555
rect 8712 16499 8780 16555
rect 8836 16499 8904 16555
rect 8960 16499 9028 16555
rect 9084 16499 9124 16555
rect 8616 16431 9124 16499
rect 8616 16375 8656 16431
rect 8712 16375 8780 16431
rect 8836 16375 8904 16431
rect 8960 16375 9028 16431
rect 9084 16375 9124 16431
rect 8616 16307 9124 16375
rect 8616 16251 8656 16307
rect 8712 16251 8780 16307
rect 8836 16251 8904 16307
rect 8960 16251 9028 16307
rect 9084 16251 9124 16307
rect 8616 16183 9124 16251
rect 8616 16127 8656 16183
rect 8712 16127 8780 16183
rect 8836 16127 8904 16183
rect 8960 16127 9028 16183
rect 9084 16127 9124 16183
rect 8616 16083 9124 16127
rect 8616 16031 8628 16083
rect 8680 16059 8736 16083
rect 8788 16059 8844 16083
rect 8712 16031 8736 16059
rect 8836 16031 8844 16059
rect 8896 16059 8952 16083
rect 9004 16059 9060 16083
rect 8896 16031 8904 16059
rect 9004 16031 9028 16059
rect 9112 16031 9124 16083
rect 8616 16003 8656 16031
rect 8712 16003 8780 16031
rect 8836 16003 8904 16031
rect 8960 16003 9028 16031
rect 9084 16003 9124 16031
rect 8616 15975 9124 16003
rect 8616 15923 8628 15975
rect 8680 15935 8736 15975
rect 8788 15935 8844 15975
rect 8712 15923 8736 15935
rect 8836 15923 8844 15935
rect 8896 15935 8952 15975
rect 9004 15935 9060 15975
rect 8896 15923 8904 15935
rect 9004 15923 9028 15935
rect 9112 15923 9124 15975
rect 8616 15879 8656 15923
rect 8712 15879 8780 15923
rect 8836 15879 8904 15923
rect 8960 15879 9028 15923
rect 9084 15879 9124 15923
rect 8616 15867 9124 15879
rect 8616 15815 8628 15867
rect 8680 15815 8736 15867
rect 8788 15815 8844 15867
rect 8896 15815 8952 15867
rect 9004 15815 9060 15867
rect 9112 15815 9124 15867
rect 8616 15811 9124 15815
rect 8616 15762 8656 15811
rect 6408 15755 6418 15762
rect 5970 15687 6418 15755
rect 5970 15631 5980 15687
rect 6036 15631 6104 15687
rect 6160 15631 6228 15687
rect 6284 15631 6352 15687
rect 6408 15631 6418 15687
rect 5970 15563 6418 15631
rect 5970 15507 5980 15563
rect 6036 15507 6104 15563
rect 6160 15507 6228 15563
rect 6284 15507 6352 15563
rect 6408 15507 6418 15563
rect 5970 15439 6418 15507
rect 5970 15383 5980 15439
rect 6036 15383 6104 15439
rect 6160 15383 6228 15439
rect 6284 15383 6352 15439
rect 6408 15383 6418 15439
rect 5970 15315 6418 15383
rect 5970 15259 5980 15315
rect 6036 15259 6104 15315
rect 6160 15259 6228 15315
rect 6284 15259 6352 15315
rect 6408 15259 6418 15315
rect 5970 15191 6418 15259
rect 5970 15135 5980 15191
rect 6036 15135 6104 15191
rect 6160 15135 6228 15191
rect 6284 15135 6352 15191
rect 6408 15135 6418 15191
rect 5970 15067 6418 15135
rect 5970 15011 5980 15067
rect 6036 15011 6104 15067
rect 6160 15011 6228 15067
rect 6284 15011 6352 15067
rect 6408 15011 6418 15067
rect 5970 14943 6418 15011
rect 5970 14887 5980 14943
rect 6036 14887 6104 14943
rect 6160 14887 6228 14943
rect 6284 14887 6352 14943
rect 6408 14887 6418 14943
rect 5970 14819 6418 14887
rect 5970 14763 5980 14819
rect 6036 14763 6104 14819
rect 6160 14763 6228 14819
rect 6284 14763 6352 14819
rect 6408 14763 6418 14819
rect 5970 14695 6418 14763
rect 5970 14639 5980 14695
rect 6036 14639 6104 14695
rect 6160 14639 6228 14695
rect 6284 14639 6352 14695
rect 6408 14639 6418 14695
rect 5970 14571 6418 14639
rect 5970 14515 5980 14571
rect 6036 14515 6104 14571
rect 6160 14515 6228 14571
rect 6284 14515 6352 14571
rect 6408 14515 6418 14571
rect 5970 14447 6418 14515
rect 5970 14391 5980 14447
rect 6036 14391 6104 14447
rect 6160 14391 6228 14447
rect 6284 14391 6352 14447
rect 6408 14391 6418 14447
rect 5970 14323 6418 14391
rect 5970 14267 5980 14323
rect 6036 14267 6104 14323
rect 6160 14267 6228 14323
rect 6284 14267 6352 14323
rect 6408 14267 6418 14323
rect 5970 14199 6418 14267
rect 5970 14143 5980 14199
rect 6036 14143 6104 14199
rect 6160 14143 6228 14199
rect 6284 14143 6352 14199
rect 6408 14143 6418 14199
rect 5970 14133 6418 14143
rect 8646 15755 8656 15762
rect 8712 15755 8780 15811
rect 8836 15755 8904 15811
rect 8960 15755 9028 15811
rect 9084 15762 9124 15811
rect 9752 56922 10260 56975
rect 9752 56866 9792 56922
rect 9848 56866 9916 56922
rect 9972 56866 10040 56922
rect 10096 56866 10164 56922
rect 10220 56866 10260 56922
rect 9752 56798 10260 56866
rect 9752 56742 9792 56798
rect 9848 56742 9916 56798
rect 9972 56742 10040 56798
rect 10096 56742 10164 56798
rect 10220 56742 10260 56798
rect 9752 56711 10260 56742
rect 9752 56659 9764 56711
rect 9816 56674 9872 56711
rect 9924 56674 9980 56711
rect 9848 56659 9872 56674
rect 9972 56659 9980 56674
rect 10032 56674 10088 56711
rect 10140 56674 10196 56711
rect 10032 56659 10040 56674
rect 10140 56659 10164 56674
rect 10248 56659 10260 56711
rect 9752 56618 9792 56659
rect 9848 56618 9916 56659
rect 9972 56618 10040 56659
rect 10096 56618 10164 56659
rect 10220 56618 10260 56659
rect 9752 56603 10260 56618
rect 9752 56551 9764 56603
rect 9816 56551 9872 56603
rect 9924 56551 9980 56603
rect 10032 56551 10088 56603
rect 10140 56551 10196 56603
rect 10248 56551 10260 56603
rect 9752 56550 10260 56551
rect 9752 56495 9792 56550
rect 9848 56495 9916 56550
rect 9972 56495 10040 56550
rect 10096 56495 10164 56550
rect 10220 56495 10260 56550
rect 9752 56443 9764 56495
rect 9848 56494 9872 56495
rect 9972 56494 9980 56495
rect 9816 56443 9872 56494
rect 9924 56443 9980 56494
rect 10032 56494 10040 56495
rect 10140 56494 10164 56495
rect 10032 56443 10088 56494
rect 10140 56443 10196 56494
rect 10248 56443 10260 56495
rect 9752 56426 10260 56443
rect 9752 56370 9792 56426
rect 9848 56370 9916 56426
rect 9972 56370 10040 56426
rect 10096 56370 10164 56426
rect 10220 56370 10260 56426
rect 9752 56302 10260 56370
rect 9752 56246 9792 56302
rect 9848 56246 9916 56302
rect 9972 56246 10040 56302
rect 10096 56246 10164 56302
rect 10220 56246 10260 56302
rect 9752 56178 10260 56246
rect 9752 56122 9792 56178
rect 9848 56122 9916 56178
rect 9972 56122 10040 56178
rect 10096 56122 10164 56178
rect 10220 56122 10260 56178
rect 9752 56054 10260 56122
rect 9752 55998 9792 56054
rect 9848 55998 9916 56054
rect 9972 55998 10040 56054
rect 10096 55998 10164 56054
rect 10220 55998 10260 56054
rect 9752 55930 10260 55998
rect 9752 55874 9792 55930
rect 9848 55874 9916 55930
rect 9972 55874 10040 55930
rect 10096 55874 10164 55930
rect 10220 55874 10260 55930
rect 9752 55806 10260 55874
rect 9752 55750 9792 55806
rect 9848 55750 9916 55806
rect 9972 55750 10040 55806
rect 10096 55750 10164 55806
rect 10220 55750 10260 55806
rect 9752 53845 10260 55750
rect 9752 53789 9792 53845
rect 9848 53789 9916 53845
rect 9972 53789 10040 53845
rect 10096 53789 10164 53845
rect 10220 53789 10260 53845
rect 9752 53721 10260 53789
rect 9752 53665 9792 53721
rect 9848 53665 9916 53721
rect 9972 53665 10040 53721
rect 10096 53665 10164 53721
rect 10220 53665 10260 53721
rect 9752 53597 10260 53665
rect 9752 53541 9792 53597
rect 9848 53541 9916 53597
rect 9972 53541 10040 53597
rect 10096 53541 10164 53597
rect 10220 53541 10260 53597
rect 9752 53473 10260 53541
rect 9752 53417 9792 53473
rect 9848 53417 9916 53473
rect 9972 53417 10040 53473
rect 10096 53417 10164 53473
rect 10220 53417 10260 53473
rect 9752 53349 10260 53417
rect 9752 53293 9792 53349
rect 9848 53293 9916 53349
rect 9972 53293 10040 53349
rect 10096 53293 10164 53349
rect 10220 53293 10260 53349
rect 9752 53225 10260 53293
rect 9752 53169 9792 53225
rect 9848 53169 9916 53225
rect 9972 53169 10040 53225
rect 10096 53169 10164 53225
rect 10220 53169 10260 53225
rect 9752 53101 10260 53169
rect 9752 53045 9792 53101
rect 9848 53045 9916 53101
rect 9972 53045 10040 53101
rect 10096 53045 10164 53101
rect 10220 53045 10260 53101
rect 9752 52996 9794 53045
rect 9846 52996 9918 53045
rect 9970 52996 10042 53045
rect 10094 52996 10166 53045
rect 10218 52996 10260 53045
rect 9752 52977 10260 52996
rect 9752 52921 9792 52977
rect 9848 52921 9916 52977
rect 9972 52921 10040 52977
rect 10096 52921 10164 52977
rect 10220 52921 10260 52977
rect 9752 52872 9794 52921
rect 9846 52872 9918 52921
rect 9970 52872 10042 52921
rect 10094 52872 10166 52921
rect 10218 52872 10260 52921
rect 9752 52853 10260 52872
rect 9752 52797 9792 52853
rect 9848 52797 9916 52853
rect 9972 52797 10040 52853
rect 10096 52797 10164 52853
rect 10220 52797 10260 52853
rect 9752 52748 9794 52797
rect 9846 52748 9918 52797
rect 9970 52748 10042 52797
rect 10094 52748 10166 52797
rect 10218 52748 10260 52797
rect 9752 52729 10260 52748
rect 9752 52673 9792 52729
rect 9848 52673 9916 52729
rect 9972 52673 10040 52729
rect 10096 52673 10164 52729
rect 10220 52673 10260 52729
rect 9752 52624 9794 52673
rect 9846 52624 9918 52673
rect 9970 52624 10042 52673
rect 10094 52624 10166 52673
rect 10218 52624 10260 52673
rect 9752 52605 10260 52624
rect 9752 52549 9792 52605
rect 9848 52549 9916 52605
rect 9972 52549 10040 52605
rect 10096 52549 10164 52605
rect 10220 52549 10260 52605
rect 9752 52500 9794 52549
rect 9846 52500 9918 52549
rect 9970 52500 10042 52549
rect 10094 52500 10166 52549
rect 10218 52500 10260 52549
rect 9752 49100 10260 52500
rect 9752 49048 9794 49100
rect 9846 49048 9918 49100
rect 9970 49048 10042 49100
rect 10094 49048 10166 49100
rect 10218 49048 10260 49100
rect 9752 49045 10260 49048
rect 9752 48989 9792 49045
rect 9848 48989 9916 49045
rect 9972 48989 10040 49045
rect 10096 48989 10164 49045
rect 10220 48989 10260 49045
rect 9752 48976 10260 48989
rect 9752 48924 9794 48976
rect 9846 48924 9918 48976
rect 9970 48924 10042 48976
rect 10094 48924 10166 48976
rect 10218 48924 10260 48976
rect 9752 48921 10260 48924
rect 9752 48865 9792 48921
rect 9848 48865 9916 48921
rect 9972 48865 10040 48921
rect 10096 48865 10164 48921
rect 10220 48865 10260 48921
rect 9752 48852 10260 48865
rect 9752 48800 9794 48852
rect 9846 48800 9918 48852
rect 9970 48800 10042 48852
rect 10094 48800 10166 48852
rect 10218 48800 10260 48852
rect 9752 48797 10260 48800
rect 9752 48741 9792 48797
rect 9848 48741 9916 48797
rect 9972 48741 10040 48797
rect 10096 48741 10164 48797
rect 10220 48741 10260 48797
rect 9752 48728 10260 48741
rect 9752 48676 9794 48728
rect 9846 48676 9918 48728
rect 9970 48676 10042 48728
rect 10094 48676 10166 48728
rect 10218 48676 10260 48728
rect 9752 48673 10260 48676
rect 9752 48617 9792 48673
rect 9848 48617 9916 48673
rect 9972 48617 10040 48673
rect 10096 48617 10164 48673
rect 10220 48617 10260 48673
rect 9752 48604 10260 48617
rect 9752 48552 9794 48604
rect 9846 48552 9918 48604
rect 9970 48552 10042 48604
rect 10094 48552 10166 48604
rect 10218 48552 10260 48604
rect 9752 48549 10260 48552
rect 9752 48493 9792 48549
rect 9848 48493 9916 48549
rect 9972 48493 10040 48549
rect 10096 48493 10164 48549
rect 10220 48493 10260 48549
rect 9752 48425 10260 48493
rect 9752 48369 9792 48425
rect 9848 48369 9916 48425
rect 9972 48369 10040 48425
rect 10096 48369 10164 48425
rect 10220 48369 10260 48425
rect 9752 48301 10260 48369
rect 9752 48245 9792 48301
rect 9848 48245 9916 48301
rect 9972 48245 10040 48301
rect 10096 48245 10164 48301
rect 10220 48245 10260 48301
rect 9752 48177 10260 48245
rect 9752 48121 9792 48177
rect 9848 48121 9916 48177
rect 9972 48121 10040 48177
rect 10096 48121 10164 48177
rect 10220 48121 10260 48177
rect 9752 48053 10260 48121
rect 9752 47997 9792 48053
rect 9848 47997 9916 48053
rect 9972 47997 10040 48053
rect 10096 47997 10164 48053
rect 10220 47997 10260 48053
rect 9752 47929 10260 47997
rect 9752 47873 9792 47929
rect 9848 47873 9916 47929
rect 9972 47873 10040 47929
rect 10096 47873 10164 47929
rect 10220 47873 10260 47929
rect 9752 47805 10260 47873
rect 9752 47749 9792 47805
rect 9848 47749 9916 47805
rect 9972 47749 10040 47805
rect 10096 47749 10164 47805
rect 10220 47749 10260 47805
rect 9752 45845 10260 47749
rect 9752 45789 9792 45845
rect 9848 45789 9916 45845
rect 9972 45789 10040 45845
rect 10096 45789 10164 45845
rect 10220 45789 10260 45845
rect 9752 45721 10260 45789
rect 9752 45665 9792 45721
rect 9848 45665 9916 45721
rect 9972 45665 10040 45721
rect 10096 45665 10164 45721
rect 10220 45665 10260 45721
rect 9752 45597 10260 45665
rect 9752 45541 9792 45597
rect 9848 45541 9916 45597
rect 9972 45541 10040 45597
rect 10096 45541 10164 45597
rect 10220 45541 10260 45597
rect 9752 45473 10260 45541
rect 9752 45417 9792 45473
rect 9848 45417 9916 45473
rect 9972 45417 10040 45473
rect 10096 45417 10164 45473
rect 10220 45417 10260 45473
rect 9752 45349 10260 45417
rect 9752 45293 9792 45349
rect 9848 45293 9916 45349
rect 9972 45293 10040 45349
rect 10096 45293 10164 45349
rect 10220 45293 10260 45349
rect 9752 45225 10260 45293
rect 9752 45169 9792 45225
rect 9848 45169 9916 45225
rect 9972 45169 10040 45225
rect 10096 45169 10164 45225
rect 10220 45169 10260 45225
rect 9752 45152 10260 45169
rect 9752 45101 9794 45152
rect 9846 45101 9918 45152
rect 9970 45101 10042 45152
rect 10094 45101 10166 45152
rect 10218 45101 10260 45152
rect 9752 45045 9792 45101
rect 9848 45045 9916 45101
rect 9972 45045 10040 45101
rect 10096 45045 10164 45101
rect 10220 45045 10260 45101
rect 9752 45028 10260 45045
rect 9752 44977 9794 45028
rect 9846 44977 9918 45028
rect 9970 44977 10042 45028
rect 10094 44977 10166 45028
rect 10218 44977 10260 45028
rect 9752 44921 9792 44977
rect 9848 44921 9916 44977
rect 9972 44921 10040 44977
rect 10096 44921 10164 44977
rect 10220 44921 10260 44977
rect 9752 44904 10260 44921
rect 9752 44853 9794 44904
rect 9846 44853 9918 44904
rect 9970 44853 10042 44904
rect 10094 44853 10166 44904
rect 10218 44853 10260 44904
rect 9752 44797 9792 44853
rect 9848 44797 9916 44853
rect 9972 44797 10040 44853
rect 10096 44797 10164 44853
rect 10220 44797 10260 44853
rect 9752 44780 10260 44797
rect 9752 44729 9794 44780
rect 9846 44729 9918 44780
rect 9970 44729 10042 44780
rect 10094 44729 10166 44780
rect 10218 44729 10260 44780
rect 9752 44673 9792 44729
rect 9848 44673 9916 44729
rect 9972 44673 10040 44729
rect 10096 44673 10164 44729
rect 10220 44673 10260 44729
rect 9752 44656 10260 44673
rect 9752 44605 9794 44656
rect 9846 44605 9918 44656
rect 9970 44605 10042 44656
rect 10094 44605 10166 44656
rect 10218 44605 10260 44656
rect 9752 44549 9792 44605
rect 9848 44549 9916 44605
rect 9972 44549 10040 44605
rect 10096 44549 10164 44605
rect 10220 44549 10260 44605
rect 9752 41204 10260 44549
rect 9752 41152 9794 41204
rect 9846 41152 9918 41204
rect 9970 41152 10042 41204
rect 10094 41152 10166 41204
rect 10218 41152 10260 41204
rect 9752 41080 10260 41152
rect 9752 41028 9794 41080
rect 9846 41028 9918 41080
rect 9970 41028 10042 41080
rect 10094 41028 10166 41080
rect 10218 41028 10260 41080
rect 9752 40956 10260 41028
rect 9752 40904 9794 40956
rect 9846 40904 9918 40956
rect 9970 40904 10042 40956
rect 10094 40904 10166 40956
rect 10218 40904 10260 40956
rect 9752 40832 10260 40904
rect 9752 40780 9794 40832
rect 9846 40780 9918 40832
rect 9970 40780 10042 40832
rect 10094 40780 10166 40832
rect 10218 40780 10260 40832
rect 9752 40708 10260 40780
rect 9752 40656 9794 40708
rect 9846 40656 9918 40708
rect 9970 40656 10042 40708
rect 10094 40656 10166 40708
rect 10218 40656 10260 40708
rect 9752 37256 10260 40656
rect 9752 37204 9794 37256
rect 9846 37204 9918 37256
rect 9970 37204 10042 37256
rect 10094 37204 10166 37256
rect 10218 37204 10260 37256
rect 9752 37132 10260 37204
rect 9752 37080 9794 37132
rect 9846 37080 9918 37132
rect 9970 37080 10042 37132
rect 10094 37080 10166 37132
rect 10218 37080 10260 37132
rect 9752 37008 10260 37080
rect 9752 36956 9794 37008
rect 9846 36956 9918 37008
rect 9970 36956 10042 37008
rect 10094 36956 10166 37008
rect 10218 36956 10260 37008
rect 9752 36884 10260 36956
rect 9752 36832 9794 36884
rect 9846 36832 9918 36884
rect 9970 36832 10042 36884
rect 10094 36832 10166 36884
rect 10218 36832 10260 36884
rect 9752 36760 10260 36832
rect 9752 36708 9794 36760
rect 9846 36708 9918 36760
rect 9970 36708 10042 36760
rect 10094 36708 10166 36760
rect 10218 36708 10260 36760
rect 9752 36251 10260 36708
rect 9752 36195 9792 36251
rect 9848 36195 9916 36251
rect 9972 36195 10040 36251
rect 10096 36195 10164 36251
rect 10220 36195 10260 36251
rect 9752 36127 10260 36195
rect 9752 36071 9792 36127
rect 9848 36071 9916 36127
rect 9972 36071 10040 36127
rect 10096 36071 10164 36127
rect 10220 36071 10260 36127
rect 9752 36003 10260 36071
rect 9752 35947 9792 36003
rect 9848 35947 9916 36003
rect 9972 35947 10040 36003
rect 10096 35947 10164 36003
rect 10220 35947 10260 36003
rect 9752 35879 10260 35947
rect 9752 35823 9792 35879
rect 9848 35823 9916 35879
rect 9972 35823 10040 35879
rect 10096 35823 10164 35879
rect 10220 35823 10260 35879
rect 9752 35755 10260 35823
rect 9752 35699 9792 35755
rect 9848 35699 9916 35755
rect 9972 35699 10040 35755
rect 10096 35699 10164 35755
rect 10220 35699 10260 35755
rect 9752 35631 10260 35699
rect 9752 35575 9792 35631
rect 9848 35575 9916 35631
rect 9972 35575 10040 35631
rect 10096 35575 10164 35631
rect 10220 35575 10260 35631
rect 9752 35507 10260 35575
rect 9752 35451 9792 35507
rect 9848 35451 9916 35507
rect 9972 35451 10040 35507
rect 10096 35451 10164 35507
rect 10220 35451 10260 35507
rect 9752 35383 10260 35451
rect 9752 35327 9792 35383
rect 9848 35327 9916 35383
rect 9972 35327 10040 35383
rect 10096 35327 10164 35383
rect 10220 35327 10260 35383
rect 9752 35259 10260 35327
rect 9752 35203 9792 35259
rect 9848 35203 9916 35259
rect 9972 35203 10040 35259
rect 10096 35203 10164 35259
rect 10220 35203 10260 35259
rect 9752 35135 10260 35203
rect 9752 35079 9792 35135
rect 9848 35079 9916 35135
rect 9972 35079 10040 35135
rect 10096 35079 10164 35135
rect 10220 35079 10260 35135
rect 9752 35011 10260 35079
rect 9752 34955 9792 35011
rect 9848 34955 9916 35011
rect 9972 34955 10040 35011
rect 10096 34955 10164 35011
rect 10220 34955 10260 35011
rect 9752 34887 10260 34955
rect 9752 34831 9792 34887
rect 9848 34831 9916 34887
rect 9972 34831 10040 34887
rect 10096 34831 10164 34887
rect 10220 34831 10260 34887
rect 9752 34763 10260 34831
rect 9752 34707 9792 34763
rect 9848 34707 9916 34763
rect 9972 34707 10040 34763
rect 10096 34707 10164 34763
rect 10220 34707 10260 34763
rect 9752 34639 10260 34707
rect 9752 34583 9792 34639
rect 9848 34583 9916 34639
rect 9972 34583 10040 34639
rect 10096 34583 10164 34639
rect 10220 34583 10260 34639
rect 9752 34515 10260 34583
rect 9752 34459 9792 34515
rect 9848 34459 9916 34515
rect 9972 34459 10040 34515
rect 10096 34459 10164 34515
rect 10220 34459 10260 34515
rect 9752 34391 10260 34459
rect 9752 34335 9792 34391
rect 9848 34335 9916 34391
rect 9972 34335 10040 34391
rect 10096 34335 10164 34391
rect 10220 34335 10260 34391
rect 9752 34267 10260 34335
rect 9752 34211 9792 34267
rect 9848 34211 9916 34267
rect 9972 34211 10040 34267
rect 10096 34211 10164 34267
rect 10220 34211 10260 34267
rect 9752 34143 10260 34211
rect 9752 34087 9792 34143
rect 9848 34087 9916 34143
rect 9972 34087 10040 34143
rect 10096 34087 10164 34143
rect 10220 34087 10260 34143
rect 9752 34019 10260 34087
rect 9752 33963 9792 34019
rect 9848 33963 9916 34019
rect 9972 33963 10040 34019
rect 10096 33963 10164 34019
rect 10220 33963 10260 34019
rect 9752 33895 10260 33963
rect 9752 33839 9792 33895
rect 9848 33839 9916 33895
rect 9972 33839 10040 33895
rect 10096 33839 10164 33895
rect 10220 33839 10260 33895
rect 9752 33771 10260 33839
rect 9752 33715 9792 33771
rect 9848 33715 9916 33771
rect 9972 33715 10040 33771
rect 10096 33715 10164 33771
rect 10220 33715 10260 33771
rect 9752 33647 10260 33715
rect 9752 33591 9792 33647
rect 9848 33591 9916 33647
rect 9972 33591 10040 33647
rect 10096 33591 10164 33647
rect 10220 33591 10260 33647
rect 9752 33523 10260 33591
rect 9752 33467 9792 33523
rect 9848 33467 9916 33523
rect 9972 33467 10040 33523
rect 10096 33467 10164 33523
rect 10220 33467 10260 33523
rect 9752 33399 10260 33467
rect 9752 33343 9792 33399
rect 9848 33343 9916 33399
rect 9972 33343 10040 33399
rect 10096 33343 10164 33399
rect 10220 33343 10260 33399
rect 9752 33308 10260 33343
rect 9752 33256 9794 33308
rect 9846 33256 9918 33308
rect 9970 33256 10042 33308
rect 10094 33256 10166 33308
rect 10218 33256 10260 33308
rect 9752 33184 10260 33256
rect 9752 33132 9794 33184
rect 9846 33132 9918 33184
rect 9970 33132 10042 33184
rect 10094 33132 10166 33184
rect 10218 33132 10260 33184
rect 9752 33060 10260 33132
rect 9752 33008 9794 33060
rect 9846 33008 9918 33060
rect 9970 33008 10042 33060
rect 10094 33008 10166 33060
rect 10218 33008 10260 33060
rect 9752 32936 10260 33008
rect 9752 32884 9794 32936
rect 9846 32884 9918 32936
rect 9970 32884 10042 32936
rect 10094 32884 10166 32936
rect 10218 32884 10260 32936
rect 9752 32812 10260 32884
rect 9752 32760 9794 32812
rect 9846 32760 9918 32812
rect 9970 32760 10042 32812
rect 10094 32760 10166 32812
rect 10218 32760 10260 32812
rect 9752 29360 10260 32760
rect 9752 29308 9794 29360
rect 9846 29308 9918 29360
rect 9970 29308 10042 29360
rect 10094 29308 10166 29360
rect 10218 29308 10260 29360
rect 9752 29236 10260 29308
rect 9752 29184 9794 29236
rect 9846 29184 9918 29236
rect 9970 29184 10042 29236
rect 10094 29184 10166 29236
rect 10218 29184 10260 29236
rect 9752 29112 10260 29184
rect 9752 29060 9794 29112
rect 9846 29060 9918 29112
rect 9970 29060 10042 29112
rect 10094 29060 10166 29112
rect 10218 29060 10260 29112
rect 9752 28988 10260 29060
rect 9752 28936 9794 28988
rect 9846 28936 9918 28988
rect 9970 28936 10042 28988
rect 10094 28936 10166 28988
rect 10218 28936 10260 28988
rect 9752 28864 10260 28936
rect 9752 28812 9794 28864
rect 9846 28812 9918 28864
rect 9970 28812 10042 28864
rect 10094 28812 10166 28864
rect 10218 28812 10260 28864
rect 9752 28245 10260 28812
rect 9752 28189 9792 28245
rect 9848 28189 9916 28245
rect 9972 28189 10040 28245
rect 10096 28189 10164 28245
rect 10220 28189 10260 28245
rect 9752 28121 10260 28189
rect 9752 28065 9792 28121
rect 9848 28065 9916 28121
rect 9972 28065 10040 28121
rect 10096 28065 10164 28121
rect 10220 28065 10260 28121
rect 9752 27997 10260 28065
rect 9752 27941 9792 27997
rect 9848 27941 9916 27997
rect 9972 27941 10040 27997
rect 10096 27941 10164 27997
rect 10220 27941 10260 27997
rect 9752 27873 10260 27941
rect 9752 27817 9792 27873
rect 9848 27817 9916 27873
rect 9972 27817 10040 27873
rect 10096 27817 10164 27873
rect 10220 27817 10260 27873
rect 9752 27749 10260 27817
rect 9752 27693 9792 27749
rect 9848 27693 9916 27749
rect 9972 27693 10040 27749
rect 10096 27693 10164 27749
rect 10220 27693 10260 27749
rect 9752 27625 10260 27693
rect 9752 27569 9792 27625
rect 9848 27569 9916 27625
rect 9972 27569 10040 27625
rect 10096 27569 10164 27625
rect 10220 27569 10260 27625
rect 9752 27501 10260 27569
rect 9752 27445 9792 27501
rect 9848 27445 9916 27501
rect 9972 27445 10040 27501
rect 10096 27445 10164 27501
rect 10220 27445 10260 27501
rect 9752 27377 10260 27445
rect 9752 27321 9792 27377
rect 9848 27321 9916 27377
rect 9972 27321 10040 27377
rect 10096 27321 10164 27377
rect 10220 27321 10260 27377
rect 9752 27253 10260 27321
rect 9752 27197 9792 27253
rect 9848 27197 9916 27253
rect 9972 27197 10040 27253
rect 10096 27197 10164 27253
rect 10220 27197 10260 27253
rect 9752 27129 10260 27197
rect 9752 27073 9792 27129
rect 9848 27073 9916 27129
rect 9972 27073 10040 27129
rect 10096 27073 10164 27129
rect 10220 27073 10260 27129
rect 9752 27005 10260 27073
rect 9752 26949 9792 27005
rect 9848 26949 9916 27005
rect 9972 26949 10040 27005
rect 10096 26949 10164 27005
rect 10220 26949 10260 27005
rect 9752 25412 10260 26949
rect 9752 25360 9794 25412
rect 9846 25360 9918 25412
rect 9970 25360 10042 25412
rect 10094 25360 10166 25412
rect 10218 25360 10260 25412
rect 9752 25288 10260 25360
rect 9752 25236 9794 25288
rect 9846 25236 9918 25288
rect 9970 25236 10042 25288
rect 10094 25236 10166 25288
rect 10218 25236 10260 25288
rect 9752 25164 10260 25236
rect 9752 25112 9794 25164
rect 9846 25112 9918 25164
rect 9970 25112 10042 25164
rect 10094 25112 10166 25164
rect 10218 25112 10260 25164
rect 9752 25040 10260 25112
rect 9752 24988 9794 25040
rect 9846 24988 9918 25040
rect 9970 24988 10042 25040
rect 10094 24988 10166 25040
rect 10218 24988 10260 25040
rect 9752 24916 10260 24988
rect 9752 24864 9794 24916
rect 9846 24864 9918 24916
rect 9970 24864 10042 24916
rect 10094 24864 10166 24916
rect 10218 24864 10260 24916
rect 9752 21469 10260 24864
rect 9752 21417 9764 21469
rect 9816 21417 9872 21469
rect 9924 21417 9980 21469
rect 10032 21417 10088 21469
rect 10140 21417 10196 21469
rect 10248 21417 10260 21469
rect 9752 21361 10260 21417
rect 9752 21309 9764 21361
rect 9816 21309 9872 21361
rect 9924 21309 9980 21361
rect 10032 21309 10088 21361
rect 10140 21309 10196 21361
rect 10248 21309 10260 21361
rect 9752 21253 10260 21309
rect 9752 21201 9764 21253
rect 9816 21201 9872 21253
rect 9924 21201 9980 21253
rect 10032 21201 10088 21253
rect 10140 21201 10196 21253
rect 10248 21201 10260 21253
rect 9752 19951 10260 21201
rect 9752 19899 9764 19951
rect 9816 19899 9872 19951
rect 9924 19899 9980 19951
rect 10032 19899 10088 19951
rect 10140 19899 10196 19951
rect 10248 19899 10260 19951
rect 9752 19843 10260 19899
rect 9752 19791 9764 19843
rect 9816 19791 9872 19843
rect 9924 19791 9980 19843
rect 10032 19791 10088 19843
rect 10140 19791 10196 19843
rect 10248 19791 10260 19843
rect 9752 19202 10260 19791
rect 9752 19150 9764 19202
rect 9816 19150 9872 19202
rect 9924 19150 9980 19202
rect 10032 19150 10088 19202
rect 10140 19150 10196 19202
rect 10248 19150 10260 19202
rect 9752 19094 10260 19150
rect 9752 19042 9764 19094
rect 9816 19042 9872 19094
rect 9924 19042 9980 19094
rect 10032 19042 10088 19094
rect 10140 19042 10196 19094
rect 10248 19042 10260 19094
rect 9752 18986 10260 19042
rect 9752 18934 9764 18986
rect 9816 18934 9872 18986
rect 9924 18934 9980 18986
rect 10032 18934 10088 18986
rect 10140 18934 10196 18986
rect 10248 18934 10260 18986
rect 9752 18330 10260 18934
rect 9752 18278 9764 18330
rect 9816 18278 9872 18330
rect 9924 18278 9980 18330
rect 10032 18278 10088 18330
rect 10140 18278 10196 18330
rect 10248 18278 10260 18330
rect 9752 18222 10260 18278
rect 9752 18170 9764 18222
rect 9816 18170 9872 18222
rect 9924 18170 9980 18222
rect 10032 18170 10088 18222
rect 10140 18170 10196 18222
rect 10248 18170 10260 18222
rect 9752 18114 10260 18170
rect 9752 18062 9764 18114
rect 9816 18062 9872 18114
rect 9924 18062 9980 18114
rect 10032 18062 10088 18114
rect 10140 18062 10196 18114
rect 10248 18062 10260 18114
rect 9752 17458 10260 18062
rect 9752 17406 9764 17458
rect 9816 17406 9872 17458
rect 9924 17406 9980 17458
rect 10032 17406 10088 17458
rect 10140 17406 10196 17458
rect 10248 17406 10260 17458
rect 9752 17350 10260 17406
rect 9752 17298 9764 17350
rect 9816 17298 9872 17350
rect 9924 17298 9980 17350
rect 10032 17298 10088 17350
rect 10140 17298 10196 17350
rect 10248 17298 10260 17350
rect 9752 17242 10260 17298
rect 9752 17190 9764 17242
rect 9816 17190 9872 17242
rect 9924 17190 9980 17242
rect 10032 17190 10088 17242
rect 10140 17190 10196 17242
rect 10248 17190 10260 17242
rect 9752 16601 10260 17190
rect 9752 16549 9764 16601
rect 9816 16549 9872 16601
rect 9924 16549 9980 16601
rect 10032 16549 10088 16601
rect 10140 16549 10196 16601
rect 10248 16549 10260 16601
rect 9752 16493 10260 16549
rect 9752 16441 9764 16493
rect 9816 16441 9872 16493
rect 9924 16441 9980 16493
rect 10032 16441 10088 16493
rect 10140 16441 10196 16493
rect 10248 16441 10260 16493
rect 9752 15762 10260 16441
rect 10888 56286 11396 56975
rect 10888 56234 11283 56286
rect 11335 56234 11396 56286
rect 10888 56178 11396 56234
rect 10888 56126 11283 56178
rect 11335 56126 11396 56178
rect 10888 56070 11396 56126
rect 10888 56018 11283 56070
rect 11335 56018 11396 56070
rect 10888 55962 11396 56018
rect 10888 55910 11283 55962
rect 11335 55910 11396 55962
rect 10888 55854 11396 55910
rect 10888 55802 11283 55854
rect 11335 55802 11396 55854
rect 10888 55746 11396 55802
rect 10888 55694 11283 55746
rect 11335 55694 11396 55746
rect 10888 55638 11396 55694
rect 10888 55586 11283 55638
rect 11335 55586 11396 55638
rect 10888 55530 11396 55586
rect 10888 55478 11283 55530
rect 11335 55478 11396 55530
rect 10888 55445 11396 55478
rect 10888 55389 10928 55445
rect 10984 55389 11052 55445
rect 11108 55389 11176 55445
rect 11232 55422 11300 55445
rect 11232 55389 11283 55422
rect 11356 55389 11396 55445
rect 10888 55370 11283 55389
rect 11335 55370 11396 55389
rect 10888 55321 11396 55370
rect 10888 55265 10928 55321
rect 10984 55265 11052 55321
rect 11108 55265 11176 55321
rect 11232 55314 11300 55321
rect 11232 55265 11283 55314
rect 11356 55265 11396 55321
rect 10888 55262 11283 55265
rect 11335 55262 11396 55265
rect 10888 55206 11396 55262
rect 10888 55197 11283 55206
rect 11335 55197 11396 55206
rect 10888 55141 10928 55197
rect 10984 55141 11052 55197
rect 11108 55141 11176 55197
rect 11232 55154 11283 55197
rect 11232 55141 11300 55154
rect 11356 55141 11396 55197
rect 10888 55098 11396 55141
rect 10888 55073 11283 55098
rect 11335 55073 11396 55098
rect 10888 55017 10928 55073
rect 10984 55017 11052 55073
rect 11108 55017 11176 55073
rect 11232 55046 11283 55073
rect 11232 55017 11300 55046
rect 11356 55017 11396 55073
rect 10888 54990 11396 55017
rect 10888 54949 11283 54990
rect 11335 54949 11396 54990
rect 10888 54893 10928 54949
rect 10984 54893 11052 54949
rect 11108 54893 11176 54949
rect 11232 54938 11283 54949
rect 11232 54893 11300 54938
rect 11356 54893 11396 54949
rect 10888 54882 11396 54893
rect 10888 54830 11283 54882
rect 11335 54830 11396 54882
rect 10888 54825 11396 54830
rect 10888 54769 10928 54825
rect 10984 54769 11052 54825
rect 11108 54769 11176 54825
rect 11232 54774 11300 54825
rect 11232 54769 11283 54774
rect 11356 54769 11396 54825
rect 10888 54722 11283 54769
rect 11335 54722 11396 54769
rect 10888 54701 11396 54722
rect 10888 54645 10928 54701
rect 10984 54645 11052 54701
rect 11108 54645 11176 54701
rect 11232 54666 11300 54701
rect 11232 54645 11283 54666
rect 11356 54645 11396 54701
rect 10888 54614 11283 54645
rect 11335 54614 11396 54645
rect 10888 54577 11396 54614
rect 10888 54521 10928 54577
rect 10984 54521 11052 54577
rect 11108 54521 11176 54577
rect 11232 54558 11300 54577
rect 11232 54521 11283 54558
rect 11356 54521 11396 54577
rect 10888 54506 11283 54521
rect 11335 54506 11396 54521
rect 10888 54453 11396 54506
rect 10888 54397 10928 54453
rect 10984 54397 11052 54453
rect 11108 54397 11176 54453
rect 11232 54450 11300 54453
rect 11232 54398 11283 54450
rect 11232 54397 11300 54398
rect 11356 54397 11396 54453
rect 10888 54342 11396 54397
rect 10888 54329 11283 54342
rect 11335 54329 11396 54342
rect 10888 54273 10928 54329
rect 10984 54273 11052 54329
rect 11108 54273 11176 54329
rect 11232 54290 11283 54329
rect 11232 54273 11300 54290
rect 11356 54273 11396 54329
rect 10888 54234 11396 54273
rect 10888 54205 11283 54234
rect 11335 54205 11396 54234
rect 10888 54149 10928 54205
rect 10984 54149 11052 54205
rect 11108 54149 11176 54205
rect 11232 54182 11283 54205
rect 11232 54149 11300 54182
rect 11356 54149 11396 54205
rect 10888 54126 11396 54149
rect 10888 54074 11283 54126
rect 11335 54074 11396 54126
rect 10888 54018 11396 54074
rect 10888 53966 11283 54018
rect 11335 53966 11396 54018
rect 10888 53910 11396 53966
rect 10888 53858 11283 53910
rect 11335 53858 11396 53910
rect 10888 53802 11396 53858
rect 10888 53750 11283 53802
rect 11335 53750 11396 53802
rect 10888 53694 11396 53750
rect 10888 53642 11283 53694
rect 11335 53642 11396 53694
rect 10888 53586 11396 53642
rect 10888 53534 11283 53586
rect 11335 53534 11396 53586
rect 10888 53478 11396 53534
rect 10888 53426 11283 53478
rect 11335 53426 11396 53478
rect 10888 53370 11396 53426
rect 10888 53318 11283 53370
rect 11335 53318 11396 53370
rect 10888 53262 11396 53318
rect 10888 53210 11283 53262
rect 11335 53210 11396 53262
rect 10888 52338 11396 53210
rect 10888 52286 11283 52338
rect 11335 52286 11396 52338
rect 10888 52230 11396 52286
rect 10888 52178 11283 52230
rect 11335 52178 11396 52230
rect 10888 52122 11396 52178
rect 10888 52070 11283 52122
rect 11335 52070 11396 52122
rect 10888 52014 11396 52070
rect 10888 51962 11283 52014
rect 11335 51962 11396 52014
rect 10888 51906 11396 51962
rect 10888 51854 11283 51906
rect 11335 51854 11396 51906
rect 10888 51798 11396 51854
rect 10888 51746 11283 51798
rect 11335 51746 11396 51798
rect 10888 51690 11396 51746
rect 10888 51638 11283 51690
rect 11335 51638 11396 51690
rect 10888 51582 11396 51638
rect 10888 51530 11283 51582
rect 11335 51530 11396 51582
rect 10888 51474 11396 51530
rect 10888 51422 11283 51474
rect 11335 51422 11396 51474
rect 10888 51366 11396 51422
rect 10888 51314 11283 51366
rect 11335 51314 11396 51366
rect 10888 51258 11396 51314
rect 10888 51206 11283 51258
rect 11335 51206 11396 51258
rect 10888 51150 11396 51206
rect 10888 51098 11283 51150
rect 11335 51098 11396 51150
rect 10888 51042 11396 51098
rect 10888 50990 11283 51042
rect 11335 50990 11396 51042
rect 10888 50934 11396 50990
rect 10888 50882 11283 50934
rect 11335 50882 11396 50934
rect 10888 50826 11396 50882
rect 10888 50774 11283 50826
rect 11335 50774 11396 50826
rect 10888 50718 11396 50774
rect 10888 50666 11283 50718
rect 11335 50666 11396 50718
rect 10888 50610 11396 50666
rect 10888 50558 11283 50610
rect 11335 50558 11396 50610
rect 10888 50502 11396 50558
rect 10888 50450 11283 50502
rect 11335 50450 11396 50502
rect 10888 50394 11396 50450
rect 10888 50342 11283 50394
rect 11335 50342 11396 50394
rect 10888 50286 11396 50342
rect 10888 50234 11283 50286
rect 11335 50234 11396 50286
rect 10888 50178 11396 50234
rect 10888 50126 11283 50178
rect 11335 50126 11396 50178
rect 10888 50070 11396 50126
rect 10888 50018 11283 50070
rect 11335 50018 11396 50070
rect 10888 49962 11396 50018
rect 10888 49910 11283 49962
rect 11335 49910 11396 49962
rect 10888 49854 11396 49910
rect 10888 49802 11283 49854
rect 11335 49802 11396 49854
rect 10888 49746 11396 49802
rect 10888 49694 11283 49746
rect 11335 49694 11396 49746
rect 10888 49638 11396 49694
rect 10888 49586 11283 49638
rect 11335 49586 11396 49638
rect 10888 49530 11396 49586
rect 10888 49478 11283 49530
rect 11335 49478 11396 49530
rect 10888 49422 11396 49478
rect 10888 49370 11283 49422
rect 11335 49370 11396 49422
rect 10888 49314 11396 49370
rect 10888 49262 11283 49314
rect 11335 49262 11396 49314
rect 10888 48390 11396 49262
rect 10888 48338 11283 48390
rect 11335 48338 11396 48390
rect 10888 48282 11396 48338
rect 10888 48230 11283 48282
rect 11335 48230 11396 48282
rect 10888 48174 11396 48230
rect 10888 48122 11283 48174
rect 11335 48122 11396 48174
rect 10888 48066 11396 48122
rect 10888 48014 11283 48066
rect 11335 48014 11396 48066
rect 10888 47958 11396 48014
rect 10888 47906 11283 47958
rect 11335 47906 11396 47958
rect 10888 47850 11396 47906
rect 10888 47798 11283 47850
rect 11335 47798 11396 47850
rect 10888 47742 11396 47798
rect 10888 47690 11283 47742
rect 11335 47690 11396 47742
rect 10888 47634 11396 47690
rect 10888 47582 11283 47634
rect 11335 47582 11396 47634
rect 10888 47526 11396 47582
rect 10888 47474 11283 47526
rect 11335 47474 11396 47526
rect 10888 47445 11396 47474
rect 10888 47389 10928 47445
rect 10984 47389 11052 47445
rect 11108 47389 11176 47445
rect 11232 47418 11300 47445
rect 11232 47389 11283 47418
rect 11356 47389 11396 47445
rect 10888 47366 11283 47389
rect 11335 47366 11396 47389
rect 10888 47321 11396 47366
rect 10888 47265 10928 47321
rect 10984 47265 11052 47321
rect 11108 47265 11176 47321
rect 11232 47310 11300 47321
rect 11232 47265 11283 47310
rect 11356 47265 11396 47321
rect 10888 47258 11283 47265
rect 11335 47258 11396 47265
rect 10888 47202 11396 47258
rect 10888 47197 11283 47202
rect 11335 47197 11396 47202
rect 10888 47141 10928 47197
rect 10984 47141 11052 47197
rect 11108 47141 11176 47197
rect 11232 47150 11283 47197
rect 11232 47141 11300 47150
rect 11356 47141 11396 47197
rect 10888 47094 11396 47141
rect 10888 47073 11283 47094
rect 11335 47073 11396 47094
rect 10888 47017 10928 47073
rect 10984 47017 11052 47073
rect 11108 47017 11176 47073
rect 11232 47042 11283 47073
rect 11232 47017 11300 47042
rect 11356 47017 11396 47073
rect 10888 46986 11396 47017
rect 10888 46949 11283 46986
rect 11335 46949 11396 46986
rect 10888 46893 10928 46949
rect 10984 46893 11052 46949
rect 11108 46893 11176 46949
rect 11232 46934 11283 46949
rect 11232 46893 11300 46934
rect 11356 46893 11396 46949
rect 10888 46878 11396 46893
rect 10888 46826 11283 46878
rect 11335 46826 11396 46878
rect 10888 46825 11396 46826
rect 10888 46769 10928 46825
rect 10984 46769 11052 46825
rect 11108 46769 11176 46825
rect 11232 46770 11300 46825
rect 11232 46769 11283 46770
rect 11356 46769 11396 46825
rect 10888 46718 11283 46769
rect 11335 46718 11396 46769
rect 10888 46701 11396 46718
rect 10888 46645 10928 46701
rect 10984 46645 11052 46701
rect 11108 46645 11176 46701
rect 11232 46662 11300 46701
rect 11232 46645 11283 46662
rect 11356 46645 11396 46701
rect 10888 46610 11283 46645
rect 11335 46610 11396 46645
rect 10888 46577 11396 46610
rect 10888 46521 10928 46577
rect 10984 46521 11052 46577
rect 11108 46521 11176 46577
rect 11232 46554 11300 46577
rect 11232 46521 11283 46554
rect 11356 46521 11396 46577
rect 10888 46502 11283 46521
rect 11335 46502 11396 46521
rect 10888 46453 11396 46502
rect 10888 46397 10928 46453
rect 10984 46397 11052 46453
rect 11108 46397 11176 46453
rect 11232 46446 11300 46453
rect 11232 46397 11283 46446
rect 11356 46397 11396 46453
rect 10888 46394 11283 46397
rect 11335 46394 11396 46397
rect 10888 46338 11396 46394
rect 10888 46329 11283 46338
rect 11335 46329 11396 46338
rect 10888 46273 10928 46329
rect 10984 46273 11052 46329
rect 11108 46273 11176 46329
rect 11232 46286 11283 46329
rect 11232 46273 11300 46286
rect 11356 46273 11396 46329
rect 10888 46230 11396 46273
rect 10888 46205 11283 46230
rect 11335 46205 11396 46230
rect 10888 46149 10928 46205
rect 10984 46149 11052 46205
rect 11108 46149 11176 46205
rect 11232 46178 11283 46205
rect 11232 46149 11300 46178
rect 11356 46149 11396 46205
rect 10888 46122 11396 46149
rect 10888 46070 11283 46122
rect 11335 46070 11396 46122
rect 10888 46014 11396 46070
rect 10888 45962 11283 46014
rect 11335 45962 11396 46014
rect 10888 45906 11396 45962
rect 10888 45854 11283 45906
rect 11335 45854 11396 45906
rect 10888 45798 11396 45854
rect 10888 45746 11283 45798
rect 11335 45746 11396 45798
rect 10888 45690 11396 45746
rect 10888 45638 11283 45690
rect 11335 45638 11396 45690
rect 10888 45582 11396 45638
rect 10888 45530 11283 45582
rect 11335 45530 11396 45582
rect 10888 45474 11396 45530
rect 10888 45422 11283 45474
rect 11335 45422 11396 45474
rect 10888 45366 11396 45422
rect 10888 45314 11283 45366
rect 11335 45314 11396 45366
rect 10888 44442 11396 45314
rect 10888 44390 11283 44442
rect 11335 44390 11396 44442
rect 10888 44334 11396 44390
rect 10888 44282 11283 44334
rect 11335 44282 11396 44334
rect 10888 44245 11396 44282
rect 10888 44189 10928 44245
rect 10984 44189 11052 44245
rect 11108 44189 11176 44245
rect 11232 44226 11300 44245
rect 11232 44189 11283 44226
rect 11356 44189 11396 44245
rect 10888 44174 11283 44189
rect 11335 44174 11396 44189
rect 10888 44121 11396 44174
rect 10888 44065 10928 44121
rect 10984 44065 11052 44121
rect 11108 44065 11176 44121
rect 11232 44118 11300 44121
rect 11232 44066 11283 44118
rect 11232 44065 11300 44066
rect 11356 44065 11396 44121
rect 10888 44010 11396 44065
rect 10888 43997 11283 44010
rect 11335 43997 11396 44010
rect 10888 43941 10928 43997
rect 10984 43941 11052 43997
rect 11108 43941 11176 43997
rect 11232 43958 11283 43997
rect 11232 43941 11300 43958
rect 11356 43941 11396 43997
rect 10888 43902 11396 43941
rect 10888 43873 11283 43902
rect 11335 43873 11396 43902
rect 10888 43817 10928 43873
rect 10984 43817 11052 43873
rect 11108 43817 11176 43873
rect 11232 43850 11283 43873
rect 11232 43817 11300 43850
rect 11356 43817 11396 43873
rect 10888 43794 11396 43817
rect 10888 43749 11283 43794
rect 11335 43749 11396 43794
rect 10888 43693 10928 43749
rect 10984 43693 11052 43749
rect 11108 43693 11176 43749
rect 11232 43742 11283 43749
rect 11232 43693 11300 43742
rect 11356 43693 11396 43749
rect 10888 43686 11396 43693
rect 10888 43634 11283 43686
rect 11335 43634 11396 43686
rect 10888 43625 11396 43634
rect 10888 43569 10928 43625
rect 10984 43569 11052 43625
rect 11108 43569 11176 43625
rect 11232 43578 11300 43625
rect 11232 43569 11283 43578
rect 11356 43569 11396 43625
rect 10888 43526 11283 43569
rect 11335 43526 11396 43569
rect 10888 43501 11396 43526
rect 10888 43445 10928 43501
rect 10984 43445 11052 43501
rect 11108 43445 11176 43501
rect 11232 43470 11300 43501
rect 11232 43445 11283 43470
rect 11356 43445 11396 43501
rect 10888 43418 11283 43445
rect 11335 43418 11396 43445
rect 10888 43377 11396 43418
rect 10888 43321 10928 43377
rect 10984 43321 11052 43377
rect 11108 43321 11176 43377
rect 11232 43362 11300 43377
rect 11232 43321 11283 43362
rect 11356 43321 11396 43377
rect 10888 43310 11283 43321
rect 11335 43310 11396 43321
rect 10888 43254 11396 43310
rect 10888 43253 11283 43254
rect 11335 43253 11396 43254
rect 10888 43197 10928 43253
rect 10984 43197 11052 43253
rect 11108 43197 11176 43253
rect 11232 43202 11283 43253
rect 11232 43197 11300 43202
rect 11356 43197 11396 43253
rect 10888 43146 11396 43197
rect 10888 43129 11283 43146
rect 11335 43129 11396 43146
rect 10888 43073 10928 43129
rect 10984 43073 11052 43129
rect 11108 43073 11176 43129
rect 11232 43094 11283 43129
rect 11232 43073 11300 43094
rect 11356 43073 11396 43129
rect 10888 43038 11396 43073
rect 10888 43005 11283 43038
rect 11335 43005 11396 43038
rect 10888 42949 10928 43005
rect 10984 42949 11052 43005
rect 11108 42949 11176 43005
rect 11232 42986 11283 43005
rect 11232 42949 11300 42986
rect 11356 42949 11396 43005
rect 10888 42930 11396 42949
rect 10888 42878 11283 42930
rect 11335 42878 11396 42930
rect 10888 42822 11396 42878
rect 10888 42770 11283 42822
rect 11335 42770 11396 42822
rect 10888 42714 11396 42770
rect 10888 42662 11283 42714
rect 11335 42662 11396 42714
rect 10888 42645 11396 42662
rect 10888 42589 10928 42645
rect 10984 42589 11052 42645
rect 11108 42589 11176 42645
rect 11232 42606 11300 42645
rect 11232 42589 11283 42606
rect 11356 42589 11396 42645
rect 10888 42554 11283 42589
rect 11335 42554 11396 42589
rect 10888 42521 11396 42554
rect 10888 42465 10928 42521
rect 10984 42465 11052 42521
rect 11108 42465 11176 42521
rect 11232 42498 11300 42521
rect 11232 42465 11283 42498
rect 11356 42465 11396 42521
rect 10888 42446 11283 42465
rect 11335 42446 11396 42465
rect 10888 42397 11396 42446
rect 10888 42341 10928 42397
rect 10984 42341 11052 42397
rect 11108 42341 11176 42397
rect 11232 42390 11300 42397
rect 11232 42341 11283 42390
rect 11356 42341 11396 42397
rect 10888 42338 11283 42341
rect 11335 42338 11396 42341
rect 10888 42282 11396 42338
rect 10888 42273 11283 42282
rect 11335 42273 11396 42282
rect 10888 42217 10928 42273
rect 10984 42217 11052 42273
rect 11108 42217 11176 42273
rect 11232 42230 11283 42273
rect 11232 42217 11300 42230
rect 11356 42217 11396 42273
rect 10888 42174 11396 42217
rect 10888 42149 11283 42174
rect 11335 42149 11396 42174
rect 10888 42093 10928 42149
rect 10984 42093 11052 42149
rect 11108 42093 11176 42149
rect 11232 42122 11283 42149
rect 11232 42093 11300 42122
rect 11356 42093 11396 42149
rect 10888 42066 11396 42093
rect 10888 42025 11283 42066
rect 11335 42025 11396 42066
rect 10888 41969 10928 42025
rect 10984 41969 11052 42025
rect 11108 41969 11176 42025
rect 11232 42014 11283 42025
rect 11232 41969 11300 42014
rect 11356 41969 11396 42025
rect 10888 41958 11396 41969
rect 10888 41906 11283 41958
rect 11335 41906 11396 41958
rect 10888 41901 11396 41906
rect 10888 41845 10928 41901
rect 10984 41845 11052 41901
rect 11108 41845 11176 41901
rect 11232 41850 11300 41901
rect 11232 41845 11283 41850
rect 11356 41845 11396 41901
rect 10888 41798 11283 41845
rect 11335 41798 11396 41845
rect 10888 41777 11396 41798
rect 10888 41721 10928 41777
rect 10984 41721 11052 41777
rect 11108 41721 11176 41777
rect 11232 41742 11300 41777
rect 11232 41721 11283 41742
rect 11356 41721 11396 41777
rect 10888 41690 11283 41721
rect 11335 41690 11396 41721
rect 10888 41653 11396 41690
rect 10888 41597 10928 41653
rect 10984 41597 11052 41653
rect 11108 41597 11176 41653
rect 11232 41634 11300 41653
rect 11232 41597 11283 41634
rect 11356 41597 11396 41653
rect 10888 41582 11283 41597
rect 11335 41582 11396 41597
rect 10888 41529 11396 41582
rect 10888 41473 10928 41529
rect 10984 41473 11052 41529
rect 11108 41473 11176 41529
rect 11232 41526 11300 41529
rect 11232 41474 11283 41526
rect 11232 41473 11300 41474
rect 11356 41473 11396 41529
rect 10888 41418 11396 41473
rect 10888 41405 11283 41418
rect 11335 41405 11396 41418
rect 10888 41349 10928 41405
rect 10984 41349 11052 41405
rect 11108 41349 11176 41405
rect 11232 41366 11283 41405
rect 11232 41349 11300 41366
rect 11356 41349 11396 41405
rect 10888 41045 11396 41349
rect 10888 40989 10928 41045
rect 10984 40989 11052 41045
rect 11108 40989 11176 41045
rect 11232 40989 11300 41045
rect 11356 40989 11396 41045
rect 10888 40921 11396 40989
rect 10888 40865 10928 40921
rect 10984 40865 11052 40921
rect 11108 40865 11176 40921
rect 11232 40865 11300 40921
rect 11356 40865 11396 40921
rect 10888 40797 11396 40865
rect 10888 40741 10928 40797
rect 10984 40741 11052 40797
rect 11108 40741 11176 40797
rect 11232 40741 11300 40797
rect 11356 40741 11396 40797
rect 10888 40673 11396 40741
rect 10888 40617 10928 40673
rect 10984 40617 11052 40673
rect 11108 40617 11176 40673
rect 11232 40617 11300 40673
rect 11356 40617 11396 40673
rect 10888 40549 11396 40617
rect 10888 40493 10928 40549
rect 10984 40493 11052 40549
rect 11108 40493 11176 40549
rect 11232 40494 11300 40549
rect 11232 40493 11283 40494
rect 11356 40493 11396 40549
rect 10888 40442 11283 40493
rect 11335 40442 11396 40493
rect 10888 40425 11396 40442
rect 10888 40369 10928 40425
rect 10984 40369 11052 40425
rect 11108 40369 11176 40425
rect 11232 40386 11300 40425
rect 11232 40369 11283 40386
rect 11356 40369 11396 40425
rect 10888 40334 11283 40369
rect 11335 40334 11396 40369
rect 10888 40301 11396 40334
rect 10888 40245 10928 40301
rect 10984 40245 11052 40301
rect 11108 40245 11176 40301
rect 11232 40278 11300 40301
rect 11232 40245 11283 40278
rect 11356 40245 11396 40301
rect 10888 40226 11283 40245
rect 11335 40226 11396 40245
rect 10888 40177 11396 40226
rect 10888 40121 10928 40177
rect 10984 40121 11052 40177
rect 11108 40121 11176 40177
rect 11232 40170 11300 40177
rect 11232 40121 11283 40170
rect 11356 40121 11396 40177
rect 10888 40118 11283 40121
rect 11335 40118 11396 40121
rect 10888 40062 11396 40118
rect 10888 40053 11283 40062
rect 11335 40053 11396 40062
rect 10888 39997 10928 40053
rect 10984 39997 11052 40053
rect 11108 39997 11176 40053
rect 11232 40010 11283 40053
rect 11232 39997 11300 40010
rect 11356 39997 11396 40053
rect 10888 39954 11396 39997
rect 10888 39929 11283 39954
rect 11335 39929 11396 39954
rect 10888 39873 10928 39929
rect 10984 39873 11052 39929
rect 11108 39873 11176 39929
rect 11232 39902 11283 39929
rect 11232 39873 11300 39902
rect 11356 39873 11396 39929
rect 10888 39846 11396 39873
rect 10888 39805 11283 39846
rect 11335 39805 11396 39846
rect 10888 39749 10928 39805
rect 10984 39749 11052 39805
rect 11108 39749 11176 39805
rect 11232 39794 11283 39805
rect 11232 39749 11300 39794
rect 11356 39749 11396 39805
rect 10888 39738 11396 39749
rect 10888 39686 11283 39738
rect 11335 39686 11396 39738
rect 10888 39630 11396 39686
rect 10888 39578 11283 39630
rect 11335 39578 11396 39630
rect 10888 39522 11396 39578
rect 10888 39470 11283 39522
rect 11335 39470 11396 39522
rect 10888 39414 11396 39470
rect 10888 39362 11283 39414
rect 11335 39362 11396 39414
rect 10888 39306 11396 39362
rect 10888 39254 11283 39306
rect 11335 39254 11396 39306
rect 10888 39198 11396 39254
rect 10888 39146 11283 39198
rect 11335 39146 11396 39198
rect 10888 39090 11396 39146
rect 10888 39038 11283 39090
rect 11335 39038 11396 39090
rect 10888 38982 11396 39038
rect 10888 38930 11283 38982
rect 11335 38930 11396 38982
rect 10888 38874 11396 38930
rect 10888 38822 11283 38874
rect 11335 38822 11396 38874
rect 10888 38766 11396 38822
rect 10888 38714 11283 38766
rect 11335 38714 11396 38766
rect 10888 38658 11396 38714
rect 10888 38606 11283 38658
rect 11335 38606 11396 38658
rect 10888 38550 11396 38606
rect 10888 38498 11283 38550
rect 11335 38498 11396 38550
rect 10888 38442 11396 38498
rect 10888 38390 11283 38442
rect 11335 38390 11396 38442
rect 10888 38334 11396 38390
rect 10888 38282 11283 38334
rect 11335 38282 11396 38334
rect 10888 38226 11396 38282
rect 10888 38174 11283 38226
rect 11335 38174 11396 38226
rect 10888 38118 11396 38174
rect 10888 38066 11283 38118
rect 11335 38066 11396 38118
rect 10888 38010 11396 38066
rect 10888 37958 11283 38010
rect 11335 37958 11396 38010
rect 10888 37902 11396 37958
rect 10888 37850 11283 37902
rect 11335 37850 11396 37902
rect 10888 37794 11396 37850
rect 10888 37742 11283 37794
rect 11335 37742 11396 37794
rect 10888 37686 11396 37742
rect 10888 37634 11283 37686
rect 11335 37634 11396 37686
rect 10888 37578 11396 37634
rect 10888 37526 11283 37578
rect 11335 37526 11396 37578
rect 10888 37470 11396 37526
rect 10888 37418 11283 37470
rect 11335 37418 11396 37470
rect 10888 36546 11396 37418
rect 10888 36494 11283 36546
rect 11335 36494 11396 36546
rect 10888 36438 11396 36494
rect 10888 36386 11283 36438
rect 11335 36386 11396 36438
rect 10888 36330 11396 36386
rect 10888 36278 11283 36330
rect 11335 36278 11396 36330
rect 10888 36222 11396 36278
rect 10888 36170 11283 36222
rect 11335 36170 11396 36222
rect 10888 36114 11396 36170
rect 10888 36062 11283 36114
rect 11335 36062 11396 36114
rect 10888 36006 11396 36062
rect 10888 35954 11283 36006
rect 11335 35954 11396 36006
rect 10888 35898 11396 35954
rect 10888 35846 11283 35898
rect 11335 35846 11396 35898
rect 10888 35790 11396 35846
rect 10888 35738 11283 35790
rect 11335 35738 11396 35790
rect 10888 35682 11396 35738
rect 10888 35630 11283 35682
rect 11335 35630 11396 35682
rect 10888 35574 11396 35630
rect 10888 35522 11283 35574
rect 11335 35522 11396 35574
rect 10888 35466 11396 35522
rect 10888 35414 11283 35466
rect 11335 35414 11396 35466
rect 10888 35358 11396 35414
rect 10888 35306 11283 35358
rect 11335 35306 11396 35358
rect 10888 35250 11396 35306
rect 10888 35198 11283 35250
rect 11335 35198 11396 35250
rect 10888 35142 11396 35198
rect 10888 35090 11283 35142
rect 11335 35090 11396 35142
rect 10888 35034 11396 35090
rect 10888 34982 11283 35034
rect 11335 34982 11396 35034
rect 10888 34926 11396 34982
rect 10888 34874 11283 34926
rect 11335 34874 11396 34926
rect 10888 34818 11396 34874
rect 10888 34766 11283 34818
rect 11335 34766 11396 34818
rect 10888 34710 11396 34766
rect 10888 34658 11283 34710
rect 11335 34658 11396 34710
rect 10888 34602 11396 34658
rect 10888 34550 11283 34602
rect 11335 34550 11396 34602
rect 10888 34494 11396 34550
rect 10888 34442 11283 34494
rect 11335 34442 11396 34494
rect 10888 34386 11396 34442
rect 10888 34334 11283 34386
rect 11335 34334 11396 34386
rect 10888 34278 11396 34334
rect 10888 34226 11283 34278
rect 11335 34226 11396 34278
rect 10888 34170 11396 34226
rect 10888 34118 11283 34170
rect 11335 34118 11396 34170
rect 10888 34062 11396 34118
rect 10888 34010 11283 34062
rect 11335 34010 11396 34062
rect 10888 33954 11396 34010
rect 10888 33902 11283 33954
rect 11335 33902 11396 33954
rect 10888 33846 11396 33902
rect 10888 33794 11283 33846
rect 11335 33794 11396 33846
rect 10888 33738 11396 33794
rect 10888 33686 11283 33738
rect 11335 33686 11396 33738
rect 10888 33630 11396 33686
rect 10888 33578 11283 33630
rect 11335 33578 11396 33630
rect 10888 33522 11396 33578
rect 10888 33470 11283 33522
rect 11335 33470 11396 33522
rect 10888 33051 11396 33470
rect 10888 32995 10928 33051
rect 10984 32995 11052 33051
rect 11108 32995 11176 33051
rect 11232 32995 11300 33051
rect 11356 32995 11396 33051
rect 10888 32927 11396 32995
rect 10888 32871 10928 32927
rect 10984 32871 11052 32927
rect 11108 32871 11176 32927
rect 11232 32871 11300 32927
rect 11356 32871 11396 32927
rect 10888 32803 11396 32871
rect 10888 32747 10928 32803
rect 10984 32747 11052 32803
rect 11108 32747 11176 32803
rect 11232 32747 11300 32803
rect 11356 32747 11396 32803
rect 10888 32679 11396 32747
rect 10888 32623 10928 32679
rect 10984 32623 11052 32679
rect 11108 32623 11176 32679
rect 11232 32623 11300 32679
rect 11356 32623 11396 32679
rect 10888 32598 11396 32623
rect 10888 32555 11283 32598
rect 11335 32555 11396 32598
rect 10888 32499 10928 32555
rect 10984 32499 11052 32555
rect 11108 32499 11176 32555
rect 11232 32546 11283 32555
rect 11232 32499 11300 32546
rect 11356 32499 11396 32555
rect 10888 32490 11396 32499
rect 10888 32438 11283 32490
rect 11335 32438 11396 32490
rect 10888 32431 11396 32438
rect 10888 32375 10928 32431
rect 10984 32375 11052 32431
rect 11108 32375 11176 32431
rect 11232 32382 11300 32431
rect 11232 32375 11283 32382
rect 11356 32375 11396 32431
rect 10888 32330 11283 32375
rect 11335 32330 11396 32375
rect 10888 32307 11396 32330
rect 10888 32251 10928 32307
rect 10984 32251 11052 32307
rect 11108 32251 11176 32307
rect 11232 32274 11300 32307
rect 11232 32251 11283 32274
rect 11356 32251 11396 32307
rect 10888 32222 11283 32251
rect 11335 32222 11396 32251
rect 10888 32183 11396 32222
rect 10888 32127 10928 32183
rect 10984 32127 11052 32183
rect 11108 32127 11176 32183
rect 11232 32166 11300 32183
rect 11232 32127 11283 32166
rect 11356 32127 11396 32183
rect 10888 32114 11283 32127
rect 11335 32114 11396 32127
rect 10888 32059 11396 32114
rect 10888 32003 10928 32059
rect 10984 32003 11052 32059
rect 11108 32003 11176 32059
rect 11232 32058 11300 32059
rect 11232 32006 11283 32058
rect 11232 32003 11300 32006
rect 11356 32003 11396 32059
rect 10888 31950 11396 32003
rect 10888 31935 11283 31950
rect 11335 31935 11396 31950
rect 10888 31879 10928 31935
rect 10984 31879 11052 31935
rect 11108 31879 11176 31935
rect 11232 31898 11283 31935
rect 11232 31879 11300 31898
rect 11356 31879 11396 31935
rect 10888 31842 11396 31879
rect 10888 31811 11283 31842
rect 11335 31811 11396 31842
rect 10888 31755 10928 31811
rect 10984 31755 11052 31811
rect 11108 31755 11176 31811
rect 11232 31790 11283 31811
rect 11232 31755 11300 31790
rect 11356 31755 11396 31811
rect 10888 31734 11396 31755
rect 10888 31687 11283 31734
rect 11335 31687 11396 31734
rect 10888 31631 10928 31687
rect 10984 31631 11052 31687
rect 11108 31631 11176 31687
rect 11232 31682 11283 31687
rect 11232 31631 11300 31682
rect 11356 31631 11396 31687
rect 10888 31626 11396 31631
rect 10888 31574 11283 31626
rect 11335 31574 11396 31626
rect 10888 31563 11396 31574
rect 10888 31507 10928 31563
rect 10984 31507 11052 31563
rect 11108 31507 11176 31563
rect 11232 31518 11300 31563
rect 11232 31507 11283 31518
rect 11356 31507 11396 31563
rect 10888 31466 11283 31507
rect 11335 31466 11396 31507
rect 10888 31439 11396 31466
rect 10888 31383 10928 31439
rect 10984 31383 11052 31439
rect 11108 31383 11176 31439
rect 11232 31410 11300 31439
rect 11232 31383 11283 31410
rect 11356 31383 11396 31439
rect 10888 31358 11283 31383
rect 11335 31358 11396 31383
rect 10888 31315 11396 31358
rect 10888 31259 10928 31315
rect 10984 31259 11052 31315
rect 11108 31259 11176 31315
rect 11232 31302 11300 31315
rect 11232 31259 11283 31302
rect 11356 31259 11396 31315
rect 10888 31250 11283 31259
rect 11335 31250 11396 31259
rect 10888 31194 11396 31250
rect 10888 31191 11283 31194
rect 11335 31191 11396 31194
rect 10888 31135 10928 31191
rect 10984 31135 11052 31191
rect 11108 31135 11176 31191
rect 11232 31142 11283 31191
rect 11232 31135 11300 31142
rect 11356 31135 11396 31191
rect 10888 31086 11396 31135
rect 10888 31067 11283 31086
rect 11335 31067 11396 31086
rect 10888 31011 10928 31067
rect 10984 31011 11052 31067
rect 11108 31011 11176 31067
rect 11232 31034 11283 31067
rect 11232 31011 11300 31034
rect 11356 31011 11396 31067
rect 10888 30978 11396 31011
rect 10888 30943 11283 30978
rect 11335 30943 11396 30978
rect 10888 30887 10928 30943
rect 10984 30887 11052 30943
rect 11108 30887 11176 30943
rect 11232 30926 11283 30943
rect 11232 30887 11300 30926
rect 11356 30887 11396 30943
rect 10888 30870 11396 30887
rect 10888 30819 11283 30870
rect 11335 30819 11396 30870
rect 10888 30763 10928 30819
rect 10984 30763 11052 30819
rect 11108 30763 11176 30819
rect 11232 30818 11283 30819
rect 11232 30763 11300 30818
rect 11356 30763 11396 30819
rect 10888 30762 11396 30763
rect 10888 30710 11283 30762
rect 11335 30710 11396 30762
rect 10888 30695 11396 30710
rect 10888 30639 10928 30695
rect 10984 30639 11052 30695
rect 11108 30639 11176 30695
rect 11232 30654 11300 30695
rect 11232 30639 11283 30654
rect 11356 30639 11396 30695
rect 10888 30602 11283 30639
rect 11335 30602 11396 30639
rect 10888 30571 11396 30602
rect 10888 30515 10928 30571
rect 10984 30515 11052 30571
rect 11108 30515 11176 30571
rect 11232 30546 11300 30571
rect 11232 30515 11283 30546
rect 11356 30515 11396 30571
rect 10888 30494 11283 30515
rect 11335 30494 11396 30515
rect 10888 30447 11396 30494
rect 10888 30391 10928 30447
rect 10984 30391 11052 30447
rect 11108 30391 11176 30447
rect 11232 30438 11300 30447
rect 11232 30391 11283 30438
rect 11356 30391 11396 30447
rect 10888 30386 11283 30391
rect 11335 30386 11396 30391
rect 10888 30330 11396 30386
rect 10888 30323 11283 30330
rect 11335 30323 11396 30330
rect 10888 30267 10928 30323
rect 10984 30267 11052 30323
rect 11108 30267 11176 30323
rect 11232 30278 11283 30323
rect 11232 30267 11300 30278
rect 11356 30267 11396 30323
rect 10888 30222 11396 30267
rect 10888 30199 11283 30222
rect 11335 30199 11396 30222
rect 10888 30143 10928 30199
rect 10984 30143 11052 30199
rect 11108 30143 11176 30199
rect 11232 30170 11283 30199
rect 11232 30143 11300 30170
rect 11356 30143 11396 30199
rect 10888 30114 11396 30143
rect 10888 30062 11283 30114
rect 11335 30062 11396 30114
rect 10888 30006 11396 30062
rect 10888 29954 11283 30006
rect 11335 29954 11396 30006
rect 10888 29898 11396 29954
rect 10888 29846 11283 29898
rect 11335 29846 11396 29898
rect 10888 29845 11396 29846
rect 10888 29789 10928 29845
rect 10984 29789 11052 29845
rect 11108 29789 11176 29845
rect 11232 29790 11300 29845
rect 11232 29789 11283 29790
rect 11356 29789 11396 29845
rect 10888 29738 11283 29789
rect 11335 29738 11396 29789
rect 10888 29721 11396 29738
rect 10888 29665 10928 29721
rect 10984 29665 11052 29721
rect 11108 29665 11176 29721
rect 11232 29682 11300 29721
rect 11232 29665 11283 29682
rect 11356 29665 11396 29721
rect 10888 29630 11283 29665
rect 11335 29630 11396 29665
rect 10888 29597 11396 29630
rect 10888 29541 10928 29597
rect 10984 29541 11052 29597
rect 11108 29541 11176 29597
rect 11232 29574 11300 29597
rect 11232 29541 11283 29574
rect 11356 29541 11396 29597
rect 10888 29522 11283 29541
rect 11335 29522 11396 29541
rect 10888 29473 11396 29522
rect 10888 29417 10928 29473
rect 10984 29417 11052 29473
rect 11108 29417 11176 29473
rect 11232 29417 11300 29473
rect 11356 29417 11396 29473
rect 10888 29349 11396 29417
rect 10888 29293 10928 29349
rect 10984 29293 11052 29349
rect 11108 29293 11176 29349
rect 11232 29293 11300 29349
rect 11356 29293 11396 29349
rect 10888 29225 11396 29293
rect 10888 29169 10928 29225
rect 10984 29169 11052 29225
rect 11108 29169 11176 29225
rect 11232 29169 11300 29225
rect 11356 29169 11396 29225
rect 10888 29101 11396 29169
rect 10888 29045 10928 29101
rect 10984 29045 11052 29101
rect 11108 29045 11176 29101
rect 11232 29045 11300 29101
rect 11356 29045 11396 29101
rect 10888 28977 11396 29045
rect 10888 28921 10928 28977
rect 10984 28921 11052 28977
rect 11108 28921 11176 28977
rect 11232 28921 11300 28977
rect 11356 28921 11396 28977
rect 10888 28853 11396 28921
rect 10888 28797 10928 28853
rect 10984 28797 11052 28853
rect 11108 28797 11176 28853
rect 11232 28797 11300 28853
rect 11356 28797 11396 28853
rect 10888 28729 11396 28797
rect 10888 28673 10928 28729
rect 10984 28673 11052 28729
rect 11108 28673 11176 28729
rect 11232 28673 11300 28729
rect 11356 28673 11396 28729
rect 10888 28650 11396 28673
rect 10888 28605 11283 28650
rect 11335 28605 11396 28650
rect 10888 28549 10928 28605
rect 10984 28549 11052 28605
rect 11108 28549 11176 28605
rect 11232 28598 11283 28605
rect 11232 28549 11300 28598
rect 11356 28549 11396 28605
rect 10888 28542 11396 28549
rect 10888 28490 11283 28542
rect 11335 28490 11396 28542
rect 10888 28434 11396 28490
rect 10888 28382 11283 28434
rect 11335 28382 11396 28434
rect 10888 28326 11396 28382
rect 10888 28274 11283 28326
rect 11335 28274 11396 28326
rect 10888 28218 11396 28274
rect 10888 28166 11283 28218
rect 11335 28166 11396 28218
rect 10888 28110 11396 28166
rect 10888 28058 11283 28110
rect 11335 28058 11396 28110
rect 10888 28002 11396 28058
rect 10888 27950 11283 28002
rect 11335 27950 11396 28002
rect 10888 27894 11396 27950
rect 10888 27842 11283 27894
rect 11335 27842 11396 27894
rect 10888 27786 11396 27842
rect 10888 27734 11283 27786
rect 11335 27734 11396 27786
rect 10888 27678 11396 27734
rect 10888 27626 11283 27678
rect 11335 27626 11396 27678
rect 10888 27570 11396 27626
rect 10888 27518 11283 27570
rect 11335 27518 11396 27570
rect 10888 27462 11396 27518
rect 10888 27410 11283 27462
rect 11335 27410 11396 27462
rect 10888 27354 11396 27410
rect 10888 27302 11283 27354
rect 11335 27302 11396 27354
rect 10888 27246 11396 27302
rect 10888 27194 11283 27246
rect 11335 27194 11396 27246
rect 10888 27138 11396 27194
rect 10888 27086 11283 27138
rect 11335 27086 11396 27138
rect 10888 27030 11396 27086
rect 10888 26978 11283 27030
rect 11335 26978 11396 27030
rect 10888 26922 11396 26978
rect 10888 26870 11283 26922
rect 11335 26870 11396 26922
rect 10888 26814 11396 26870
rect 10888 26762 11283 26814
rect 11335 26762 11396 26814
rect 10888 26706 11396 26762
rect 10888 26654 11283 26706
rect 11335 26654 11396 26706
rect 10888 26651 11396 26654
rect 10888 26595 10928 26651
rect 10984 26595 11052 26651
rect 11108 26595 11176 26651
rect 11232 26598 11300 26651
rect 11232 26595 11283 26598
rect 11356 26595 11396 26651
rect 10888 26546 11283 26595
rect 11335 26546 11396 26595
rect 10888 26527 11396 26546
rect 10888 26471 10928 26527
rect 10984 26471 11052 26527
rect 11108 26471 11176 26527
rect 11232 26490 11300 26527
rect 11232 26471 11283 26490
rect 11356 26471 11396 26527
rect 10888 26438 11283 26471
rect 11335 26438 11396 26471
rect 10888 26403 11396 26438
rect 10888 26347 10928 26403
rect 10984 26347 11052 26403
rect 11108 26347 11176 26403
rect 11232 26382 11300 26403
rect 11232 26347 11283 26382
rect 11356 26347 11396 26403
rect 10888 26330 11283 26347
rect 11335 26330 11396 26347
rect 10888 26279 11396 26330
rect 10888 26223 10928 26279
rect 10984 26223 11052 26279
rect 11108 26223 11176 26279
rect 11232 26274 11300 26279
rect 11232 26223 11283 26274
rect 11356 26223 11396 26279
rect 10888 26222 11283 26223
rect 11335 26222 11396 26223
rect 10888 26166 11396 26222
rect 10888 26155 11283 26166
rect 11335 26155 11396 26166
rect 10888 26099 10928 26155
rect 10984 26099 11052 26155
rect 11108 26099 11176 26155
rect 11232 26114 11283 26155
rect 11232 26099 11300 26114
rect 11356 26099 11396 26155
rect 10888 26058 11396 26099
rect 10888 26031 11283 26058
rect 11335 26031 11396 26058
rect 10888 25975 10928 26031
rect 10984 25975 11052 26031
rect 11108 25975 11176 26031
rect 11232 26006 11283 26031
rect 11232 25975 11300 26006
rect 11356 25975 11396 26031
rect 10888 25950 11396 25975
rect 10888 25907 11283 25950
rect 11335 25907 11396 25950
rect 10888 25851 10928 25907
rect 10984 25851 11052 25907
rect 11108 25851 11176 25907
rect 11232 25898 11283 25907
rect 11232 25851 11300 25898
rect 11356 25851 11396 25907
rect 10888 25842 11396 25851
rect 10888 25790 11283 25842
rect 11335 25790 11396 25842
rect 10888 25783 11396 25790
rect 10888 25727 10928 25783
rect 10984 25727 11052 25783
rect 11108 25727 11176 25783
rect 11232 25734 11300 25783
rect 11232 25727 11283 25734
rect 11356 25727 11396 25783
rect 10888 25682 11283 25727
rect 11335 25682 11396 25727
rect 10888 25659 11396 25682
rect 10888 25603 10928 25659
rect 10984 25603 11052 25659
rect 11108 25603 11176 25659
rect 11232 25626 11300 25659
rect 11232 25603 11283 25626
rect 11356 25603 11396 25659
rect 10888 25574 11283 25603
rect 11335 25574 11396 25603
rect 10888 25535 11396 25574
rect 10888 25479 10928 25535
rect 10984 25479 11052 25535
rect 11108 25479 11176 25535
rect 11232 25479 11300 25535
rect 11356 25479 11396 25535
rect 10888 25411 11396 25479
rect 10888 25355 10928 25411
rect 10984 25355 11052 25411
rect 11108 25355 11176 25411
rect 11232 25355 11300 25411
rect 11356 25355 11396 25411
rect 10888 25287 11396 25355
rect 10888 25231 10928 25287
rect 10984 25231 11052 25287
rect 11108 25231 11176 25287
rect 11232 25231 11300 25287
rect 11356 25231 11396 25287
rect 10888 25163 11396 25231
rect 10888 25107 10928 25163
rect 10984 25107 11052 25163
rect 11108 25107 11176 25163
rect 11232 25107 11300 25163
rect 11356 25107 11396 25163
rect 10888 25039 11396 25107
rect 10888 24983 10928 25039
rect 10984 24983 11052 25039
rect 11108 24983 11176 25039
rect 11232 24983 11300 25039
rect 11356 24983 11396 25039
rect 10888 24915 11396 24983
rect 10888 24859 10928 24915
rect 10984 24859 11052 24915
rect 11108 24859 11176 24915
rect 11232 24859 11300 24915
rect 11356 24859 11396 24915
rect 10888 24791 11396 24859
rect 10888 24735 10928 24791
rect 10984 24735 11052 24791
rect 11108 24735 11176 24791
rect 11232 24735 11300 24791
rect 11356 24735 11396 24791
rect 10888 24702 11396 24735
rect 10888 24667 11283 24702
rect 11335 24667 11396 24702
rect 10888 24611 10928 24667
rect 10984 24611 11052 24667
rect 11108 24611 11176 24667
rect 11232 24650 11283 24667
rect 11232 24611 11300 24650
rect 11356 24611 11396 24667
rect 10888 24594 11396 24611
rect 10888 24543 11283 24594
rect 11335 24543 11396 24594
rect 10888 24487 10928 24543
rect 10984 24487 11052 24543
rect 11108 24487 11176 24543
rect 11232 24542 11283 24543
rect 11232 24487 11300 24542
rect 11356 24487 11396 24543
rect 10888 24486 11396 24487
rect 10888 24434 11283 24486
rect 11335 24434 11396 24486
rect 10888 24419 11396 24434
rect 10888 24363 10928 24419
rect 10984 24363 11052 24419
rect 11108 24363 11176 24419
rect 11232 24378 11300 24419
rect 11232 24363 11283 24378
rect 11356 24363 11396 24419
rect 10888 24326 11283 24363
rect 11335 24326 11396 24363
rect 10888 24295 11396 24326
rect 10888 24239 10928 24295
rect 10984 24239 11052 24295
rect 11108 24239 11176 24295
rect 11232 24270 11300 24295
rect 11232 24239 11283 24270
rect 11356 24239 11396 24295
rect 10888 24218 11283 24239
rect 11335 24218 11396 24239
rect 10888 24171 11396 24218
rect 10888 24115 10928 24171
rect 10984 24115 11052 24171
rect 11108 24115 11176 24171
rect 11232 24162 11300 24171
rect 11232 24115 11283 24162
rect 11356 24115 11396 24171
rect 10888 24110 11283 24115
rect 11335 24110 11396 24115
rect 10888 24054 11396 24110
rect 10888 24047 11283 24054
rect 11335 24047 11396 24054
rect 10888 23991 10928 24047
rect 10984 23991 11052 24047
rect 11108 23991 11176 24047
rect 11232 24002 11283 24047
rect 11232 23991 11300 24002
rect 11356 23991 11396 24047
rect 10888 23946 11396 23991
rect 10888 23923 11283 23946
rect 11335 23923 11396 23946
rect 10888 23867 10928 23923
rect 10984 23867 11052 23923
rect 11108 23867 11176 23923
rect 11232 23894 11283 23923
rect 11232 23867 11300 23894
rect 11356 23867 11396 23923
rect 10888 23838 11396 23867
rect 10888 23799 11283 23838
rect 11335 23799 11396 23838
rect 10888 23743 10928 23799
rect 10984 23743 11052 23799
rect 11108 23743 11176 23799
rect 11232 23786 11283 23799
rect 11232 23743 11300 23786
rect 11356 23743 11396 23799
rect 10888 23730 11396 23743
rect 10888 23678 11283 23730
rect 11335 23678 11396 23730
rect 10888 23622 11396 23678
rect 10888 23570 11283 23622
rect 11335 23570 11396 23622
rect 10888 23514 11396 23570
rect 10888 23462 11283 23514
rect 11335 23462 11396 23514
rect 10888 23451 11396 23462
rect 10888 23395 10928 23451
rect 10984 23395 11052 23451
rect 11108 23395 11176 23451
rect 11232 23406 11300 23451
rect 11232 23395 11283 23406
rect 11356 23395 11396 23451
rect 10888 23354 11283 23395
rect 11335 23354 11396 23395
rect 10888 23327 11396 23354
rect 10888 23271 10928 23327
rect 10984 23271 11052 23327
rect 11108 23271 11176 23327
rect 11232 23298 11300 23327
rect 11232 23271 11283 23298
rect 11356 23271 11396 23327
rect 10888 23246 11283 23271
rect 11335 23246 11396 23271
rect 10888 23203 11396 23246
rect 10888 23147 10928 23203
rect 10984 23147 11052 23203
rect 11108 23147 11176 23203
rect 11232 23190 11300 23203
rect 11232 23147 11283 23190
rect 11356 23147 11396 23203
rect 10888 23138 11283 23147
rect 11335 23138 11396 23147
rect 10888 23082 11396 23138
rect 10888 23079 11283 23082
rect 11335 23079 11396 23082
rect 10888 23023 10928 23079
rect 10984 23023 11052 23079
rect 11108 23023 11176 23079
rect 11232 23030 11283 23079
rect 11232 23023 11300 23030
rect 11356 23023 11396 23079
rect 10888 22974 11396 23023
rect 10888 22955 11283 22974
rect 11335 22955 11396 22974
rect 10888 22899 10928 22955
rect 10984 22899 11052 22955
rect 11108 22899 11176 22955
rect 11232 22922 11283 22955
rect 11232 22899 11300 22922
rect 11356 22899 11396 22955
rect 10888 22866 11396 22899
rect 10888 22831 11283 22866
rect 11335 22831 11396 22866
rect 10888 22775 10928 22831
rect 10984 22775 11052 22831
rect 11108 22775 11176 22831
rect 11232 22814 11283 22831
rect 11232 22775 11300 22814
rect 11356 22775 11396 22831
rect 10888 22758 11396 22775
rect 10888 22707 11283 22758
rect 11335 22707 11396 22758
rect 10888 22651 10928 22707
rect 10984 22651 11052 22707
rect 11108 22651 11176 22707
rect 11232 22706 11283 22707
rect 11232 22651 11300 22706
rect 11356 22651 11396 22707
rect 10888 22650 11396 22651
rect 10888 22598 11283 22650
rect 11335 22598 11396 22650
rect 10888 22583 11396 22598
rect 10888 22527 10928 22583
rect 10984 22527 11052 22583
rect 11108 22527 11176 22583
rect 11232 22542 11300 22583
rect 11232 22527 11283 22542
rect 11356 22527 11396 22583
rect 10888 22490 11283 22527
rect 11335 22490 11396 22527
rect 10888 22459 11396 22490
rect 10888 22403 10928 22459
rect 10984 22403 11052 22459
rect 11108 22403 11176 22459
rect 11232 22434 11300 22459
rect 11232 22403 11283 22434
rect 11356 22403 11396 22459
rect 10888 22382 11283 22403
rect 11335 22382 11396 22403
rect 10888 22335 11396 22382
rect 10888 22279 10928 22335
rect 10984 22279 11052 22335
rect 11108 22279 11176 22335
rect 11232 22326 11300 22335
rect 11232 22279 11283 22326
rect 11356 22279 11396 22335
rect 10888 22274 11283 22279
rect 11335 22274 11396 22279
rect 10888 22218 11396 22274
rect 10888 22211 11283 22218
rect 11335 22211 11396 22218
rect 10888 22155 10928 22211
rect 10984 22155 11052 22211
rect 11108 22155 11176 22211
rect 11232 22166 11283 22211
rect 11232 22155 11300 22166
rect 11356 22155 11396 22211
rect 10888 22110 11396 22155
rect 10888 22087 11283 22110
rect 11335 22087 11396 22110
rect 10888 22031 10928 22087
rect 10984 22031 11052 22087
rect 11108 22031 11176 22087
rect 11232 22058 11283 22087
rect 11232 22031 11300 22058
rect 11356 22031 11396 22087
rect 10888 22002 11396 22031
rect 10888 21963 11283 22002
rect 11335 21963 11396 22002
rect 10888 21907 10928 21963
rect 10984 21907 11052 21963
rect 11108 21907 11176 21963
rect 11232 21950 11283 21963
rect 11232 21907 11300 21950
rect 11356 21907 11396 21963
rect 10888 21894 11396 21907
rect 10888 21842 11283 21894
rect 11335 21842 11396 21894
rect 10888 21839 11396 21842
rect 10888 21783 10928 21839
rect 10984 21783 11052 21839
rect 11108 21783 11176 21839
rect 11232 21786 11300 21839
rect 11232 21783 11283 21786
rect 11356 21783 11396 21839
rect 10888 21734 11283 21783
rect 11335 21734 11396 21783
rect 10888 21715 11396 21734
rect 10888 21659 10928 21715
rect 10984 21659 11052 21715
rect 11108 21659 11176 21715
rect 11232 21678 11300 21715
rect 11232 21659 11283 21678
rect 11356 21659 11396 21715
rect 10888 21626 11283 21659
rect 11335 21626 11396 21659
rect 10888 21591 11396 21626
rect 10888 21535 10928 21591
rect 10984 21535 11052 21591
rect 11108 21535 11176 21591
rect 11232 21535 11300 21591
rect 11356 21535 11396 21591
rect 10888 21467 11396 21535
rect 10888 21411 10928 21467
rect 10984 21411 11052 21467
rect 11108 21411 11176 21467
rect 11232 21411 11300 21467
rect 11356 21411 11396 21467
rect 10888 21343 11396 21411
rect 10888 21287 10928 21343
rect 10984 21287 11052 21343
rect 11108 21287 11176 21343
rect 11232 21287 11300 21343
rect 11356 21287 11396 21343
rect 10888 21219 11396 21287
rect 10888 21163 10928 21219
rect 10984 21163 11052 21219
rect 11108 21163 11176 21219
rect 11232 21163 11300 21219
rect 11356 21163 11396 21219
rect 10888 21095 11396 21163
rect 10888 21039 10928 21095
rect 10984 21039 11052 21095
rect 11108 21039 11176 21095
rect 11232 21039 11300 21095
rect 11356 21039 11396 21095
rect 10888 20971 11396 21039
rect 10888 20915 10928 20971
rect 10984 20915 11052 20971
rect 11108 20915 11176 20971
rect 11232 20915 11300 20971
rect 11356 20915 11396 20971
rect 10888 20847 11396 20915
rect 10888 20791 10928 20847
rect 10984 20791 11052 20847
rect 11108 20791 11176 20847
rect 11232 20791 11300 20847
rect 11356 20791 11396 20847
rect 10888 20723 11396 20791
rect 10888 20667 10928 20723
rect 10984 20667 11052 20723
rect 11108 20667 11176 20723
rect 11232 20667 11300 20723
rect 11356 20667 11396 20723
rect 10888 20599 11396 20667
rect 10888 20577 10928 20599
rect 10984 20577 11052 20599
rect 11108 20577 11176 20599
rect 11232 20577 11300 20599
rect 11356 20577 11396 20599
rect 10888 20525 10900 20577
rect 10984 20543 11008 20577
rect 11108 20543 11116 20577
rect 10952 20525 11008 20543
rect 11060 20525 11116 20543
rect 11168 20543 11176 20577
rect 11276 20543 11300 20577
rect 11168 20525 11224 20543
rect 11276 20525 11332 20543
rect 11384 20525 11396 20577
rect 10888 20469 11396 20525
rect 10888 20417 10900 20469
rect 10952 20417 11008 20469
rect 11060 20417 11116 20469
rect 11168 20417 11224 20469
rect 11276 20417 11332 20469
rect 11384 20417 11396 20469
rect 10888 20361 11396 20417
rect 10888 20309 10900 20361
rect 10952 20309 11008 20361
rect 11060 20309 11116 20361
rect 11168 20309 11224 20361
rect 11276 20309 11332 20361
rect 11384 20309 11396 20361
rect 10888 20251 11396 20309
rect 10888 20195 10928 20251
rect 10984 20195 11052 20251
rect 11108 20195 11176 20251
rect 11232 20195 11300 20251
rect 11356 20195 11396 20251
rect 10888 20127 11396 20195
rect 10888 20071 10928 20127
rect 10984 20071 11052 20127
rect 11108 20071 11176 20127
rect 11232 20071 11300 20127
rect 11356 20071 11396 20127
rect 10888 20003 11396 20071
rect 10888 19947 10928 20003
rect 10984 19947 11052 20003
rect 11108 19947 11176 20003
rect 11232 19947 11300 20003
rect 11356 19947 11396 20003
rect 10888 19879 11396 19947
rect 10888 19823 10928 19879
rect 10984 19823 11052 19879
rect 11108 19823 11176 19879
rect 11232 19823 11300 19879
rect 11356 19823 11396 19879
rect 10888 19755 11396 19823
rect 10888 19699 10928 19755
rect 10984 19699 11052 19755
rect 11108 19699 11176 19755
rect 11232 19699 11300 19755
rect 11356 19699 11396 19755
rect 10888 19631 11396 19699
rect 10888 19584 10928 19631
rect 10984 19584 11052 19631
rect 11108 19584 11176 19631
rect 11232 19584 11300 19631
rect 11356 19584 11396 19631
rect 10888 19532 10900 19584
rect 10984 19575 11008 19584
rect 11108 19575 11116 19584
rect 10952 19532 11008 19575
rect 11060 19532 11116 19575
rect 11168 19575 11176 19584
rect 11276 19575 11300 19584
rect 11168 19532 11224 19575
rect 11276 19532 11332 19575
rect 11384 19532 11396 19584
rect 10888 19507 11396 19532
rect 10888 19476 10928 19507
rect 10984 19476 11052 19507
rect 11108 19476 11176 19507
rect 11232 19476 11300 19507
rect 11356 19476 11396 19507
rect 10888 19424 10900 19476
rect 10984 19451 11008 19476
rect 11108 19451 11116 19476
rect 10952 19424 11008 19451
rect 11060 19424 11116 19451
rect 11168 19451 11176 19476
rect 11276 19451 11300 19476
rect 11168 19424 11224 19451
rect 11276 19424 11332 19451
rect 11384 19424 11396 19476
rect 10888 19383 11396 19424
rect 10888 19327 10928 19383
rect 10984 19327 11052 19383
rect 11108 19327 11176 19383
rect 11232 19327 11300 19383
rect 11356 19327 11396 19383
rect 10888 19259 11396 19327
rect 10888 19203 10928 19259
rect 10984 19203 11052 19259
rect 11108 19203 11176 19259
rect 11232 19203 11300 19259
rect 11356 19203 11396 19259
rect 10888 19135 11396 19203
rect 10888 19079 10928 19135
rect 10984 19079 11052 19135
rect 11108 19079 11176 19135
rect 11232 19079 11300 19135
rect 11356 19079 11396 19135
rect 10888 19011 11396 19079
rect 10888 18955 10928 19011
rect 10984 18955 11052 19011
rect 11108 18955 11176 19011
rect 11232 18955 11300 19011
rect 11356 18955 11396 19011
rect 10888 18887 11396 18955
rect 10888 18831 10928 18887
rect 10984 18831 11052 18887
rect 11108 18831 11176 18887
rect 11232 18831 11300 18887
rect 11356 18831 11396 18887
rect 10888 18763 11396 18831
rect 10888 18712 10928 18763
rect 10984 18712 11052 18763
rect 11108 18712 11176 18763
rect 11232 18712 11300 18763
rect 11356 18712 11396 18763
rect 10888 18660 10900 18712
rect 10984 18707 11008 18712
rect 11108 18707 11116 18712
rect 10952 18660 11008 18707
rect 11060 18660 11116 18707
rect 11168 18707 11176 18712
rect 11276 18707 11300 18712
rect 11168 18660 11224 18707
rect 11276 18660 11332 18707
rect 11384 18660 11396 18712
rect 10888 18639 11396 18660
rect 10888 18604 10928 18639
rect 10984 18604 11052 18639
rect 11108 18604 11176 18639
rect 11232 18604 11300 18639
rect 11356 18604 11396 18639
rect 10888 18552 10900 18604
rect 10984 18583 11008 18604
rect 11108 18583 11116 18604
rect 10952 18552 11008 18583
rect 11060 18552 11116 18583
rect 11168 18583 11176 18604
rect 11276 18583 11300 18604
rect 11168 18552 11224 18583
rect 11276 18552 11332 18583
rect 11384 18552 11396 18604
rect 10888 18515 11396 18552
rect 10888 18459 10928 18515
rect 10984 18459 11052 18515
rect 11108 18459 11176 18515
rect 11232 18459 11300 18515
rect 11356 18459 11396 18515
rect 10888 18391 11396 18459
rect 10888 18335 10928 18391
rect 10984 18335 11052 18391
rect 11108 18335 11176 18391
rect 11232 18335 11300 18391
rect 11356 18335 11396 18391
rect 10888 18267 11396 18335
rect 10888 18211 10928 18267
rect 10984 18211 11052 18267
rect 11108 18211 11176 18267
rect 11232 18211 11300 18267
rect 11356 18211 11396 18267
rect 10888 18143 11396 18211
rect 10888 18087 10928 18143
rect 10984 18087 11052 18143
rect 11108 18087 11176 18143
rect 11232 18087 11300 18143
rect 11356 18087 11396 18143
rect 10888 18019 11396 18087
rect 10888 17963 10928 18019
rect 10984 17963 11052 18019
rect 11108 17963 11176 18019
rect 11232 17963 11300 18019
rect 11356 17963 11396 18019
rect 10888 17895 11396 17963
rect 10888 17840 10928 17895
rect 10984 17840 11052 17895
rect 11108 17840 11176 17895
rect 11232 17840 11300 17895
rect 11356 17840 11396 17895
rect 10888 17788 10900 17840
rect 10984 17839 11008 17840
rect 11108 17839 11116 17840
rect 10952 17788 11008 17839
rect 11060 17788 11116 17839
rect 11168 17839 11176 17840
rect 11276 17839 11300 17840
rect 11168 17788 11224 17839
rect 11276 17788 11332 17839
rect 11384 17788 11396 17840
rect 10888 17771 11396 17788
rect 10888 17732 10928 17771
rect 10984 17732 11052 17771
rect 11108 17732 11176 17771
rect 11232 17732 11300 17771
rect 11356 17732 11396 17771
rect 10888 17680 10900 17732
rect 10984 17715 11008 17732
rect 11108 17715 11116 17732
rect 10952 17680 11008 17715
rect 11060 17680 11116 17715
rect 11168 17715 11176 17732
rect 11276 17715 11300 17732
rect 11168 17680 11224 17715
rect 11276 17680 11332 17715
rect 11384 17680 11396 17732
rect 10888 17647 11396 17680
rect 10888 17591 10928 17647
rect 10984 17591 11052 17647
rect 11108 17591 11176 17647
rect 11232 17591 11300 17647
rect 11356 17591 11396 17647
rect 10888 17523 11396 17591
rect 10888 17467 10928 17523
rect 10984 17467 11052 17523
rect 11108 17467 11176 17523
rect 11232 17467 11300 17523
rect 11356 17467 11396 17523
rect 10888 17399 11396 17467
rect 10888 17343 10928 17399
rect 10984 17343 11052 17399
rect 11108 17343 11176 17399
rect 11232 17343 11300 17399
rect 11356 17343 11396 17399
rect 10888 17051 11396 17343
rect 10888 16995 10928 17051
rect 10984 16995 11052 17051
rect 11108 16995 11176 17051
rect 11232 16995 11300 17051
rect 11356 16995 11396 17051
rect 10888 16968 11396 16995
rect 10888 16916 10900 16968
rect 10952 16927 11008 16968
rect 11060 16927 11116 16968
rect 10984 16916 11008 16927
rect 11108 16916 11116 16927
rect 11168 16927 11224 16968
rect 11276 16927 11332 16968
rect 11168 16916 11176 16927
rect 11276 16916 11300 16927
rect 11384 16916 11396 16968
rect 10888 16871 10928 16916
rect 10984 16871 11052 16916
rect 11108 16871 11176 16916
rect 11232 16871 11300 16916
rect 11356 16871 11396 16916
rect 10888 16860 11396 16871
rect 10888 16808 10900 16860
rect 10952 16808 11008 16860
rect 11060 16808 11116 16860
rect 11168 16808 11224 16860
rect 11276 16808 11332 16860
rect 11384 16808 11396 16860
rect 10888 16803 11396 16808
rect 10888 16747 10928 16803
rect 10984 16747 11052 16803
rect 11108 16747 11176 16803
rect 11232 16747 11300 16803
rect 11356 16747 11396 16803
rect 10888 16679 11396 16747
rect 10888 16623 10928 16679
rect 10984 16623 11052 16679
rect 11108 16623 11176 16679
rect 11232 16623 11300 16679
rect 11356 16623 11396 16679
rect 10888 16555 11396 16623
rect 10888 16499 10928 16555
rect 10984 16499 11052 16555
rect 11108 16499 11176 16555
rect 11232 16499 11300 16555
rect 11356 16499 11396 16555
rect 10888 16431 11396 16499
rect 10888 16375 10928 16431
rect 10984 16375 11052 16431
rect 11108 16375 11176 16431
rect 11232 16375 11300 16431
rect 11356 16375 11396 16431
rect 10888 16307 11396 16375
rect 10888 16251 10928 16307
rect 10984 16251 11052 16307
rect 11108 16251 11176 16307
rect 11232 16251 11300 16307
rect 11356 16251 11396 16307
rect 10888 16183 11396 16251
rect 10888 16127 10928 16183
rect 10984 16127 11052 16183
rect 11108 16127 11176 16183
rect 11232 16127 11300 16183
rect 11356 16127 11396 16183
rect 10888 16083 11396 16127
rect 10888 16031 10900 16083
rect 10952 16059 11008 16083
rect 11060 16059 11116 16083
rect 10984 16031 11008 16059
rect 11108 16031 11116 16059
rect 11168 16059 11224 16083
rect 11276 16059 11332 16083
rect 11168 16031 11176 16059
rect 11276 16031 11300 16059
rect 11384 16031 11396 16083
rect 10888 16003 10928 16031
rect 10984 16003 11052 16031
rect 11108 16003 11176 16031
rect 11232 16003 11300 16031
rect 11356 16003 11396 16031
rect 10888 15975 11396 16003
rect 10888 15923 10900 15975
rect 10952 15935 11008 15975
rect 11060 15935 11116 15975
rect 10984 15923 11008 15935
rect 11108 15923 11116 15935
rect 11168 15935 11224 15975
rect 11276 15935 11332 15975
rect 11168 15923 11176 15935
rect 11276 15923 11300 15935
rect 11384 15923 11396 15975
rect 10888 15879 10928 15923
rect 10984 15879 11052 15923
rect 11108 15879 11176 15923
rect 11232 15879 11300 15923
rect 11356 15879 11396 15923
rect 10888 15867 11396 15879
rect 10888 15815 10900 15867
rect 10952 15815 11008 15867
rect 11060 15815 11116 15867
rect 11168 15815 11224 15867
rect 11276 15815 11332 15867
rect 11384 15815 11396 15867
rect 10888 15811 11396 15815
rect 10888 15762 10928 15811
rect 9084 15755 9094 15762
rect 8646 15687 9094 15755
rect 8646 15631 8656 15687
rect 8712 15631 8780 15687
rect 8836 15631 8904 15687
rect 8960 15631 9028 15687
rect 9084 15631 9094 15687
rect 8646 15563 9094 15631
rect 8646 15507 8656 15563
rect 8712 15507 8780 15563
rect 8836 15507 8904 15563
rect 8960 15507 9028 15563
rect 9084 15507 9094 15563
rect 8646 15439 9094 15507
rect 8646 15383 8656 15439
rect 8712 15383 8780 15439
rect 8836 15383 8904 15439
rect 8960 15383 9028 15439
rect 9084 15383 9094 15439
rect 8646 15315 9094 15383
rect 8646 15259 8656 15315
rect 8712 15259 8780 15315
rect 8836 15259 8904 15315
rect 8960 15259 9028 15315
rect 9084 15259 9094 15315
rect 8646 15191 9094 15259
rect 8646 15135 8656 15191
rect 8712 15135 8780 15191
rect 8836 15135 8904 15191
rect 8960 15135 9028 15191
rect 9084 15135 9094 15191
rect 8646 15067 9094 15135
rect 8646 15011 8656 15067
rect 8712 15011 8780 15067
rect 8836 15011 8904 15067
rect 8960 15011 9028 15067
rect 9084 15011 9094 15067
rect 8646 14943 9094 15011
rect 8646 14887 8656 14943
rect 8712 14887 8780 14943
rect 8836 14887 8904 14943
rect 8960 14887 9028 14943
rect 9084 14887 9094 14943
rect 8646 14819 9094 14887
rect 8646 14763 8656 14819
rect 8712 14763 8780 14819
rect 8836 14763 8904 14819
rect 8960 14763 9028 14819
rect 9084 14763 9094 14819
rect 8646 14695 9094 14763
rect 8646 14639 8656 14695
rect 8712 14639 8780 14695
rect 8836 14639 8904 14695
rect 8960 14639 9028 14695
rect 9084 14639 9094 14695
rect 8646 14571 9094 14639
rect 8646 14515 8656 14571
rect 8712 14515 8780 14571
rect 8836 14515 8904 14571
rect 8960 14515 9028 14571
rect 9084 14515 9094 14571
rect 8646 14447 9094 14515
rect 8646 14391 8656 14447
rect 8712 14391 8780 14447
rect 8836 14391 8904 14447
rect 8960 14391 9028 14447
rect 9084 14391 9094 14447
rect 8646 14323 9094 14391
rect 8646 14267 8656 14323
rect 8712 14267 8780 14323
rect 8836 14267 8904 14323
rect 8960 14267 9028 14323
rect 9084 14267 9094 14323
rect 8646 14199 9094 14267
rect 8646 14143 8656 14199
rect 8712 14143 8780 14199
rect 8836 14143 8904 14199
rect 8960 14143 9028 14199
rect 9084 14143 9094 14199
rect 8646 14133 9094 14143
rect 10918 15755 10928 15762
rect 10984 15755 11052 15811
rect 11108 15755 11176 15811
rect 11232 15755 11300 15811
rect 11356 15762 11396 15811
rect 12024 56922 12532 56975
rect 12024 56866 12064 56922
rect 12120 56866 12188 56922
rect 12244 56866 12312 56922
rect 12368 56866 12436 56922
rect 12492 56866 12532 56922
rect 12024 56798 12532 56866
rect 12024 56742 12064 56798
rect 12120 56742 12188 56798
rect 12244 56742 12312 56798
rect 12368 56742 12436 56798
rect 12492 56742 12532 56798
rect 12024 56711 12532 56742
rect 12024 56659 12036 56711
rect 12088 56674 12144 56711
rect 12196 56674 12252 56711
rect 12120 56659 12144 56674
rect 12244 56659 12252 56674
rect 12304 56674 12360 56711
rect 12412 56674 12468 56711
rect 12304 56659 12312 56674
rect 12412 56659 12436 56674
rect 12520 56659 12532 56711
rect 12024 56618 12064 56659
rect 12120 56618 12188 56659
rect 12244 56618 12312 56659
rect 12368 56618 12436 56659
rect 12492 56618 12532 56659
rect 12024 56603 12532 56618
rect 12024 56551 12036 56603
rect 12088 56551 12144 56603
rect 12196 56551 12252 56603
rect 12304 56551 12360 56603
rect 12412 56551 12468 56603
rect 12520 56551 12532 56603
rect 12024 56550 12532 56551
rect 12024 56495 12064 56550
rect 12120 56495 12188 56550
rect 12244 56495 12312 56550
rect 12368 56495 12436 56550
rect 12492 56495 12532 56550
rect 12024 56443 12036 56495
rect 12120 56494 12144 56495
rect 12244 56494 12252 56495
rect 12088 56443 12144 56494
rect 12196 56443 12252 56494
rect 12304 56494 12312 56495
rect 12412 56494 12436 56495
rect 12304 56443 12360 56494
rect 12412 56443 12468 56494
rect 12520 56443 12532 56495
rect 12024 56426 12532 56443
rect 12024 56370 12064 56426
rect 12120 56370 12188 56426
rect 12244 56370 12312 56426
rect 12368 56370 12436 56426
rect 12492 56370 12532 56426
rect 12024 56302 12532 56370
rect 12024 56246 12064 56302
rect 12120 56246 12188 56302
rect 12244 56246 12312 56302
rect 12368 56246 12436 56302
rect 12492 56246 12532 56302
rect 12024 56178 12532 56246
rect 12024 56122 12064 56178
rect 12120 56122 12188 56178
rect 12244 56122 12312 56178
rect 12368 56122 12436 56178
rect 12492 56122 12532 56178
rect 12024 56054 12532 56122
rect 12024 55998 12064 56054
rect 12120 55998 12188 56054
rect 12244 55998 12312 56054
rect 12368 55998 12436 56054
rect 12492 55998 12532 56054
rect 12024 55930 12532 55998
rect 12024 55874 12064 55930
rect 12120 55874 12188 55930
rect 12244 55874 12312 55930
rect 12368 55874 12436 55930
rect 12492 55874 12532 55930
rect 12024 55806 12532 55874
rect 12024 55750 12064 55806
rect 12120 55750 12188 55806
rect 12244 55750 12312 55806
rect 12368 55750 12436 55806
rect 12492 55750 12532 55806
rect 12024 53845 12532 55750
rect 12024 53789 12064 53845
rect 12120 53789 12188 53845
rect 12244 53789 12312 53845
rect 12368 53789 12436 53845
rect 12492 53789 12532 53845
rect 12024 53721 12532 53789
rect 12024 53665 12064 53721
rect 12120 53665 12188 53721
rect 12244 53665 12312 53721
rect 12368 53665 12436 53721
rect 12492 53665 12532 53721
rect 12024 53597 12532 53665
rect 12024 53541 12064 53597
rect 12120 53541 12188 53597
rect 12244 53541 12312 53597
rect 12368 53541 12436 53597
rect 12492 53541 12532 53597
rect 12024 53473 12532 53541
rect 12024 53417 12064 53473
rect 12120 53417 12188 53473
rect 12244 53417 12312 53473
rect 12368 53417 12436 53473
rect 12492 53417 12532 53473
rect 12024 53349 12532 53417
rect 12024 53293 12064 53349
rect 12120 53293 12188 53349
rect 12244 53293 12312 53349
rect 12368 53293 12436 53349
rect 12492 53293 12532 53349
rect 12024 53225 12532 53293
rect 12024 53169 12064 53225
rect 12120 53169 12188 53225
rect 12244 53169 12312 53225
rect 12368 53169 12436 53225
rect 12492 53169 12532 53225
rect 12024 53101 12532 53169
rect 12024 53045 12064 53101
rect 12120 53045 12188 53101
rect 12244 53045 12312 53101
rect 12368 53045 12436 53101
rect 12492 53045 12532 53101
rect 12024 52996 12066 53045
rect 12118 52996 12190 53045
rect 12242 52996 12314 53045
rect 12366 52996 12438 53045
rect 12490 52996 12532 53045
rect 12024 52977 12532 52996
rect 12024 52921 12064 52977
rect 12120 52921 12188 52977
rect 12244 52921 12312 52977
rect 12368 52921 12436 52977
rect 12492 52921 12532 52977
rect 12024 52872 12066 52921
rect 12118 52872 12190 52921
rect 12242 52872 12314 52921
rect 12366 52872 12438 52921
rect 12490 52872 12532 52921
rect 12024 52853 12532 52872
rect 12024 52797 12064 52853
rect 12120 52797 12188 52853
rect 12244 52797 12312 52853
rect 12368 52797 12436 52853
rect 12492 52797 12532 52853
rect 12024 52748 12066 52797
rect 12118 52748 12190 52797
rect 12242 52748 12314 52797
rect 12366 52748 12438 52797
rect 12490 52748 12532 52797
rect 12024 52729 12532 52748
rect 12024 52673 12064 52729
rect 12120 52673 12188 52729
rect 12244 52673 12312 52729
rect 12368 52673 12436 52729
rect 12492 52673 12532 52729
rect 12024 52624 12066 52673
rect 12118 52624 12190 52673
rect 12242 52624 12314 52673
rect 12366 52624 12438 52673
rect 12490 52624 12532 52673
rect 12024 52605 12532 52624
rect 12024 52549 12064 52605
rect 12120 52549 12188 52605
rect 12244 52549 12312 52605
rect 12368 52549 12436 52605
rect 12492 52549 12532 52605
rect 12024 52500 12066 52549
rect 12118 52500 12190 52549
rect 12242 52500 12314 52549
rect 12366 52500 12438 52549
rect 12490 52500 12532 52549
rect 12024 49100 12532 52500
rect 12024 49048 12066 49100
rect 12118 49048 12190 49100
rect 12242 49048 12314 49100
rect 12366 49048 12438 49100
rect 12490 49048 12532 49100
rect 12024 49045 12532 49048
rect 12024 48989 12064 49045
rect 12120 48989 12188 49045
rect 12244 48989 12312 49045
rect 12368 48989 12436 49045
rect 12492 48989 12532 49045
rect 12024 48976 12532 48989
rect 12024 48924 12066 48976
rect 12118 48924 12190 48976
rect 12242 48924 12314 48976
rect 12366 48924 12438 48976
rect 12490 48924 12532 48976
rect 12024 48921 12532 48924
rect 12024 48865 12064 48921
rect 12120 48865 12188 48921
rect 12244 48865 12312 48921
rect 12368 48865 12436 48921
rect 12492 48865 12532 48921
rect 12024 48852 12532 48865
rect 12024 48800 12066 48852
rect 12118 48800 12190 48852
rect 12242 48800 12314 48852
rect 12366 48800 12438 48852
rect 12490 48800 12532 48852
rect 12024 48797 12532 48800
rect 12024 48741 12064 48797
rect 12120 48741 12188 48797
rect 12244 48741 12312 48797
rect 12368 48741 12436 48797
rect 12492 48741 12532 48797
rect 12024 48728 12532 48741
rect 12024 48676 12066 48728
rect 12118 48676 12190 48728
rect 12242 48676 12314 48728
rect 12366 48676 12438 48728
rect 12490 48676 12532 48728
rect 12024 48673 12532 48676
rect 12024 48617 12064 48673
rect 12120 48617 12188 48673
rect 12244 48617 12312 48673
rect 12368 48617 12436 48673
rect 12492 48617 12532 48673
rect 12024 48604 12532 48617
rect 12024 48552 12066 48604
rect 12118 48552 12190 48604
rect 12242 48552 12314 48604
rect 12366 48552 12438 48604
rect 12490 48552 12532 48604
rect 12024 48549 12532 48552
rect 12024 48493 12064 48549
rect 12120 48493 12188 48549
rect 12244 48493 12312 48549
rect 12368 48493 12436 48549
rect 12492 48493 12532 48549
rect 12024 48425 12532 48493
rect 12024 48369 12064 48425
rect 12120 48369 12188 48425
rect 12244 48369 12312 48425
rect 12368 48369 12436 48425
rect 12492 48369 12532 48425
rect 12024 48301 12532 48369
rect 12024 48245 12064 48301
rect 12120 48245 12188 48301
rect 12244 48245 12312 48301
rect 12368 48245 12436 48301
rect 12492 48245 12532 48301
rect 12024 48177 12532 48245
rect 12024 48121 12064 48177
rect 12120 48121 12188 48177
rect 12244 48121 12312 48177
rect 12368 48121 12436 48177
rect 12492 48121 12532 48177
rect 12024 48053 12532 48121
rect 12024 47997 12064 48053
rect 12120 47997 12188 48053
rect 12244 47997 12312 48053
rect 12368 47997 12436 48053
rect 12492 47997 12532 48053
rect 12024 47929 12532 47997
rect 12024 47873 12064 47929
rect 12120 47873 12188 47929
rect 12244 47873 12312 47929
rect 12368 47873 12436 47929
rect 12492 47873 12532 47929
rect 12024 47805 12532 47873
rect 12024 47749 12064 47805
rect 12120 47749 12188 47805
rect 12244 47749 12312 47805
rect 12368 47749 12436 47805
rect 12492 47749 12532 47805
rect 12024 45845 12532 47749
rect 12024 45789 12064 45845
rect 12120 45789 12188 45845
rect 12244 45789 12312 45845
rect 12368 45789 12436 45845
rect 12492 45789 12532 45845
rect 12024 45721 12532 45789
rect 12024 45665 12064 45721
rect 12120 45665 12188 45721
rect 12244 45665 12312 45721
rect 12368 45665 12436 45721
rect 12492 45665 12532 45721
rect 12024 45597 12532 45665
rect 12024 45541 12064 45597
rect 12120 45541 12188 45597
rect 12244 45541 12312 45597
rect 12368 45541 12436 45597
rect 12492 45541 12532 45597
rect 12024 45473 12532 45541
rect 12024 45417 12064 45473
rect 12120 45417 12188 45473
rect 12244 45417 12312 45473
rect 12368 45417 12436 45473
rect 12492 45417 12532 45473
rect 12024 45349 12532 45417
rect 12024 45293 12064 45349
rect 12120 45293 12188 45349
rect 12244 45293 12312 45349
rect 12368 45293 12436 45349
rect 12492 45293 12532 45349
rect 12024 45225 12532 45293
rect 12024 45169 12064 45225
rect 12120 45169 12188 45225
rect 12244 45169 12312 45225
rect 12368 45169 12436 45225
rect 12492 45169 12532 45225
rect 12024 45152 12532 45169
rect 12024 45101 12066 45152
rect 12118 45101 12190 45152
rect 12242 45101 12314 45152
rect 12366 45101 12438 45152
rect 12490 45101 12532 45152
rect 12024 45045 12064 45101
rect 12120 45045 12188 45101
rect 12244 45045 12312 45101
rect 12368 45045 12436 45101
rect 12492 45045 12532 45101
rect 12024 45028 12532 45045
rect 12024 44977 12066 45028
rect 12118 44977 12190 45028
rect 12242 44977 12314 45028
rect 12366 44977 12438 45028
rect 12490 44977 12532 45028
rect 12024 44921 12064 44977
rect 12120 44921 12188 44977
rect 12244 44921 12312 44977
rect 12368 44921 12436 44977
rect 12492 44921 12532 44977
rect 12024 44904 12532 44921
rect 12024 44853 12066 44904
rect 12118 44853 12190 44904
rect 12242 44853 12314 44904
rect 12366 44853 12438 44904
rect 12490 44853 12532 44904
rect 12024 44797 12064 44853
rect 12120 44797 12188 44853
rect 12244 44797 12312 44853
rect 12368 44797 12436 44853
rect 12492 44797 12532 44853
rect 12024 44780 12532 44797
rect 12024 44729 12066 44780
rect 12118 44729 12190 44780
rect 12242 44729 12314 44780
rect 12366 44729 12438 44780
rect 12490 44729 12532 44780
rect 12024 44673 12064 44729
rect 12120 44673 12188 44729
rect 12244 44673 12312 44729
rect 12368 44673 12436 44729
rect 12492 44673 12532 44729
rect 12024 44656 12532 44673
rect 12024 44605 12066 44656
rect 12118 44605 12190 44656
rect 12242 44605 12314 44656
rect 12366 44605 12438 44656
rect 12490 44605 12532 44656
rect 12024 44549 12064 44605
rect 12120 44549 12188 44605
rect 12244 44549 12312 44605
rect 12368 44549 12436 44605
rect 12492 44549 12532 44605
rect 12024 41204 12532 44549
rect 12024 41152 12066 41204
rect 12118 41152 12190 41204
rect 12242 41152 12314 41204
rect 12366 41152 12438 41204
rect 12490 41152 12532 41204
rect 12024 41080 12532 41152
rect 12024 41028 12066 41080
rect 12118 41028 12190 41080
rect 12242 41028 12314 41080
rect 12366 41028 12438 41080
rect 12490 41028 12532 41080
rect 12024 40956 12532 41028
rect 12024 40904 12066 40956
rect 12118 40904 12190 40956
rect 12242 40904 12314 40956
rect 12366 40904 12438 40956
rect 12490 40904 12532 40956
rect 12024 40832 12532 40904
rect 12024 40780 12066 40832
rect 12118 40780 12190 40832
rect 12242 40780 12314 40832
rect 12366 40780 12438 40832
rect 12490 40780 12532 40832
rect 12024 40708 12532 40780
rect 12024 40656 12066 40708
rect 12118 40656 12190 40708
rect 12242 40656 12314 40708
rect 12366 40656 12438 40708
rect 12490 40656 12532 40708
rect 12024 37256 12532 40656
rect 12024 37204 12066 37256
rect 12118 37204 12190 37256
rect 12242 37204 12314 37256
rect 12366 37204 12438 37256
rect 12490 37204 12532 37256
rect 12024 37132 12532 37204
rect 12024 37080 12066 37132
rect 12118 37080 12190 37132
rect 12242 37080 12314 37132
rect 12366 37080 12438 37132
rect 12490 37080 12532 37132
rect 12024 37008 12532 37080
rect 12024 36956 12066 37008
rect 12118 36956 12190 37008
rect 12242 36956 12314 37008
rect 12366 36956 12438 37008
rect 12490 36956 12532 37008
rect 12024 36884 12532 36956
rect 12024 36832 12066 36884
rect 12118 36832 12190 36884
rect 12242 36832 12314 36884
rect 12366 36832 12438 36884
rect 12490 36832 12532 36884
rect 12024 36760 12532 36832
rect 12024 36708 12066 36760
rect 12118 36708 12190 36760
rect 12242 36708 12314 36760
rect 12366 36708 12438 36760
rect 12490 36708 12532 36760
rect 12024 36251 12532 36708
rect 12024 36195 12064 36251
rect 12120 36195 12188 36251
rect 12244 36195 12312 36251
rect 12368 36195 12436 36251
rect 12492 36195 12532 36251
rect 12024 36127 12532 36195
rect 12024 36071 12064 36127
rect 12120 36071 12188 36127
rect 12244 36071 12312 36127
rect 12368 36071 12436 36127
rect 12492 36071 12532 36127
rect 12024 36003 12532 36071
rect 12024 35947 12064 36003
rect 12120 35947 12188 36003
rect 12244 35947 12312 36003
rect 12368 35947 12436 36003
rect 12492 35947 12532 36003
rect 12024 35879 12532 35947
rect 12024 35823 12064 35879
rect 12120 35823 12188 35879
rect 12244 35823 12312 35879
rect 12368 35823 12436 35879
rect 12492 35823 12532 35879
rect 12024 35755 12532 35823
rect 12024 35699 12064 35755
rect 12120 35699 12188 35755
rect 12244 35699 12312 35755
rect 12368 35699 12436 35755
rect 12492 35699 12532 35755
rect 12024 35631 12532 35699
rect 12024 35575 12064 35631
rect 12120 35575 12188 35631
rect 12244 35575 12312 35631
rect 12368 35575 12436 35631
rect 12492 35575 12532 35631
rect 12024 35507 12532 35575
rect 12024 35451 12064 35507
rect 12120 35451 12188 35507
rect 12244 35451 12312 35507
rect 12368 35451 12436 35507
rect 12492 35451 12532 35507
rect 12024 35383 12532 35451
rect 12024 35327 12064 35383
rect 12120 35327 12188 35383
rect 12244 35327 12312 35383
rect 12368 35327 12436 35383
rect 12492 35327 12532 35383
rect 12024 35259 12532 35327
rect 12024 35203 12064 35259
rect 12120 35203 12188 35259
rect 12244 35203 12312 35259
rect 12368 35203 12436 35259
rect 12492 35203 12532 35259
rect 12024 35135 12532 35203
rect 12024 35079 12064 35135
rect 12120 35079 12188 35135
rect 12244 35079 12312 35135
rect 12368 35079 12436 35135
rect 12492 35079 12532 35135
rect 12024 35011 12532 35079
rect 12024 34955 12064 35011
rect 12120 34955 12188 35011
rect 12244 34955 12312 35011
rect 12368 34955 12436 35011
rect 12492 34955 12532 35011
rect 12024 34887 12532 34955
rect 12024 34831 12064 34887
rect 12120 34831 12188 34887
rect 12244 34831 12312 34887
rect 12368 34831 12436 34887
rect 12492 34831 12532 34887
rect 12024 34763 12532 34831
rect 12024 34707 12064 34763
rect 12120 34707 12188 34763
rect 12244 34707 12312 34763
rect 12368 34707 12436 34763
rect 12492 34707 12532 34763
rect 12024 34639 12532 34707
rect 12024 34583 12064 34639
rect 12120 34583 12188 34639
rect 12244 34583 12312 34639
rect 12368 34583 12436 34639
rect 12492 34583 12532 34639
rect 12024 34515 12532 34583
rect 12024 34459 12064 34515
rect 12120 34459 12188 34515
rect 12244 34459 12312 34515
rect 12368 34459 12436 34515
rect 12492 34459 12532 34515
rect 12024 34391 12532 34459
rect 12024 34335 12064 34391
rect 12120 34335 12188 34391
rect 12244 34335 12312 34391
rect 12368 34335 12436 34391
rect 12492 34335 12532 34391
rect 12024 34267 12532 34335
rect 12024 34211 12064 34267
rect 12120 34211 12188 34267
rect 12244 34211 12312 34267
rect 12368 34211 12436 34267
rect 12492 34211 12532 34267
rect 12024 34143 12532 34211
rect 12024 34087 12064 34143
rect 12120 34087 12188 34143
rect 12244 34087 12312 34143
rect 12368 34087 12436 34143
rect 12492 34087 12532 34143
rect 12024 34019 12532 34087
rect 12024 33963 12064 34019
rect 12120 33963 12188 34019
rect 12244 33963 12312 34019
rect 12368 33963 12436 34019
rect 12492 33963 12532 34019
rect 12024 33895 12532 33963
rect 12024 33839 12064 33895
rect 12120 33839 12188 33895
rect 12244 33839 12312 33895
rect 12368 33839 12436 33895
rect 12492 33839 12532 33895
rect 12024 33771 12532 33839
rect 12024 33715 12064 33771
rect 12120 33715 12188 33771
rect 12244 33715 12312 33771
rect 12368 33715 12436 33771
rect 12492 33715 12532 33771
rect 12024 33647 12532 33715
rect 12024 33591 12064 33647
rect 12120 33591 12188 33647
rect 12244 33591 12312 33647
rect 12368 33591 12436 33647
rect 12492 33591 12532 33647
rect 12024 33523 12532 33591
rect 12024 33467 12064 33523
rect 12120 33467 12188 33523
rect 12244 33467 12312 33523
rect 12368 33467 12436 33523
rect 12492 33467 12532 33523
rect 12024 33399 12532 33467
rect 12024 33343 12064 33399
rect 12120 33343 12188 33399
rect 12244 33343 12312 33399
rect 12368 33343 12436 33399
rect 12492 33343 12532 33399
rect 12024 33308 12532 33343
rect 12024 33256 12066 33308
rect 12118 33256 12190 33308
rect 12242 33256 12314 33308
rect 12366 33256 12438 33308
rect 12490 33256 12532 33308
rect 12024 33184 12532 33256
rect 12024 33132 12066 33184
rect 12118 33132 12190 33184
rect 12242 33132 12314 33184
rect 12366 33132 12438 33184
rect 12490 33132 12532 33184
rect 12024 33060 12532 33132
rect 12024 33008 12066 33060
rect 12118 33008 12190 33060
rect 12242 33008 12314 33060
rect 12366 33008 12438 33060
rect 12490 33008 12532 33060
rect 12024 32936 12532 33008
rect 12024 32884 12066 32936
rect 12118 32884 12190 32936
rect 12242 32884 12314 32936
rect 12366 32884 12438 32936
rect 12490 32884 12532 32936
rect 12024 32812 12532 32884
rect 12024 32760 12066 32812
rect 12118 32760 12190 32812
rect 12242 32760 12314 32812
rect 12366 32760 12438 32812
rect 12490 32760 12532 32812
rect 12024 29360 12532 32760
rect 12024 29308 12066 29360
rect 12118 29308 12190 29360
rect 12242 29308 12314 29360
rect 12366 29308 12438 29360
rect 12490 29308 12532 29360
rect 12024 29236 12532 29308
rect 12024 29184 12066 29236
rect 12118 29184 12190 29236
rect 12242 29184 12314 29236
rect 12366 29184 12438 29236
rect 12490 29184 12532 29236
rect 12024 29112 12532 29184
rect 12024 29060 12066 29112
rect 12118 29060 12190 29112
rect 12242 29060 12314 29112
rect 12366 29060 12438 29112
rect 12490 29060 12532 29112
rect 12024 28988 12532 29060
rect 12024 28936 12066 28988
rect 12118 28936 12190 28988
rect 12242 28936 12314 28988
rect 12366 28936 12438 28988
rect 12490 28936 12532 28988
rect 12024 28864 12532 28936
rect 12024 28812 12066 28864
rect 12118 28812 12190 28864
rect 12242 28812 12314 28864
rect 12366 28812 12438 28864
rect 12490 28812 12532 28864
rect 12024 28245 12532 28812
rect 12024 28189 12064 28245
rect 12120 28189 12188 28245
rect 12244 28189 12312 28245
rect 12368 28189 12436 28245
rect 12492 28189 12532 28245
rect 12024 28121 12532 28189
rect 12024 28065 12064 28121
rect 12120 28065 12188 28121
rect 12244 28065 12312 28121
rect 12368 28065 12436 28121
rect 12492 28065 12532 28121
rect 12024 27997 12532 28065
rect 12024 27941 12064 27997
rect 12120 27941 12188 27997
rect 12244 27941 12312 27997
rect 12368 27941 12436 27997
rect 12492 27941 12532 27997
rect 12024 27873 12532 27941
rect 12024 27817 12064 27873
rect 12120 27817 12188 27873
rect 12244 27817 12312 27873
rect 12368 27817 12436 27873
rect 12492 27817 12532 27873
rect 12024 27749 12532 27817
rect 12024 27693 12064 27749
rect 12120 27693 12188 27749
rect 12244 27693 12312 27749
rect 12368 27693 12436 27749
rect 12492 27693 12532 27749
rect 12024 27625 12532 27693
rect 12024 27569 12064 27625
rect 12120 27569 12188 27625
rect 12244 27569 12312 27625
rect 12368 27569 12436 27625
rect 12492 27569 12532 27625
rect 12024 27501 12532 27569
rect 12024 27445 12064 27501
rect 12120 27445 12188 27501
rect 12244 27445 12312 27501
rect 12368 27445 12436 27501
rect 12492 27445 12532 27501
rect 12024 27377 12532 27445
rect 12024 27321 12064 27377
rect 12120 27321 12188 27377
rect 12244 27321 12312 27377
rect 12368 27321 12436 27377
rect 12492 27321 12532 27377
rect 12024 27253 12532 27321
rect 12024 27197 12064 27253
rect 12120 27197 12188 27253
rect 12244 27197 12312 27253
rect 12368 27197 12436 27253
rect 12492 27197 12532 27253
rect 12024 27129 12532 27197
rect 12024 27073 12064 27129
rect 12120 27073 12188 27129
rect 12244 27073 12312 27129
rect 12368 27073 12436 27129
rect 12492 27073 12532 27129
rect 12024 27005 12532 27073
rect 12024 26949 12064 27005
rect 12120 26949 12188 27005
rect 12244 26949 12312 27005
rect 12368 26949 12436 27005
rect 12492 26949 12532 27005
rect 12024 25412 12532 26949
rect 12024 25360 12066 25412
rect 12118 25360 12190 25412
rect 12242 25360 12314 25412
rect 12366 25360 12438 25412
rect 12490 25360 12532 25412
rect 12024 25288 12532 25360
rect 12024 25236 12066 25288
rect 12118 25236 12190 25288
rect 12242 25236 12314 25288
rect 12366 25236 12438 25288
rect 12490 25236 12532 25288
rect 12024 25164 12532 25236
rect 12024 25112 12066 25164
rect 12118 25112 12190 25164
rect 12242 25112 12314 25164
rect 12366 25112 12438 25164
rect 12490 25112 12532 25164
rect 12024 25040 12532 25112
rect 12024 24988 12066 25040
rect 12118 24988 12190 25040
rect 12242 24988 12314 25040
rect 12366 24988 12438 25040
rect 12490 24988 12532 25040
rect 12024 24916 12532 24988
rect 12024 24864 12066 24916
rect 12118 24864 12190 24916
rect 12242 24864 12314 24916
rect 12366 24864 12438 24916
rect 12490 24864 12532 24916
rect 12024 21469 12532 24864
rect 12024 21417 12036 21469
rect 12088 21417 12144 21469
rect 12196 21417 12252 21469
rect 12304 21417 12360 21469
rect 12412 21417 12468 21469
rect 12520 21417 12532 21469
rect 12024 21361 12532 21417
rect 12024 21309 12036 21361
rect 12088 21309 12144 21361
rect 12196 21309 12252 21361
rect 12304 21309 12360 21361
rect 12412 21309 12468 21361
rect 12520 21309 12532 21361
rect 12024 21253 12532 21309
rect 12024 21201 12036 21253
rect 12088 21201 12144 21253
rect 12196 21201 12252 21253
rect 12304 21201 12360 21253
rect 12412 21201 12468 21253
rect 12520 21201 12532 21253
rect 12024 15762 12532 21201
rect 12592 55445 13100 56975
rect 12592 55389 12632 55445
rect 12688 55389 12756 55445
rect 12812 55389 12880 55445
rect 12936 55389 13004 55445
rect 13060 55389 13100 55445
rect 12592 55321 13100 55389
rect 12592 55265 12632 55321
rect 12688 55265 12756 55321
rect 12812 55265 12880 55321
rect 12936 55265 13004 55321
rect 13060 55265 13100 55321
rect 12592 55197 13100 55265
rect 12592 55141 12632 55197
rect 12688 55141 12756 55197
rect 12812 55141 12880 55197
rect 12936 55141 13004 55197
rect 13060 55141 13100 55197
rect 12592 55073 13100 55141
rect 12592 55017 12632 55073
rect 12688 55017 12756 55073
rect 12812 55017 12880 55073
rect 12936 55017 13004 55073
rect 13060 55017 13100 55073
rect 12592 54949 13100 55017
rect 12592 54893 12632 54949
rect 12688 54893 12756 54949
rect 12812 54893 12880 54949
rect 12936 54893 13004 54949
rect 13060 54893 13100 54949
rect 12592 54825 13100 54893
rect 12592 54769 12632 54825
rect 12688 54769 12756 54825
rect 12812 54769 12880 54825
rect 12936 54769 13004 54825
rect 13060 54769 13100 54825
rect 12592 54701 13100 54769
rect 12592 54645 12632 54701
rect 12688 54645 12756 54701
rect 12812 54645 12880 54701
rect 12936 54645 13004 54701
rect 13060 54645 13100 54701
rect 12592 54577 13100 54645
rect 12592 54521 12632 54577
rect 12688 54521 12756 54577
rect 12812 54521 12880 54577
rect 12936 54521 13004 54577
rect 13060 54521 13100 54577
rect 12592 54453 13100 54521
rect 12592 54397 12632 54453
rect 12688 54397 12756 54453
rect 12812 54397 12880 54453
rect 12936 54397 13004 54453
rect 13060 54397 13100 54453
rect 12592 54329 13100 54397
rect 12592 54273 12632 54329
rect 12688 54273 12756 54329
rect 12812 54273 12880 54329
rect 12936 54273 13004 54329
rect 13060 54273 13100 54329
rect 12592 54205 13100 54273
rect 12592 54149 12632 54205
rect 12688 54149 12756 54205
rect 12812 54149 12880 54205
rect 12936 54149 13004 54205
rect 13060 54149 13100 54205
rect 12592 47445 13100 54149
rect 13160 56922 13668 56975
rect 13160 56866 13200 56922
rect 13256 56866 13324 56922
rect 13380 56866 13448 56922
rect 13504 56866 13572 56922
rect 13628 56866 13668 56922
rect 13160 56798 13668 56866
rect 13160 56742 13200 56798
rect 13256 56742 13324 56798
rect 13380 56742 13448 56798
rect 13504 56742 13572 56798
rect 13628 56742 13668 56798
rect 13160 56711 13668 56742
rect 13160 56659 13172 56711
rect 13224 56674 13280 56711
rect 13332 56674 13388 56711
rect 13256 56659 13280 56674
rect 13380 56659 13388 56674
rect 13440 56674 13496 56711
rect 13548 56674 13604 56711
rect 13440 56659 13448 56674
rect 13548 56659 13572 56674
rect 13656 56659 13668 56711
rect 13160 56618 13200 56659
rect 13256 56618 13324 56659
rect 13380 56618 13448 56659
rect 13504 56618 13572 56659
rect 13628 56618 13668 56659
rect 13160 56603 13668 56618
rect 13160 56551 13172 56603
rect 13224 56551 13280 56603
rect 13332 56551 13388 56603
rect 13440 56551 13496 56603
rect 13548 56551 13604 56603
rect 13656 56551 13668 56603
rect 13160 56550 13668 56551
rect 13160 56495 13200 56550
rect 13256 56495 13324 56550
rect 13380 56495 13448 56550
rect 13504 56495 13572 56550
rect 13628 56495 13668 56550
rect 13160 56443 13172 56495
rect 13256 56494 13280 56495
rect 13380 56494 13388 56495
rect 13224 56443 13280 56494
rect 13332 56443 13388 56494
rect 13440 56494 13448 56495
rect 13548 56494 13572 56495
rect 13440 56443 13496 56494
rect 13548 56443 13604 56494
rect 13656 56443 13668 56495
rect 13160 56426 13668 56443
rect 13160 56370 13200 56426
rect 13256 56370 13324 56426
rect 13380 56370 13448 56426
rect 13504 56370 13572 56426
rect 13628 56370 13668 56426
rect 13160 56302 13668 56370
rect 13160 56246 13200 56302
rect 13256 56246 13324 56302
rect 13380 56246 13448 56302
rect 13504 56246 13572 56302
rect 13628 56246 13668 56302
rect 13160 56178 13668 56246
rect 13160 56122 13200 56178
rect 13256 56122 13324 56178
rect 13380 56122 13448 56178
rect 13504 56122 13572 56178
rect 13628 56122 13668 56178
rect 13160 56054 13668 56122
rect 13160 55998 13200 56054
rect 13256 55998 13324 56054
rect 13380 55998 13448 56054
rect 13504 55998 13572 56054
rect 13628 55998 13668 56054
rect 13160 55930 13668 55998
rect 13160 55874 13200 55930
rect 13256 55874 13324 55930
rect 13380 55874 13448 55930
rect 13504 55874 13572 55930
rect 13628 55874 13668 55930
rect 13160 55806 13668 55874
rect 13160 55750 13200 55806
rect 13256 55750 13324 55806
rect 13380 55750 13448 55806
rect 13504 55750 13572 55806
rect 13628 55750 13668 55806
rect 13160 53845 13668 55750
rect 13160 53789 13200 53845
rect 13256 53789 13324 53845
rect 13380 53789 13448 53845
rect 13504 53789 13572 53845
rect 13628 53789 13668 53845
rect 13160 53721 13668 53789
rect 13160 53665 13200 53721
rect 13256 53665 13324 53721
rect 13380 53665 13448 53721
rect 13504 53665 13572 53721
rect 13628 53665 13668 53721
rect 13160 53597 13668 53665
rect 13160 53541 13200 53597
rect 13256 53541 13324 53597
rect 13380 53541 13448 53597
rect 13504 53541 13572 53597
rect 13628 53541 13668 53597
rect 13160 53473 13668 53541
rect 13160 53417 13200 53473
rect 13256 53417 13324 53473
rect 13380 53417 13448 53473
rect 13504 53417 13572 53473
rect 13628 53417 13668 53473
rect 13160 53349 13668 53417
rect 13160 53293 13200 53349
rect 13256 53293 13324 53349
rect 13380 53293 13448 53349
rect 13504 53293 13572 53349
rect 13628 53293 13668 53349
rect 13160 53225 13668 53293
rect 13160 53169 13200 53225
rect 13256 53169 13324 53225
rect 13380 53169 13448 53225
rect 13504 53169 13572 53225
rect 13628 53169 13668 53225
rect 13160 53101 13668 53169
rect 13160 53045 13200 53101
rect 13256 53045 13324 53101
rect 13380 53045 13448 53101
rect 13504 53045 13572 53101
rect 13628 53045 13668 53101
rect 13160 52996 13202 53045
rect 13254 52996 13326 53045
rect 13378 52996 13450 53045
rect 13502 52996 13574 53045
rect 13626 52996 13668 53045
rect 13160 52977 13668 52996
rect 13160 52921 13200 52977
rect 13256 52921 13324 52977
rect 13380 52921 13448 52977
rect 13504 52921 13572 52977
rect 13628 52921 13668 52977
rect 13160 52872 13202 52921
rect 13254 52872 13326 52921
rect 13378 52872 13450 52921
rect 13502 52872 13574 52921
rect 13626 52872 13668 52921
rect 13160 52853 13668 52872
rect 13160 52797 13200 52853
rect 13256 52797 13324 52853
rect 13380 52797 13448 52853
rect 13504 52797 13572 52853
rect 13628 52797 13668 52853
rect 13160 52748 13202 52797
rect 13254 52748 13326 52797
rect 13378 52748 13450 52797
rect 13502 52748 13574 52797
rect 13626 52748 13668 52797
rect 13160 52729 13668 52748
rect 13160 52673 13200 52729
rect 13256 52673 13324 52729
rect 13380 52673 13448 52729
rect 13504 52673 13572 52729
rect 13628 52673 13668 52729
rect 13160 52624 13202 52673
rect 13254 52624 13326 52673
rect 13378 52624 13450 52673
rect 13502 52624 13574 52673
rect 13626 52624 13668 52673
rect 13160 52605 13668 52624
rect 13160 52549 13200 52605
rect 13256 52549 13324 52605
rect 13380 52549 13448 52605
rect 13504 52549 13572 52605
rect 13628 52549 13668 52605
rect 13160 52500 13202 52549
rect 13254 52500 13326 52549
rect 13378 52500 13450 52549
rect 13502 52500 13574 52549
rect 13626 52500 13668 52549
rect 13160 52427 13668 52500
rect 12592 47389 12632 47445
rect 12688 47389 12756 47445
rect 12812 47389 12880 47445
rect 12936 47389 13004 47445
rect 13060 47389 13100 47445
rect 12592 47321 13100 47389
rect 12592 47265 12632 47321
rect 12688 47265 12756 47321
rect 12812 47265 12880 47321
rect 12936 47265 13004 47321
rect 13060 47265 13100 47321
rect 12592 47197 13100 47265
rect 12592 47141 12632 47197
rect 12688 47141 12756 47197
rect 12812 47141 12880 47197
rect 12936 47141 13004 47197
rect 13060 47141 13100 47197
rect 12592 47073 13100 47141
rect 12592 47017 12632 47073
rect 12688 47017 12756 47073
rect 12812 47017 12880 47073
rect 12936 47017 13004 47073
rect 13060 47017 13100 47073
rect 12592 46949 13100 47017
rect 12592 46893 12632 46949
rect 12688 46893 12756 46949
rect 12812 46893 12880 46949
rect 12936 46893 13004 46949
rect 13060 46893 13100 46949
rect 12592 46825 13100 46893
rect 12592 46769 12632 46825
rect 12688 46769 12756 46825
rect 12812 46769 12880 46825
rect 12936 46769 13004 46825
rect 13060 46769 13100 46825
rect 12592 46701 13100 46769
rect 12592 46645 12632 46701
rect 12688 46645 12756 46701
rect 12812 46645 12880 46701
rect 12936 46645 13004 46701
rect 13060 46645 13100 46701
rect 12592 46577 13100 46645
rect 12592 46521 12632 46577
rect 12688 46521 12756 46577
rect 12812 46521 12880 46577
rect 12936 46521 13004 46577
rect 13060 46521 13100 46577
rect 12592 46453 13100 46521
rect 12592 46397 12632 46453
rect 12688 46397 12756 46453
rect 12812 46397 12880 46453
rect 12936 46397 13004 46453
rect 13060 46397 13100 46453
rect 12592 46329 13100 46397
rect 12592 46273 12632 46329
rect 12688 46273 12756 46329
rect 12812 46273 12880 46329
rect 12936 46273 13004 46329
rect 13060 46273 13100 46329
rect 12592 46205 13100 46273
rect 12592 46149 12632 46205
rect 12688 46149 12756 46205
rect 12812 46149 12880 46205
rect 12936 46149 13004 46205
rect 13060 46149 13100 46205
rect 12592 44245 13100 46149
rect 12592 44189 12632 44245
rect 12688 44189 12756 44245
rect 12812 44189 12880 44245
rect 12936 44189 13004 44245
rect 13060 44189 13100 44245
rect 12592 44121 13100 44189
rect 12592 44065 12632 44121
rect 12688 44065 12756 44121
rect 12812 44065 12880 44121
rect 12936 44065 13004 44121
rect 13060 44065 13100 44121
rect 12592 43997 13100 44065
rect 12592 43941 12632 43997
rect 12688 43941 12756 43997
rect 12812 43941 12880 43997
rect 12936 43941 13004 43997
rect 13060 43941 13100 43997
rect 12592 43873 13100 43941
rect 12592 43817 12632 43873
rect 12688 43817 12756 43873
rect 12812 43817 12880 43873
rect 12936 43817 13004 43873
rect 13060 43817 13100 43873
rect 12592 43749 13100 43817
rect 12592 43693 12632 43749
rect 12688 43693 12756 43749
rect 12812 43693 12880 43749
rect 12936 43693 13004 43749
rect 13060 43693 13100 43749
rect 12592 43625 13100 43693
rect 12592 43569 12632 43625
rect 12688 43569 12756 43625
rect 12812 43569 12880 43625
rect 12936 43569 13004 43625
rect 13060 43569 13100 43625
rect 12592 43501 13100 43569
rect 12592 43445 12632 43501
rect 12688 43445 12756 43501
rect 12812 43445 12880 43501
rect 12936 43445 13004 43501
rect 13060 43445 13100 43501
rect 12592 43377 13100 43445
rect 12592 43321 12632 43377
rect 12688 43321 12756 43377
rect 12812 43321 12880 43377
rect 12936 43321 13004 43377
rect 13060 43321 13100 43377
rect 12592 43253 13100 43321
rect 12592 43197 12632 43253
rect 12688 43197 12756 43253
rect 12812 43197 12880 43253
rect 12936 43197 13004 43253
rect 13060 43197 13100 43253
rect 12592 43129 13100 43197
rect 12592 43073 12632 43129
rect 12688 43073 12756 43129
rect 12812 43073 12880 43129
rect 12936 43073 13004 43129
rect 13060 43073 13100 43129
rect 12592 43005 13100 43073
rect 12592 42949 12632 43005
rect 12688 42949 12756 43005
rect 12812 42949 12880 43005
rect 12936 42949 13004 43005
rect 13060 42949 13100 43005
rect 12592 42645 13100 42949
rect 12592 42589 12632 42645
rect 12688 42589 12756 42645
rect 12812 42589 12880 42645
rect 12936 42589 13004 42645
rect 13060 42589 13100 42645
rect 12592 42521 13100 42589
rect 12592 42465 12632 42521
rect 12688 42465 12756 42521
rect 12812 42465 12880 42521
rect 12936 42465 13004 42521
rect 13060 42465 13100 42521
rect 12592 42397 13100 42465
rect 12592 42341 12632 42397
rect 12688 42341 12756 42397
rect 12812 42341 12880 42397
rect 12936 42341 13004 42397
rect 13060 42341 13100 42397
rect 12592 42273 13100 42341
rect 12592 42217 12632 42273
rect 12688 42217 12756 42273
rect 12812 42217 12880 42273
rect 12936 42217 13004 42273
rect 13060 42217 13100 42273
rect 12592 42149 13100 42217
rect 12592 42093 12632 42149
rect 12688 42093 12756 42149
rect 12812 42093 12880 42149
rect 12936 42093 13004 42149
rect 13060 42093 13100 42149
rect 12592 42025 13100 42093
rect 12592 41969 12632 42025
rect 12688 41969 12756 42025
rect 12812 41969 12880 42025
rect 12936 41969 13004 42025
rect 13060 41969 13100 42025
rect 12592 41901 13100 41969
rect 12592 41845 12632 41901
rect 12688 41845 12756 41901
rect 12812 41845 12880 41901
rect 12936 41845 13004 41901
rect 13060 41845 13100 41901
rect 12592 41777 13100 41845
rect 12592 41721 12632 41777
rect 12688 41721 12756 41777
rect 12812 41721 12880 41777
rect 12936 41721 13004 41777
rect 13060 41721 13100 41777
rect 12592 41653 13100 41721
rect 12592 41597 12632 41653
rect 12688 41597 12756 41653
rect 12812 41597 12880 41653
rect 12936 41597 13004 41653
rect 13060 41597 13100 41653
rect 12592 41529 13100 41597
rect 12592 41473 12632 41529
rect 12688 41473 12756 41529
rect 12812 41473 12880 41529
rect 12936 41473 13004 41529
rect 13060 41473 13100 41529
rect 12592 41405 13100 41473
rect 12592 41349 12632 41405
rect 12688 41349 12756 41405
rect 12812 41349 12880 41405
rect 12936 41349 13004 41405
rect 13060 41349 13100 41405
rect 12592 41045 13100 41349
rect 12592 40989 12632 41045
rect 12688 40989 12756 41045
rect 12812 40989 12880 41045
rect 12936 40989 13004 41045
rect 13060 40989 13100 41045
rect 12592 40921 13100 40989
rect 12592 40865 12632 40921
rect 12688 40865 12756 40921
rect 12812 40865 12880 40921
rect 12936 40865 13004 40921
rect 13060 40865 13100 40921
rect 12592 40797 13100 40865
rect 12592 40741 12632 40797
rect 12688 40741 12756 40797
rect 12812 40741 12880 40797
rect 12936 40741 13004 40797
rect 13060 40741 13100 40797
rect 12592 40673 13100 40741
rect 12592 40617 12632 40673
rect 12688 40617 12756 40673
rect 12812 40617 12880 40673
rect 12936 40617 13004 40673
rect 13060 40617 13100 40673
rect 12592 40549 13100 40617
rect 12592 40493 12632 40549
rect 12688 40493 12756 40549
rect 12812 40493 12880 40549
rect 12936 40493 13004 40549
rect 13060 40493 13100 40549
rect 12592 40425 13100 40493
rect 12592 40369 12632 40425
rect 12688 40369 12756 40425
rect 12812 40369 12880 40425
rect 12936 40369 13004 40425
rect 13060 40369 13100 40425
rect 12592 40301 13100 40369
rect 12592 40245 12632 40301
rect 12688 40245 12756 40301
rect 12812 40245 12880 40301
rect 12936 40245 13004 40301
rect 13060 40245 13100 40301
rect 12592 40177 13100 40245
rect 12592 40121 12632 40177
rect 12688 40121 12756 40177
rect 12812 40121 12880 40177
rect 12936 40121 13004 40177
rect 13060 40121 13100 40177
rect 12592 40053 13100 40121
rect 12592 39997 12632 40053
rect 12688 39997 12756 40053
rect 12812 39997 12880 40053
rect 12936 39997 13004 40053
rect 13060 39997 13100 40053
rect 12592 39929 13100 39997
rect 12592 39873 12632 39929
rect 12688 39873 12756 39929
rect 12812 39873 12880 39929
rect 12936 39873 13004 39929
rect 13060 39873 13100 39929
rect 12592 39805 13100 39873
rect 12592 39749 12632 39805
rect 12688 39749 12756 39805
rect 12812 39749 12880 39805
rect 12936 39749 13004 39805
rect 13060 39749 13100 39805
rect 12592 33051 13100 39749
rect 13160 52245 13360 52297
rect 13160 52189 13170 52245
rect 13226 52189 13294 52245
rect 13350 52189 13360 52245
rect 13160 52121 13360 52189
rect 13160 52065 13170 52121
rect 13226 52065 13294 52121
rect 13350 52065 13360 52121
rect 13160 51997 13360 52065
rect 13160 51941 13170 51997
rect 13226 51941 13294 51997
rect 13350 51941 13360 51997
rect 13160 51873 13360 51941
rect 13160 51817 13170 51873
rect 13226 51817 13294 51873
rect 13350 51817 13360 51873
rect 13160 51749 13360 51817
rect 13160 51693 13170 51749
rect 13226 51693 13294 51749
rect 13350 51693 13360 51749
rect 13160 51625 13360 51693
rect 13160 51569 13170 51625
rect 13226 51569 13294 51625
rect 13350 51569 13360 51625
rect 13160 51501 13360 51569
rect 13160 51445 13170 51501
rect 13226 51445 13294 51501
rect 13350 51445 13360 51501
rect 13160 51377 13360 51445
rect 13160 51321 13170 51377
rect 13226 51321 13294 51377
rect 13350 51321 13360 51377
rect 13160 51253 13360 51321
rect 13160 51197 13170 51253
rect 13226 51197 13294 51253
rect 13350 51197 13360 51253
rect 13160 51129 13360 51197
rect 13160 51073 13170 51129
rect 13226 51073 13294 51129
rect 13350 51073 13360 51129
rect 13160 51005 13360 51073
rect 13160 50949 13170 51005
rect 13226 50949 13294 51005
rect 13350 50949 13360 51005
rect 13160 37845 13360 50949
rect 13160 37789 13170 37845
rect 13226 37789 13294 37845
rect 13350 37789 13360 37845
rect 13160 37721 13360 37789
rect 13160 37665 13170 37721
rect 13226 37665 13294 37721
rect 13350 37665 13360 37721
rect 13160 37597 13360 37665
rect 13160 37541 13170 37597
rect 13226 37541 13294 37597
rect 13350 37541 13360 37597
rect 13160 37473 13360 37541
rect 13160 37417 13170 37473
rect 13226 37417 13294 37473
rect 13350 37417 13360 37473
rect 13160 37349 13360 37417
rect 13160 37293 13170 37349
rect 13226 37293 13294 37349
rect 13350 37293 13360 37349
rect 13160 37225 13360 37293
rect 13160 37169 13170 37225
rect 13226 37169 13294 37225
rect 13350 37169 13360 37225
rect 13160 37101 13360 37169
rect 13160 37045 13170 37101
rect 13226 37045 13294 37101
rect 13350 37045 13360 37101
rect 13160 36977 13360 37045
rect 13160 36921 13170 36977
rect 13226 36921 13294 36977
rect 13350 36921 13360 36977
rect 13160 36853 13360 36921
rect 13160 36797 13170 36853
rect 13226 36797 13294 36853
rect 13350 36797 13360 36853
rect 13160 36729 13360 36797
rect 13160 36673 13170 36729
rect 13226 36673 13294 36729
rect 13350 36673 13360 36729
rect 13160 36605 13360 36673
rect 13160 36549 13170 36605
rect 13226 36549 13294 36605
rect 13350 36549 13360 36605
rect 13160 36497 13360 36549
rect 13468 49100 13668 52427
rect 13468 49048 13480 49100
rect 13532 49048 13604 49100
rect 13656 49048 13668 49100
rect 13468 49045 13668 49048
rect 13468 48989 13478 49045
rect 13534 48989 13602 49045
rect 13658 48989 13668 49045
rect 13468 48976 13668 48989
rect 13468 48924 13480 48976
rect 13532 48924 13604 48976
rect 13656 48924 13668 48976
rect 13468 48921 13668 48924
rect 13468 48865 13478 48921
rect 13534 48865 13602 48921
rect 13658 48865 13668 48921
rect 13468 48852 13668 48865
rect 13468 48800 13480 48852
rect 13532 48800 13604 48852
rect 13656 48800 13668 48852
rect 13468 48797 13668 48800
rect 13468 48741 13478 48797
rect 13534 48741 13602 48797
rect 13658 48741 13668 48797
rect 13468 48728 13668 48741
rect 13468 48676 13480 48728
rect 13532 48676 13604 48728
rect 13656 48676 13668 48728
rect 13468 48673 13668 48676
rect 13468 48617 13478 48673
rect 13534 48617 13602 48673
rect 13658 48617 13668 48673
rect 13468 48604 13668 48617
rect 13468 48552 13480 48604
rect 13532 48552 13604 48604
rect 13656 48552 13668 48604
rect 13468 48549 13668 48552
rect 13468 48493 13478 48549
rect 13534 48493 13602 48549
rect 13658 48493 13668 48549
rect 13468 48425 13668 48493
rect 13468 48369 13478 48425
rect 13534 48369 13602 48425
rect 13658 48369 13668 48425
rect 13468 48301 13668 48369
rect 13468 48245 13478 48301
rect 13534 48245 13602 48301
rect 13658 48245 13668 48301
rect 13468 48177 13668 48245
rect 13468 48121 13478 48177
rect 13534 48121 13602 48177
rect 13658 48121 13668 48177
rect 13468 48053 13668 48121
rect 13468 47997 13478 48053
rect 13534 47997 13602 48053
rect 13658 47997 13668 48053
rect 13468 47929 13668 47997
rect 13468 47873 13478 47929
rect 13534 47873 13602 47929
rect 13658 47873 13668 47929
rect 13468 47805 13668 47873
rect 13468 47749 13478 47805
rect 13534 47749 13602 47805
rect 13658 47749 13668 47805
rect 13468 45845 13668 47749
rect 13468 45789 13478 45845
rect 13534 45789 13602 45845
rect 13658 45789 13668 45845
rect 13468 45721 13668 45789
rect 13468 45665 13478 45721
rect 13534 45665 13602 45721
rect 13658 45665 13668 45721
rect 13468 45597 13668 45665
rect 13468 45541 13478 45597
rect 13534 45541 13602 45597
rect 13658 45541 13668 45597
rect 13468 45473 13668 45541
rect 13468 45417 13478 45473
rect 13534 45417 13602 45473
rect 13658 45417 13668 45473
rect 13468 45349 13668 45417
rect 13468 45293 13478 45349
rect 13534 45293 13602 45349
rect 13658 45293 13668 45349
rect 13468 45225 13668 45293
rect 13468 45169 13478 45225
rect 13534 45169 13602 45225
rect 13658 45169 13668 45225
rect 13468 45152 13668 45169
rect 13468 45101 13480 45152
rect 13532 45101 13604 45152
rect 13656 45101 13668 45152
rect 13468 45045 13478 45101
rect 13534 45045 13602 45101
rect 13658 45045 13668 45101
rect 13468 45028 13668 45045
rect 13468 44977 13480 45028
rect 13532 44977 13604 45028
rect 13656 44977 13668 45028
rect 13468 44921 13478 44977
rect 13534 44921 13602 44977
rect 13658 44921 13668 44977
rect 13468 44904 13668 44921
rect 13468 44853 13480 44904
rect 13532 44853 13604 44904
rect 13656 44853 13668 44904
rect 13468 44797 13478 44853
rect 13534 44797 13602 44853
rect 13658 44797 13668 44853
rect 13468 44780 13668 44797
rect 13468 44729 13480 44780
rect 13532 44729 13604 44780
rect 13656 44729 13668 44780
rect 13468 44673 13478 44729
rect 13534 44673 13602 44729
rect 13658 44673 13668 44729
rect 13468 44656 13668 44673
rect 13468 44605 13480 44656
rect 13532 44605 13604 44656
rect 13656 44605 13668 44656
rect 13468 44549 13478 44605
rect 13534 44549 13602 44605
rect 13658 44549 13668 44605
rect 13468 41204 13668 44549
rect 13468 41152 13480 41204
rect 13532 41152 13604 41204
rect 13656 41152 13668 41204
rect 13468 41080 13668 41152
rect 13468 41028 13480 41080
rect 13532 41028 13604 41080
rect 13656 41028 13668 41080
rect 13468 40956 13668 41028
rect 13468 40904 13480 40956
rect 13532 40904 13604 40956
rect 13656 40904 13668 40956
rect 13468 40832 13668 40904
rect 13468 40780 13480 40832
rect 13532 40780 13604 40832
rect 13656 40780 13668 40832
rect 13468 40708 13668 40780
rect 13468 40656 13480 40708
rect 13532 40656 13604 40708
rect 13656 40656 13668 40708
rect 13468 37256 13668 40656
rect 13468 37204 13480 37256
rect 13532 37204 13604 37256
rect 13656 37204 13668 37256
rect 13468 37132 13668 37204
rect 13468 37080 13480 37132
rect 13532 37080 13604 37132
rect 13656 37080 13668 37132
rect 13468 37008 13668 37080
rect 13468 36956 13480 37008
rect 13532 36956 13604 37008
rect 13656 36956 13668 37008
rect 13468 36884 13668 36956
rect 13468 36832 13480 36884
rect 13532 36832 13604 36884
rect 13656 36832 13668 36884
rect 13468 36760 13668 36832
rect 13468 36708 13480 36760
rect 13532 36708 13604 36760
rect 13656 36708 13668 36760
rect 13468 36261 13668 36708
rect 13190 36260 13668 36261
rect 12592 32995 12632 33051
rect 12688 32995 12756 33051
rect 12812 32995 12880 33051
rect 12936 32995 13004 33051
rect 13060 32995 13100 33051
rect 12592 32927 13100 32995
rect 12592 32871 12632 32927
rect 12688 32871 12756 32927
rect 12812 32871 12880 32927
rect 12936 32871 13004 32927
rect 13060 32871 13100 32927
rect 12592 32803 13100 32871
rect 12592 32747 12632 32803
rect 12688 32747 12756 32803
rect 12812 32747 12880 32803
rect 12936 32747 13004 32803
rect 13060 32747 13100 32803
rect 12592 32679 13100 32747
rect 12592 32623 12632 32679
rect 12688 32623 12756 32679
rect 12812 32623 12880 32679
rect 12936 32623 13004 32679
rect 13060 32623 13100 32679
rect 12592 32555 13100 32623
rect 12592 32499 12632 32555
rect 12688 32499 12756 32555
rect 12812 32499 12880 32555
rect 12936 32499 13004 32555
rect 13060 32499 13100 32555
rect 12592 32431 13100 32499
rect 12592 32375 12632 32431
rect 12688 32375 12756 32431
rect 12812 32375 12880 32431
rect 12936 32375 13004 32431
rect 13060 32375 13100 32431
rect 12592 32307 13100 32375
rect 12592 32251 12632 32307
rect 12688 32251 12756 32307
rect 12812 32251 12880 32307
rect 12936 32251 13004 32307
rect 13060 32251 13100 32307
rect 12592 32183 13100 32251
rect 12592 32127 12632 32183
rect 12688 32127 12756 32183
rect 12812 32127 12880 32183
rect 12936 32127 13004 32183
rect 13060 32127 13100 32183
rect 12592 32059 13100 32127
rect 12592 32003 12632 32059
rect 12688 32003 12756 32059
rect 12812 32003 12880 32059
rect 12936 32003 13004 32059
rect 13060 32003 13100 32059
rect 12592 31935 13100 32003
rect 12592 31879 12632 31935
rect 12688 31879 12756 31935
rect 12812 31879 12880 31935
rect 12936 31879 13004 31935
rect 13060 31879 13100 31935
rect 12592 31811 13100 31879
rect 12592 31755 12632 31811
rect 12688 31755 12756 31811
rect 12812 31755 12880 31811
rect 12936 31755 13004 31811
rect 13060 31755 13100 31811
rect 12592 31687 13100 31755
rect 12592 31631 12632 31687
rect 12688 31631 12756 31687
rect 12812 31631 12880 31687
rect 12936 31631 13004 31687
rect 13060 31631 13100 31687
rect 12592 31563 13100 31631
rect 12592 31507 12632 31563
rect 12688 31507 12756 31563
rect 12812 31507 12880 31563
rect 12936 31507 13004 31563
rect 13060 31507 13100 31563
rect 12592 31439 13100 31507
rect 12592 31383 12632 31439
rect 12688 31383 12756 31439
rect 12812 31383 12880 31439
rect 12936 31383 13004 31439
rect 13060 31383 13100 31439
rect 12592 31315 13100 31383
rect 12592 31259 12632 31315
rect 12688 31259 12756 31315
rect 12812 31259 12880 31315
rect 12936 31259 13004 31315
rect 13060 31259 13100 31315
rect 12592 31191 13100 31259
rect 12592 31135 12632 31191
rect 12688 31135 12756 31191
rect 12812 31135 12880 31191
rect 12936 31135 13004 31191
rect 13060 31135 13100 31191
rect 12592 31067 13100 31135
rect 12592 31011 12632 31067
rect 12688 31011 12756 31067
rect 12812 31011 12880 31067
rect 12936 31011 13004 31067
rect 13060 31011 13100 31067
rect 12592 30943 13100 31011
rect 12592 30887 12632 30943
rect 12688 30887 12756 30943
rect 12812 30887 12880 30943
rect 12936 30887 13004 30943
rect 13060 30887 13100 30943
rect 12592 30819 13100 30887
rect 12592 30763 12632 30819
rect 12688 30763 12756 30819
rect 12812 30763 12880 30819
rect 12936 30763 13004 30819
rect 13060 30763 13100 30819
rect 12592 30695 13100 30763
rect 12592 30639 12632 30695
rect 12688 30639 12756 30695
rect 12812 30639 12880 30695
rect 12936 30639 13004 30695
rect 13060 30639 13100 30695
rect 12592 30571 13100 30639
rect 12592 30515 12632 30571
rect 12688 30515 12756 30571
rect 12812 30515 12880 30571
rect 12936 30515 13004 30571
rect 13060 30515 13100 30571
rect 12592 30447 13100 30515
rect 12592 30391 12632 30447
rect 12688 30391 12756 30447
rect 12812 30391 12880 30447
rect 12936 30391 13004 30447
rect 13060 30391 13100 30447
rect 12592 30323 13100 30391
rect 12592 30267 12632 30323
rect 12688 30267 12756 30323
rect 12812 30267 12880 30323
rect 12936 30267 13004 30323
rect 13060 30267 13100 30323
rect 12592 30199 13100 30267
rect 12592 30143 12632 30199
rect 12688 30143 12756 30199
rect 12812 30143 12880 30199
rect 12936 30143 13004 30199
rect 13060 30143 13100 30199
rect 12592 29845 13100 30143
rect 12592 29789 12632 29845
rect 12688 29789 12756 29845
rect 12812 29789 12880 29845
rect 12936 29789 13004 29845
rect 13060 29789 13100 29845
rect 12592 29721 13100 29789
rect 12592 29665 12632 29721
rect 12688 29665 12756 29721
rect 12812 29665 12880 29721
rect 12936 29665 13004 29721
rect 13060 29665 13100 29721
rect 12592 29597 13100 29665
rect 12592 29541 12632 29597
rect 12688 29541 12756 29597
rect 12812 29541 12880 29597
rect 12936 29541 13004 29597
rect 13060 29541 13100 29597
rect 12592 29473 13100 29541
rect 12592 29417 12632 29473
rect 12688 29417 12756 29473
rect 12812 29417 12880 29473
rect 12936 29417 13004 29473
rect 13060 29417 13100 29473
rect 12592 29349 13100 29417
rect 12592 29293 12632 29349
rect 12688 29293 12756 29349
rect 12812 29293 12880 29349
rect 12936 29293 13004 29349
rect 13060 29293 13100 29349
rect 12592 29225 13100 29293
rect 12592 29169 12632 29225
rect 12688 29169 12756 29225
rect 12812 29169 12880 29225
rect 12936 29169 13004 29225
rect 13060 29169 13100 29225
rect 12592 29101 13100 29169
rect 12592 29045 12632 29101
rect 12688 29045 12756 29101
rect 12812 29045 12880 29101
rect 12936 29045 13004 29101
rect 13060 29045 13100 29101
rect 12592 28977 13100 29045
rect 12592 28921 12632 28977
rect 12688 28921 12756 28977
rect 12812 28921 12880 28977
rect 12936 28921 13004 28977
rect 13060 28921 13100 28977
rect 12592 28853 13100 28921
rect 12592 28797 12632 28853
rect 12688 28797 12756 28853
rect 12812 28797 12880 28853
rect 12936 28797 13004 28853
rect 13060 28797 13100 28853
rect 12592 28729 13100 28797
rect 12592 28673 12632 28729
rect 12688 28673 12756 28729
rect 12812 28673 12880 28729
rect 12936 28673 13004 28729
rect 13060 28673 13100 28729
rect 12592 28605 13100 28673
rect 12592 28549 12632 28605
rect 12688 28549 12756 28605
rect 12812 28549 12880 28605
rect 12936 28549 13004 28605
rect 13060 28549 13100 28605
rect 12592 26651 13100 28549
rect 12592 26595 12632 26651
rect 12688 26595 12756 26651
rect 12812 26595 12880 26651
rect 12936 26595 13004 26651
rect 13060 26595 13100 26651
rect 12592 26527 13100 26595
rect 12592 26471 12632 26527
rect 12688 26471 12756 26527
rect 12812 26471 12880 26527
rect 12936 26471 13004 26527
rect 13060 26471 13100 26527
rect 12592 26403 13100 26471
rect 12592 26347 12632 26403
rect 12688 26347 12756 26403
rect 12812 26347 12880 26403
rect 12936 26347 13004 26403
rect 13060 26347 13100 26403
rect 12592 26279 13100 26347
rect 12592 26223 12632 26279
rect 12688 26223 12756 26279
rect 12812 26223 12880 26279
rect 12936 26223 13004 26279
rect 13060 26223 13100 26279
rect 12592 26155 13100 26223
rect 12592 26099 12632 26155
rect 12688 26099 12756 26155
rect 12812 26099 12880 26155
rect 12936 26099 13004 26155
rect 13060 26099 13100 26155
rect 12592 26031 13100 26099
rect 12592 25975 12632 26031
rect 12688 25975 12756 26031
rect 12812 25975 12880 26031
rect 12936 25975 13004 26031
rect 13060 25975 13100 26031
rect 12592 25907 13100 25975
rect 12592 25851 12632 25907
rect 12688 25851 12756 25907
rect 12812 25851 12880 25907
rect 12936 25851 13004 25907
rect 13060 25851 13100 25907
rect 12592 25783 13100 25851
rect 12592 25727 12632 25783
rect 12688 25727 12756 25783
rect 12812 25727 12880 25783
rect 12936 25727 13004 25783
rect 13060 25727 13100 25783
rect 12592 25659 13100 25727
rect 12592 25603 12632 25659
rect 12688 25603 12756 25659
rect 12812 25603 12880 25659
rect 12936 25603 13004 25659
rect 13060 25603 13100 25659
rect 12592 25535 13100 25603
rect 12592 25479 12632 25535
rect 12688 25479 12756 25535
rect 12812 25479 12880 25535
rect 12936 25479 13004 25535
rect 13060 25479 13100 25535
rect 12592 25411 13100 25479
rect 12592 25355 12632 25411
rect 12688 25355 12756 25411
rect 12812 25355 12880 25411
rect 12936 25355 13004 25411
rect 13060 25355 13100 25411
rect 12592 25287 13100 25355
rect 12592 25231 12632 25287
rect 12688 25231 12756 25287
rect 12812 25231 12880 25287
rect 12936 25231 13004 25287
rect 13060 25231 13100 25287
rect 12592 25163 13100 25231
rect 12592 25107 12632 25163
rect 12688 25107 12756 25163
rect 12812 25107 12880 25163
rect 12936 25107 13004 25163
rect 13060 25107 13100 25163
rect 12592 25039 13100 25107
rect 12592 24983 12632 25039
rect 12688 24983 12756 25039
rect 12812 24983 12880 25039
rect 12936 24983 13004 25039
rect 13060 24983 13100 25039
rect 12592 24915 13100 24983
rect 12592 24859 12632 24915
rect 12688 24859 12756 24915
rect 12812 24859 12880 24915
rect 12936 24859 13004 24915
rect 13060 24859 13100 24915
rect 12592 24791 13100 24859
rect 12592 24735 12632 24791
rect 12688 24735 12756 24791
rect 12812 24735 12880 24791
rect 12936 24735 13004 24791
rect 13060 24735 13100 24791
rect 12592 24667 13100 24735
rect 12592 24611 12632 24667
rect 12688 24611 12756 24667
rect 12812 24611 12880 24667
rect 12936 24611 13004 24667
rect 13060 24611 13100 24667
rect 12592 24543 13100 24611
rect 12592 24487 12632 24543
rect 12688 24487 12756 24543
rect 12812 24487 12880 24543
rect 12936 24487 13004 24543
rect 13060 24487 13100 24543
rect 12592 24419 13100 24487
rect 12592 24363 12632 24419
rect 12688 24363 12756 24419
rect 12812 24363 12880 24419
rect 12936 24363 13004 24419
rect 13060 24363 13100 24419
rect 12592 24295 13100 24363
rect 12592 24239 12632 24295
rect 12688 24239 12756 24295
rect 12812 24239 12880 24295
rect 12936 24239 13004 24295
rect 13060 24239 13100 24295
rect 12592 24171 13100 24239
rect 12592 24115 12632 24171
rect 12688 24115 12756 24171
rect 12812 24115 12880 24171
rect 12936 24115 13004 24171
rect 13060 24115 13100 24171
rect 12592 24047 13100 24115
rect 12592 23991 12632 24047
rect 12688 23991 12756 24047
rect 12812 23991 12880 24047
rect 12936 23991 13004 24047
rect 13060 23991 13100 24047
rect 12592 23923 13100 23991
rect 12592 23867 12632 23923
rect 12688 23867 12756 23923
rect 12812 23867 12880 23923
rect 12936 23867 13004 23923
rect 13060 23867 13100 23923
rect 12592 23799 13100 23867
rect 12592 23743 12632 23799
rect 12688 23743 12756 23799
rect 12812 23743 12880 23799
rect 12936 23743 13004 23799
rect 13060 23743 13100 23799
rect 12592 23451 13100 23743
rect 12592 23395 12632 23451
rect 12688 23395 12756 23451
rect 12812 23395 12880 23451
rect 12936 23395 13004 23451
rect 13060 23395 13100 23451
rect 12592 23327 13100 23395
rect 12592 23271 12632 23327
rect 12688 23271 12756 23327
rect 12812 23271 12880 23327
rect 12936 23271 13004 23327
rect 13060 23271 13100 23327
rect 12592 23203 13100 23271
rect 12592 23147 12632 23203
rect 12688 23147 12756 23203
rect 12812 23147 12880 23203
rect 12936 23147 13004 23203
rect 13060 23147 13100 23203
rect 12592 23079 13100 23147
rect 12592 23023 12632 23079
rect 12688 23023 12756 23079
rect 12812 23023 12880 23079
rect 12936 23023 13004 23079
rect 13060 23023 13100 23079
rect 12592 22955 13100 23023
rect 12592 22899 12632 22955
rect 12688 22899 12756 22955
rect 12812 22899 12880 22955
rect 12936 22899 13004 22955
rect 13060 22899 13100 22955
rect 12592 22831 13100 22899
rect 12592 22775 12632 22831
rect 12688 22775 12756 22831
rect 12812 22775 12880 22831
rect 12936 22775 13004 22831
rect 13060 22775 13100 22831
rect 12592 22707 13100 22775
rect 12592 22651 12632 22707
rect 12688 22651 12756 22707
rect 12812 22651 12880 22707
rect 12936 22651 13004 22707
rect 13060 22651 13100 22707
rect 12592 22583 13100 22651
rect 12592 22527 12632 22583
rect 12688 22527 12756 22583
rect 12812 22527 12880 22583
rect 12936 22527 13004 22583
rect 13060 22527 13100 22583
rect 12592 22459 13100 22527
rect 12592 22403 12632 22459
rect 12688 22403 12756 22459
rect 12812 22403 12880 22459
rect 12936 22403 13004 22459
rect 13060 22403 13100 22459
rect 12592 22335 13100 22403
rect 12592 22279 12632 22335
rect 12688 22279 12756 22335
rect 12812 22279 12880 22335
rect 12936 22279 13004 22335
rect 13060 22279 13100 22335
rect 12592 22211 13100 22279
rect 12592 22155 12632 22211
rect 12688 22155 12756 22211
rect 12812 22155 12880 22211
rect 12936 22155 13004 22211
rect 13060 22155 13100 22211
rect 12592 22087 13100 22155
rect 12592 22031 12632 22087
rect 12688 22031 12756 22087
rect 12812 22031 12880 22087
rect 12936 22031 13004 22087
rect 13060 22031 13100 22087
rect 12592 21963 13100 22031
rect 12592 21907 12632 21963
rect 12688 21907 12756 21963
rect 12812 21907 12880 21963
rect 12936 21907 13004 21963
rect 13060 21907 13100 21963
rect 12592 21839 13100 21907
rect 12592 21783 12632 21839
rect 12688 21783 12756 21839
rect 12812 21783 12880 21839
rect 12936 21783 13004 21839
rect 13060 21783 13100 21839
rect 12592 21715 13100 21783
rect 12592 21659 12632 21715
rect 12688 21659 12756 21715
rect 12812 21659 12880 21715
rect 12936 21659 13004 21715
rect 13060 21659 13100 21715
rect 12592 21591 13100 21659
rect 12592 21535 12632 21591
rect 12688 21535 12756 21591
rect 12812 21535 12880 21591
rect 12936 21535 13004 21591
rect 13060 21535 13100 21591
rect 12592 21467 13100 21535
rect 12592 21411 12632 21467
rect 12688 21411 12756 21467
rect 12812 21411 12880 21467
rect 12936 21411 13004 21467
rect 13060 21411 13100 21467
rect 12592 21343 13100 21411
rect 12592 21287 12632 21343
rect 12688 21287 12756 21343
rect 12812 21287 12880 21343
rect 12936 21287 13004 21343
rect 13060 21287 13100 21343
rect 12592 21219 13100 21287
rect 12592 21163 12632 21219
rect 12688 21163 12756 21219
rect 12812 21163 12880 21219
rect 12936 21163 13004 21219
rect 13060 21163 13100 21219
rect 12592 21095 13100 21163
rect 12592 21039 12632 21095
rect 12688 21039 12756 21095
rect 12812 21039 12880 21095
rect 12936 21039 13004 21095
rect 13060 21039 13100 21095
rect 12592 20971 13100 21039
rect 12592 20915 12632 20971
rect 12688 20915 12756 20971
rect 12812 20915 12880 20971
rect 12936 20915 13004 20971
rect 13060 20915 13100 20971
rect 12592 20847 13100 20915
rect 12592 20791 12632 20847
rect 12688 20791 12756 20847
rect 12812 20791 12880 20847
rect 12936 20791 13004 20847
rect 13060 20791 13100 20847
rect 12592 20723 13100 20791
rect 12592 20667 12632 20723
rect 12688 20667 12756 20723
rect 12812 20667 12880 20723
rect 12936 20667 13004 20723
rect 13060 20667 13100 20723
rect 12592 20599 13100 20667
rect 12592 20543 12632 20599
rect 12688 20543 12756 20599
rect 12812 20543 12880 20599
rect 12936 20543 13004 20599
rect 13060 20543 13100 20599
rect 12592 20251 13100 20543
rect 12592 20195 12632 20251
rect 12688 20195 12756 20251
rect 12812 20195 12880 20251
rect 12936 20195 13004 20251
rect 13060 20195 13100 20251
rect 12592 20127 13100 20195
rect 12592 20071 12632 20127
rect 12688 20071 12756 20127
rect 12812 20071 12880 20127
rect 12936 20071 13004 20127
rect 13060 20071 13100 20127
rect 12592 20003 13100 20071
rect 12592 19947 12632 20003
rect 12688 19947 12756 20003
rect 12812 19947 12880 20003
rect 12936 19947 13004 20003
rect 13060 19947 13100 20003
rect 12592 19879 13100 19947
rect 12592 19823 12632 19879
rect 12688 19823 12756 19879
rect 12812 19823 12880 19879
rect 12936 19823 13004 19879
rect 13060 19823 13100 19879
rect 12592 19755 13100 19823
rect 12592 19699 12632 19755
rect 12688 19699 12756 19755
rect 12812 19699 12880 19755
rect 12936 19699 13004 19755
rect 13060 19699 13100 19755
rect 12592 19631 13100 19699
rect 12592 19575 12632 19631
rect 12688 19575 12756 19631
rect 12812 19575 12880 19631
rect 12936 19575 13004 19631
rect 13060 19575 13100 19631
rect 12592 19507 13100 19575
rect 12592 19451 12632 19507
rect 12688 19451 12756 19507
rect 12812 19451 12880 19507
rect 12936 19451 13004 19507
rect 13060 19451 13100 19507
rect 12592 19383 13100 19451
rect 12592 19327 12632 19383
rect 12688 19327 12756 19383
rect 12812 19327 12880 19383
rect 12936 19327 13004 19383
rect 13060 19327 13100 19383
rect 12592 19259 13100 19327
rect 12592 19203 12632 19259
rect 12688 19203 12756 19259
rect 12812 19203 12880 19259
rect 12936 19203 13004 19259
rect 13060 19203 13100 19259
rect 12592 19135 13100 19203
rect 12592 19079 12632 19135
rect 12688 19079 12756 19135
rect 12812 19079 12880 19135
rect 12936 19079 13004 19135
rect 13060 19079 13100 19135
rect 12592 19011 13100 19079
rect 12592 18955 12632 19011
rect 12688 18955 12756 19011
rect 12812 18955 12880 19011
rect 12936 18955 13004 19011
rect 13060 18955 13100 19011
rect 12592 18887 13100 18955
rect 12592 18831 12632 18887
rect 12688 18831 12756 18887
rect 12812 18831 12880 18887
rect 12936 18831 13004 18887
rect 13060 18831 13100 18887
rect 12592 18763 13100 18831
rect 12592 18707 12632 18763
rect 12688 18707 12756 18763
rect 12812 18707 12880 18763
rect 12936 18707 13004 18763
rect 13060 18707 13100 18763
rect 12592 18639 13100 18707
rect 12592 18583 12632 18639
rect 12688 18583 12756 18639
rect 12812 18583 12880 18639
rect 12936 18583 13004 18639
rect 13060 18583 13100 18639
rect 12592 18515 13100 18583
rect 12592 18459 12632 18515
rect 12688 18459 12756 18515
rect 12812 18459 12880 18515
rect 12936 18459 13004 18515
rect 13060 18459 13100 18515
rect 12592 18391 13100 18459
rect 12592 18335 12632 18391
rect 12688 18335 12756 18391
rect 12812 18335 12880 18391
rect 12936 18335 13004 18391
rect 13060 18335 13100 18391
rect 12592 18267 13100 18335
rect 12592 18211 12632 18267
rect 12688 18211 12756 18267
rect 12812 18211 12880 18267
rect 12936 18211 13004 18267
rect 13060 18211 13100 18267
rect 12592 18143 13100 18211
rect 12592 18087 12632 18143
rect 12688 18087 12756 18143
rect 12812 18087 12880 18143
rect 12936 18087 13004 18143
rect 13060 18087 13100 18143
rect 12592 18019 13100 18087
rect 12592 17963 12632 18019
rect 12688 17963 12756 18019
rect 12812 17963 12880 18019
rect 12936 17963 13004 18019
rect 13060 17963 13100 18019
rect 12592 17895 13100 17963
rect 12592 17839 12632 17895
rect 12688 17839 12756 17895
rect 12812 17839 12880 17895
rect 12936 17839 13004 17895
rect 13060 17839 13100 17895
rect 12592 17771 13100 17839
rect 12592 17715 12632 17771
rect 12688 17715 12756 17771
rect 12812 17715 12880 17771
rect 12936 17715 13004 17771
rect 13060 17715 13100 17771
rect 12592 17647 13100 17715
rect 12592 17591 12632 17647
rect 12688 17591 12756 17647
rect 12812 17591 12880 17647
rect 12936 17591 13004 17647
rect 13060 17591 13100 17647
rect 12592 17523 13100 17591
rect 12592 17467 12632 17523
rect 12688 17467 12756 17523
rect 12812 17467 12880 17523
rect 12936 17467 13004 17523
rect 13060 17467 13100 17523
rect 12592 17399 13100 17467
rect 12592 17343 12632 17399
rect 12688 17343 12756 17399
rect 12812 17343 12880 17399
rect 12936 17343 13004 17399
rect 13060 17343 13100 17399
rect 12592 17051 13100 17343
rect 12592 16995 12632 17051
rect 12688 16995 12756 17051
rect 12812 16995 12880 17051
rect 12936 16995 13004 17051
rect 13060 16995 13100 17051
rect 12592 16927 13100 16995
rect 12592 16871 12632 16927
rect 12688 16871 12756 16927
rect 12812 16871 12880 16927
rect 12936 16871 13004 16927
rect 13060 16871 13100 16927
rect 12592 16803 13100 16871
rect 12592 16747 12632 16803
rect 12688 16747 12756 16803
rect 12812 16747 12880 16803
rect 12936 16747 13004 16803
rect 13060 16747 13100 16803
rect 12592 16679 13100 16747
rect 12592 16623 12632 16679
rect 12688 16623 12756 16679
rect 12812 16623 12880 16679
rect 12936 16623 13004 16679
rect 13060 16623 13100 16679
rect 12592 16555 13100 16623
rect 12592 16499 12632 16555
rect 12688 16499 12756 16555
rect 12812 16499 12880 16555
rect 12936 16499 13004 16555
rect 13060 16499 13100 16555
rect 12592 16431 13100 16499
rect 12592 16375 12632 16431
rect 12688 16375 12756 16431
rect 12812 16375 12880 16431
rect 12936 16375 13004 16431
rect 13060 16375 13100 16431
rect 12592 16307 13100 16375
rect 12592 16251 12632 16307
rect 12688 16251 12756 16307
rect 12812 16251 12880 16307
rect 12936 16251 13004 16307
rect 13060 16251 13100 16307
rect 12592 16183 13100 16251
rect 12592 16127 12632 16183
rect 12688 16127 12756 16183
rect 12812 16127 12880 16183
rect 12936 16127 13004 16183
rect 13060 16127 13100 16183
rect 12592 16059 13100 16127
rect 12592 16003 12632 16059
rect 12688 16003 12756 16059
rect 12812 16003 12880 16059
rect 12936 16003 13004 16059
rect 13060 16003 13100 16059
rect 12592 15935 13100 16003
rect 12592 15879 12632 15935
rect 12688 15879 12756 15935
rect 12812 15879 12880 15935
rect 12936 15879 13004 15935
rect 13060 15879 13100 15935
rect 12592 15811 13100 15879
rect 12592 15762 12632 15811
rect 11356 15755 11366 15762
rect 10918 15687 11366 15755
rect 10918 15631 10928 15687
rect 10984 15631 11052 15687
rect 11108 15631 11176 15687
rect 11232 15631 11300 15687
rect 11356 15631 11366 15687
rect 10918 15563 11366 15631
rect 10918 15507 10928 15563
rect 10984 15507 11052 15563
rect 11108 15507 11176 15563
rect 11232 15507 11300 15563
rect 11356 15507 11366 15563
rect 10918 15439 11366 15507
rect 10918 15383 10928 15439
rect 10984 15383 11052 15439
rect 11108 15383 11176 15439
rect 11232 15383 11300 15439
rect 11356 15383 11366 15439
rect 10918 15315 11366 15383
rect 10918 15259 10928 15315
rect 10984 15259 11052 15315
rect 11108 15259 11176 15315
rect 11232 15259 11300 15315
rect 11356 15259 11366 15315
rect 10918 15191 11366 15259
rect 10918 15135 10928 15191
rect 10984 15135 11052 15191
rect 11108 15135 11176 15191
rect 11232 15135 11300 15191
rect 11356 15135 11366 15191
rect 10918 15067 11366 15135
rect 10918 15011 10928 15067
rect 10984 15011 11052 15067
rect 11108 15011 11176 15067
rect 11232 15011 11300 15067
rect 11356 15011 11366 15067
rect 10918 14943 11366 15011
rect 10918 14887 10928 14943
rect 10984 14887 11052 14943
rect 11108 14887 11176 14943
rect 11232 14887 11300 14943
rect 11356 14887 11366 14943
rect 10918 14819 11366 14887
rect 10918 14763 10928 14819
rect 10984 14763 11052 14819
rect 11108 14763 11176 14819
rect 11232 14763 11300 14819
rect 11356 14763 11366 14819
rect 10918 14695 11366 14763
rect 10918 14639 10928 14695
rect 10984 14639 11052 14695
rect 11108 14639 11176 14695
rect 11232 14639 11300 14695
rect 11356 14639 11366 14695
rect 10918 14571 11366 14639
rect 10918 14515 10928 14571
rect 10984 14515 11052 14571
rect 11108 14515 11176 14571
rect 11232 14515 11300 14571
rect 11356 14515 11366 14571
rect 10918 14447 11366 14515
rect 10918 14391 10928 14447
rect 10984 14391 11052 14447
rect 11108 14391 11176 14447
rect 11232 14391 11300 14447
rect 11356 14391 11366 14447
rect 10918 14323 11366 14391
rect 10918 14267 10928 14323
rect 10984 14267 11052 14323
rect 11108 14267 11176 14323
rect 11232 14267 11300 14323
rect 11356 14267 11366 14323
rect 10918 14199 11366 14267
rect 10918 14143 10928 14199
rect 10984 14143 11052 14199
rect 11108 14143 11176 14199
rect 11232 14143 11300 14199
rect 11356 14143 11366 14199
rect 10918 14133 11366 14143
rect 12622 15755 12632 15762
rect 12688 15755 12756 15811
rect 12812 15755 12880 15811
rect 12936 15755 13004 15811
rect 13060 15762 13100 15811
rect 13160 36251 13668 36260
rect 13160 36195 13200 36251
rect 13256 36195 13324 36251
rect 13380 36195 13448 36251
rect 13504 36195 13572 36251
rect 13628 36195 13668 36251
rect 13160 36127 13668 36195
rect 13160 36071 13200 36127
rect 13256 36071 13324 36127
rect 13380 36071 13448 36127
rect 13504 36071 13572 36127
rect 13628 36071 13668 36127
rect 13160 36003 13668 36071
rect 13160 35947 13200 36003
rect 13256 35947 13324 36003
rect 13380 35947 13448 36003
rect 13504 35947 13572 36003
rect 13628 35947 13668 36003
rect 13160 35879 13668 35947
rect 13160 35823 13200 35879
rect 13256 35823 13324 35879
rect 13380 35823 13448 35879
rect 13504 35823 13572 35879
rect 13628 35823 13668 35879
rect 13160 35755 13668 35823
rect 13160 35699 13200 35755
rect 13256 35699 13324 35755
rect 13380 35699 13448 35755
rect 13504 35699 13572 35755
rect 13628 35699 13668 35755
rect 13160 35631 13668 35699
rect 13160 35575 13200 35631
rect 13256 35575 13324 35631
rect 13380 35575 13448 35631
rect 13504 35575 13572 35631
rect 13628 35575 13668 35631
rect 13160 35507 13668 35575
rect 13160 35451 13200 35507
rect 13256 35451 13324 35507
rect 13380 35451 13448 35507
rect 13504 35451 13572 35507
rect 13628 35451 13668 35507
rect 13160 35383 13668 35451
rect 13160 35327 13200 35383
rect 13256 35327 13324 35383
rect 13380 35327 13448 35383
rect 13504 35327 13572 35383
rect 13628 35327 13668 35383
rect 13160 35259 13668 35327
rect 13160 35203 13200 35259
rect 13256 35203 13324 35259
rect 13380 35203 13448 35259
rect 13504 35203 13572 35259
rect 13628 35203 13668 35259
rect 13160 35135 13668 35203
rect 13160 35079 13200 35135
rect 13256 35079 13324 35135
rect 13380 35079 13448 35135
rect 13504 35079 13572 35135
rect 13628 35079 13668 35135
rect 13160 35011 13668 35079
rect 13160 34955 13200 35011
rect 13256 34955 13324 35011
rect 13380 34955 13448 35011
rect 13504 34955 13572 35011
rect 13628 34955 13668 35011
rect 13160 34887 13668 34955
rect 13160 34831 13200 34887
rect 13256 34831 13324 34887
rect 13380 34831 13448 34887
rect 13504 34831 13572 34887
rect 13628 34831 13668 34887
rect 13160 34763 13668 34831
rect 13160 34707 13200 34763
rect 13256 34707 13324 34763
rect 13380 34707 13448 34763
rect 13504 34707 13572 34763
rect 13628 34707 13668 34763
rect 13160 34639 13668 34707
rect 13160 34583 13200 34639
rect 13256 34583 13324 34639
rect 13380 34583 13448 34639
rect 13504 34583 13572 34639
rect 13628 34583 13668 34639
rect 13160 34515 13668 34583
rect 13160 34459 13200 34515
rect 13256 34459 13324 34515
rect 13380 34459 13448 34515
rect 13504 34459 13572 34515
rect 13628 34459 13668 34515
rect 13160 34391 13668 34459
rect 13160 34335 13200 34391
rect 13256 34335 13324 34391
rect 13380 34335 13448 34391
rect 13504 34335 13572 34391
rect 13628 34335 13668 34391
rect 13160 34267 13668 34335
rect 13160 34211 13200 34267
rect 13256 34211 13324 34267
rect 13380 34211 13448 34267
rect 13504 34211 13572 34267
rect 13628 34211 13668 34267
rect 13160 34143 13668 34211
rect 13160 34087 13200 34143
rect 13256 34087 13324 34143
rect 13380 34087 13448 34143
rect 13504 34087 13572 34143
rect 13628 34087 13668 34143
rect 13160 34019 13668 34087
rect 13160 33963 13200 34019
rect 13256 33963 13324 34019
rect 13380 33963 13448 34019
rect 13504 33963 13572 34019
rect 13628 33963 13668 34019
rect 13160 33895 13668 33963
rect 13160 33839 13200 33895
rect 13256 33839 13324 33895
rect 13380 33839 13448 33895
rect 13504 33839 13572 33895
rect 13628 33839 13668 33895
rect 13160 33771 13668 33839
rect 13160 33715 13200 33771
rect 13256 33715 13324 33771
rect 13380 33715 13448 33771
rect 13504 33715 13572 33771
rect 13628 33715 13668 33771
rect 13160 33647 13668 33715
rect 13160 33591 13200 33647
rect 13256 33591 13324 33647
rect 13380 33591 13448 33647
rect 13504 33591 13572 33647
rect 13628 33591 13668 33647
rect 13160 33523 13668 33591
rect 13160 33467 13200 33523
rect 13256 33467 13324 33523
rect 13380 33467 13448 33523
rect 13504 33467 13572 33523
rect 13628 33467 13668 33523
rect 13160 33399 13668 33467
rect 13160 33343 13200 33399
rect 13256 33343 13324 33399
rect 13380 33343 13448 33399
rect 13504 33343 13572 33399
rect 13628 33343 13668 33399
rect 13160 33308 13668 33343
rect 13160 33256 13202 33308
rect 13254 33256 13326 33308
rect 13378 33256 13450 33308
rect 13502 33256 13574 33308
rect 13626 33256 13668 33308
rect 13160 33184 13668 33256
rect 13160 33132 13202 33184
rect 13254 33132 13326 33184
rect 13378 33132 13450 33184
rect 13502 33132 13574 33184
rect 13626 33132 13668 33184
rect 13160 33060 13668 33132
rect 13160 33008 13202 33060
rect 13254 33008 13326 33060
rect 13378 33008 13450 33060
rect 13502 33008 13574 33060
rect 13626 33008 13668 33060
rect 13160 32936 13668 33008
rect 13160 32884 13202 32936
rect 13254 32884 13326 32936
rect 13378 32884 13450 32936
rect 13502 32884 13574 32936
rect 13626 32884 13668 32936
rect 13160 32812 13668 32884
rect 13160 32760 13202 32812
rect 13254 32760 13326 32812
rect 13378 32760 13450 32812
rect 13502 32760 13574 32812
rect 13626 32760 13668 32812
rect 13160 29360 13668 32760
rect 13160 29308 13202 29360
rect 13254 29308 13326 29360
rect 13378 29308 13450 29360
rect 13502 29308 13574 29360
rect 13626 29308 13668 29360
rect 13160 29236 13668 29308
rect 13160 29184 13202 29236
rect 13254 29184 13326 29236
rect 13378 29184 13450 29236
rect 13502 29184 13574 29236
rect 13626 29184 13668 29236
rect 13160 29112 13668 29184
rect 13160 29060 13202 29112
rect 13254 29060 13326 29112
rect 13378 29060 13450 29112
rect 13502 29060 13574 29112
rect 13626 29060 13668 29112
rect 13160 28988 13668 29060
rect 13160 28936 13202 28988
rect 13254 28936 13326 28988
rect 13378 28936 13450 28988
rect 13502 28936 13574 28988
rect 13626 28936 13668 28988
rect 13160 28864 13668 28936
rect 13160 28812 13202 28864
rect 13254 28812 13326 28864
rect 13378 28812 13450 28864
rect 13502 28812 13574 28864
rect 13626 28812 13668 28864
rect 13160 28245 13668 28812
rect 13160 28189 13200 28245
rect 13256 28189 13324 28245
rect 13380 28189 13448 28245
rect 13504 28189 13572 28245
rect 13628 28189 13668 28245
rect 13160 28121 13668 28189
rect 13160 28065 13200 28121
rect 13256 28065 13324 28121
rect 13380 28065 13448 28121
rect 13504 28065 13572 28121
rect 13628 28065 13668 28121
rect 13160 27997 13668 28065
rect 13160 27941 13200 27997
rect 13256 27941 13324 27997
rect 13380 27941 13448 27997
rect 13504 27941 13572 27997
rect 13628 27941 13668 27997
rect 13160 27873 13668 27941
rect 13160 27817 13200 27873
rect 13256 27817 13324 27873
rect 13380 27817 13448 27873
rect 13504 27817 13572 27873
rect 13628 27817 13668 27873
rect 13160 27749 13668 27817
rect 13160 27693 13200 27749
rect 13256 27693 13324 27749
rect 13380 27693 13448 27749
rect 13504 27693 13572 27749
rect 13628 27693 13668 27749
rect 13160 27625 13668 27693
rect 13160 27569 13200 27625
rect 13256 27569 13324 27625
rect 13380 27569 13448 27625
rect 13504 27569 13572 27625
rect 13628 27569 13668 27625
rect 13160 27501 13668 27569
rect 13160 27445 13200 27501
rect 13256 27445 13324 27501
rect 13380 27445 13448 27501
rect 13504 27445 13572 27501
rect 13628 27445 13668 27501
rect 13160 27377 13668 27445
rect 13160 27321 13200 27377
rect 13256 27321 13324 27377
rect 13380 27321 13448 27377
rect 13504 27321 13572 27377
rect 13628 27321 13668 27377
rect 13160 27253 13668 27321
rect 13160 27197 13200 27253
rect 13256 27197 13324 27253
rect 13380 27197 13448 27253
rect 13504 27197 13572 27253
rect 13628 27197 13668 27253
rect 13160 27129 13668 27197
rect 13160 27073 13200 27129
rect 13256 27073 13324 27129
rect 13380 27073 13448 27129
rect 13504 27073 13572 27129
rect 13628 27073 13668 27129
rect 13160 27005 13668 27073
rect 13160 26949 13200 27005
rect 13256 26949 13324 27005
rect 13380 26949 13448 27005
rect 13504 26949 13572 27005
rect 13628 26949 13668 27005
rect 13160 25412 13668 26949
rect 13160 25360 13202 25412
rect 13254 25360 13326 25412
rect 13378 25360 13450 25412
rect 13502 25360 13574 25412
rect 13626 25360 13668 25412
rect 13160 25288 13668 25360
rect 13160 25236 13202 25288
rect 13254 25236 13326 25288
rect 13378 25236 13450 25288
rect 13502 25236 13574 25288
rect 13626 25236 13668 25288
rect 13160 25164 13668 25236
rect 13160 25112 13202 25164
rect 13254 25112 13326 25164
rect 13378 25112 13450 25164
rect 13502 25112 13574 25164
rect 13626 25112 13668 25164
rect 13160 25040 13668 25112
rect 13160 24988 13202 25040
rect 13254 24988 13326 25040
rect 13378 24988 13450 25040
rect 13502 24988 13574 25040
rect 13626 24988 13668 25040
rect 13160 24916 13668 24988
rect 13160 24864 13202 24916
rect 13254 24864 13326 24916
rect 13378 24864 13450 24916
rect 13502 24864 13574 24916
rect 13626 24864 13668 24916
rect 13160 21469 13668 24864
rect 13160 21417 13172 21469
rect 13224 21417 13280 21469
rect 13332 21417 13388 21469
rect 13440 21417 13496 21469
rect 13548 21417 13604 21469
rect 13656 21417 13668 21469
rect 13160 21361 13668 21417
rect 13160 21309 13172 21361
rect 13224 21309 13280 21361
rect 13332 21309 13388 21361
rect 13440 21309 13496 21361
rect 13548 21309 13604 21361
rect 13656 21309 13668 21361
rect 13160 21253 13668 21309
rect 13160 21201 13172 21253
rect 13224 21201 13280 21253
rect 13332 21201 13388 21253
rect 13440 21201 13496 21253
rect 13548 21201 13604 21253
rect 13656 21201 13668 21253
rect 13160 15762 13668 21201
rect 13728 56324 14236 56975
rect 13728 56272 13786 56324
rect 13838 56272 13910 56324
rect 13962 56272 14034 56324
rect 14086 56272 14236 56324
rect 13728 56200 14236 56272
rect 13728 56148 13786 56200
rect 13838 56148 13910 56200
rect 13962 56148 14034 56200
rect 14086 56148 14236 56200
rect 13728 56076 14236 56148
rect 13728 56024 13786 56076
rect 13838 56024 13910 56076
rect 13962 56024 14034 56076
rect 14086 56024 14236 56076
rect 13728 55952 14236 56024
rect 13728 55900 13786 55952
rect 13838 55900 13910 55952
rect 13962 55900 14034 55952
rect 14086 55900 14236 55952
rect 13728 55828 14236 55900
rect 13728 55776 13786 55828
rect 13838 55776 13910 55828
rect 13962 55776 14034 55828
rect 14086 55776 14236 55828
rect 13728 55704 14236 55776
rect 13728 55652 13786 55704
rect 13838 55652 13910 55704
rect 13962 55652 14034 55704
rect 14086 55652 14236 55704
rect 13728 55580 14236 55652
rect 13728 55528 13786 55580
rect 13838 55528 13910 55580
rect 13962 55528 14034 55580
rect 14086 55528 14236 55580
rect 13728 55456 14236 55528
rect 13728 55445 13786 55456
rect 13838 55445 13910 55456
rect 13962 55445 14034 55456
rect 14086 55445 14236 55456
rect 13728 55389 13768 55445
rect 13838 55404 13892 55445
rect 13962 55404 14016 55445
rect 14086 55404 14140 55445
rect 13824 55389 13892 55404
rect 13948 55389 14016 55404
rect 14072 55389 14140 55404
rect 14196 55389 14236 55445
rect 13728 55332 14236 55389
rect 13728 55321 13786 55332
rect 13838 55321 13910 55332
rect 13962 55321 14034 55332
rect 14086 55321 14236 55332
rect 13728 55265 13768 55321
rect 13838 55280 13892 55321
rect 13962 55280 14016 55321
rect 14086 55280 14140 55321
rect 13824 55265 13892 55280
rect 13948 55265 14016 55280
rect 14072 55265 14140 55280
rect 14196 55265 14236 55321
rect 13728 55208 14236 55265
rect 13728 55197 13786 55208
rect 13838 55197 13910 55208
rect 13962 55197 14034 55208
rect 14086 55197 14236 55208
rect 13728 55141 13768 55197
rect 13838 55156 13892 55197
rect 13962 55156 14016 55197
rect 14086 55156 14140 55197
rect 13824 55141 13892 55156
rect 13948 55141 14016 55156
rect 14072 55141 14140 55156
rect 14196 55141 14236 55197
rect 13728 55084 14236 55141
rect 13728 55073 13786 55084
rect 13838 55073 13910 55084
rect 13962 55073 14034 55084
rect 14086 55073 14236 55084
rect 13728 55017 13768 55073
rect 13838 55032 13892 55073
rect 13962 55032 14016 55073
rect 14086 55032 14140 55073
rect 13824 55017 13892 55032
rect 13948 55017 14016 55032
rect 14072 55017 14140 55032
rect 14196 55017 14236 55073
rect 13728 54960 14236 55017
rect 13728 54949 13786 54960
rect 13838 54949 13910 54960
rect 13962 54949 14034 54960
rect 14086 54949 14236 54960
rect 13728 54893 13768 54949
rect 13838 54908 13892 54949
rect 13962 54908 14016 54949
rect 14086 54908 14140 54949
rect 13824 54893 13892 54908
rect 13948 54893 14016 54908
rect 14072 54893 14140 54908
rect 14196 54893 14236 54949
rect 13728 54836 14236 54893
rect 13728 54825 13786 54836
rect 13838 54825 13910 54836
rect 13962 54825 14034 54836
rect 14086 54825 14236 54836
rect 13728 54769 13768 54825
rect 13838 54784 13892 54825
rect 13962 54784 14016 54825
rect 14086 54784 14140 54825
rect 13824 54769 13892 54784
rect 13948 54769 14016 54784
rect 14072 54769 14140 54784
rect 14196 54769 14236 54825
rect 13728 54712 14236 54769
rect 13728 54701 13786 54712
rect 13838 54701 13910 54712
rect 13962 54701 14034 54712
rect 14086 54701 14236 54712
rect 13728 54645 13768 54701
rect 13838 54660 13892 54701
rect 13962 54660 14016 54701
rect 14086 54660 14140 54701
rect 13824 54645 13892 54660
rect 13948 54645 14016 54660
rect 14072 54645 14140 54660
rect 14196 54645 14236 54701
rect 13728 54588 14236 54645
rect 13728 54577 13786 54588
rect 13838 54577 13910 54588
rect 13962 54577 14034 54588
rect 14086 54577 14236 54588
rect 13728 54521 13768 54577
rect 13838 54536 13892 54577
rect 13962 54536 14016 54577
rect 14086 54536 14140 54577
rect 13824 54521 13892 54536
rect 13948 54521 14016 54536
rect 14072 54521 14140 54536
rect 14196 54521 14236 54577
rect 13728 54464 14236 54521
rect 13728 54453 13786 54464
rect 13838 54453 13910 54464
rect 13962 54453 14034 54464
rect 14086 54453 14236 54464
rect 13728 54397 13768 54453
rect 13838 54412 13892 54453
rect 13962 54412 14016 54453
rect 14086 54412 14140 54453
rect 13824 54397 13892 54412
rect 13948 54397 14016 54412
rect 14072 54397 14140 54412
rect 14196 54397 14236 54453
rect 13728 54340 14236 54397
rect 13728 54329 13786 54340
rect 13838 54329 13910 54340
rect 13962 54329 14034 54340
rect 14086 54329 14236 54340
rect 13728 54273 13768 54329
rect 13838 54288 13892 54329
rect 13962 54288 14016 54329
rect 14086 54288 14140 54329
rect 13824 54273 13892 54288
rect 13948 54273 14016 54288
rect 14072 54273 14140 54288
rect 14196 54273 14236 54329
rect 13728 54216 14236 54273
rect 13728 54205 13786 54216
rect 13838 54205 13910 54216
rect 13962 54205 14034 54216
rect 14086 54205 14236 54216
rect 13728 54149 13768 54205
rect 13838 54164 13892 54205
rect 13962 54164 14016 54205
rect 14086 54164 14140 54205
rect 13824 54149 13892 54164
rect 13948 54149 14016 54164
rect 14072 54149 14140 54164
rect 14196 54149 14236 54205
rect 13728 54092 14236 54149
rect 13728 54040 13786 54092
rect 13838 54040 13910 54092
rect 13962 54040 14034 54092
rect 14086 54040 14236 54092
rect 13728 53968 14236 54040
rect 13728 53916 13786 53968
rect 13838 53916 13910 53968
rect 13962 53916 14034 53968
rect 14086 53916 14236 53968
rect 13728 53844 14236 53916
rect 13728 53792 13786 53844
rect 13838 53792 13910 53844
rect 13962 53792 14034 53844
rect 14086 53792 14236 53844
rect 13728 53720 14236 53792
rect 13728 53668 13786 53720
rect 13838 53668 13910 53720
rect 13962 53668 14034 53720
rect 14086 53668 14236 53720
rect 13728 53596 14236 53668
rect 13728 53544 13786 53596
rect 13838 53544 13910 53596
rect 13962 53544 14034 53596
rect 14086 53544 14236 53596
rect 13728 53472 14236 53544
rect 13728 53420 13786 53472
rect 13838 53420 13910 53472
rect 13962 53420 14034 53472
rect 14086 53420 14236 53472
rect 13728 53348 14236 53420
rect 13728 53296 13786 53348
rect 13838 53296 13910 53348
rect 13962 53296 14034 53348
rect 14086 53296 14236 53348
rect 13728 53224 14236 53296
rect 13728 53172 13786 53224
rect 13838 53172 13910 53224
rect 13962 53172 14034 53224
rect 14086 53172 14236 53224
rect 13728 52376 14236 53172
rect 13728 52324 13786 52376
rect 13838 52324 13910 52376
rect 13962 52324 14034 52376
rect 14086 52324 14236 52376
rect 13728 52252 14236 52324
rect 13728 52200 13786 52252
rect 13838 52200 13910 52252
rect 13962 52200 14034 52252
rect 14086 52200 14236 52252
rect 13728 52128 14236 52200
rect 13728 52076 13786 52128
rect 13838 52076 13910 52128
rect 13962 52076 14034 52128
rect 14086 52076 14236 52128
rect 13728 52004 14236 52076
rect 13728 51952 13786 52004
rect 13838 51952 13910 52004
rect 13962 51952 14034 52004
rect 14086 51952 14236 52004
rect 13728 51880 14236 51952
rect 13728 51828 13786 51880
rect 13838 51828 13910 51880
rect 13962 51828 14034 51880
rect 14086 51828 14236 51880
rect 13728 51756 14236 51828
rect 13728 51704 13786 51756
rect 13838 51704 13910 51756
rect 13962 51704 14034 51756
rect 14086 51704 14236 51756
rect 13728 51632 14236 51704
rect 13728 51580 13786 51632
rect 13838 51580 13910 51632
rect 13962 51580 14034 51632
rect 14086 51580 14236 51632
rect 13728 51508 14236 51580
rect 13728 51456 13786 51508
rect 13838 51456 13910 51508
rect 13962 51456 14034 51508
rect 14086 51456 14236 51508
rect 13728 51384 14236 51456
rect 13728 51332 13786 51384
rect 13838 51332 13910 51384
rect 13962 51332 14034 51384
rect 14086 51332 14236 51384
rect 13728 51260 14236 51332
rect 13728 51208 13786 51260
rect 13838 51208 13910 51260
rect 13962 51208 14034 51260
rect 14086 51208 14236 51260
rect 13728 51136 14236 51208
rect 13728 51084 13786 51136
rect 13838 51084 13910 51136
rect 13962 51084 14034 51136
rect 14086 51084 14236 51136
rect 13728 51012 14236 51084
rect 13728 50960 13786 51012
rect 13838 50960 13910 51012
rect 13962 50960 14034 51012
rect 14086 50960 14236 51012
rect 13728 50888 14236 50960
rect 13728 50836 13786 50888
rect 13838 50836 13910 50888
rect 13962 50836 14034 50888
rect 14086 50836 14236 50888
rect 13728 50764 14236 50836
rect 13728 50712 13786 50764
rect 13838 50712 13910 50764
rect 13962 50712 14034 50764
rect 14086 50712 14236 50764
rect 13728 50640 14236 50712
rect 13728 50588 13786 50640
rect 13838 50588 13910 50640
rect 13962 50588 14034 50640
rect 14086 50588 14236 50640
rect 13728 50516 14236 50588
rect 13728 50464 13786 50516
rect 13838 50464 13910 50516
rect 13962 50464 14034 50516
rect 14086 50464 14236 50516
rect 13728 50392 14236 50464
rect 13728 50340 13786 50392
rect 13838 50340 13910 50392
rect 13962 50340 14034 50392
rect 14086 50340 14236 50392
rect 13728 50268 14236 50340
rect 13728 50216 13786 50268
rect 13838 50216 13910 50268
rect 13962 50216 14034 50268
rect 14086 50216 14236 50268
rect 13728 50144 14236 50216
rect 13728 50092 13786 50144
rect 13838 50092 13910 50144
rect 13962 50092 14034 50144
rect 14086 50092 14236 50144
rect 13728 50020 14236 50092
rect 13728 49968 13786 50020
rect 13838 49968 13910 50020
rect 13962 49968 14034 50020
rect 14086 49968 14236 50020
rect 13728 49896 14236 49968
rect 13728 49844 13786 49896
rect 13838 49844 13910 49896
rect 13962 49844 14034 49896
rect 14086 49844 14236 49896
rect 13728 49772 14236 49844
rect 13728 49720 13786 49772
rect 13838 49720 13910 49772
rect 13962 49720 14034 49772
rect 14086 49720 14236 49772
rect 13728 49648 14236 49720
rect 13728 49596 13786 49648
rect 13838 49596 13910 49648
rect 13962 49596 14034 49648
rect 14086 49596 14236 49648
rect 13728 49524 14236 49596
rect 13728 49472 13786 49524
rect 13838 49472 13910 49524
rect 13962 49472 14034 49524
rect 14086 49472 14236 49524
rect 13728 49400 14236 49472
rect 13728 49348 13786 49400
rect 13838 49348 13910 49400
rect 13962 49348 14034 49400
rect 14086 49348 14236 49400
rect 13728 49276 14236 49348
rect 13728 49224 13786 49276
rect 13838 49224 13910 49276
rect 13962 49224 14034 49276
rect 14086 49224 14236 49276
rect 13728 48428 14236 49224
rect 13728 48376 13786 48428
rect 13838 48376 13910 48428
rect 13962 48376 14034 48428
rect 14086 48376 14236 48428
rect 13728 48304 14236 48376
rect 13728 48252 13786 48304
rect 13838 48252 13910 48304
rect 13962 48252 14034 48304
rect 14086 48252 14236 48304
rect 13728 48180 14236 48252
rect 13728 48128 13786 48180
rect 13838 48128 13910 48180
rect 13962 48128 14034 48180
rect 14086 48128 14236 48180
rect 13728 48056 14236 48128
rect 13728 48004 13786 48056
rect 13838 48004 13910 48056
rect 13962 48004 14034 48056
rect 14086 48004 14236 48056
rect 13728 47932 14236 48004
rect 13728 47880 13786 47932
rect 13838 47880 13910 47932
rect 13962 47880 14034 47932
rect 14086 47880 14236 47932
rect 13728 47808 14236 47880
rect 13728 47756 13786 47808
rect 13838 47756 13910 47808
rect 13962 47756 14034 47808
rect 14086 47756 14236 47808
rect 13728 47684 14236 47756
rect 13728 47632 13786 47684
rect 13838 47632 13910 47684
rect 13962 47632 14034 47684
rect 14086 47632 14236 47684
rect 13728 47560 14236 47632
rect 13728 47508 13786 47560
rect 13838 47508 13910 47560
rect 13962 47508 14034 47560
rect 14086 47508 14236 47560
rect 13728 47445 14236 47508
rect 13728 47389 13768 47445
rect 13824 47436 13892 47445
rect 13948 47436 14016 47445
rect 14072 47436 14140 47445
rect 13838 47389 13892 47436
rect 13962 47389 14016 47436
rect 14086 47389 14140 47436
rect 14196 47389 14236 47445
rect 13728 47384 13786 47389
rect 13838 47384 13910 47389
rect 13962 47384 14034 47389
rect 14086 47384 14236 47389
rect 13728 47321 14236 47384
rect 13728 47265 13768 47321
rect 13824 47312 13892 47321
rect 13948 47312 14016 47321
rect 14072 47312 14140 47321
rect 13838 47265 13892 47312
rect 13962 47265 14016 47312
rect 14086 47265 14140 47312
rect 14196 47265 14236 47321
rect 13728 47260 13786 47265
rect 13838 47260 13910 47265
rect 13962 47260 14034 47265
rect 14086 47260 14236 47265
rect 13728 47197 14236 47260
rect 13728 47141 13768 47197
rect 13824 47188 13892 47197
rect 13948 47188 14016 47197
rect 14072 47188 14140 47197
rect 13838 47141 13892 47188
rect 13962 47141 14016 47188
rect 14086 47141 14140 47188
rect 14196 47141 14236 47197
rect 13728 47136 13786 47141
rect 13838 47136 13910 47141
rect 13962 47136 14034 47141
rect 14086 47136 14236 47141
rect 13728 47073 14236 47136
rect 13728 47017 13768 47073
rect 13824 47064 13892 47073
rect 13948 47064 14016 47073
rect 14072 47064 14140 47073
rect 13838 47017 13892 47064
rect 13962 47017 14016 47064
rect 14086 47017 14140 47064
rect 14196 47017 14236 47073
rect 13728 47012 13786 47017
rect 13838 47012 13910 47017
rect 13962 47012 14034 47017
rect 14086 47012 14236 47017
rect 13728 46949 14236 47012
rect 13728 46893 13768 46949
rect 13824 46940 13892 46949
rect 13948 46940 14016 46949
rect 14072 46940 14140 46949
rect 13838 46893 13892 46940
rect 13962 46893 14016 46940
rect 14086 46893 14140 46940
rect 14196 46893 14236 46949
rect 13728 46888 13786 46893
rect 13838 46888 13910 46893
rect 13962 46888 14034 46893
rect 14086 46888 14236 46893
rect 13728 46825 14236 46888
rect 13728 46769 13768 46825
rect 13824 46816 13892 46825
rect 13948 46816 14016 46825
rect 14072 46816 14140 46825
rect 13838 46769 13892 46816
rect 13962 46769 14016 46816
rect 14086 46769 14140 46816
rect 14196 46769 14236 46825
rect 13728 46764 13786 46769
rect 13838 46764 13910 46769
rect 13962 46764 14034 46769
rect 14086 46764 14236 46769
rect 13728 46701 14236 46764
rect 13728 46645 13768 46701
rect 13824 46692 13892 46701
rect 13948 46692 14016 46701
rect 14072 46692 14140 46701
rect 13838 46645 13892 46692
rect 13962 46645 14016 46692
rect 14086 46645 14140 46692
rect 14196 46645 14236 46701
rect 13728 46640 13786 46645
rect 13838 46640 13910 46645
rect 13962 46640 14034 46645
rect 14086 46640 14236 46645
rect 13728 46577 14236 46640
rect 13728 46521 13768 46577
rect 13824 46568 13892 46577
rect 13948 46568 14016 46577
rect 14072 46568 14140 46577
rect 13838 46521 13892 46568
rect 13962 46521 14016 46568
rect 14086 46521 14140 46568
rect 14196 46521 14236 46577
rect 13728 46516 13786 46521
rect 13838 46516 13910 46521
rect 13962 46516 14034 46521
rect 14086 46516 14236 46521
rect 13728 46453 14236 46516
rect 13728 46397 13768 46453
rect 13824 46444 13892 46453
rect 13948 46444 14016 46453
rect 14072 46444 14140 46453
rect 13838 46397 13892 46444
rect 13962 46397 14016 46444
rect 14086 46397 14140 46444
rect 14196 46397 14236 46453
rect 13728 46392 13786 46397
rect 13838 46392 13910 46397
rect 13962 46392 14034 46397
rect 14086 46392 14236 46397
rect 13728 46329 14236 46392
rect 13728 46273 13768 46329
rect 13824 46320 13892 46329
rect 13948 46320 14016 46329
rect 14072 46320 14140 46329
rect 13838 46273 13892 46320
rect 13962 46273 14016 46320
rect 14086 46273 14140 46320
rect 14196 46273 14236 46329
rect 13728 46268 13786 46273
rect 13838 46268 13910 46273
rect 13962 46268 14034 46273
rect 14086 46268 14236 46273
rect 13728 46205 14236 46268
rect 13728 46149 13768 46205
rect 13824 46196 13892 46205
rect 13948 46196 14016 46205
rect 14072 46196 14140 46205
rect 13838 46149 13892 46196
rect 13962 46149 14016 46196
rect 14086 46149 14140 46196
rect 14196 46149 14236 46205
rect 13728 46144 13786 46149
rect 13838 46144 13910 46149
rect 13962 46144 14034 46149
rect 14086 46144 14236 46149
rect 13728 46072 14236 46144
rect 13728 46020 13786 46072
rect 13838 46020 13910 46072
rect 13962 46020 14034 46072
rect 14086 46020 14236 46072
rect 13728 45948 14236 46020
rect 13728 45896 13786 45948
rect 13838 45896 13910 45948
rect 13962 45896 14034 45948
rect 14086 45896 14236 45948
rect 13728 45824 14236 45896
rect 13728 45772 13786 45824
rect 13838 45772 13910 45824
rect 13962 45772 14034 45824
rect 14086 45772 14236 45824
rect 13728 45700 14236 45772
rect 13728 45648 13786 45700
rect 13838 45648 13910 45700
rect 13962 45648 14034 45700
rect 14086 45648 14236 45700
rect 13728 45576 14236 45648
rect 13728 45524 13786 45576
rect 13838 45524 13910 45576
rect 13962 45524 14034 45576
rect 14086 45524 14236 45576
rect 13728 45452 14236 45524
rect 13728 45400 13786 45452
rect 13838 45400 13910 45452
rect 13962 45400 14034 45452
rect 14086 45400 14236 45452
rect 13728 45328 14236 45400
rect 13728 45276 13786 45328
rect 13838 45276 13910 45328
rect 13962 45276 14034 45328
rect 14086 45276 14236 45328
rect 13728 44480 14236 45276
rect 13728 44428 13786 44480
rect 13838 44428 13910 44480
rect 13962 44428 14034 44480
rect 14086 44428 14236 44480
rect 13728 44356 14236 44428
rect 13728 44304 13786 44356
rect 13838 44304 13910 44356
rect 13962 44304 14034 44356
rect 14086 44304 14236 44356
rect 13728 44245 14236 44304
rect 13728 44189 13768 44245
rect 13824 44232 13892 44245
rect 13948 44232 14016 44245
rect 14072 44232 14140 44245
rect 13838 44189 13892 44232
rect 13962 44189 14016 44232
rect 14086 44189 14140 44232
rect 14196 44189 14236 44245
rect 13728 44180 13786 44189
rect 13838 44180 13910 44189
rect 13962 44180 14034 44189
rect 14086 44180 14236 44189
rect 13728 44121 14236 44180
rect 13728 44065 13768 44121
rect 13824 44108 13892 44121
rect 13948 44108 14016 44121
rect 14072 44108 14140 44121
rect 13838 44065 13892 44108
rect 13962 44065 14016 44108
rect 14086 44065 14140 44108
rect 14196 44065 14236 44121
rect 13728 44056 13786 44065
rect 13838 44056 13910 44065
rect 13962 44056 14034 44065
rect 14086 44056 14236 44065
rect 13728 43997 14236 44056
rect 13728 43941 13768 43997
rect 13824 43984 13892 43997
rect 13948 43984 14016 43997
rect 14072 43984 14140 43997
rect 13838 43941 13892 43984
rect 13962 43941 14016 43984
rect 14086 43941 14140 43984
rect 14196 43941 14236 43997
rect 13728 43932 13786 43941
rect 13838 43932 13910 43941
rect 13962 43932 14034 43941
rect 14086 43932 14236 43941
rect 13728 43873 14236 43932
rect 13728 43817 13768 43873
rect 13824 43860 13892 43873
rect 13948 43860 14016 43873
rect 14072 43860 14140 43873
rect 13838 43817 13892 43860
rect 13962 43817 14016 43860
rect 14086 43817 14140 43860
rect 14196 43817 14236 43873
rect 13728 43808 13786 43817
rect 13838 43808 13910 43817
rect 13962 43808 14034 43817
rect 14086 43808 14236 43817
rect 13728 43749 14236 43808
rect 13728 43693 13768 43749
rect 13824 43736 13892 43749
rect 13948 43736 14016 43749
rect 14072 43736 14140 43749
rect 13838 43693 13892 43736
rect 13962 43693 14016 43736
rect 14086 43693 14140 43736
rect 14196 43693 14236 43749
rect 13728 43684 13786 43693
rect 13838 43684 13910 43693
rect 13962 43684 14034 43693
rect 14086 43684 14236 43693
rect 13728 43625 14236 43684
rect 13728 43569 13768 43625
rect 13824 43612 13892 43625
rect 13948 43612 14016 43625
rect 14072 43612 14140 43625
rect 13838 43569 13892 43612
rect 13962 43569 14016 43612
rect 14086 43569 14140 43612
rect 14196 43569 14236 43625
rect 13728 43560 13786 43569
rect 13838 43560 13910 43569
rect 13962 43560 14034 43569
rect 14086 43560 14236 43569
rect 13728 43501 14236 43560
rect 13728 43445 13768 43501
rect 13824 43488 13892 43501
rect 13948 43488 14016 43501
rect 14072 43488 14140 43501
rect 13838 43445 13892 43488
rect 13962 43445 14016 43488
rect 14086 43445 14140 43488
rect 14196 43445 14236 43501
rect 13728 43436 13786 43445
rect 13838 43436 13910 43445
rect 13962 43436 14034 43445
rect 14086 43436 14236 43445
rect 13728 43377 14236 43436
rect 13728 43321 13768 43377
rect 13824 43364 13892 43377
rect 13948 43364 14016 43377
rect 14072 43364 14140 43377
rect 13838 43321 13892 43364
rect 13962 43321 14016 43364
rect 14086 43321 14140 43364
rect 14196 43321 14236 43377
rect 13728 43312 13786 43321
rect 13838 43312 13910 43321
rect 13962 43312 14034 43321
rect 14086 43312 14236 43321
rect 13728 43253 14236 43312
rect 13728 43197 13768 43253
rect 13824 43240 13892 43253
rect 13948 43240 14016 43253
rect 14072 43240 14140 43253
rect 13838 43197 13892 43240
rect 13962 43197 14016 43240
rect 14086 43197 14140 43240
rect 14196 43197 14236 43253
rect 13728 43188 13786 43197
rect 13838 43188 13910 43197
rect 13962 43188 14034 43197
rect 14086 43188 14236 43197
rect 13728 43129 14236 43188
rect 13728 43073 13768 43129
rect 13824 43116 13892 43129
rect 13948 43116 14016 43129
rect 14072 43116 14140 43129
rect 13838 43073 13892 43116
rect 13962 43073 14016 43116
rect 14086 43073 14140 43116
rect 14196 43073 14236 43129
rect 13728 43064 13786 43073
rect 13838 43064 13910 43073
rect 13962 43064 14034 43073
rect 14086 43064 14236 43073
rect 13728 43005 14236 43064
rect 13728 42949 13768 43005
rect 13824 42992 13892 43005
rect 13948 42992 14016 43005
rect 14072 42992 14140 43005
rect 13838 42949 13892 42992
rect 13962 42949 14016 42992
rect 14086 42949 14140 42992
rect 14196 42949 14236 43005
rect 13728 42940 13786 42949
rect 13838 42940 13910 42949
rect 13962 42940 14034 42949
rect 14086 42940 14236 42949
rect 13728 42868 14236 42940
rect 13728 42816 13786 42868
rect 13838 42816 13910 42868
rect 13962 42816 14034 42868
rect 14086 42816 14236 42868
rect 13728 42744 14236 42816
rect 13728 42692 13786 42744
rect 13838 42692 13910 42744
rect 13962 42692 14034 42744
rect 14086 42692 14236 42744
rect 13728 42645 14236 42692
rect 13728 42589 13768 42645
rect 13824 42620 13892 42645
rect 13948 42620 14016 42645
rect 14072 42620 14140 42645
rect 13838 42589 13892 42620
rect 13962 42589 14016 42620
rect 14086 42589 14140 42620
rect 14196 42589 14236 42645
rect 13728 42568 13786 42589
rect 13838 42568 13910 42589
rect 13962 42568 14034 42589
rect 14086 42568 14236 42589
rect 13728 42521 14236 42568
rect 13728 42465 13768 42521
rect 13824 42496 13892 42521
rect 13948 42496 14016 42521
rect 14072 42496 14140 42521
rect 13838 42465 13892 42496
rect 13962 42465 14016 42496
rect 14086 42465 14140 42496
rect 14196 42465 14236 42521
rect 13728 42444 13786 42465
rect 13838 42444 13910 42465
rect 13962 42444 14034 42465
rect 14086 42444 14236 42465
rect 13728 42397 14236 42444
rect 13728 42341 13768 42397
rect 13824 42372 13892 42397
rect 13948 42372 14016 42397
rect 14072 42372 14140 42397
rect 13838 42341 13892 42372
rect 13962 42341 14016 42372
rect 14086 42341 14140 42372
rect 14196 42341 14236 42397
rect 13728 42320 13786 42341
rect 13838 42320 13910 42341
rect 13962 42320 14034 42341
rect 14086 42320 14236 42341
rect 13728 42273 14236 42320
rect 13728 42217 13768 42273
rect 13824 42248 13892 42273
rect 13948 42248 14016 42273
rect 14072 42248 14140 42273
rect 13838 42217 13892 42248
rect 13962 42217 14016 42248
rect 14086 42217 14140 42248
rect 14196 42217 14236 42273
rect 13728 42196 13786 42217
rect 13838 42196 13910 42217
rect 13962 42196 14034 42217
rect 14086 42196 14236 42217
rect 13728 42149 14236 42196
rect 13728 42093 13768 42149
rect 13824 42124 13892 42149
rect 13948 42124 14016 42149
rect 14072 42124 14140 42149
rect 13838 42093 13892 42124
rect 13962 42093 14016 42124
rect 14086 42093 14140 42124
rect 14196 42093 14236 42149
rect 13728 42072 13786 42093
rect 13838 42072 13910 42093
rect 13962 42072 14034 42093
rect 14086 42072 14236 42093
rect 13728 42025 14236 42072
rect 13728 41969 13768 42025
rect 13824 42000 13892 42025
rect 13948 42000 14016 42025
rect 14072 42000 14140 42025
rect 13838 41969 13892 42000
rect 13962 41969 14016 42000
rect 14086 41969 14140 42000
rect 14196 41969 14236 42025
rect 13728 41948 13786 41969
rect 13838 41948 13910 41969
rect 13962 41948 14034 41969
rect 14086 41948 14236 41969
rect 13728 41901 14236 41948
rect 13728 41845 13768 41901
rect 13824 41876 13892 41901
rect 13948 41876 14016 41901
rect 14072 41876 14140 41901
rect 13838 41845 13892 41876
rect 13962 41845 14016 41876
rect 14086 41845 14140 41876
rect 14196 41845 14236 41901
rect 13728 41824 13786 41845
rect 13838 41824 13910 41845
rect 13962 41824 14034 41845
rect 14086 41824 14236 41845
rect 13728 41777 14236 41824
rect 13728 41721 13768 41777
rect 13824 41752 13892 41777
rect 13948 41752 14016 41777
rect 14072 41752 14140 41777
rect 13838 41721 13892 41752
rect 13962 41721 14016 41752
rect 14086 41721 14140 41752
rect 14196 41721 14236 41777
rect 13728 41700 13786 41721
rect 13838 41700 13910 41721
rect 13962 41700 14034 41721
rect 14086 41700 14236 41721
rect 13728 41653 14236 41700
rect 13728 41597 13768 41653
rect 13824 41628 13892 41653
rect 13948 41628 14016 41653
rect 14072 41628 14140 41653
rect 13838 41597 13892 41628
rect 13962 41597 14016 41628
rect 14086 41597 14140 41628
rect 14196 41597 14236 41653
rect 13728 41576 13786 41597
rect 13838 41576 13910 41597
rect 13962 41576 14034 41597
rect 14086 41576 14236 41597
rect 13728 41529 14236 41576
rect 13728 41473 13768 41529
rect 13824 41504 13892 41529
rect 13948 41504 14016 41529
rect 14072 41504 14140 41529
rect 13838 41473 13892 41504
rect 13962 41473 14016 41504
rect 14086 41473 14140 41504
rect 14196 41473 14236 41529
rect 13728 41452 13786 41473
rect 13838 41452 13910 41473
rect 13962 41452 14034 41473
rect 14086 41452 14236 41473
rect 13728 41405 14236 41452
rect 13728 41349 13768 41405
rect 13824 41380 13892 41405
rect 13948 41380 14016 41405
rect 14072 41380 14140 41405
rect 13838 41349 13892 41380
rect 13962 41349 14016 41380
rect 14086 41349 14140 41380
rect 14196 41349 14236 41405
rect 13728 41328 13786 41349
rect 13838 41328 13910 41349
rect 13962 41328 14034 41349
rect 14086 41328 14236 41349
rect 13728 41045 14236 41328
rect 13728 40989 13768 41045
rect 13824 40989 13892 41045
rect 13948 40989 14016 41045
rect 14072 40989 14140 41045
rect 14196 40989 14236 41045
rect 13728 40921 14236 40989
rect 13728 40865 13768 40921
rect 13824 40865 13892 40921
rect 13948 40865 14016 40921
rect 14072 40865 14140 40921
rect 14196 40865 14236 40921
rect 13728 40797 14236 40865
rect 13728 40741 13768 40797
rect 13824 40741 13892 40797
rect 13948 40741 14016 40797
rect 14072 40741 14140 40797
rect 14196 40741 14236 40797
rect 13728 40673 14236 40741
rect 13728 40617 13768 40673
rect 13824 40617 13892 40673
rect 13948 40617 14016 40673
rect 14072 40617 14140 40673
rect 14196 40617 14236 40673
rect 13728 40549 14236 40617
rect 13728 40493 13768 40549
rect 13824 40532 13892 40549
rect 13948 40532 14016 40549
rect 14072 40532 14140 40549
rect 13838 40493 13892 40532
rect 13962 40493 14016 40532
rect 14086 40493 14140 40532
rect 14196 40493 14236 40549
rect 13728 40480 13786 40493
rect 13838 40480 13910 40493
rect 13962 40480 14034 40493
rect 14086 40480 14236 40493
rect 13728 40425 14236 40480
rect 13728 40369 13768 40425
rect 13824 40408 13892 40425
rect 13948 40408 14016 40425
rect 14072 40408 14140 40425
rect 13838 40369 13892 40408
rect 13962 40369 14016 40408
rect 14086 40369 14140 40408
rect 14196 40369 14236 40425
rect 13728 40356 13786 40369
rect 13838 40356 13910 40369
rect 13962 40356 14034 40369
rect 14086 40356 14236 40369
rect 13728 40301 14236 40356
rect 13728 40245 13768 40301
rect 13824 40284 13892 40301
rect 13948 40284 14016 40301
rect 14072 40284 14140 40301
rect 13838 40245 13892 40284
rect 13962 40245 14016 40284
rect 14086 40245 14140 40284
rect 14196 40245 14236 40301
rect 13728 40232 13786 40245
rect 13838 40232 13910 40245
rect 13962 40232 14034 40245
rect 14086 40232 14236 40245
rect 13728 40177 14236 40232
rect 13728 40121 13768 40177
rect 13824 40160 13892 40177
rect 13948 40160 14016 40177
rect 14072 40160 14140 40177
rect 13838 40121 13892 40160
rect 13962 40121 14016 40160
rect 14086 40121 14140 40160
rect 14196 40121 14236 40177
rect 13728 40108 13786 40121
rect 13838 40108 13910 40121
rect 13962 40108 14034 40121
rect 14086 40108 14236 40121
rect 13728 40053 14236 40108
rect 13728 39997 13768 40053
rect 13824 40036 13892 40053
rect 13948 40036 14016 40053
rect 14072 40036 14140 40053
rect 13838 39997 13892 40036
rect 13962 39997 14016 40036
rect 14086 39997 14140 40036
rect 14196 39997 14236 40053
rect 13728 39984 13786 39997
rect 13838 39984 13910 39997
rect 13962 39984 14034 39997
rect 14086 39984 14236 39997
rect 13728 39929 14236 39984
rect 13728 39873 13768 39929
rect 13824 39912 13892 39929
rect 13948 39912 14016 39929
rect 14072 39912 14140 39929
rect 13838 39873 13892 39912
rect 13962 39873 14016 39912
rect 14086 39873 14140 39912
rect 14196 39873 14236 39929
rect 13728 39860 13786 39873
rect 13838 39860 13910 39873
rect 13962 39860 14034 39873
rect 14086 39860 14236 39873
rect 13728 39805 14236 39860
rect 13728 39749 13768 39805
rect 13824 39788 13892 39805
rect 13948 39788 14016 39805
rect 14072 39788 14140 39805
rect 13838 39749 13892 39788
rect 13962 39749 14016 39788
rect 14086 39749 14140 39788
rect 14196 39749 14236 39805
rect 13728 39736 13786 39749
rect 13838 39736 13910 39749
rect 13962 39736 14034 39749
rect 14086 39736 14236 39749
rect 13728 39664 14236 39736
rect 13728 39612 13786 39664
rect 13838 39612 13910 39664
rect 13962 39612 14034 39664
rect 14086 39612 14236 39664
rect 13728 39540 14236 39612
rect 13728 39488 13786 39540
rect 13838 39488 13910 39540
rect 13962 39488 14034 39540
rect 14086 39488 14236 39540
rect 13728 39416 14236 39488
rect 13728 39364 13786 39416
rect 13838 39364 13910 39416
rect 13962 39364 14034 39416
rect 14086 39364 14236 39416
rect 13728 39292 14236 39364
rect 13728 39240 13786 39292
rect 13838 39240 13910 39292
rect 13962 39240 14034 39292
rect 14086 39240 14236 39292
rect 13728 39168 14236 39240
rect 13728 39116 13786 39168
rect 13838 39116 13910 39168
rect 13962 39116 14034 39168
rect 14086 39116 14236 39168
rect 13728 39044 14236 39116
rect 13728 38992 13786 39044
rect 13838 38992 13910 39044
rect 13962 38992 14034 39044
rect 14086 38992 14236 39044
rect 13728 38920 14236 38992
rect 13728 38868 13786 38920
rect 13838 38868 13910 38920
rect 13962 38868 14034 38920
rect 14086 38868 14236 38920
rect 13728 38796 14236 38868
rect 13728 38744 13786 38796
rect 13838 38744 13910 38796
rect 13962 38744 14034 38796
rect 14086 38744 14236 38796
rect 13728 38672 14236 38744
rect 13728 38620 13786 38672
rect 13838 38620 13910 38672
rect 13962 38620 14034 38672
rect 14086 38620 14236 38672
rect 13728 38548 14236 38620
rect 13728 38496 13786 38548
rect 13838 38496 13910 38548
rect 13962 38496 14034 38548
rect 14086 38496 14236 38548
rect 13728 38424 14236 38496
rect 13728 38372 13786 38424
rect 13838 38372 13910 38424
rect 13962 38372 14034 38424
rect 14086 38372 14236 38424
rect 13728 38300 14236 38372
rect 13728 38248 13786 38300
rect 13838 38248 13910 38300
rect 13962 38248 14034 38300
rect 14086 38248 14236 38300
rect 13728 38176 14236 38248
rect 13728 38124 13786 38176
rect 13838 38124 13910 38176
rect 13962 38124 14034 38176
rect 14086 38124 14236 38176
rect 13728 38052 14236 38124
rect 13728 38000 13786 38052
rect 13838 38000 13910 38052
rect 13962 38000 14034 38052
rect 14086 38000 14236 38052
rect 13728 37928 14236 38000
rect 13728 37876 13786 37928
rect 13838 37876 13910 37928
rect 13962 37876 14034 37928
rect 14086 37876 14236 37928
rect 13728 37804 14236 37876
rect 13728 37752 13786 37804
rect 13838 37752 13910 37804
rect 13962 37752 14034 37804
rect 14086 37752 14236 37804
rect 13728 37680 14236 37752
rect 13728 37628 13786 37680
rect 13838 37628 13910 37680
rect 13962 37628 14034 37680
rect 14086 37628 14236 37680
rect 13728 37556 14236 37628
rect 13728 37504 13786 37556
rect 13838 37504 13910 37556
rect 13962 37504 14034 37556
rect 14086 37504 14236 37556
rect 13728 37432 14236 37504
rect 13728 37380 13786 37432
rect 13838 37380 13910 37432
rect 13962 37380 14034 37432
rect 14086 37380 14236 37432
rect 13728 36584 14236 37380
rect 13728 36532 13786 36584
rect 13838 36532 13910 36584
rect 13962 36532 14034 36584
rect 14086 36532 14236 36584
rect 13728 36460 14236 36532
rect 13728 36408 13786 36460
rect 13838 36408 13910 36460
rect 13962 36408 14034 36460
rect 14086 36408 14236 36460
rect 13728 36336 14236 36408
rect 13728 36284 13786 36336
rect 13838 36284 13910 36336
rect 13962 36284 14034 36336
rect 14086 36284 14236 36336
rect 13728 36212 14236 36284
rect 13728 36160 13786 36212
rect 13838 36160 13910 36212
rect 13962 36160 14034 36212
rect 14086 36160 14236 36212
rect 13728 36088 14236 36160
rect 13728 36036 13786 36088
rect 13838 36036 13910 36088
rect 13962 36036 14034 36088
rect 14086 36036 14236 36088
rect 13728 35964 14236 36036
rect 13728 35912 13786 35964
rect 13838 35912 13910 35964
rect 13962 35912 14034 35964
rect 14086 35912 14236 35964
rect 13728 35840 14236 35912
rect 13728 35788 13786 35840
rect 13838 35788 13910 35840
rect 13962 35788 14034 35840
rect 14086 35788 14236 35840
rect 13728 35716 14236 35788
rect 13728 35664 13786 35716
rect 13838 35664 13910 35716
rect 13962 35664 14034 35716
rect 14086 35664 14236 35716
rect 13728 35592 14236 35664
rect 13728 35540 13786 35592
rect 13838 35540 13910 35592
rect 13962 35540 14034 35592
rect 14086 35540 14236 35592
rect 13728 35468 14236 35540
rect 13728 35416 13786 35468
rect 13838 35416 13910 35468
rect 13962 35416 14034 35468
rect 14086 35416 14236 35468
rect 13728 35344 14236 35416
rect 13728 35292 13786 35344
rect 13838 35292 13910 35344
rect 13962 35292 14034 35344
rect 14086 35292 14236 35344
rect 13728 35220 14236 35292
rect 13728 35168 13786 35220
rect 13838 35168 13910 35220
rect 13962 35168 14034 35220
rect 14086 35168 14236 35220
rect 13728 35096 14236 35168
rect 13728 35044 13786 35096
rect 13838 35044 13910 35096
rect 13962 35044 14034 35096
rect 14086 35044 14236 35096
rect 13728 34972 14236 35044
rect 13728 34920 13786 34972
rect 13838 34920 13910 34972
rect 13962 34920 14034 34972
rect 14086 34920 14236 34972
rect 13728 34848 14236 34920
rect 13728 34796 13786 34848
rect 13838 34796 13910 34848
rect 13962 34796 14034 34848
rect 14086 34796 14236 34848
rect 13728 34724 14236 34796
rect 13728 34672 13786 34724
rect 13838 34672 13910 34724
rect 13962 34672 14034 34724
rect 14086 34672 14236 34724
rect 13728 34600 14236 34672
rect 13728 34548 13786 34600
rect 13838 34548 13910 34600
rect 13962 34548 14034 34600
rect 14086 34548 14236 34600
rect 13728 34476 14236 34548
rect 13728 34424 13786 34476
rect 13838 34424 13910 34476
rect 13962 34424 14034 34476
rect 14086 34424 14236 34476
rect 13728 34352 14236 34424
rect 13728 34300 13786 34352
rect 13838 34300 13910 34352
rect 13962 34300 14034 34352
rect 14086 34300 14236 34352
rect 13728 34228 14236 34300
rect 13728 34176 13786 34228
rect 13838 34176 13910 34228
rect 13962 34176 14034 34228
rect 14086 34176 14236 34228
rect 13728 34104 14236 34176
rect 13728 34052 13786 34104
rect 13838 34052 13910 34104
rect 13962 34052 14034 34104
rect 14086 34052 14236 34104
rect 13728 33980 14236 34052
rect 13728 33928 13786 33980
rect 13838 33928 13910 33980
rect 13962 33928 14034 33980
rect 14086 33928 14236 33980
rect 13728 33856 14236 33928
rect 13728 33804 13786 33856
rect 13838 33804 13910 33856
rect 13962 33804 14034 33856
rect 14086 33804 14236 33856
rect 13728 33732 14236 33804
rect 13728 33680 13786 33732
rect 13838 33680 13910 33732
rect 13962 33680 14034 33732
rect 14086 33680 14236 33732
rect 13728 33608 14236 33680
rect 13728 33556 13786 33608
rect 13838 33556 13910 33608
rect 13962 33556 14034 33608
rect 14086 33556 14236 33608
rect 13728 33484 14236 33556
rect 13728 33432 13786 33484
rect 13838 33432 13910 33484
rect 13962 33432 14034 33484
rect 14086 33432 14236 33484
rect 13728 33051 14236 33432
rect 13728 32995 13768 33051
rect 13824 32995 13892 33051
rect 13948 32995 14016 33051
rect 14072 32995 14140 33051
rect 14196 32995 14236 33051
rect 13728 32927 14236 32995
rect 13728 32871 13768 32927
rect 13824 32871 13892 32927
rect 13948 32871 14016 32927
rect 14072 32871 14140 32927
rect 14196 32871 14236 32927
rect 13728 32803 14236 32871
rect 13728 32747 13768 32803
rect 13824 32747 13892 32803
rect 13948 32747 14016 32803
rect 14072 32747 14140 32803
rect 14196 32747 14236 32803
rect 13728 32679 14236 32747
rect 13728 32623 13768 32679
rect 13824 32636 13892 32679
rect 13948 32636 14016 32679
rect 14072 32636 14140 32679
rect 13838 32623 13892 32636
rect 13962 32623 14016 32636
rect 14086 32623 14140 32636
rect 14196 32623 14236 32679
rect 13728 32584 13786 32623
rect 13838 32584 13910 32623
rect 13962 32584 14034 32623
rect 14086 32584 14236 32623
rect 13728 32555 14236 32584
rect 13728 32499 13768 32555
rect 13824 32512 13892 32555
rect 13948 32512 14016 32555
rect 14072 32512 14140 32555
rect 13838 32499 13892 32512
rect 13962 32499 14016 32512
rect 14086 32499 14140 32512
rect 14196 32499 14236 32555
rect 13728 32460 13786 32499
rect 13838 32460 13910 32499
rect 13962 32460 14034 32499
rect 14086 32460 14236 32499
rect 13728 32431 14236 32460
rect 13728 32375 13768 32431
rect 13824 32388 13892 32431
rect 13948 32388 14016 32431
rect 14072 32388 14140 32431
rect 13838 32375 13892 32388
rect 13962 32375 14016 32388
rect 14086 32375 14140 32388
rect 14196 32375 14236 32431
rect 13728 32336 13786 32375
rect 13838 32336 13910 32375
rect 13962 32336 14034 32375
rect 14086 32336 14236 32375
rect 13728 32307 14236 32336
rect 13728 32251 13768 32307
rect 13824 32264 13892 32307
rect 13948 32264 14016 32307
rect 14072 32264 14140 32307
rect 13838 32251 13892 32264
rect 13962 32251 14016 32264
rect 14086 32251 14140 32264
rect 14196 32251 14236 32307
rect 13728 32212 13786 32251
rect 13838 32212 13910 32251
rect 13962 32212 14034 32251
rect 14086 32212 14236 32251
rect 13728 32183 14236 32212
rect 13728 32127 13768 32183
rect 13824 32140 13892 32183
rect 13948 32140 14016 32183
rect 14072 32140 14140 32183
rect 13838 32127 13892 32140
rect 13962 32127 14016 32140
rect 14086 32127 14140 32140
rect 14196 32127 14236 32183
rect 13728 32088 13786 32127
rect 13838 32088 13910 32127
rect 13962 32088 14034 32127
rect 14086 32088 14236 32127
rect 13728 32059 14236 32088
rect 13728 32003 13768 32059
rect 13824 32016 13892 32059
rect 13948 32016 14016 32059
rect 14072 32016 14140 32059
rect 13838 32003 13892 32016
rect 13962 32003 14016 32016
rect 14086 32003 14140 32016
rect 14196 32003 14236 32059
rect 13728 31964 13786 32003
rect 13838 31964 13910 32003
rect 13962 31964 14034 32003
rect 14086 31964 14236 32003
rect 13728 31935 14236 31964
rect 13728 31879 13768 31935
rect 13824 31892 13892 31935
rect 13948 31892 14016 31935
rect 14072 31892 14140 31935
rect 13838 31879 13892 31892
rect 13962 31879 14016 31892
rect 14086 31879 14140 31892
rect 14196 31879 14236 31935
rect 13728 31840 13786 31879
rect 13838 31840 13910 31879
rect 13962 31840 14034 31879
rect 14086 31840 14236 31879
rect 13728 31811 14236 31840
rect 13728 31755 13768 31811
rect 13824 31768 13892 31811
rect 13948 31768 14016 31811
rect 14072 31768 14140 31811
rect 13838 31755 13892 31768
rect 13962 31755 14016 31768
rect 14086 31755 14140 31768
rect 14196 31755 14236 31811
rect 13728 31716 13786 31755
rect 13838 31716 13910 31755
rect 13962 31716 14034 31755
rect 14086 31716 14236 31755
rect 13728 31687 14236 31716
rect 13728 31631 13768 31687
rect 13824 31644 13892 31687
rect 13948 31644 14016 31687
rect 14072 31644 14140 31687
rect 13838 31631 13892 31644
rect 13962 31631 14016 31644
rect 14086 31631 14140 31644
rect 14196 31631 14236 31687
rect 13728 31592 13786 31631
rect 13838 31592 13910 31631
rect 13962 31592 14034 31631
rect 14086 31592 14236 31631
rect 13728 31563 14236 31592
rect 13728 31507 13768 31563
rect 13824 31520 13892 31563
rect 13948 31520 14016 31563
rect 14072 31520 14140 31563
rect 13838 31507 13892 31520
rect 13962 31507 14016 31520
rect 14086 31507 14140 31520
rect 14196 31507 14236 31563
rect 13728 31468 13786 31507
rect 13838 31468 13910 31507
rect 13962 31468 14034 31507
rect 14086 31468 14236 31507
rect 13728 31439 14236 31468
rect 13728 31383 13768 31439
rect 13824 31396 13892 31439
rect 13948 31396 14016 31439
rect 14072 31396 14140 31439
rect 13838 31383 13892 31396
rect 13962 31383 14016 31396
rect 14086 31383 14140 31396
rect 14196 31383 14236 31439
rect 13728 31344 13786 31383
rect 13838 31344 13910 31383
rect 13962 31344 14034 31383
rect 14086 31344 14236 31383
rect 13728 31315 14236 31344
rect 13728 31259 13768 31315
rect 13824 31272 13892 31315
rect 13948 31272 14016 31315
rect 14072 31272 14140 31315
rect 13838 31259 13892 31272
rect 13962 31259 14016 31272
rect 14086 31259 14140 31272
rect 14196 31259 14236 31315
rect 13728 31220 13786 31259
rect 13838 31220 13910 31259
rect 13962 31220 14034 31259
rect 14086 31220 14236 31259
rect 13728 31191 14236 31220
rect 13728 31135 13768 31191
rect 13824 31148 13892 31191
rect 13948 31148 14016 31191
rect 14072 31148 14140 31191
rect 13838 31135 13892 31148
rect 13962 31135 14016 31148
rect 14086 31135 14140 31148
rect 14196 31135 14236 31191
rect 13728 31096 13786 31135
rect 13838 31096 13910 31135
rect 13962 31096 14034 31135
rect 14086 31096 14236 31135
rect 13728 31067 14236 31096
rect 13728 31011 13768 31067
rect 13824 31024 13892 31067
rect 13948 31024 14016 31067
rect 14072 31024 14140 31067
rect 13838 31011 13892 31024
rect 13962 31011 14016 31024
rect 14086 31011 14140 31024
rect 14196 31011 14236 31067
rect 13728 30972 13786 31011
rect 13838 30972 13910 31011
rect 13962 30972 14034 31011
rect 14086 30972 14236 31011
rect 13728 30943 14236 30972
rect 13728 30887 13768 30943
rect 13824 30900 13892 30943
rect 13948 30900 14016 30943
rect 14072 30900 14140 30943
rect 13838 30887 13892 30900
rect 13962 30887 14016 30900
rect 14086 30887 14140 30900
rect 14196 30887 14236 30943
rect 13728 30848 13786 30887
rect 13838 30848 13910 30887
rect 13962 30848 14034 30887
rect 14086 30848 14236 30887
rect 13728 30819 14236 30848
rect 13728 30763 13768 30819
rect 13824 30776 13892 30819
rect 13948 30776 14016 30819
rect 14072 30776 14140 30819
rect 13838 30763 13892 30776
rect 13962 30763 14016 30776
rect 14086 30763 14140 30776
rect 14196 30763 14236 30819
rect 13728 30724 13786 30763
rect 13838 30724 13910 30763
rect 13962 30724 14034 30763
rect 14086 30724 14236 30763
rect 13728 30695 14236 30724
rect 13728 30639 13768 30695
rect 13824 30652 13892 30695
rect 13948 30652 14016 30695
rect 14072 30652 14140 30695
rect 13838 30639 13892 30652
rect 13962 30639 14016 30652
rect 14086 30639 14140 30652
rect 14196 30639 14236 30695
rect 13728 30600 13786 30639
rect 13838 30600 13910 30639
rect 13962 30600 14034 30639
rect 14086 30600 14236 30639
rect 13728 30571 14236 30600
rect 13728 30515 13768 30571
rect 13824 30528 13892 30571
rect 13948 30528 14016 30571
rect 14072 30528 14140 30571
rect 13838 30515 13892 30528
rect 13962 30515 14016 30528
rect 14086 30515 14140 30528
rect 14196 30515 14236 30571
rect 13728 30476 13786 30515
rect 13838 30476 13910 30515
rect 13962 30476 14034 30515
rect 14086 30476 14236 30515
rect 13728 30447 14236 30476
rect 13728 30391 13768 30447
rect 13824 30404 13892 30447
rect 13948 30404 14016 30447
rect 14072 30404 14140 30447
rect 13838 30391 13892 30404
rect 13962 30391 14016 30404
rect 14086 30391 14140 30404
rect 14196 30391 14236 30447
rect 13728 30352 13786 30391
rect 13838 30352 13910 30391
rect 13962 30352 14034 30391
rect 14086 30352 14236 30391
rect 13728 30323 14236 30352
rect 13728 30267 13768 30323
rect 13824 30280 13892 30323
rect 13948 30280 14016 30323
rect 14072 30280 14140 30323
rect 13838 30267 13892 30280
rect 13962 30267 14016 30280
rect 14086 30267 14140 30280
rect 14196 30267 14236 30323
rect 13728 30228 13786 30267
rect 13838 30228 13910 30267
rect 13962 30228 14034 30267
rect 14086 30228 14236 30267
rect 13728 30199 14236 30228
rect 13728 30143 13768 30199
rect 13824 30156 13892 30199
rect 13948 30156 14016 30199
rect 14072 30156 14140 30199
rect 13838 30143 13892 30156
rect 13962 30143 14016 30156
rect 14086 30143 14140 30156
rect 14196 30143 14236 30199
rect 13728 30104 13786 30143
rect 13838 30104 13910 30143
rect 13962 30104 14034 30143
rect 14086 30104 14236 30143
rect 13728 30032 14236 30104
rect 13728 29980 13786 30032
rect 13838 29980 13910 30032
rect 13962 29980 14034 30032
rect 14086 29980 14236 30032
rect 13728 29908 14236 29980
rect 13728 29856 13786 29908
rect 13838 29856 13910 29908
rect 13962 29856 14034 29908
rect 14086 29856 14236 29908
rect 13728 29845 14236 29856
rect 13728 29789 13768 29845
rect 13824 29789 13892 29845
rect 13948 29789 14016 29845
rect 14072 29789 14140 29845
rect 14196 29789 14236 29845
rect 13728 29784 14236 29789
rect 13728 29732 13786 29784
rect 13838 29732 13910 29784
rect 13962 29732 14034 29784
rect 14086 29732 14236 29784
rect 13728 29721 14236 29732
rect 13728 29665 13768 29721
rect 13824 29665 13892 29721
rect 13948 29665 14016 29721
rect 14072 29665 14140 29721
rect 14196 29665 14236 29721
rect 13728 29660 14236 29665
rect 13728 29608 13786 29660
rect 13838 29608 13910 29660
rect 13962 29608 14034 29660
rect 14086 29608 14236 29660
rect 13728 29597 14236 29608
rect 13728 29541 13768 29597
rect 13824 29541 13892 29597
rect 13948 29541 14016 29597
rect 14072 29541 14140 29597
rect 14196 29541 14236 29597
rect 13728 29536 14236 29541
rect 13728 29484 13786 29536
rect 13838 29484 13910 29536
rect 13962 29484 14034 29536
rect 14086 29484 14236 29536
rect 13728 29473 14236 29484
rect 13728 29417 13768 29473
rect 13824 29417 13892 29473
rect 13948 29417 14016 29473
rect 14072 29417 14140 29473
rect 14196 29417 14236 29473
rect 13728 29349 14236 29417
rect 13728 29293 13768 29349
rect 13824 29293 13892 29349
rect 13948 29293 14016 29349
rect 14072 29293 14140 29349
rect 14196 29293 14236 29349
rect 13728 29225 14236 29293
rect 13728 29169 13768 29225
rect 13824 29169 13892 29225
rect 13948 29169 14016 29225
rect 14072 29169 14140 29225
rect 14196 29169 14236 29225
rect 13728 29101 14236 29169
rect 13728 29045 13768 29101
rect 13824 29045 13892 29101
rect 13948 29045 14016 29101
rect 14072 29045 14140 29101
rect 14196 29045 14236 29101
rect 13728 28977 14236 29045
rect 13728 28921 13768 28977
rect 13824 28921 13892 28977
rect 13948 28921 14016 28977
rect 14072 28921 14140 28977
rect 14196 28921 14236 28977
rect 13728 28853 14236 28921
rect 13728 28797 13768 28853
rect 13824 28797 13892 28853
rect 13948 28797 14016 28853
rect 14072 28797 14140 28853
rect 14196 28797 14236 28853
rect 13728 28729 14236 28797
rect 13728 28673 13768 28729
rect 13824 28688 13892 28729
rect 13948 28688 14016 28729
rect 14072 28688 14140 28729
rect 13838 28673 13892 28688
rect 13962 28673 14016 28688
rect 14086 28673 14140 28688
rect 14196 28673 14236 28729
rect 13728 28636 13786 28673
rect 13838 28636 13910 28673
rect 13962 28636 14034 28673
rect 14086 28636 14236 28673
rect 13728 28605 14236 28636
rect 13728 28549 13768 28605
rect 13824 28564 13892 28605
rect 13948 28564 14016 28605
rect 14072 28564 14140 28605
rect 13838 28549 13892 28564
rect 13962 28549 14016 28564
rect 14086 28549 14140 28564
rect 14196 28549 14236 28605
rect 13728 28512 13786 28549
rect 13838 28512 13910 28549
rect 13962 28512 14034 28549
rect 14086 28512 14236 28549
rect 13728 28440 14236 28512
rect 13728 28388 13786 28440
rect 13838 28388 13910 28440
rect 13962 28388 14034 28440
rect 14086 28388 14236 28440
rect 13728 28316 14236 28388
rect 13728 28264 13786 28316
rect 13838 28264 13910 28316
rect 13962 28264 14034 28316
rect 14086 28264 14236 28316
rect 13728 28192 14236 28264
rect 13728 28140 13786 28192
rect 13838 28140 13910 28192
rect 13962 28140 14034 28192
rect 14086 28140 14236 28192
rect 13728 28068 14236 28140
rect 13728 28016 13786 28068
rect 13838 28016 13910 28068
rect 13962 28016 14034 28068
rect 14086 28016 14236 28068
rect 13728 27944 14236 28016
rect 13728 27892 13786 27944
rect 13838 27892 13910 27944
rect 13962 27892 14034 27944
rect 14086 27892 14236 27944
rect 13728 27820 14236 27892
rect 13728 27768 13786 27820
rect 13838 27768 13910 27820
rect 13962 27768 14034 27820
rect 14086 27768 14236 27820
rect 13728 27696 14236 27768
rect 13728 27644 13786 27696
rect 13838 27644 13910 27696
rect 13962 27644 14034 27696
rect 14086 27644 14236 27696
rect 13728 27572 14236 27644
rect 13728 27520 13786 27572
rect 13838 27520 13910 27572
rect 13962 27520 14034 27572
rect 14086 27520 14236 27572
rect 13728 27448 14236 27520
rect 13728 27396 13786 27448
rect 13838 27396 13910 27448
rect 13962 27396 14034 27448
rect 14086 27396 14236 27448
rect 13728 27324 14236 27396
rect 13728 27272 13786 27324
rect 13838 27272 13910 27324
rect 13962 27272 14034 27324
rect 14086 27272 14236 27324
rect 13728 27200 14236 27272
rect 13728 27148 13786 27200
rect 13838 27148 13910 27200
rect 13962 27148 14034 27200
rect 14086 27148 14236 27200
rect 13728 27076 14236 27148
rect 13728 27024 13786 27076
rect 13838 27024 13910 27076
rect 13962 27024 14034 27076
rect 14086 27024 14236 27076
rect 13728 26952 14236 27024
rect 13728 26900 13786 26952
rect 13838 26900 13910 26952
rect 13962 26900 14034 26952
rect 14086 26900 14236 26952
rect 13728 26828 14236 26900
rect 13728 26776 13786 26828
rect 13838 26776 13910 26828
rect 13962 26776 14034 26828
rect 14086 26776 14236 26828
rect 13728 26704 14236 26776
rect 13728 26652 13786 26704
rect 13838 26652 13910 26704
rect 13962 26652 14034 26704
rect 14086 26652 14236 26704
rect 13728 26651 14236 26652
rect 13728 26595 13768 26651
rect 13824 26595 13892 26651
rect 13948 26595 14016 26651
rect 14072 26595 14140 26651
rect 14196 26595 14236 26651
rect 13728 26580 14236 26595
rect 13728 26528 13786 26580
rect 13838 26528 13910 26580
rect 13962 26528 14034 26580
rect 14086 26528 14236 26580
rect 13728 26527 14236 26528
rect 13728 26471 13768 26527
rect 13824 26471 13892 26527
rect 13948 26471 14016 26527
rect 14072 26471 14140 26527
rect 14196 26471 14236 26527
rect 13728 26456 14236 26471
rect 13728 26404 13786 26456
rect 13838 26404 13910 26456
rect 13962 26404 14034 26456
rect 14086 26404 14236 26456
rect 13728 26403 14236 26404
rect 13728 26347 13768 26403
rect 13824 26347 13892 26403
rect 13948 26347 14016 26403
rect 14072 26347 14140 26403
rect 14196 26347 14236 26403
rect 13728 26332 14236 26347
rect 13728 26280 13786 26332
rect 13838 26280 13910 26332
rect 13962 26280 14034 26332
rect 14086 26280 14236 26332
rect 13728 26279 14236 26280
rect 13728 26223 13768 26279
rect 13824 26223 13892 26279
rect 13948 26223 14016 26279
rect 14072 26223 14140 26279
rect 14196 26223 14236 26279
rect 13728 26208 14236 26223
rect 13728 26156 13786 26208
rect 13838 26156 13910 26208
rect 13962 26156 14034 26208
rect 14086 26156 14236 26208
rect 13728 26155 14236 26156
rect 13728 26099 13768 26155
rect 13824 26099 13892 26155
rect 13948 26099 14016 26155
rect 14072 26099 14140 26155
rect 14196 26099 14236 26155
rect 13728 26084 14236 26099
rect 13728 26032 13786 26084
rect 13838 26032 13910 26084
rect 13962 26032 14034 26084
rect 14086 26032 14236 26084
rect 13728 26031 14236 26032
rect 13728 25975 13768 26031
rect 13824 25975 13892 26031
rect 13948 25975 14016 26031
rect 14072 25975 14140 26031
rect 14196 25975 14236 26031
rect 13728 25960 14236 25975
rect 13728 25908 13786 25960
rect 13838 25908 13910 25960
rect 13962 25908 14034 25960
rect 14086 25908 14236 25960
rect 13728 25907 14236 25908
rect 13728 25851 13768 25907
rect 13824 25851 13892 25907
rect 13948 25851 14016 25907
rect 14072 25851 14140 25907
rect 14196 25851 14236 25907
rect 13728 25836 14236 25851
rect 13728 25784 13786 25836
rect 13838 25784 13910 25836
rect 13962 25784 14034 25836
rect 14086 25784 14236 25836
rect 13728 25783 14236 25784
rect 13728 25727 13768 25783
rect 13824 25727 13892 25783
rect 13948 25727 14016 25783
rect 14072 25727 14140 25783
rect 14196 25727 14236 25783
rect 13728 25712 14236 25727
rect 13728 25660 13786 25712
rect 13838 25660 13910 25712
rect 13962 25660 14034 25712
rect 14086 25660 14236 25712
rect 13728 25659 14236 25660
rect 13728 25603 13768 25659
rect 13824 25603 13892 25659
rect 13948 25603 14016 25659
rect 14072 25603 14140 25659
rect 14196 25603 14236 25659
rect 13728 25588 14236 25603
rect 13728 25536 13786 25588
rect 13838 25536 13910 25588
rect 13962 25536 14034 25588
rect 14086 25536 14236 25588
rect 13728 25535 14236 25536
rect 13728 25479 13768 25535
rect 13824 25479 13892 25535
rect 13948 25479 14016 25535
rect 14072 25479 14140 25535
rect 14196 25479 14236 25535
rect 13728 25411 14236 25479
rect 13728 25355 13768 25411
rect 13824 25355 13892 25411
rect 13948 25355 14016 25411
rect 14072 25355 14140 25411
rect 14196 25355 14236 25411
rect 13728 25287 14236 25355
rect 13728 25231 13768 25287
rect 13824 25231 13892 25287
rect 13948 25231 14016 25287
rect 14072 25231 14140 25287
rect 14196 25231 14236 25287
rect 13728 25163 14236 25231
rect 13728 25107 13768 25163
rect 13824 25107 13892 25163
rect 13948 25107 14016 25163
rect 14072 25107 14140 25163
rect 14196 25107 14236 25163
rect 13728 25039 14236 25107
rect 13728 24983 13768 25039
rect 13824 24983 13892 25039
rect 13948 24983 14016 25039
rect 14072 24983 14140 25039
rect 14196 24983 14236 25039
rect 13728 24915 14236 24983
rect 13728 24859 13768 24915
rect 13824 24859 13892 24915
rect 13948 24859 14016 24915
rect 14072 24859 14140 24915
rect 14196 24859 14236 24915
rect 13728 24791 14236 24859
rect 13728 24735 13768 24791
rect 13824 24740 13892 24791
rect 13948 24740 14016 24791
rect 14072 24740 14140 24791
rect 13838 24735 13892 24740
rect 13962 24735 14016 24740
rect 14086 24735 14140 24740
rect 14196 24735 14236 24791
rect 13728 24688 13786 24735
rect 13838 24688 13910 24735
rect 13962 24688 14034 24735
rect 14086 24688 14236 24735
rect 13728 24667 14236 24688
rect 13728 24611 13768 24667
rect 13824 24616 13892 24667
rect 13948 24616 14016 24667
rect 14072 24616 14140 24667
rect 13838 24611 13892 24616
rect 13962 24611 14016 24616
rect 14086 24611 14140 24616
rect 14196 24611 14236 24667
rect 13728 24564 13786 24611
rect 13838 24564 13910 24611
rect 13962 24564 14034 24611
rect 14086 24564 14236 24611
rect 13728 24543 14236 24564
rect 13728 24487 13768 24543
rect 13824 24492 13892 24543
rect 13948 24492 14016 24543
rect 14072 24492 14140 24543
rect 13838 24487 13892 24492
rect 13962 24487 14016 24492
rect 14086 24487 14140 24492
rect 14196 24487 14236 24543
rect 13728 24440 13786 24487
rect 13838 24440 13910 24487
rect 13962 24440 14034 24487
rect 14086 24440 14236 24487
rect 13728 24419 14236 24440
rect 13728 24363 13768 24419
rect 13824 24368 13892 24419
rect 13948 24368 14016 24419
rect 14072 24368 14140 24419
rect 13838 24363 13892 24368
rect 13962 24363 14016 24368
rect 14086 24363 14140 24368
rect 14196 24363 14236 24419
rect 13728 24316 13786 24363
rect 13838 24316 13910 24363
rect 13962 24316 14034 24363
rect 14086 24316 14236 24363
rect 13728 24295 14236 24316
rect 13728 24239 13768 24295
rect 13824 24244 13892 24295
rect 13948 24244 14016 24295
rect 14072 24244 14140 24295
rect 13838 24239 13892 24244
rect 13962 24239 14016 24244
rect 14086 24239 14140 24244
rect 14196 24239 14236 24295
rect 13728 24192 13786 24239
rect 13838 24192 13910 24239
rect 13962 24192 14034 24239
rect 14086 24192 14236 24239
rect 13728 24171 14236 24192
rect 13728 24115 13768 24171
rect 13824 24120 13892 24171
rect 13948 24120 14016 24171
rect 14072 24120 14140 24171
rect 13838 24115 13892 24120
rect 13962 24115 14016 24120
rect 14086 24115 14140 24120
rect 14196 24115 14236 24171
rect 13728 24068 13786 24115
rect 13838 24068 13910 24115
rect 13962 24068 14034 24115
rect 14086 24068 14236 24115
rect 13728 24047 14236 24068
rect 13728 23991 13768 24047
rect 13824 23996 13892 24047
rect 13948 23996 14016 24047
rect 14072 23996 14140 24047
rect 13838 23991 13892 23996
rect 13962 23991 14016 23996
rect 14086 23991 14140 23996
rect 14196 23991 14236 24047
rect 13728 23944 13786 23991
rect 13838 23944 13910 23991
rect 13962 23944 14034 23991
rect 14086 23944 14236 23991
rect 13728 23923 14236 23944
rect 13728 23867 13768 23923
rect 13824 23872 13892 23923
rect 13948 23872 14016 23923
rect 14072 23872 14140 23923
rect 13838 23867 13892 23872
rect 13962 23867 14016 23872
rect 14086 23867 14140 23872
rect 14196 23867 14236 23923
rect 13728 23820 13786 23867
rect 13838 23820 13910 23867
rect 13962 23820 14034 23867
rect 14086 23820 14236 23867
rect 13728 23799 14236 23820
rect 13728 23743 13768 23799
rect 13824 23748 13892 23799
rect 13948 23748 14016 23799
rect 14072 23748 14140 23799
rect 13838 23743 13892 23748
rect 13962 23743 14016 23748
rect 14086 23743 14140 23748
rect 14196 23743 14236 23799
rect 13728 23696 13786 23743
rect 13838 23696 13910 23743
rect 13962 23696 14034 23743
rect 14086 23696 14236 23743
rect 13728 23624 14236 23696
rect 13728 23572 13786 23624
rect 13838 23572 13910 23624
rect 13962 23572 14034 23624
rect 14086 23572 14236 23624
rect 13728 23500 14236 23572
rect 13728 23451 13786 23500
rect 13838 23451 13910 23500
rect 13962 23451 14034 23500
rect 14086 23451 14236 23500
rect 13728 23395 13768 23451
rect 13838 23448 13892 23451
rect 13962 23448 14016 23451
rect 14086 23448 14140 23451
rect 13824 23395 13892 23448
rect 13948 23395 14016 23448
rect 14072 23395 14140 23448
rect 14196 23395 14236 23451
rect 13728 23376 14236 23395
rect 13728 23327 13786 23376
rect 13838 23327 13910 23376
rect 13962 23327 14034 23376
rect 14086 23327 14236 23376
rect 13728 23271 13768 23327
rect 13838 23324 13892 23327
rect 13962 23324 14016 23327
rect 14086 23324 14140 23327
rect 13824 23271 13892 23324
rect 13948 23271 14016 23324
rect 14072 23271 14140 23324
rect 14196 23271 14236 23327
rect 13728 23252 14236 23271
rect 13728 23203 13786 23252
rect 13838 23203 13910 23252
rect 13962 23203 14034 23252
rect 14086 23203 14236 23252
rect 13728 23147 13768 23203
rect 13838 23200 13892 23203
rect 13962 23200 14016 23203
rect 14086 23200 14140 23203
rect 13824 23147 13892 23200
rect 13948 23147 14016 23200
rect 14072 23147 14140 23200
rect 14196 23147 14236 23203
rect 13728 23128 14236 23147
rect 13728 23079 13786 23128
rect 13838 23079 13910 23128
rect 13962 23079 14034 23128
rect 14086 23079 14236 23128
rect 13728 23023 13768 23079
rect 13838 23076 13892 23079
rect 13962 23076 14016 23079
rect 14086 23076 14140 23079
rect 13824 23023 13892 23076
rect 13948 23023 14016 23076
rect 14072 23023 14140 23076
rect 14196 23023 14236 23079
rect 13728 23004 14236 23023
rect 13728 22955 13786 23004
rect 13838 22955 13910 23004
rect 13962 22955 14034 23004
rect 14086 22955 14236 23004
rect 13728 22899 13768 22955
rect 13838 22952 13892 22955
rect 13962 22952 14016 22955
rect 14086 22952 14140 22955
rect 13824 22899 13892 22952
rect 13948 22899 14016 22952
rect 14072 22899 14140 22952
rect 14196 22899 14236 22955
rect 13728 22880 14236 22899
rect 13728 22831 13786 22880
rect 13838 22831 13910 22880
rect 13962 22831 14034 22880
rect 14086 22831 14236 22880
rect 13728 22775 13768 22831
rect 13838 22828 13892 22831
rect 13962 22828 14016 22831
rect 14086 22828 14140 22831
rect 13824 22775 13892 22828
rect 13948 22775 14016 22828
rect 14072 22775 14140 22828
rect 14196 22775 14236 22831
rect 13728 22756 14236 22775
rect 13728 22707 13786 22756
rect 13838 22707 13910 22756
rect 13962 22707 14034 22756
rect 14086 22707 14236 22756
rect 13728 22651 13768 22707
rect 13838 22704 13892 22707
rect 13962 22704 14016 22707
rect 14086 22704 14140 22707
rect 13824 22651 13892 22704
rect 13948 22651 14016 22704
rect 14072 22651 14140 22704
rect 14196 22651 14236 22707
rect 13728 22632 14236 22651
rect 13728 22583 13786 22632
rect 13838 22583 13910 22632
rect 13962 22583 14034 22632
rect 14086 22583 14236 22632
rect 13728 22527 13768 22583
rect 13838 22580 13892 22583
rect 13962 22580 14016 22583
rect 14086 22580 14140 22583
rect 13824 22527 13892 22580
rect 13948 22527 14016 22580
rect 14072 22527 14140 22580
rect 14196 22527 14236 22583
rect 13728 22508 14236 22527
rect 13728 22459 13786 22508
rect 13838 22459 13910 22508
rect 13962 22459 14034 22508
rect 14086 22459 14236 22508
rect 13728 22403 13768 22459
rect 13838 22456 13892 22459
rect 13962 22456 14016 22459
rect 14086 22456 14140 22459
rect 13824 22403 13892 22456
rect 13948 22403 14016 22456
rect 14072 22403 14140 22456
rect 14196 22403 14236 22459
rect 13728 22384 14236 22403
rect 13728 22335 13786 22384
rect 13838 22335 13910 22384
rect 13962 22335 14034 22384
rect 14086 22335 14236 22384
rect 13728 22279 13768 22335
rect 13838 22332 13892 22335
rect 13962 22332 14016 22335
rect 14086 22332 14140 22335
rect 13824 22279 13892 22332
rect 13948 22279 14016 22332
rect 14072 22279 14140 22332
rect 14196 22279 14236 22335
rect 13728 22260 14236 22279
rect 13728 22211 13786 22260
rect 13838 22211 13910 22260
rect 13962 22211 14034 22260
rect 14086 22211 14236 22260
rect 13728 22155 13768 22211
rect 13838 22208 13892 22211
rect 13962 22208 14016 22211
rect 14086 22208 14140 22211
rect 13824 22155 13892 22208
rect 13948 22155 14016 22208
rect 14072 22155 14140 22208
rect 14196 22155 14236 22211
rect 13728 22136 14236 22155
rect 13728 22087 13786 22136
rect 13838 22087 13910 22136
rect 13962 22087 14034 22136
rect 14086 22087 14236 22136
rect 13728 22031 13768 22087
rect 13838 22084 13892 22087
rect 13962 22084 14016 22087
rect 14086 22084 14140 22087
rect 13824 22031 13892 22084
rect 13948 22031 14016 22084
rect 14072 22031 14140 22084
rect 14196 22031 14236 22087
rect 13728 22012 14236 22031
rect 13728 21963 13786 22012
rect 13838 21963 13910 22012
rect 13962 21963 14034 22012
rect 14086 21963 14236 22012
rect 13728 21907 13768 21963
rect 13838 21960 13892 21963
rect 13962 21960 14016 21963
rect 14086 21960 14140 21963
rect 13824 21907 13892 21960
rect 13948 21907 14016 21960
rect 14072 21907 14140 21960
rect 14196 21907 14236 21963
rect 13728 21888 14236 21907
rect 13728 21839 13786 21888
rect 13838 21839 13910 21888
rect 13962 21839 14034 21888
rect 14086 21839 14236 21888
rect 13728 21783 13768 21839
rect 13838 21836 13892 21839
rect 13962 21836 14016 21839
rect 14086 21836 14140 21839
rect 13824 21783 13892 21836
rect 13948 21783 14016 21836
rect 14072 21783 14140 21836
rect 14196 21783 14236 21839
rect 13728 21764 14236 21783
rect 13728 21715 13786 21764
rect 13838 21715 13910 21764
rect 13962 21715 14034 21764
rect 14086 21715 14236 21764
rect 13728 21659 13768 21715
rect 13838 21712 13892 21715
rect 13962 21712 14016 21715
rect 14086 21712 14140 21715
rect 13824 21659 13892 21712
rect 13948 21659 14016 21712
rect 14072 21659 14140 21712
rect 14196 21659 14236 21715
rect 13728 21640 14236 21659
rect 13728 21591 13786 21640
rect 13838 21591 13910 21640
rect 13962 21591 14034 21640
rect 14086 21591 14236 21640
rect 13728 21535 13768 21591
rect 13838 21588 13892 21591
rect 13962 21588 14016 21591
rect 14086 21588 14140 21591
rect 13824 21535 13892 21588
rect 13948 21535 14016 21588
rect 14072 21535 14140 21588
rect 14196 21535 14236 21591
rect 13728 21467 14236 21535
rect 13728 21411 13768 21467
rect 13824 21411 13892 21467
rect 13948 21411 14016 21467
rect 14072 21411 14140 21467
rect 14196 21411 14236 21467
rect 13728 21343 14236 21411
rect 13728 21287 13768 21343
rect 13824 21287 13892 21343
rect 13948 21287 14016 21343
rect 14072 21287 14140 21343
rect 14196 21287 14236 21343
rect 13728 21219 14236 21287
rect 13728 21163 13768 21219
rect 13824 21163 13892 21219
rect 13948 21163 14016 21219
rect 14072 21163 14140 21219
rect 14196 21163 14236 21219
rect 13728 21095 14236 21163
rect 13728 21039 13768 21095
rect 13824 21039 13892 21095
rect 13948 21039 14016 21095
rect 14072 21039 14140 21095
rect 14196 21039 14236 21095
rect 13728 20971 14236 21039
rect 13728 20915 13768 20971
rect 13824 20915 13892 20971
rect 13948 20915 14016 20971
rect 14072 20915 14140 20971
rect 14196 20915 14236 20971
rect 13728 20847 14236 20915
rect 13728 20791 13768 20847
rect 13824 20791 13892 20847
rect 13948 20791 14016 20847
rect 14072 20791 14140 20847
rect 14196 20791 14236 20847
rect 13728 20723 14236 20791
rect 13728 20667 13768 20723
rect 13824 20667 13892 20723
rect 13948 20667 14016 20723
rect 14072 20667 14140 20723
rect 14196 20667 14236 20723
rect 13728 20599 14236 20667
rect 13728 20543 13768 20599
rect 13824 20543 13892 20599
rect 13948 20543 14016 20599
rect 14072 20543 14140 20599
rect 14196 20543 14236 20599
rect 13728 20251 14236 20543
rect 13728 20195 13768 20251
rect 13824 20195 13892 20251
rect 13948 20195 14016 20251
rect 14072 20195 14140 20251
rect 14196 20195 14236 20251
rect 13728 20127 14236 20195
rect 13728 20071 13768 20127
rect 13824 20071 13892 20127
rect 13948 20071 14016 20127
rect 14072 20071 14140 20127
rect 14196 20071 14236 20127
rect 13728 20003 14236 20071
rect 13728 19947 13768 20003
rect 13824 19947 13892 20003
rect 13948 19947 14016 20003
rect 14072 19947 14140 20003
rect 14196 19947 14236 20003
rect 13728 19879 14236 19947
rect 13728 19823 13768 19879
rect 13824 19823 13892 19879
rect 13948 19823 14016 19879
rect 14072 19823 14140 19879
rect 14196 19823 14236 19879
rect 13728 19755 14236 19823
rect 13728 19699 13768 19755
rect 13824 19699 13892 19755
rect 13948 19699 14016 19755
rect 14072 19699 14140 19755
rect 14196 19699 14236 19755
rect 13728 19631 14236 19699
rect 13728 19575 13768 19631
rect 13824 19575 13892 19631
rect 13948 19575 14016 19631
rect 14072 19575 14140 19631
rect 14196 19575 14236 19631
rect 13728 19507 14236 19575
rect 13728 19451 13768 19507
rect 13824 19451 13892 19507
rect 13948 19451 14016 19507
rect 14072 19451 14140 19507
rect 14196 19451 14236 19507
rect 13728 19383 14236 19451
rect 13728 19327 13768 19383
rect 13824 19327 13892 19383
rect 13948 19327 14016 19383
rect 14072 19327 14140 19383
rect 14196 19327 14236 19383
rect 13728 19259 14236 19327
rect 13728 19203 13768 19259
rect 13824 19203 13892 19259
rect 13948 19203 14016 19259
rect 14072 19203 14140 19259
rect 14196 19203 14236 19259
rect 13728 19135 14236 19203
rect 13728 19079 13768 19135
rect 13824 19079 13892 19135
rect 13948 19079 14016 19135
rect 14072 19079 14140 19135
rect 14196 19079 14236 19135
rect 13728 19011 14236 19079
rect 13728 18955 13768 19011
rect 13824 18955 13892 19011
rect 13948 18955 14016 19011
rect 14072 18955 14140 19011
rect 14196 18955 14236 19011
rect 13728 18887 14236 18955
rect 13728 18831 13768 18887
rect 13824 18831 13892 18887
rect 13948 18831 14016 18887
rect 14072 18831 14140 18887
rect 14196 18831 14236 18887
rect 13728 18763 14236 18831
rect 13728 18707 13768 18763
rect 13824 18707 13892 18763
rect 13948 18707 14016 18763
rect 14072 18707 14140 18763
rect 14196 18707 14236 18763
rect 13728 18639 14236 18707
rect 13728 18583 13768 18639
rect 13824 18583 13892 18639
rect 13948 18583 14016 18639
rect 14072 18583 14140 18639
rect 14196 18583 14236 18639
rect 13728 18515 14236 18583
rect 13728 18459 13768 18515
rect 13824 18459 13892 18515
rect 13948 18459 14016 18515
rect 14072 18459 14140 18515
rect 14196 18459 14236 18515
rect 13728 18391 14236 18459
rect 13728 18335 13768 18391
rect 13824 18335 13892 18391
rect 13948 18335 14016 18391
rect 14072 18335 14140 18391
rect 14196 18335 14236 18391
rect 13728 18267 14236 18335
rect 13728 18211 13768 18267
rect 13824 18211 13892 18267
rect 13948 18211 14016 18267
rect 14072 18211 14140 18267
rect 14196 18211 14236 18267
rect 13728 18143 14236 18211
rect 13728 18087 13768 18143
rect 13824 18087 13892 18143
rect 13948 18087 14016 18143
rect 14072 18087 14140 18143
rect 14196 18087 14236 18143
rect 13728 18019 14236 18087
rect 13728 17963 13768 18019
rect 13824 17963 13892 18019
rect 13948 17963 14016 18019
rect 14072 17963 14140 18019
rect 14196 17963 14236 18019
rect 13728 17895 14236 17963
rect 13728 17839 13768 17895
rect 13824 17839 13892 17895
rect 13948 17839 14016 17895
rect 14072 17839 14140 17895
rect 14196 17839 14236 17895
rect 13728 17771 14236 17839
rect 13728 17715 13768 17771
rect 13824 17715 13892 17771
rect 13948 17715 14016 17771
rect 14072 17715 14140 17771
rect 14196 17715 14236 17771
rect 13728 17647 14236 17715
rect 13728 17591 13768 17647
rect 13824 17591 13892 17647
rect 13948 17591 14016 17647
rect 14072 17591 14140 17647
rect 14196 17591 14236 17647
rect 13728 17523 14236 17591
rect 13728 17467 13768 17523
rect 13824 17467 13892 17523
rect 13948 17467 14016 17523
rect 14072 17467 14140 17523
rect 14196 17467 14236 17523
rect 13728 17399 14236 17467
rect 13728 17343 13768 17399
rect 13824 17343 13892 17399
rect 13948 17343 14016 17399
rect 14072 17343 14140 17399
rect 14196 17343 14236 17399
rect 13728 17051 14236 17343
rect 13728 16995 13768 17051
rect 13824 16995 13892 17051
rect 13948 16995 14016 17051
rect 14072 16995 14140 17051
rect 14196 16995 14236 17051
rect 13728 16927 14236 16995
rect 13728 16871 13768 16927
rect 13824 16871 13892 16927
rect 13948 16871 14016 16927
rect 14072 16871 14140 16927
rect 14196 16871 14236 16927
rect 13728 16803 14236 16871
rect 13728 16747 13768 16803
rect 13824 16747 13892 16803
rect 13948 16747 14016 16803
rect 14072 16747 14140 16803
rect 14196 16747 14236 16803
rect 13728 16679 14236 16747
rect 13728 16623 13768 16679
rect 13824 16623 13892 16679
rect 13948 16623 14016 16679
rect 14072 16623 14140 16679
rect 14196 16623 14236 16679
rect 13728 16555 14236 16623
rect 13728 16499 13768 16555
rect 13824 16499 13892 16555
rect 13948 16499 14016 16555
rect 14072 16499 14140 16555
rect 14196 16499 14236 16555
rect 13728 16431 14236 16499
rect 13728 16375 13768 16431
rect 13824 16375 13892 16431
rect 13948 16375 14016 16431
rect 14072 16375 14140 16431
rect 14196 16375 14236 16431
rect 13728 16307 14236 16375
rect 13728 16251 13768 16307
rect 13824 16251 13892 16307
rect 13948 16251 14016 16307
rect 14072 16251 14140 16307
rect 14196 16251 14236 16307
rect 13728 16183 14236 16251
rect 13728 16127 13768 16183
rect 13824 16127 13892 16183
rect 13948 16127 14016 16183
rect 14072 16127 14140 16183
rect 14196 16127 14236 16183
rect 13728 16059 14236 16127
rect 13728 16003 13768 16059
rect 13824 16003 13892 16059
rect 13948 16003 14016 16059
rect 14072 16003 14140 16059
rect 14196 16003 14236 16059
rect 13728 15935 14236 16003
rect 13728 15879 13768 15935
rect 13824 15879 13892 15935
rect 13948 15879 14016 15935
rect 14072 15879 14140 15935
rect 14196 15879 14236 15935
rect 13728 15811 14236 15879
rect 13060 15755 13070 15762
rect 12622 15687 13070 15755
rect 12622 15631 12632 15687
rect 12688 15631 12756 15687
rect 12812 15631 12880 15687
rect 12936 15631 13004 15687
rect 13060 15631 13070 15687
rect 12622 15563 13070 15631
rect 12622 15507 12632 15563
rect 12688 15507 12756 15563
rect 12812 15507 12880 15563
rect 12936 15507 13004 15563
rect 13060 15507 13070 15563
rect 12622 15439 13070 15507
rect 12622 15383 12632 15439
rect 12688 15383 12756 15439
rect 12812 15383 12880 15439
rect 12936 15383 13004 15439
rect 13060 15383 13070 15439
rect 12622 15315 13070 15383
rect 12622 15259 12632 15315
rect 12688 15259 12756 15315
rect 12812 15259 12880 15315
rect 12936 15259 13004 15315
rect 13060 15259 13070 15315
rect 12622 15191 13070 15259
rect 12622 15135 12632 15191
rect 12688 15135 12756 15191
rect 12812 15135 12880 15191
rect 12936 15135 13004 15191
rect 13060 15135 13070 15191
rect 12622 15067 13070 15135
rect 12622 15011 12632 15067
rect 12688 15011 12756 15067
rect 12812 15011 12880 15067
rect 12936 15011 13004 15067
rect 13060 15011 13070 15067
rect 12622 14943 13070 15011
rect 12622 14887 12632 14943
rect 12688 14887 12756 14943
rect 12812 14887 12880 14943
rect 12936 14887 13004 14943
rect 13060 14887 13070 14943
rect 12622 14819 13070 14887
rect 12622 14763 12632 14819
rect 12688 14763 12756 14819
rect 12812 14763 12880 14819
rect 12936 14763 13004 14819
rect 13060 14763 13070 14819
rect 12622 14695 13070 14763
rect 12622 14639 12632 14695
rect 12688 14639 12756 14695
rect 12812 14639 12880 14695
rect 12936 14639 13004 14695
rect 13060 14639 13070 14695
rect 12622 14571 13070 14639
rect 12622 14515 12632 14571
rect 12688 14515 12756 14571
rect 12812 14515 12880 14571
rect 12936 14515 13004 14571
rect 13060 14515 13070 14571
rect 12622 14447 13070 14515
rect 12622 14391 12632 14447
rect 12688 14391 12756 14447
rect 12812 14391 12880 14447
rect 12936 14391 13004 14447
rect 13060 14391 13070 14447
rect 12622 14323 13070 14391
rect 12622 14267 12632 14323
rect 12688 14267 12756 14323
rect 12812 14267 12880 14323
rect 12936 14267 13004 14323
rect 13060 14267 13070 14323
rect 12622 14199 13070 14267
rect 12622 14143 12632 14199
rect 12688 14143 12756 14199
rect 12812 14143 12880 14199
rect 12936 14143 13004 14199
rect 13060 14143 13070 14199
rect 12622 14133 13070 14143
rect 13728 15755 13768 15811
rect 13824 15755 13892 15811
rect 13948 15755 14016 15811
rect 14072 15755 14140 15811
rect 14196 15755 14236 15811
rect 13728 15687 14236 15755
rect 13728 15631 13768 15687
rect 13824 15631 13892 15687
rect 13948 15631 14016 15687
rect 14072 15631 14140 15687
rect 14196 15631 14236 15687
rect 13728 15563 14236 15631
rect 13728 15507 13768 15563
rect 13824 15507 13892 15563
rect 13948 15507 14016 15563
rect 14072 15507 14140 15563
rect 14196 15507 14236 15563
rect 13728 15439 14236 15507
rect 13728 15383 13768 15439
rect 13824 15383 13892 15439
rect 13948 15383 14016 15439
rect 14072 15383 14140 15439
rect 14196 15383 14236 15439
rect 13728 15315 14236 15383
rect 13728 15259 13768 15315
rect 13824 15259 13892 15315
rect 13948 15259 14016 15315
rect 14072 15259 14140 15315
rect 14196 15259 14236 15315
rect 13728 15191 14236 15259
rect 13728 15135 13768 15191
rect 13824 15135 13892 15191
rect 13948 15135 14016 15191
rect 14072 15135 14140 15191
rect 14196 15135 14236 15191
rect 13728 15067 14236 15135
rect 13728 15011 13768 15067
rect 13824 15011 13892 15067
rect 13948 15011 14016 15067
rect 14072 15011 14140 15067
rect 14196 15011 14236 15067
rect 13728 14943 14236 15011
rect 13728 14887 13768 14943
rect 13824 14887 13892 14943
rect 13948 14887 14016 14943
rect 14072 14887 14140 14943
rect 14196 14887 14236 14943
rect 13728 14819 14236 14887
rect 13728 14763 13768 14819
rect 13824 14763 13892 14819
rect 13948 14763 14016 14819
rect 14072 14763 14140 14819
rect 14196 14763 14236 14819
rect 13728 14695 14236 14763
rect 13728 14639 13768 14695
rect 13824 14639 13892 14695
rect 13948 14639 14016 14695
rect 14072 14639 14140 14695
rect 14196 14639 14236 14695
rect 13728 14571 14236 14639
rect 13728 14515 13768 14571
rect 13824 14515 13892 14571
rect 13948 14515 14016 14571
rect 14072 14515 14140 14571
rect 14196 14515 14236 14571
rect 13728 14447 14236 14515
rect 13728 14391 13768 14447
rect 13824 14391 13892 14447
rect 13948 14391 14016 14447
rect 14072 14391 14140 14447
rect 14196 14391 14236 14447
rect 13728 14323 14236 14391
rect 13728 14267 13768 14323
rect 13824 14267 13892 14323
rect 13948 14267 14016 14323
rect 14072 14267 14140 14323
rect 14196 14267 14236 14323
rect 13728 14199 14236 14267
rect 13728 14143 13768 14199
rect 13824 14143 13892 14199
rect 13948 14143 14016 14199
rect 14072 14143 14140 14199
rect 14196 14143 14236 14199
rect 260 13789 300 13845
rect 356 13789 424 13845
rect 480 13789 548 13845
rect 604 13789 672 13845
rect 728 13789 768 13845
rect 260 13721 768 13789
rect 260 13665 300 13721
rect 356 13665 424 13721
rect 480 13665 548 13721
rect 604 13665 672 13721
rect 728 13665 768 13721
rect 260 13597 768 13665
rect 260 13541 300 13597
rect 356 13541 424 13597
rect 480 13541 548 13597
rect 604 13541 672 13597
rect 728 13541 768 13597
rect 260 13473 768 13541
rect 260 13417 300 13473
rect 356 13417 424 13473
rect 480 13417 548 13473
rect 604 13417 672 13473
rect 728 13417 768 13473
rect 260 13349 768 13417
rect 260 13293 300 13349
rect 356 13293 424 13349
rect 480 13293 548 13349
rect 604 13293 672 13349
rect 728 13293 768 13349
rect 260 13225 768 13293
rect 260 13169 300 13225
rect 356 13169 424 13225
rect 480 13169 548 13225
rect 604 13169 672 13225
rect 728 13169 768 13225
rect 260 13101 768 13169
rect 260 13045 300 13101
rect 356 13045 424 13101
rect 480 13045 548 13101
rect 604 13045 672 13101
rect 728 13045 768 13101
rect 260 12977 768 13045
rect 260 12921 300 12977
rect 356 12921 424 12977
rect 480 12921 548 12977
rect 604 12921 672 12977
rect 728 12921 768 12977
rect 260 12853 768 12921
rect 260 12797 300 12853
rect 356 12797 424 12853
rect 480 12797 548 12853
rect 604 12797 672 12853
rect 728 12797 768 12853
rect 260 12729 768 12797
rect 260 12673 300 12729
rect 356 12673 424 12729
rect 480 12673 548 12729
rect 604 12673 672 12729
rect 728 12673 768 12729
rect 260 12605 768 12673
rect 260 12549 300 12605
rect 356 12549 424 12605
rect 480 12549 548 12605
rect 604 12549 672 12605
rect 728 12549 768 12605
rect 260 10651 768 12549
rect 1136 12255 1336 14133
rect 1426 13845 1874 13855
rect 1426 13789 1436 13845
rect 1492 13789 1560 13845
rect 1616 13789 1684 13845
rect 1740 13789 1808 13845
rect 1864 13789 1874 13845
rect 1426 13721 1874 13789
rect 1426 13665 1436 13721
rect 1492 13665 1560 13721
rect 1616 13665 1684 13721
rect 1740 13665 1808 13721
rect 1864 13665 1874 13721
rect 1426 13597 1874 13665
rect 1426 13541 1436 13597
rect 1492 13541 1560 13597
rect 1616 13541 1684 13597
rect 1740 13541 1808 13597
rect 1864 13541 1874 13597
rect 1426 13473 1874 13541
rect 1426 13417 1436 13473
rect 1492 13417 1560 13473
rect 1616 13417 1684 13473
rect 1740 13417 1808 13473
rect 1864 13417 1874 13473
rect 1426 13349 1874 13417
rect 1426 13293 1436 13349
rect 1492 13293 1560 13349
rect 1616 13293 1684 13349
rect 1740 13293 1808 13349
rect 1864 13293 1874 13349
rect 1426 13225 1874 13293
rect 1426 13169 1436 13225
rect 1492 13169 1560 13225
rect 1616 13169 1684 13225
rect 1740 13169 1808 13225
rect 1864 13169 1874 13225
rect 1426 13101 1874 13169
rect 1426 13045 1436 13101
rect 1492 13045 1560 13101
rect 1616 13045 1684 13101
rect 1740 13045 1808 13101
rect 1864 13045 1874 13101
rect 1426 12977 1874 13045
rect 1426 12921 1436 12977
rect 1492 12921 1560 12977
rect 1616 12921 1684 12977
rect 1740 12921 1808 12977
rect 1864 12921 1874 12977
rect 1426 12853 1874 12921
rect 1426 12797 1436 12853
rect 1492 12797 1560 12853
rect 1616 12797 1684 12853
rect 1740 12797 1808 12853
rect 1864 12797 1874 12853
rect 1426 12729 1874 12797
rect 1426 12673 1436 12729
rect 1492 12673 1560 12729
rect 1616 12673 1684 12729
rect 1740 12673 1808 12729
rect 1864 12673 1874 12729
rect 1426 12605 1874 12673
rect 1426 12549 1436 12605
rect 1492 12549 1560 12605
rect 1616 12549 1684 12605
rect 1740 12549 1808 12605
rect 1864 12549 1874 12605
rect 1426 12539 1874 12549
rect 2562 13845 3010 13855
rect 2562 13789 2572 13845
rect 2628 13789 2696 13845
rect 2752 13789 2820 13845
rect 2876 13789 2944 13845
rect 3000 13789 3010 13845
rect 2562 13721 3010 13789
rect 2562 13665 2572 13721
rect 2628 13665 2696 13721
rect 2752 13665 2820 13721
rect 2876 13665 2944 13721
rect 3000 13665 3010 13721
rect 2562 13597 3010 13665
rect 2562 13541 2572 13597
rect 2628 13541 2696 13597
rect 2752 13541 2820 13597
rect 2876 13541 2944 13597
rect 3000 13541 3010 13597
rect 2562 13473 3010 13541
rect 2562 13417 2572 13473
rect 2628 13417 2696 13473
rect 2752 13417 2820 13473
rect 2876 13417 2944 13473
rect 3000 13417 3010 13473
rect 2562 13349 3010 13417
rect 2562 13293 2572 13349
rect 2628 13293 2696 13349
rect 2752 13293 2820 13349
rect 2876 13293 2944 13349
rect 3000 13293 3010 13349
rect 2562 13225 3010 13293
rect 2562 13169 2572 13225
rect 2628 13169 2696 13225
rect 2752 13169 2820 13225
rect 2876 13169 2944 13225
rect 3000 13169 3010 13225
rect 2562 13101 3010 13169
rect 2562 13045 2572 13101
rect 2628 13045 2696 13101
rect 2752 13045 2820 13101
rect 2876 13045 2944 13101
rect 3000 13045 3010 13101
rect 2562 12977 3010 13045
rect 2562 12921 2572 12977
rect 2628 12921 2696 12977
rect 2752 12921 2820 12977
rect 2876 12921 2944 12977
rect 3000 12921 3010 12977
rect 2562 12853 3010 12921
rect 2562 12797 2572 12853
rect 2628 12797 2696 12853
rect 2752 12797 2820 12853
rect 2876 12797 2944 12853
rect 3000 12797 3010 12853
rect 2562 12729 3010 12797
rect 2562 12673 2572 12729
rect 2628 12673 2696 12729
rect 2752 12673 2820 12729
rect 2876 12673 2944 12729
rect 3000 12673 3010 12729
rect 2562 12605 3010 12673
rect 2562 12549 2572 12605
rect 2628 12549 2696 12605
rect 2752 12549 2820 12605
rect 2876 12549 2944 12605
rect 3000 12549 3010 12605
rect 2562 12539 3010 12549
rect 4834 13845 5282 13855
rect 4834 13789 4844 13845
rect 4900 13789 4968 13845
rect 5024 13789 5092 13845
rect 5148 13789 5216 13845
rect 5272 13789 5282 13845
rect 4834 13721 5282 13789
rect 4834 13665 4844 13721
rect 4900 13665 4968 13721
rect 5024 13665 5092 13721
rect 5148 13665 5216 13721
rect 5272 13665 5282 13721
rect 4834 13597 5282 13665
rect 4834 13541 4844 13597
rect 4900 13541 4968 13597
rect 5024 13541 5092 13597
rect 5148 13541 5216 13597
rect 5272 13541 5282 13597
rect 4834 13473 5282 13541
rect 4834 13417 4844 13473
rect 4900 13417 4968 13473
rect 5024 13417 5092 13473
rect 5148 13417 5216 13473
rect 5272 13417 5282 13473
rect 4834 13349 5282 13417
rect 4834 13293 4844 13349
rect 4900 13293 4968 13349
rect 5024 13293 5092 13349
rect 5148 13293 5216 13349
rect 5272 13293 5282 13349
rect 4834 13225 5282 13293
rect 4834 13169 4844 13225
rect 4900 13169 4968 13225
rect 5024 13169 5092 13225
rect 5148 13169 5216 13225
rect 5272 13169 5282 13225
rect 4834 13101 5282 13169
rect 4834 13045 4844 13101
rect 4900 13045 4968 13101
rect 5024 13045 5092 13101
rect 5148 13045 5216 13101
rect 5272 13045 5282 13101
rect 4834 12977 5282 13045
rect 4834 12921 4844 12977
rect 4900 12921 4968 12977
rect 5024 12921 5092 12977
rect 5148 12921 5216 12977
rect 5272 12921 5282 12977
rect 4834 12853 5282 12921
rect 4834 12797 4844 12853
rect 4900 12797 4968 12853
rect 5024 12797 5092 12853
rect 5148 12797 5216 12853
rect 5272 12797 5282 12853
rect 4834 12729 5282 12797
rect 4834 12673 4844 12729
rect 4900 12673 4968 12729
rect 5024 12673 5092 12729
rect 5148 12673 5216 12729
rect 5272 12673 5282 12729
rect 4834 12605 5282 12673
rect 4834 12549 4844 12605
rect 4900 12549 4968 12605
rect 5024 12549 5092 12605
rect 5148 12549 5216 12605
rect 5272 12549 5282 12605
rect 4834 12539 5282 12549
rect 7127 13845 7451 13855
rect 7127 13789 7137 13845
rect 7193 13789 7261 13845
rect 7317 13789 7385 13845
rect 7441 13789 7451 13845
rect 7127 13721 7451 13789
rect 7127 13665 7137 13721
rect 7193 13665 7261 13721
rect 7317 13665 7385 13721
rect 7441 13665 7451 13721
rect 7127 13597 7451 13665
rect 7127 13541 7137 13597
rect 7193 13541 7261 13597
rect 7317 13541 7385 13597
rect 7441 13541 7451 13597
rect 7127 13473 7451 13541
rect 7127 13417 7137 13473
rect 7193 13417 7261 13473
rect 7317 13417 7385 13473
rect 7441 13417 7451 13473
rect 7127 13349 7451 13417
rect 7127 13293 7137 13349
rect 7193 13293 7261 13349
rect 7317 13293 7385 13349
rect 7441 13293 7451 13349
rect 7127 13225 7451 13293
rect 7127 13169 7137 13225
rect 7193 13169 7261 13225
rect 7317 13169 7385 13225
rect 7441 13169 7451 13225
rect 7127 13101 7451 13169
rect 7127 13045 7137 13101
rect 7193 13045 7261 13101
rect 7317 13045 7385 13101
rect 7441 13045 7451 13101
rect 7127 12977 7451 13045
rect 7127 12921 7137 12977
rect 7193 12921 7261 12977
rect 7317 12921 7385 12977
rect 7441 12921 7451 12977
rect 7127 12853 7451 12921
rect 7127 12797 7137 12853
rect 7193 12797 7261 12853
rect 7317 12797 7385 12853
rect 7441 12797 7451 12853
rect 7127 12729 7451 12797
rect 7127 12673 7137 12729
rect 7193 12673 7261 12729
rect 7317 12673 7385 12729
rect 7441 12673 7451 12729
rect 7127 12605 7451 12673
rect 7127 12549 7137 12605
rect 7193 12549 7261 12605
rect 7317 12549 7385 12605
rect 7441 12549 7451 12605
rect 7127 12539 7451 12549
rect 7613 13845 7937 13855
rect 7613 13789 7623 13845
rect 7679 13789 7747 13845
rect 7803 13789 7871 13845
rect 7927 13789 7937 13845
rect 7613 13721 7937 13789
rect 7613 13665 7623 13721
rect 7679 13665 7747 13721
rect 7803 13665 7871 13721
rect 7927 13665 7937 13721
rect 7613 13597 7937 13665
rect 7613 13541 7623 13597
rect 7679 13541 7747 13597
rect 7803 13541 7871 13597
rect 7927 13541 7937 13597
rect 7613 13473 7937 13541
rect 7613 13417 7623 13473
rect 7679 13417 7747 13473
rect 7803 13417 7871 13473
rect 7927 13417 7937 13473
rect 7613 13349 7937 13417
rect 7613 13293 7623 13349
rect 7679 13293 7747 13349
rect 7803 13293 7871 13349
rect 7927 13293 7937 13349
rect 7613 13225 7937 13293
rect 7613 13169 7623 13225
rect 7679 13169 7747 13225
rect 7803 13169 7871 13225
rect 7927 13169 7937 13225
rect 7613 13101 7937 13169
rect 7613 13045 7623 13101
rect 7679 13045 7747 13101
rect 7803 13045 7871 13101
rect 7927 13045 7937 13101
rect 7613 12977 7937 13045
rect 7613 12921 7623 12977
rect 7679 12921 7747 12977
rect 7803 12921 7871 12977
rect 7927 12921 7937 12977
rect 7613 12853 7937 12921
rect 7613 12797 7623 12853
rect 7679 12797 7747 12853
rect 7803 12797 7871 12853
rect 7927 12797 7937 12853
rect 7613 12729 7937 12797
rect 7613 12673 7623 12729
rect 7679 12673 7747 12729
rect 7803 12673 7871 12729
rect 7927 12673 7937 12729
rect 7613 12605 7937 12673
rect 7613 12549 7623 12605
rect 7679 12549 7747 12605
rect 7803 12549 7871 12605
rect 7927 12549 7937 12605
rect 7613 12539 7937 12549
rect 9782 13845 10230 13855
rect 9782 13789 9792 13845
rect 9848 13789 9916 13845
rect 9972 13789 10040 13845
rect 10096 13789 10164 13845
rect 10220 13789 10230 13845
rect 9782 13721 10230 13789
rect 9782 13665 9792 13721
rect 9848 13665 9916 13721
rect 9972 13665 10040 13721
rect 10096 13665 10164 13721
rect 10220 13665 10230 13721
rect 9782 13597 10230 13665
rect 9782 13541 9792 13597
rect 9848 13541 9916 13597
rect 9972 13541 10040 13597
rect 10096 13541 10164 13597
rect 10220 13541 10230 13597
rect 9782 13473 10230 13541
rect 9782 13417 9792 13473
rect 9848 13417 9916 13473
rect 9972 13417 10040 13473
rect 10096 13417 10164 13473
rect 10220 13417 10230 13473
rect 9782 13349 10230 13417
rect 9782 13293 9792 13349
rect 9848 13293 9916 13349
rect 9972 13293 10040 13349
rect 10096 13293 10164 13349
rect 10220 13293 10230 13349
rect 9782 13225 10230 13293
rect 9782 13169 9792 13225
rect 9848 13169 9916 13225
rect 9972 13169 10040 13225
rect 10096 13169 10164 13225
rect 10220 13169 10230 13225
rect 9782 13101 10230 13169
rect 9782 13045 9792 13101
rect 9848 13045 9916 13101
rect 9972 13045 10040 13101
rect 10096 13045 10164 13101
rect 10220 13045 10230 13101
rect 9782 12977 10230 13045
rect 9782 12921 9792 12977
rect 9848 12921 9916 12977
rect 9972 12921 10040 12977
rect 10096 12921 10164 12977
rect 10220 12921 10230 12977
rect 9782 12853 10230 12921
rect 9782 12797 9792 12853
rect 9848 12797 9916 12853
rect 9972 12797 10040 12853
rect 10096 12797 10164 12853
rect 10220 12797 10230 12853
rect 9782 12729 10230 12797
rect 9782 12673 9792 12729
rect 9848 12673 9916 12729
rect 9972 12673 10040 12729
rect 10096 12673 10164 12729
rect 10220 12673 10230 12729
rect 9782 12605 10230 12673
rect 9782 12549 9792 12605
rect 9848 12549 9916 12605
rect 9972 12549 10040 12605
rect 10096 12549 10164 12605
rect 10220 12549 10230 12605
rect 9782 12539 10230 12549
rect 12054 13845 12502 13855
rect 12054 13789 12064 13845
rect 12120 13789 12188 13845
rect 12244 13789 12312 13845
rect 12368 13789 12436 13845
rect 12492 13789 12502 13845
rect 12054 13721 12502 13789
rect 12054 13665 12064 13721
rect 12120 13665 12188 13721
rect 12244 13665 12312 13721
rect 12368 13665 12436 13721
rect 12492 13665 12502 13721
rect 12054 13597 12502 13665
rect 12054 13541 12064 13597
rect 12120 13541 12188 13597
rect 12244 13541 12312 13597
rect 12368 13541 12436 13597
rect 12492 13541 12502 13597
rect 12054 13473 12502 13541
rect 12054 13417 12064 13473
rect 12120 13417 12188 13473
rect 12244 13417 12312 13473
rect 12368 13417 12436 13473
rect 12492 13417 12502 13473
rect 12054 13349 12502 13417
rect 12054 13293 12064 13349
rect 12120 13293 12188 13349
rect 12244 13293 12312 13349
rect 12368 13293 12436 13349
rect 12492 13293 12502 13349
rect 12054 13225 12502 13293
rect 12054 13169 12064 13225
rect 12120 13169 12188 13225
rect 12244 13169 12312 13225
rect 12368 13169 12436 13225
rect 12492 13169 12502 13225
rect 12054 13101 12502 13169
rect 12054 13045 12064 13101
rect 12120 13045 12188 13101
rect 12244 13045 12312 13101
rect 12368 13045 12436 13101
rect 12492 13045 12502 13101
rect 12054 12977 12502 13045
rect 12054 12921 12064 12977
rect 12120 12921 12188 12977
rect 12244 12921 12312 12977
rect 12368 12921 12436 12977
rect 12492 12921 12502 12977
rect 12054 12853 12502 12921
rect 12054 12797 12064 12853
rect 12120 12797 12188 12853
rect 12244 12797 12312 12853
rect 12368 12797 12436 12853
rect 12492 12797 12502 12853
rect 12054 12729 12502 12797
rect 12054 12673 12064 12729
rect 12120 12673 12188 12729
rect 12244 12673 12312 12729
rect 12368 12673 12436 12729
rect 12492 12673 12502 12729
rect 12054 12605 12502 12673
rect 12054 12549 12064 12605
rect 12120 12549 12188 12605
rect 12244 12549 12312 12605
rect 12368 12549 12436 12605
rect 12492 12549 12502 12605
rect 12054 12539 12502 12549
rect 13190 13845 13638 13855
rect 13190 13789 13200 13845
rect 13256 13789 13324 13845
rect 13380 13789 13448 13845
rect 13504 13789 13572 13845
rect 13628 13789 13638 13845
rect 13190 13721 13638 13789
rect 13190 13665 13200 13721
rect 13256 13665 13324 13721
rect 13380 13665 13448 13721
rect 13504 13665 13572 13721
rect 13628 13665 13638 13721
rect 13190 13597 13638 13665
rect 13190 13541 13200 13597
rect 13256 13541 13324 13597
rect 13380 13541 13448 13597
rect 13504 13541 13572 13597
rect 13628 13541 13638 13597
rect 13190 13473 13638 13541
rect 13190 13417 13200 13473
rect 13256 13417 13324 13473
rect 13380 13417 13448 13473
rect 13504 13417 13572 13473
rect 13628 13417 13638 13473
rect 13190 13349 13638 13417
rect 13190 13293 13200 13349
rect 13256 13293 13324 13349
rect 13380 13293 13448 13349
rect 13504 13293 13572 13349
rect 13628 13293 13638 13349
rect 13190 13225 13638 13293
rect 13190 13169 13200 13225
rect 13256 13169 13324 13225
rect 13380 13169 13448 13225
rect 13504 13169 13572 13225
rect 13628 13169 13638 13225
rect 13190 13101 13638 13169
rect 13190 13045 13200 13101
rect 13256 13045 13324 13101
rect 13380 13045 13448 13101
rect 13504 13045 13572 13101
rect 13628 13045 13638 13101
rect 13190 12977 13638 13045
rect 13190 12921 13200 12977
rect 13256 12921 13324 12977
rect 13380 12921 13448 12977
rect 13504 12921 13572 12977
rect 13628 12921 13638 12977
rect 13190 12853 13638 12921
rect 13190 12797 13200 12853
rect 13256 12797 13324 12853
rect 13380 12797 13448 12853
rect 13504 12797 13572 12853
rect 13628 12797 13638 12853
rect 13190 12729 13638 12797
rect 13190 12673 13200 12729
rect 13256 12673 13324 12729
rect 13380 12673 13448 12729
rect 13504 12673 13572 12729
rect 13628 12673 13638 12729
rect 13190 12605 13638 12673
rect 13190 12549 13200 12605
rect 13256 12549 13324 12605
rect 13380 12549 13448 12605
rect 13504 12549 13572 12605
rect 13628 12549 13638 12605
rect 13190 12539 13638 12549
rect 858 12245 1336 12255
rect 858 12189 868 12245
rect 924 12189 992 12245
rect 1048 12189 1116 12245
rect 1172 12189 1240 12245
rect 1296 12189 1336 12245
rect 858 12121 1336 12189
rect 858 12065 868 12121
rect 924 12065 992 12121
rect 1048 12065 1116 12121
rect 1172 12065 1240 12121
rect 1296 12065 1336 12121
rect 858 11997 1336 12065
rect 858 11941 868 11997
rect 924 11941 992 11997
rect 1048 11941 1116 11997
rect 1172 11941 1240 11997
rect 1296 11941 1336 11997
rect 858 11873 1336 11941
rect 858 11817 868 11873
rect 924 11817 992 11873
rect 1048 11817 1116 11873
rect 1172 11817 1240 11873
rect 1296 11817 1336 11873
rect 858 11749 1336 11817
rect 858 11693 868 11749
rect 924 11693 992 11749
rect 1048 11693 1116 11749
rect 1172 11693 1240 11749
rect 1296 11693 1336 11749
rect 858 11625 1336 11693
rect 858 11569 868 11625
rect 924 11569 992 11625
rect 1048 11569 1116 11625
rect 1172 11569 1240 11625
rect 1296 11569 1336 11625
rect 858 11501 1336 11569
rect 858 11445 868 11501
rect 924 11445 992 11501
rect 1048 11445 1116 11501
rect 1172 11445 1240 11501
rect 1296 11445 1336 11501
rect 858 11377 1336 11445
rect 858 11321 868 11377
rect 924 11321 992 11377
rect 1048 11321 1116 11377
rect 1172 11321 1240 11377
rect 1296 11321 1336 11377
rect 858 11253 1336 11321
rect 858 11197 868 11253
rect 924 11197 992 11253
rect 1048 11197 1116 11253
rect 1172 11197 1240 11253
rect 1296 11197 1336 11253
rect 858 11129 1336 11197
rect 858 11073 868 11129
rect 924 11073 992 11129
rect 1048 11073 1116 11129
rect 1172 11073 1240 11129
rect 1296 11073 1336 11129
rect 858 11005 1336 11073
rect 858 10949 868 11005
rect 924 10949 992 11005
rect 1048 10949 1116 11005
rect 1172 10949 1240 11005
rect 1296 10949 1336 11005
rect 858 10939 1336 10949
rect 1994 12245 2442 12255
rect 1994 12189 2004 12245
rect 2060 12189 2128 12245
rect 2184 12189 2252 12245
rect 2308 12189 2376 12245
rect 2432 12189 2442 12245
rect 1994 12121 2442 12189
rect 1994 12065 2004 12121
rect 2060 12065 2128 12121
rect 2184 12065 2252 12121
rect 2308 12065 2376 12121
rect 2432 12065 2442 12121
rect 1994 11997 2442 12065
rect 1994 11941 2004 11997
rect 2060 11941 2128 11997
rect 2184 11941 2252 11997
rect 2308 11941 2376 11997
rect 2432 11941 2442 11997
rect 1994 11873 2442 11941
rect 1994 11817 2004 11873
rect 2060 11817 2128 11873
rect 2184 11817 2252 11873
rect 2308 11817 2376 11873
rect 2432 11817 2442 11873
rect 1994 11749 2442 11817
rect 1994 11693 2004 11749
rect 2060 11693 2128 11749
rect 2184 11693 2252 11749
rect 2308 11693 2376 11749
rect 2432 11693 2442 11749
rect 1994 11625 2442 11693
rect 1994 11569 2004 11625
rect 2060 11569 2128 11625
rect 2184 11569 2252 11625
rect 2308 11569 2376 11625
rect 2432 11569 2442 11625
rect 1994 11501 2442 11569
rect 1994 11445 2004 11501
rect 2060 11445 2128 11501
rect 2184 11445 2252 11501
rect 2308 11445 2376 11501
rect 2432 11445 2442 11501
rect 1994 11377 2442 11445
rect 1994 11321 2004 11377
rect 2060 11321 2128 11377
rect 2184 11321 2252 11377
rect 2308 11321 2376 11377
rect 2432 11321 2442 11377
rect 1994 11253 2442 11321
rect 1994 11197 2004 11253
rect 2060 11197 2128 11253
rect 2184 11197 2252 11253
rect 2308 11197 2376 11253
rect 2432 11197 2442 11253
rect 1994 11129 2442 11197
rect 1994 11073 2004 11129
rect 2060 11073 2128 11129
rect 2184 11073 2252 11129
rect 2308 11073 2376 11129
rect 2432 11073 2442 11129
rect 1994 11005 2442 11073
rect 1994 10949 2004 11005
rect 2060 10949 2128 11005
rect 2184 10949 2252 11005
rect 2308 10949 2376 11005
rect 2432 10949 2442 11005
rect 1994 10939 2442 10949
rect 3698 12245 4146 12255
rect 3698 12189 3708 12245
rect 3764 12189 3832 12245
rect 3888 12189 3956 12245
rect 4012 12189 4080 12245
rect 4136 12189 4146 12245
rect 3698 12121 4146 12189
rect 3698 12065 3708 12121
rect 3764 12065 3832 12121
rect 3888 12065 3956 12121
rect 4012 12065 4080 12121
rect 4136 12065 4146 12121
rect 3698 11997 4146 12065
rect 3698 11941 3708 11997
rect 3764 11941 3832 11997
rect 3888 11941 3956 11997
rect 4012 11941 4080 11997
rect 4136 11941 4146 11997
rect 3698 11873 4146 11941
rect 3698 11817 3708 11873
rect 3764 11817 3832 11873
rect 3888 11817 3956 11873
rect 4012 11817 4080 11873
rect 4136 11817 4146 11873
rect 3698 11749 4146 11817
rect 3698 11693 3708 11749
rect 3764 11693 3832 11749
rect 3888 11693 3956 11749
rect 4012 11693 4080 11749
rect 4136 11693 4146 11749
rect 3698 11625 4146 11693
rect 3698 11569 3708 11625
rect 3764 11569 3832 11625
rect 3888 11569 3956 11625
rect 4012 11569 4080 11625
rect 4136 11569 4146 11625
rect 3698 11501 4146 11569
rect 3698 11445 3708 11501
rect 3764 11445 3832 11501
rect 3888 11445 3956 11501
rect 4012 11445 4080 11501
rect 4136 11445 4146 11501
rect 3698 11377 4146 11445
rect 3698 11321 3708 11377
rect 3764 11321 3832 11377
rect 3888 11321 3956 11377
rect 4012 11321 4080 11377
rect 4136 11321 4146 11377
rect 3698 11253 4146 11321
rect 3698 11197 3708 11253
rect 3764 11197 3832 11253
rect 3888 11197 3956 11253
rect 4012 11197 4080 11253
rect 4136 11197 4146 11253
rect 3698 11129 4146 11197
rect 3698 11073 3708 11129
rect 3764 11073 3832 11129
rect 3888 11073 3956 11129
rect 4012 11073 4080 11129
rect 4136 11073 4146 11129
rect 3698 11005 4146 11073
rect 3698 10949 3708 11005
rect 3764 10949 3832 11005
rect 3888 10949 3956 11005
rect 4012 10949 4080 11005
rect 4136 10949 4146 11005
rect 3698 10939 4146 10949
rect 5970 12245 6418 12255
rect 5970 12189 5980 12245
rect 6036 12189 6104 12245
rect 6160 12189 6228 12245
rect 6284 12189 6352 12245
rect 6408 12189 6418 12245
rect 5970 12121 6418 12189
rect 5970 12065 5980 12121
rect 6036 12065 6104 12121
rect 6160 12065 6228 12121
rect 6284 12065 6352 12121
rect 6408 12065 6418 12121
rect 5970 11997 6418 12065
rect 5970 11941 5980 11997
rect 6036 11941 6104 11997
rect 6160 11941 6228 11997
rect 6284 11941 6352 11997
rect 6408 11941 6418 11997
rect 5970 11873 6418 11941
rect 5970 11817 5980 11873
rect 6036 11817 6104 11873
rect 6160 11817 6228 11873
rect 6284 11817 6352 11873
rect 6408 11817 6418 11873
rect 5970 11749 6418 11817
rect 5970 11693 5980 11749
rect 6036 11693 6104 11749
rect 6160 11693 6228 11749
rect 6284 11693 6352 11749
rect 6408 11693 6418 11749
rect 5970 11625 6418 11693
rect 5970 11569 5980 11625
rect 6036 11569 6104 11625
rect 6160 11569 6228 11625
rect 6284 11569 6352 11625
rect 6408 11569 6418 11625
rect 5970 11501 6418 11569
rect 5970 11445 5980 11501
rect 6036 11445 6104 11501
rect 6160 11445 6228 11501
rect 6284 11445 6352 11501
rect 6408 11445 6418 11501
rect 5970 11377 6418 11445
rect 5970 11321 5980 11377
rect 6036 11321 6104 11377
rect 6160 11321 6228 11377
rect 6284 11321 6352 11377
rect 6408 11321 6418 11377
rect 5970 11253 6418 11321
rect 5970 11197 5980 11253
rect 6036 11197 6104 11253
rect 6160 11197 6228 11253
rect 6284 11197 6352 11253
rect 6408 11197 6418 11253
rect 5970 11129 6418 11197
rect 5970 11073 5980 11129
rect 6036 11073 6104 11129
rect 6160 11073 6228 11129
rect 6284 11073 6352 11129
rect 6408 11073 6418 11129
rect 5970 11005 6418 11073
rect 5970 10949 5980 11005
rect 6036 10949 6104 11005
rect 6160 10949 6228 11005
rect 6284 10949 6352 11005
rect 6408 10949 6418 11005
rect 5970 10939 6418 10949
rect 8646 12245 9094 12255
rect 8646 12189 8656 12245
rect 8712 12189 8780 12245
rect 8836 12189 8904 12245
rect 8960 12189 9028 12245
rect 9084 12189 9094 12245
rect 8646 12121 9094 12189
rect 8646 12065 8656 12121
rect 8712 12065 8780 12121
rect 8836 12065 8904 12121
rect 8960 12065 9028 12121
rect 9084 12065 9094 12121
rect 8646 11997 9094 12065
rect 8646 11941 8656 11997
rect 8712 11941 8780 11997
rect 8836 11941 8904 11997
rect 8960 11941 9028 11997
rect 9084 11941 9094 11997
rect 8646 11873 9094 11941
rect 8646 11817 8656 11873
rect 8712 11817 8780 11873
rect 8836 11817 8904 11873
rect 8960 11817 9028 11873
rect 9084 11817 9094 11873
rect 8646 11749 9094 11817
rect 8646 11693 8656 11749
rect 8712 11693 8780 11749
rect 8836 11693 8904 11749
rect 8960 11693 9028 11749
rect 9084 11693 9094 11749
rect 8646 11625 9094 11693
rect 8646 11569 8656 11625
rect 8712 11569 8780 11625
rect 8836 11569 8904 11625
rect 8960 11569 9028 11625
rect 9084 11569 9094 11625
rect 8646 11501 9094 11569
rect 8646 11445 8656 11501
rect 8712 11445 8780 11501
rect 8836 11445 8904 11501
rect 8960 11445 9028 11501
rect 9084 11445 9094 11501
rect 8646 11377 9094 11445
rect 8646 11321 8656 11377
rect 8712 11321 8780 11377
rect 8836 11321 8904 11377
rect 8960 11321 9028 11377
rect 9084 11321 9094 11377
rect 8646 11253 9094 11321
rect 8646 11197 8656 11253
rect 8712 11197 8780 11253
rect 8836 11197 8904 11253
rect 8960 11197 9028 11253
rect 9084 11197 9094 11253
rect 8646 11129 9094 11197
rect 8646 11073 8656 11129
rect 8712 11073 8780 11129
rect 8836 11073 8904 11129
rect 8960 11073 9028 11129
rect 9084 11073 9094 11129
rect 8646 11005 9094 11073
rect 8646 10949 8656 11005
rect 8712 10949 8780 11005
rect 8836 10949 8904 11005
rect 8960 10949 9028 11005
rect 9084 10949 9094 11005
rect 8646 10939 9094 10949
rect 10918 12245 11366 12255
rect 10918 12189 10928 12245
rect 10984 12189 11052 12245
rect 11108 12189 11176 12245
rect 11232 12189 11300 12245
rect 11356 12189 11366 12245
rect 10918 12121 11366 12189
rect 10918 12065 10928 12121
rect 10984 12065 11052 12121
rect 11108 12065 11176 12121
rect 11232 12065 11300 12121
rect 11356 12065 11366 12121
rect 10918 11997 11366 12065
rect 10918 11941 10928 11997
rect 10984 11941 11052 11997
rect 11108 11941 11176 11997
rect 11232 11941 11300 11997
rect 11356 11941 11366 11997
rect 10918 11873 11366 11941
rect 10918 11817 10928 11873
rect 10984 11817 11052 11873
rect 11108 11817 11176 11873
rect 11232 11817 11300 11873
rect 11356 11817 11366 11873
rect 10918 11749 11366 11817
rect 10918 11693 10928 11749
rect 10984 11693 11052 11749
rect 11108 11693 11176 11749
rect 11232 11693 11300 11749
rect 11356 11693 11366 11749
rect 10918 11625 11366 11693
rect 10918 11569 10928 11625
rect 10984 11569 11052 11625
rect 11108 11569 11176 11625
rect 11232 11569 11300 11625
rect 11356 11569 11366 11625
rect 10918 11501 11366 11569
rect 10918 11445 10928 11501
rect 10984 11445 11052 11501
rect 11108 11445 11176 11501
rect 11232 11445 11300 11501
rect 11356 11445 11366 11501
rect 10918 11377 11366 11445
rect 10918 11321 10928 11377
rect 10984 11321 11052 11377
rect 11108 11321 11176 11377
rect 11232 11321 11300 11377
rect 11356 11321 11366 11377
rect 10918 11253 11366 11321
rect 10918 11197 10928 11253
rect 10984 11197 11052 11253
rect 11108 11197 11176 11253
rect 11232 11197 11300 11253
rect 11356 11197 11366 11253
rect 10918 11129 11366 11197
rect 10918 11073 10928 11129
rect 10984 11073 11052 11129
rect 11108 11073 11176 11129
rect 11232 11073 11300 11129
rect 11356 11073 11366 11129
rect 10918 11005 11366 11073
rect 10918 10949 10928 11005
rect 10984 10949 11052 11005
rect 11108 10949 11176 11005
rect 11232 10949 11300 11005
rect 11356 10949 11366 11005
rect 10918 10939 11366 10949
rect 12622 12245 13070 12255
rect 12622 12189 12632 12245
rect 12688 12189 12756 12245
rect 12812 12189 12880 12245
rect 12936 12189 13004 12245
rect 13060 12189 13070 12245
rect 12622 12121 13070 12189
rect 12622 12065 12632 12121
rect 12688 12065 12756 12121
rect 12812 12065 12880 12121
rect 12936 12065 13004 12121
rect 13060 12065 13070 12121
rect 12622 11997 13070 12065
rect 12622 11941 12632 11997
rect 12688 11941 12756 11997
rect 12812 11941 12880 11997
rect 12936 11941 13004 11997
rect 13060 11941 13070 11997
rect 12622 11873 13070 11941
rect 12622 11817 12632 11873
rect 12688 11817 12756 11873
rect 12812 11817 12880 11873
rect 12936 11817 13004 11873
rect 13060 11817 13070 11873
rect 12622 11749 13070 11817
rect 12622 11693 12632 11749
rect 12688 11693 12756 11749
rect 12812 11693 12880 11749
rect 12936 11693 13004 11749
rect 13060 11693 13070 11749
rect 12622 11625 13070 11693
rect 12622 11569 12632 11625
rect 12688 11569 12756 11625
rect 12812 11569 12880 11625
rect 12936 11569 13004 11625
rect 13060 11569 13070 11625
rect 12622 11501 13070 11569
rect 12622 11445 12632 11501
rect 12688 11445 12756 11501
rect 12812 11445 12880 11501
rect 12936 11445 13004 11501
rect 13060 11445 13070 11501
rect 12622 11377 13070 11445
rect 12622 11321 12632 11377
rect 12688 11321 12756 11377
rect 12812 11321 12880 11377
rect 12936 11321 13004 11377
rect 13060 11321 13070 11377
rect 12622 11253 13070 11321
rect 12622 11197 12632 11253
rect 12688 11197 12756 11253
rect 12812 11197 12880 11253
rect 12936 11197 13004 11253
rect 13060 11197 13070 11253
rect 12622 11129 13070 11197
rect 12622 11073 12632 11129
rect 12688 11073 12756 11129
rect 12812 11073 12880 11129
rect 12936 11073 13004 11129
rect 13060 11073 13070 11129
rect 12622 11005 13070 11073
rect 12622 10949 12632 11005
rect 12688 10949 12756 11005
rect 12812 10949 12880 11005
rect 12936 10949 13004 11005
rect 13060 10949 13070 11005
rect 12622 10939 13070 10949
rect 13728 12245 14236 14143
rect 13728 12189 13768 12245
rect 13824 12189 13892 12245
rect 13948 12189 14016 12245
rect 14072 12189 14140 12245
rect 14196 12189 14236 12245
rect 13728 12121 14236 12189
rect 13728 12065 13768 12121
rect 13824 12065 13892 12121
rect 13948 12065 14016 12121
rect 14072 12065 14140 12121
rect 14196 12065 14236 12121
rect 13728 11997 14236 12065
rect 13728 11941 13768 11997
rect 13824 11941 13892 11997
rect 13948 11941 14016 11997
rect 14072 11941 14140 11997
rect 14196 11941 14236 11997
rect 13728 11873 14236 11941
rect 13728 11817 13768 11873
rect 13824 11817 13892 11873
rect 13948 11817 14016 11873
rect 14072 11817 14140 11873
rect 14196 11817 14236 11873
rect 13728 11749 14236 11817
rect 13728 11693 13768 11749
rect 13824 11693 13892 11749
rect 13948 11693 14016 11749
rect 14072 11693 14140 11749
rect 14196 11693 14236 11749
rect 13728 11625 14236 11693
rect 13728 11569 13768 11625
rect 13824 11569 13892 11625
rect 13948 11569 14016 11625
rect 14072 11569 14140 11625
rect 14196 11569 14236 11625
rect 13728 11501 14236 11569
rect 13728 11445 13768 11501
rect 13824 11445 13892 11501
rect 13948 11445 14016 11501
rect 14072 11445 14140 11501
rect 14196 11445 14236 11501
rect 13728 11377 14236 11445
rect 13728 11321 13768 11377
rect 13824 11321 13892 11377
rect 13948 11321 14016 11377
rect 14072 11321 14140 11377
rect 14196 11321 14236 11377
rect 13728 11253 14236 11321
rect 13728 11197 13768 11253
rect 13824 11197 13892 11253
rect 13948 11197 14016 11253
rect 14072 11197 14140 11253
rect 14196 11197 14236 11253
rect 13728 11129 14236 11197
rect 13728 11073 13768 11129
rect 13824 11073 13892 11129
rect 13948 11073 14016 11129
rect 14072 11073 14140 11129
rect 14196 11073 14236 11129
rect 13728 11005 14236 11073
rect 13728 10949 13768 11005
rect 13824 10949 13892 11005
rect 13948 10949 14016 11005
rect 14072 10949 14140 11005
rect 14196 10949 14236 11005
rect 260 10595 300 10651
rect 356 10595 424 10651
rect 480 10595 548 10651
rect 604 10595 672 10651
rect 728 10595 768 10651
rect 260 10527 768 10595
rect 260 10471 300 10527
rect 356 10471 424 10527
rect 480 10471 548 10527
rect 604 10471 672 10527
rect 728 10471 768 10527
rect 260 10403 768 10471
rect 260 10347 300 10403
rect 356 10347 424 10403
rect 480 10347 548 10403
rect 604 10347 672 10403
rect 728 10347 768 10403
rect 260 10279 768 10347
rect 260 10223 300 10279
rect 356 10223 424 10279
rect 480 10223 548 10279
rect 604 10223 672 10279
rect 728 10223 768 10279
rect 260 10155 768 10223
rect 260 10099 300 10155
rect 356 10099 424 10155
rect 480 10099 548 10155
rect 604 10099 672 10155
rect 728 10099 768 10155
rect 260 10031 768 10099
rect 260 9975 300 10031
rect 356 9975 424 10031
rect 480 9975 548 10031
rect 604 9975 672 10031
rect 728 9975 768 10031
rect 260 9907 768 9975
rect 260 9851 300 9907
rect 356 9851 424 9907
rect 480 9851 548 9907
rect 604 9851 672 9907
rect 728 9851 768 9907
rect 260 9783 768 9851
rect 260 9727 300 9783
rect 356 9727 424 9783
rect 480 9727 548 9783
rect 604 9727 672 9783
rect 728 9727 768 9783
rect 260 9659 768 9727
rect 260 9603 300 9659
rect 356 9603 424 9659
rect 480 9603 548 9659
rect 604 9603 672 9659
rect 728 9603 768 9659
rect 260 9535 768 9603
rect 260 9479 300 9535
rect 356 9479 424 9535
rect 480 9479 548 9535
rect 604 9479 672 9535
rect 728 9479 768 9535
rect 260 9411 768 9479
rect 260 9355 300 9411
rect 356 9355 424 9411
rect 480 9355 548 9411
rect 604 9355 672 9411
rect 728 9355 768 9411
rect 260 9287 768 9355
rect 260 9231 300 9287
rect 356 9231 424 9287
rect 480 9231 548 9287
rect 604 9231 672 9287
rect 728 9231 768 9287
rect 260 9163 768 9231
rect 260 9107 300 9163
rect 356 9107 424 9163
rect 480 9107 548 9163
rect 604 9107 672 9163
rect 728 9107 768 9163
rect 260 9039 768 9107
rect 260 8983 300 9039
rect 356 8983 424 9039
rect 480 8983 548 9039
rect 604 8983 672 9039
rect 728 8983 768 9039
rect 260 8915 768 8983
rect 260 8859 300 8915
rect 356 8859 424 8915
rect 480 8859 548 8915
rect 604 8859 672 8915
rect 728 8859 768 8915
rect 260 8791 768 8859
rect 260 8735 300 8791
rect 356 8735 424 8791
rect 480 8735 548 8791
rect 604 8735 672 8791
rect 728 8735 768 8791
rect 260 8667 768 8735
rect 260 8611 300 8667
rect 356 8611 424 8667
rect 480 8611 548 8667
rect 604 8611 672 8667
rect 728 8611 768 8667
rect 260 8543 768 8611
rect 260 8487 300 8543
rect 356 8487 424 8543
rect 480 8487 548 8543
rect 604 8487 672 8543
rect 728 8487 768 8543
rect 260 8419 768 8487
rect 260 8363 300 8419
rect 356 8363 424 8419
rect 480 8363 548 8419
rect 604 8363 672 8419
rect 728 8363 768 8419
rect 260 8295 768 8363
rect 260 8239 300 8295
rect 356 8239 424 8295
rect 480 8239 548 8295
rect 604 8239 672 8295
rect 728 8239 768 8295
rect 260 8171 768 8239
rect 260 8115 300 8171
rect 356 8115 424 8171
rect 480 8115 548 8171
rect 604 8115 672 8171
rect 728 8115 768 8171
rect 260 8047 768 8115
rect 260 7991 300 8047
rect 356 7991 424 8047
rect 480 7991 548 8047
rect 604 7991 672 8047
rect 728 7991 768 8047
rect 260 7923 768 7991
rect 260 7867 300 7923
rect 356 7867 424 7923
rect 480 7867 548 7923
rect 604 7867 672 7923
rect 728 7867 768 7923
rect 260 7799 768 7867
rect 260 7743 300 7799
rect 356 7743 424 7799
rect 480 7743 548 7799
rect 604 7743 672 7799
rect 728 7743 768 7799
rect 260 7451 768 7743
rect 260 7395 300 7451
rect 356 7395 424 7451
rect 480 7395 548 7451
rect 604 7395 672 7451
rect 728 7395 768 7451
rect 260 7327 768 7395
rect 260 7271 300 7327
rect 356 7271 424 7327
rect 480 7271 548 7327
rect 604 7271 672 7327
rect 728 7271 768 7327
rect 260 7203 768 7271
rect 260 7147 300 7203
rect 356 7147 424 7203
rect 480 7147 548 7203
rect 604 7147 672 7203
rect 728 7147 768 7203
rect 260 7079 768 7147
rect 260 7023 300 7079
rect 356 7023 424 7079
rect 480 7023 548 7079
rect 604 7023 672 7079
rect 728 7023 768 7079
rect 260 6955 768 7023
rect 260 6899 300 6955
rect 356 6899 424 6955
rect 480 6899 548 6955
rect 604 6899 672 6955
rect 728 6899 768 6955
rect 260 6831 768 6899
rect 260 6775 300 6831
rect 356 6775 424 6831
rect 480 6775 548 6831
rect 604 6775 672 6831
rect 728 6775 768 6831
rect 260 6707 768 6775
rect 260 6651 300 6707
rect 356 6651 424 6707
rect 480 6651 548 6707
rect 604 6651 672 6707
rect 728 6651 768 6707
rect 260 6583 768 6651
rect 260 6527 300 6583
rect 356 6527 424 6583
rect 480 6527 548 6583
rect 604 6527 672 6583
rect 728 6527 768 6583
rect 260 6459 768 6527
rect 260 6403 300 6459
rect 356 6403 424 6459
rect 480 6403 548 6459
rect 604 6403 672 6459
rect 728 6403 768 6459
rect 260 6335 768 6403
rect 260 6279 300 6335
rect 356 6279 424 6335
rect 480 6279 548 6335
rect 604 6279 672 6335
rect 728 6279 768 6335
rect 260 6211 768 6279
rect 260 6155 300 6211
rect 356 6155 424 6211
rect 480 6155 548 6211
rect 604 6155 672 6211
rect 728 6155 768 6211
rect 260 6087 768 6155
rect 260 6031 300 6087
rect 356 6031 424 6087
rect 480 6031 548 6087
rect 604 6031 672 6087
rect 728 6031 768 6087
rect 260 5963 768 6031
rect 260 5907 300 5963
rect 356 5907 424 5963
rect 480 5907 548 5963
rect 604 5907 672 5963
rect 728 5907 768 5963
rect 260 5839 768 5907
rect 260 5783 300 5839
rect 356 5783 424 5839
rect 480 5783 548 5839
rect 604 5783 672 5839
rect 728 5783 768 5839
rect 260 5715 768 5783
rect 260 5659 300 5715
rect 356 5659 424 5715
rect 480 5659 548 5715
rect 604 5659 672 5715
rect 728 5659 768 5715
rect 260 5591 768 5659
rect 260 5535 300 5591
rect 356 5535 424 5591
rect 480 5535 548 5591
rect 604 5535 672 5591
rect 728 5535 768 5591
rect 260 5467 768 5535
rect 260 5411 300 5467
rect 356 5411 424 5467
rect 480 5411 548 5467
rect 604 5411 672 5467
rect 728 5411 768 5467
rect 260 5343 768 5411
rect 260 5287 300 5343
rect 356 5287 424 5343
rect 480 5287 548 5343
rect 604 5287 672 5343
rect 728 5287 768 5343
rect 260 5219 768 5287
rect 260 5163 300 5219
rect 356 5163 424 5219
rect 480 5163 548 5219
rect 604 5163 672 5219
rect 728 5163 768 5219
rect 260 5095 768 5163
rect 260 5039 300 5095
rect 356 5039 424 5095
rect 480 5039 548 5095
rect 604 5039 672 5095
rect 728 5039 768 5095
rect 260 4971 768 5039
rect 260 4915 300 4971
rect 356 4915 424 4971
rect 480 4915 548 4971
rect 604 4915 672 4971
rect 728 4915 768 4971
rect 260 4847 768 4915
rect 260 4791 300 4847
rect 356 4791 424 4847
rect 480 4791 548 4847
rect 604 4791 672 4847
rect 728 4791 768 4847
rect 260 4723 768 4791
rect 260 4667 300 4723
rect 356 4667 424 4723
rect 480 4667 548 4723
rect 604 4667 672 4723
rect 728 4667 768 4723
rect 260 4599 768 4667
rect 260 4543 300 4599
rect 356 4543 424 4599
rect 480 4543 548 4599
rect 604 4543 672 4599
rect 728 4543 768 4599
rect 260 4251 768 4543
rect 260 4195 300 4251
rect 356 4195 424 4251
rect 480 4195 548 4251
rect 604 4195 672 4251
rect 728 4195 768 4251
rect 260 4127 768 4195
rect 260 4071 300 4127
rect 356 4071 424 4127
rect 480 4071 548 4127
rect 604 4071 672 4127
rect 728 4071 768 4127
rect 260 4003 768 4071
rect 260 3947 300 4003
rect 356 3947 424 4003
rect 480 3947 548 4003
rect 604 3947 672 4003
rect 728 3947 768 4003
rect 260 3879 768 3947
rect 260 3823 300 3879
rect 356 3823 424 3879
rect 480 3823 548 3879
rect 604 3823 672 3879
rect 728 3823 768 3879
rect 260 3755 768 3823
rect 260 3699 300 3755
rect 356 3699 424 3755
rect 480 3699 548 3755
rect 604 3699 672 3755
rect 728 3699 768 3755
rect 260 3631 768 3699
rect 260 3575 300 3631
rect 356 3575 424 3631
rect 480 3575 548 3631
rect 604 3575 672 3631
rect 728 3575 768 3631
rect 260 3507 768 3575
rect 260 3451 300 3507
rect 356 3451 424 3507
rect 480 3451 548 3507
rect 604 3451 672 3507
rect 728 3451 768 3507
rect 260 3383 768 3451
rect 260 3327 300 3383
rect 356 3327 424 3383
rect 480 3327 548 3383
rect 604 3327 672 3383
rect 728 3327 768 3383
rect 260 3259 768 3327
rect 260 3203 300 3259
rect 356 3203 424 3259
rect 480 3203 548 3259
rect 604 3203 672 3259
rect 728 3203 768 3259
rect 260 3135 768 3203
rect 260 3079 300 3135
rect 356 3079 424 3135
rect 480 3079 548 3135
rect 604 3079 672 3135
rect 728 3079 768 3135
rect 260 3011 768 3079
rect 260 2955 300 3011
rect 356 2955 424 3011
rect 480 2955 548 3011
rect 604 2955 672 3011
rect 728 2955 768 3011
rect 260 2887 768 2955
rect 260 2831 300 2887
rect 356 2831 424 2887
rect 480 2831 548 2887
rect 604 2831 672 2887
rect 728 2831 768 2887
rect 260 2763 768 2831
rect 260 2707 300 2763
rect 356 2707 424 2763
rect 480 2707 548 2763
rect 604 2707 672 2763
rect 728 2707 768 2763
rect 260 2639 768 2707
rect 260 2583 300 2639
rect 356 2583 424 2639
rect 480 2583 548 2639
rect 604 2583 672 2639
rect 728 2583 768 2639
rect 260 2515 768 2583
rect 260 2459 300 2515
rect 356 2459 424 2515
rect 480 2459 548 2515
rect 604 2459 672 2515
rect 728 2459 768 2515
rect 260 2391 768 2459
rect 260 2335 300 2391
rect 356 2335 424 2391
rect 480 2335 548 2391
rect 604 2335 672 2391
rect 728 2335 768 2391
rect 260 2267 768 2335
rect 260 2211 300 2267
rect 356 2211 424 2267
rect 480 2211 548 2267
rect 604 2211 672 2267
rect 728 2211 768 2267
rect 260 2143 768 2211
rect 260 2087 300 2143
rect 356 2087 424 2143
rect 480 2087 548 2143
rect 604 2087 672 2143
rect 728 2087 768 2143
rect 260 2019 768 2087
rect 260 1963 300 2019
rect 356 1963 424 2019
rect 480 1963 548 2019
rect 604 1963 672 2019
rect 728 1963 768 2019
rect 260 1895 768 1963
rect 260 1839 300 1895
rect 356 1839 424 1895
rect 480 1839 548 1895
rect 604 1839 672 1895
rect 728 1839 768 1895
rect 260 1771 768 1839
rect 260 1715 300 1771
rect 356 1715 424 1771
rect 480 1715 548 1771
rect 604 1715 672 1771
rect 728 1715 768 1771
rect 260 1647 768 1715
rect 260 1591 300 1647
rect 356 1591 424 1647
rect 480 1591 548 1647
rect 604 1591 672 1647
rect 728 1591 768 1647
rect 260 1523 768 1591
rect 260 1467 300 1523
rect 356 1467 424 1523
rect 480 1467 548 1523
rect 604 1467 672 1523
rect 728 1467 768 1523
rect 260 1399 768 1467
rect 260 1343 300 1399
rect 356 1343 424 1399
rect 480 1343 548 1399
rect 604 1343 672 1399
rect 728 1343 768 1399
rect 260 900 768 1343
rect 1136 900 1336 10939
rect 1426 10651 1874 10661
rect 1426 10595 1436 10651
rect 1492 10595 1560 10651
rect 1616 10595 1684 10651
rect 1740 10595 1808 10651
rect 1864 10595 1874 10651
rect 1426 10527 1874 10595
rect 1426 10471 1436 10527
rect 1492 10471 1560 10527
rect 1616 10471 1684 10527
rect 1740 10471 1808 10527
rect 1864 10471 1874 10527
rect 1426 10403 1874 10471
rect 1426 10347 1436 10403
rect 1492 10347 1560 10403
rect 1616 10347 1684 10403
rect 1740 10347 1808 10403
rect 1864 10347 1874 10403
rect 1426 10279 1874 10347
rect 1426 10223 1436 10279
rect 1492 10223 1560 10279
rect 1616 10223 1684 10279
rect 1740 10223 1808 10279
rect 1864 10223 1874 10279
rect 1426 10155 1874 10223
rect 1426 10099 1436 10155
rect 1492 10099 1560 10155
rect 1616 10099 1684 10155
rect 1740 10099 1808 10155
rect 1864 10099 1874 10155
rect 1426 10031 1874 10099
rect 1426 9975 1436 10031
rect 1492 9975 1560 10031
rect 1616 9975 1684 10031
rect 1740 9975 1808 10031
rect 1864 9975 1874 10031
rect 1426 9907 1874 9975
rect 1426 9851 1436 9907
rect 1492 9851 1560 9907
rect 1616 9851 1684 9907
rect 1740 9851 1808 9907
rect 1864 9851 1874 9907
rect 1426 9783 1874 9851
rect 1426 9727 1436 9783
rect 1492 9727 1560 9783
rect 1616 9727 1684 9783
rect 1740 9727 1808 9783
rect 1864 9727 1874 9783
rect 1426 9659 1874 9727
rect 1426 9603 1436 9659
rect 1492 9603 1560 9659
rect 1616 9603 1684 9659
rect 1740 9603 1808 9659
rect 1864 9603 1874 9659
rect 1426 9535 1874 9603
rect 1426 9479 1436 9535
rect 1492 9479 1560 9535
rect 1616 9479 1684 9535
rect 1740 9479 1808 9535
rect 1864 9479 1874 9535
rect 1426 9411 1874 9479
rect 1426 9355 1436 9411
rect 1492 9355 1560 9411
rect 1616 9355 1684 9411
rect 1740 9355 1808 9411
rect 1864 9355 1874 9411
rect 1426 9287 1874 9355
rect 1426 9231 1436 9287
rect 1492 9231 1560 9287
rect 1616 9231 1684 9287
rect 1740 9231 1808 9287
rect 1864 9231 1874 9287
rect 1426 9163 1874 9231
rect 1426 9107 1436 9163
rect 1492 9107 1560 9163
rect 1616 9107 1684 9163
rect 1740 9107 1808 9163
rect 1864 9107 1874 9163
rect 1426 9039 1874 9107
rect 1426 8983 1436 9039
rect 1492 8983 1560 9039
rect 1616 8983 1684 9039
rect 1740 8983 1808 9039
rect 1864 8983 1874 9039
rect 1426 8915 1874 8983
rect 1426 8859 1436 8915
rect 1492 8859 1560 8915
rect 1616 8859 1684 8915
rect 1740 8859 1808 8915
rect 1864 8859 1874 8915
rect 1426 8791 1874 8859
rect 1426 8735 1436 8791
rect 1492 8735 1560 8791
rect 1616 8735 1684 8791
rect 1740 8735 1808 8791
rect 1864 8735 1874 8791
rect 1426 8667 1874 8735
rect 1426 8611 1436 8667
rect 1492 8611 1560 8667
rect 1616 8611 1684 8667
rect 1740 8611 1808 8667
rect 1864 8611 1874 8667
rect 1426 8543 1874 8611
rect 1426 8487 1436 8543
rect 1492 8487 1560 8543
rect 1616 8487 1684 8543
rect 1740 8487 1808 8543
rect 1864 8487 1874 8543
rect 1426 8419 1874 8487
rect 1426 8363 1436 8419
rect 1492 8363 1560 8419
rect 1616 8363 1684 8419
rect 1740 8363 1808 8419
rect 1864 8363 1874 8419
rect 1426 8295 1874 8363
rect 1426 8239 1436 8295
rect 1492 8239 1560 8295
rect 1616 8239 1684 8295
rect 1740 8239 1808 8295
rect 1864 8239 1874 8295
rect 1426 8171 1874 8239
rect 1426 8115 1436 8171
rect 1492 8115 1560 8171
rect 1616 8115 1684 8171
rect 1740 8115 1808 8171
rect 1864 8115 1874 8171
rect 1426 8047 1874 8115
rect 1426 7991 1436 8047
rect 1492 7991 1560 8047
rect 1616 7991 1684 8047
rect 1740 7991 1808 8047
rect 1864 7991 1874 8047
rect 1426 7923 1874 7991
rect 1426 7867 1436 7923
rect 1492 7867 1560 7923
rect 1616 7867 1684 7923
rect 1740 7867 1808 7923
rect 1864 7867 1874 7923
rect 1426 7799 1874 7867
rect 1426 7743 1436 7799
rect 1492 7743 1560 7799
rect 1616 7743 1684 7799
rect 1740 7743 1808 7799
rect 1864 7743 1874 7799
rect 1426 7733 1874 7743
rect 2562 10651 3010 10661
rect 2562 10595 2572 10651
rect 2628 10595 2696 10651
rect 2752 10595 2820 10651
rect 2876 10595 2944 10651
rect 3000 10595 3010 10651
rect 2562 10527 3010 10595
rect 2562 10471 2572 10527
rect 2628 10471 2696 10527
rect 2752 10471 2820 10527
rect 2876 10471 2944 10527
rect 3000 10471 3010 10527
rect 2562 10403 3010 10471
rect 2562 10347 2572 10403
rect 2628 10347 2696 10403
rect 2752 10347 2820 10403
rect 2876 10347 2944 10403
rect 3000 10347 3010 10403
rect 2562 10279 3010 10347
rect 2562 10223 2572 10279
rect 2628 10223 2696 10279
rect 2752 10223 2820 10279
rect 2876 10223 2944 10279
rect 3000 10223 3010 10279
rect 2562 10155 3010 10223
rect 2562 10099 2572 10155
rect 2628 10099 2696 10155
rect 2752 10099 2820 10155
rect 2876 10099 2944 10155
rect 3000 10099 3010 10155
rect 2562 10031 3010 10099
rect 2562 9975 2572 10031
rect 2628 9975 2696 10031
rect 2752 9975 2820 10031
rect 2876 9975 2944 10031
rect 3000 9975 3010 10031
rect 2562 9907 3010 9975
rect 2562 9851 2572 9907
rect 2628 9851 2696 9907
rect 2752 9851 2820 9907
rect 2876 9851 2944 9907
rect 3000 9851 3010 9907
rect 2562 9783 3010 9851
rect 2562 9727 2572 9783
rect 2628 9727 2696 9783
rect 2752 9727 2820 9783
rect 2876 9727 2944 9783
rect 3000 9727 3010 9783
rect 2562 9659 3010 9727
rect 2562 9603 2572 9659
rect 2628 9603 2696 9659
rect 2752 9603 2820 9659
rect 2876 9603 2944 9659
rect 3000 9603 3010 9659
rect 2562 9535 3010 9603
rect 2562 9479 2572 9535
rect 2628 9479 2696 9535
rect 2752 9479 2820 9535
rect 2876 9479 2944 9535
rect 3000 9479 3010 9535
rect 2562 9411 3010 9479
rect 2562 9355 2572 9411
rect 2628 9355 2696 9411
rect 2752 9355 2820 9411
rect 2876 9355 2944 9411
rect 3000 9355 3010 9411
rect 2562 9287 3010 9355
rect 2562 9231 2572 9287
rect 2628 9231 2696 9287
rect 2752 9231 2820 9287
rect 2876 9231 2944 9287
rect 3000 9231 3010 9287
rect 2562 9163 3010 9231
rect 2562 9107 2572 9163
rect 2628 9107 2696 9163
rect 2752 9107 2820 9163
rect 2876 9107 2944 9163
rect 3000 9107 3010 9163
rect 2562 9039 3010 9107
rect 2562 8983 2572 9039
rect 2628 8983 2696 9039
rect 2752 8983 2820 9039
rect 2876 8983 2944 9039
rect 3000 8983 3010 9039
rect 2562 8915 3010 8983
rect 2562 8859 2572 8915
rect 2628 8859 2696 8915
rect 2752 8859 2820 8915
rect 2876 8859 2944 8915
rect 3000 8859 3010 8915
rect 2562 8791 3010 8859
rect 2562 8735 2572 8791
rect 2628 8735 2696 8791
rect 2752 8735 2820 8791
rect 2876 8735 2944 8791
rect 3000 8735 3010 8791
rect 2562 8667 3010 8735
rect 2562 8611 2572 8667
rect 2628 8611 2696 8667
rect 2752 8611 2820 8667
rect 2876 8611 2944 8667
rect 3000 8611 3010 8667
rect 2562 8543 3010 8611
rect 2562 8487 2572 8543
rect 2628 8487 2696 8543
rect 2752 8487 2820 8543
rect 2876 8487 2944 8543
rect 3000 8487 3010 8543
rect 2562 8419 3010 8487
rect 2562 8363 2572 8419
rect 2628 8363 2696 8419
rect 2752 8363 2820 8419
rect 2876 8363 2944 8419
rect 3000 8363 3010 8419
rect 2562 8295 3010 8363
rect 2562 8239 2572 8295
rect 2628 8239 2696 8295
rect 2752 8239 2820 8295
rect 2876 8239 2944 8295
rect 3000 8239 3010 8295
rect 2562 8171 3010 8239
rect 2562 8115 2572 8171
rect 2628 8115 2696 8171
rect 2752 8115 2820 8171
rect 2876 8115 2944 8171
rect 3000 8115 3010 8171
rect 2562 8047 3010 8115
rect 2562 7991 2572 8047
rect 2628 7991 2696 8047
rect 2752 7991 2820 8047
rect 2876 7991 2944 8047
rect 3000 7991 3010 8047
rect 2562 7923 3010 7991
rect 2562 7867 2572 7923
rect 2628 7867 2696 7923
rect 2752 7867 2820 7923
rect 2876 7867 2944 7923
rect 3000 7867 3010 7923
rect 2562 7799 3010 7867
rect 2562 7743 2572 7799
rect 2628 7743 2696 7799
rect 2752 7743 2820 7799
rect 2876 7743 2944 7799
rect 3000 7743 3010 7799
rect 2562 7733 3010 7743
rect 4834 10651 5282 10661
rect 4834 10595 4844 10651
rect 4900 10595 4968 10651
rect 5024 10595 5092 10651
rect 5148 10595 5216 10651
rect 5272 10595 5282 10651
rect 4834 10527 5282 10595
rect 4834 10471 4844 10527
rect 4900 10471 4968 10527
rect 5024 10471 5092 10527
rect 5148 10471 5216 10527
rect 5272 10471 5282 10527
rect 4834 10403 5282 10471
rect 4834 10347 4844 10403
rect 4900 10347 4968 10403
rect 5024 10347 5092 10403
rect 5148 10347 5216 10403
rect 5272 10347 5282 10403
rect 4834 10279 5282 10347
rect 4834 10223 4844 10279
rect 4900 10223 4968 10279
rect 5024 10223 5092 10279
rect 5148 10223 5216 10279
rect 5272 10223 5282 10279
rect 4834 10155 5282 10223
rect 4834 10099 4844 10155
rect 4900 10099 4968 10155
rect 5024 10099 5092 10155
rect 5148 10099 5216 10155
rect 5272 10099 5282 10155
rect 4834 10031 5282 10099
rect 4834 9975 4844 10031
rect 4900 9975 4968 10031
rect 5024 9975 5092 10031
rect 5148 9975 5216 10031
rect 5272 9975 5282 10031
rect 4834 9907 5282 9975
rect 4834 9851 4844 9907
rect 4900 9851 4968 9907
rect 5024 9851 5092 9907
rect 5148 9851 5216 9907
rect 5272 9851 5282 9907
rect 4834 9783 5282 9851
rect 4834 9727 4844 9783
rect 4900 9727 4968 9783
rect 5024 9727 5092 9783
rect 5148 9727 5216 9783
rect 5272 9727 5282 9783
rect 4834 9659 5282 9727
rect 4834 9603 4844 9659
rect 4900 9603 4968 9659
rect 5024 9603 5092 9659
rect 5148 9603 5216 9659
rect 5272 9603 5282 9659
rect 4834 9535 5282 9603
rect 4834 9479 4844 9535
rect 4900 9479 4968 9535
rect 5024 9479 5092 9535
rect 5148 9479 5216 9535
rect 5272 9479 5282 9535
rect 4834 9411 5282 9479
rect 4834 9355 4844 9411
rect 4900 9355 4968 9411
rect 5024 9355 5092 9411
rect 5148 9355 5216 9411
rect 5272 9355 5282 9411
rect 4834 9287 5282 9355
rect 4834 9231 4844 9287
rect 4900 9231 4968 9287
rect 5024 9231 5092 9287
rect 5148 9231 5216 9287
rect 5272 9231 5282 9287
rect 4834 9163 5282 9231
rect 4834 9107 4844 9163
rect 4900 9107 4968 9163
rect 5024 9107 5092 9163
rect 5148 9107 5216 9163
rect 5272 9107 5282 9163
rect 4834 9039 5282 9107
rect 4834 8983 4844 9039
rect 4900 8983 4968 9039
rect 5024 8983 5092 9039
rect 5148 8983 5216 9039
rect 5272 8983 5282 9039
rect 4834 8915 5282 8983
rect 4834 8859 4844 8915
rect 4900 8859 4968 8915
rect 5024 8859 5092 8915
rect 5148 8859 5216 8915
rect 5272 8859 5282 8915
rect 4834 8791 5282 8859
rect 4834 8735 4844 8791
rect 4900 8735 4968 8791
rect 5024 8735 5092 8791
rect 5148 8735 5216 8791
rect 5272 8735 5282 8791
rect 4834 8667 5282 8735
rect 4834 8611 4844 8667
rect 4900 8611 4968 8667
rect 5024 8611 5092 8667
rect 5148 8611 5216 8667
rect 5272 8611 5282 8667
rect 4834 8543 5282 8611
rect 4834 8487 4844 8543
rect 4900 8487 4968 8543
rect 5024 8487 5092 8543
rect 5148 8487 5216 8543
rect 5272 8487 5282 8543
rect 4834 8419 5282 8487
rect 4834 8363 4844 8419
rect 4900 8363 4968 8419
rect 5024 8363 5092 8419
rect 5148 8363 5216 8419
rect 5272 8363 5282 8419
rect 4834 8295 5282 8363
rect 4834 8239 4844 8295
rect 4900 8239 4968 8295
rect 5024 8239 5092 8295
rect 5148 8239 5216 8295
rect 5272 8239 5282 8295
rect 4834 8171 5282 8239
rect 4834 8115 4844 8171
rect 4900 8115 4968 8171
rect 5024 8115 5092 8171
rect 5148 8115 5216 8171
rect 5272 8115 5282 8171
rect 4834 8047 5282 8115
rect 4834 7991 4844 8047
rect 4900 7991 4968 8047
rect 5024 7991 5092 8047
rect 5148 7991 5216 8047
rect 5272 7991 5282 8047
rect 4834 7923 5282 7991
rect 4834 7867 4844 7923
rect 4900 7867 4968 7923
rect 5024 7867 5092 7923
rect 5148 7867 5216 7923
rect 5272 7867 5282 7923
rect 4834 7799 5282 7867
rect 4834 7743 4844 7799
rect 4900 7743 4968 7799
rect 5024 7743 5092 7799
rect 5148 7743 5216 7799
rect 5272 7743 5282 7799
rect 4834 7733 5282 7743
rect 7127 10651 7451 10661
rect 7127 10595 7137 10651
rect 7193 10595 7261 10651
rect 7317 10595 7385 10651
rect 7441 10595 7451 10651
rect 7127 10527 7451 10595
rect 7127 10471 7137 10527
rect 7193 10471 7261 10527
rect 7317 10471 7385 10527
rect 7441 10471 7451 10527
rect 7127 10403 7451 10471
rect 7127 10347 7137 10403
rect 7193 10347 7261 10403
rect 7317 10347 7385 10403
rect 7441 10347 7451 10403
rect 7127 10279 7451 10347
rect 7127 10223 7137 10279
rect 7193 10223 7261 10279
rect 7317 10223 7385 10279
rect 7441 10223 7451 10279
rect 7127 10155 7451 10223
rect 7127 10099 7137 10155
rect 7193 10099 7261 10155
rect 7317 10099 7385 10155
rect 7441 10099 7451 10155
rect 7127 10031 7451 10099
rect 7127 9975 7137 10031
rect 7193 9975 7261 10031
rect 7317 9975 7385 10031
rect 7441 9975 7451 10031
rect 7127 9907 7451 9975
rect 7127 9851 7137 9907
rect 7193 9851 7261 9907
rect 7317 9851 7385 9907
rect 7441 9851 7451 9907
rect 7127 9783 7451 9851
rect 7127 9727 7137 9783
rect 7193 9727 7261 9783
rect 7317 9727 7385 9783
rect 7441 9727 7451 9783
rect 7127 9659 7451 9727
rect 7127 9603 7137 9659
rect 7193 9603 7261 9659
rect 7317 9603 7385 9659
rect 7441 9603 7451 9659
rect 7127 9535 7451 9603
rect 7127 9479 7137 9535
rect 7193 9479 7261 9535
rect 7317 9479 7385 9535
rect 7441 9479 7451 9535
rect 7127 9411 7451 9479
rect 7127 9355 7137 9411
rect 7193 9355 7261 9411
rect 7317 9355 7385 9411
rect 7441 9355 7451 9411
rect 7127 9287 7451 9355
rect 7127 9231 7137 9287
rect 7193 9231 7261 9287
rect 7317 9231 7385 9287
rect 7441 9231 7451 9287
rect 7127 9163 7451 9231
rect 7127 9107 7137 9163
rect 7193 9107 7261 9163
rect 7317 9107 7385 9163
rect 7441 9107 7451 9163
rect 7127 9039 7451 9107
rect 7127 8983 7137 9039
rect 7193 8983 7261 9039
rect 7317 8983 7385 9039
rect 7441 8983 7451 9039
rect 7127 8915 7451 8983
rect 7127 8859 7137 8915
rect 7193 8859 7261 8915
rect 7317 8859 7385 8915
rect 7441 8859 7451 8915
rect 7127 8791 7451 8859
rect 7127 8735 7137 8791
rect 7193 8735 7261 8791
rect 7317 8735 7385 8791
rect 7441 8735 7451 8791
rect 7127 8667 7451 8735
rect 7127 8611 7137 8667
rect 7193 8611 7261 8667
rect 7317 8611 7385 8667
rect 7441 8611 7451 8667
rect 7127 8543 7451 8611
rect 7127 8487 7137 8543
rect 7193 8487 7261 8543
rect 7317 8487 7385 8543
rect 7441 8487 7451 8543
rect 7127 8419 7451 8487
rect 7127 8363 7137 8419
rect 7193 8363 7261 8419
rect 7317 8363 7385 8419
rect 7441 8363 7451 8419
rect 7127 8295 7451 8363
rect 7127 8239 7137 8295
rect 7193 8239 7261 8295
rect 7317 8239 7385 8295
rect 7441 8239 7451 8295
rect 7127 8171 7451 8239
rect 7127 8115 7137 8171
rect 7193 8115 7261 8171
rect 7317 8115 7385 8171
rect 7441 8115 7451 8171
rect 7127 8047 7451 8115
rect 7127 7991 7137 8047
rect 7193 7991 7261 8047
rect 7317 7991 7385 8047
rect 7441 7991 7451 8047
rect 7127 7923 7451 7991
rect 7127 7867 7137 7923
rect 7193 7867 7261 7923
rect 7317 7867 7385 7923
rect 7441 7867 7451 7923
rect 7127 7799 7451 7867
rect 7127 7743 7137 7799
rect 7193 7743 7261 7799
rect 7317 7743 7385 7799
rect 7441 7743 7451 7799
rect 7127 7733 7451 7743
rect 7613 10651 7937 10661
rect 7613 10595 7623 10651
rect 7679 10595 7747 10651
rect 7803 10595 7871 10651
rect 7927 10595 7937 10651
rect 7613 10527 7937 10595
rect 7613 10471 7623 10527
rect 7679 10471 7747 10527
rect 7803 10471 7871 10527
rect 7927 10471 7937 10527
rect 7613 10403 7937 10471
rect 7613 10347 7623 10403
rect 7679 10347 7747 10403
rect 7803 10347 7871 10403
rect 7927 10347 7937 10403
rect 7613 10279 7937 10347
rect 7613 10223 7623 10279
rect 7679 10223 7747 10279
rect 7803 10223 7871 10279
rect 7927 10223 7937 10279
rect 7613 10155 7937 10223
rect 7613 10099 7623 10155
rect 7679 10099 7747 10155
rect 7803 10099 7871 10155
rect 7927 10099 7937 10155
rect 7613 10031 7937 10099
rect 7613 9975 7623 10031
rect 7679 9975 7747 10031
rect 7803 9975 7871 10031
rect 7927 9975 7937 10031
rect 7613 9907 7937 9975
rect 7613 9851 7623 9907
rect 7679 9851 7747 9907
rect 7803 9851 7871 9907
rect 7927 9851 7937 9907
rect 7613 9783 7937 9851
rect 7613 9727 7623 9783
rect 7679 9727 7747 9783
rect 7803 9727 7871 9783
rect 7927 9727 7937 9783
rect 7613 9659 7937 9727
rect 7613 9603 7623 9659
rect 7679 9603 7747 9659
rect 7803 9603 7871 9659
rect 7927 9603 7937 9659
rect 7613 9535 7937 9603
rect 7613 9479 7623 9535
rect 7679 9479 7747 9535
rect 7803 9479 7871 9535
rect 7927 9479 7937 9535
rect 7613 9411 7937 9479
rect 7613 9355 7623 9411
rect 7679 9355 7747 9411
rect 7803 9355 7871 9411
rect 7927 9355 7937 9411
rect 7613 9287 7937 9355
rect 7613 9231 7623 9287
rect 7679 9231 7747 9287
rect 7803 9231 7871 9287
rect 7927 9231 7937 9287
rect 7613 9163 7937 9231
rect 7613 9107 7623 9163
rect 7679 9107 7747 9163
rect 7803 9107 7871 9163
rect 7927 9107 7937 9163
rect 7613 9039 7937 9107
rect 7613 8983 7623 9039
rect 7679 8983 7747 9039
rect 7803 8983 7871 9039
rect 7927 8983 7937 9039
rect 7613 8915 7937 8983
rect 7613 8859 7623 8915
rect 7679 8859 7747 8915
rect 7803 8859 7871 8915
rect 7927 8859 7937 8915
rect 7613 8791 7937 8859
rect 7613 8735 7623 8791
rect 7679 8735 7747 8791
rect 7803 8735 7871 8791
rect 7927 8735 7937 8791
rect 7613 8667 7937 8735
rect 7613 8611 7623 8667
rect 7679 8611 7747 8667
rect 7803 8611 7871 8667
rect 7927 8611 7937 8667
rect 7613 8543 7937 8611
rect 7613 8487 7623 8543
rect 7679 8487 7747 8543
rect 7803 8487 7871 8543
rect 7927 8487 7937 8543
rect 7613 8419 7937 8487
rect 7613 8363 7623 8419
rect 7679 8363 7747 8419
rect 7803 8363 7871 8419
rect 7927 8363 7937 8419
rect 7613 8295 7937 8363
rect 7613 8239 7623 8295
rect 7679 8239 7747 8295
rect 7803 8239 7871 8295
rect 7927 8239 7937 8295
rect 7613 8171 7937 8239
rect 7613 8115 7623 8171
rect 7679 8115 7747 8171
rect 7803 8115 7871 8171
rect 7927 8115 7937 8171
rect 7613 8047 7937 8115
rect 7613 7991 7623 8047
rect 7679 7991 7747 8047
rect 7803 7991 7871 8047
rect 7927 7991 7937 8047
rect 7613 7923 7937 7991
rect 7613 7867 7623 7923
rect 7679 7867 7747 7923
rect 7803 7867 7871 7923
rect 7927 7867 7937 7923
rect 7613 7799 7937 7867
rect 7613 7743 7623 7799
rect 7679 7743 7747 7799
rect 7803 7743 7871 7799
rect 7927 7743 7937 7799
rect 7613 7733 7937 7743
rect 9782 10651 10230 10661
rect 9782 10595 9792 10651
rect 9848 10595 9916 10651
rect 9972 10595 10040 10651
rect 10096 10595 10164 10651
rect 10220 10595 10230 10651
rect 9782 10527 10230 10595
rect 9782 10471 9792 10527
rect 9848 10471 9916 10527
rect 9972 10471 10040 10527
rect 10096 10471 10164 10527
rect 10220 10471 10230 10527
rect 9782 10403 10230 10471
rect 9782 10347 9792 10403
rect 9848 10347 9916 10403
rect 9972 10347 10040 10403
rect 10096 10347 10164 10403
rect 10220 10347 10230 10403
rect 9782 10279 10230 10347
rect 9782 10223 9792 10279
rect 9848 10223 9916 10279
rect 9972 10223 10040 10279
rect 10096 10223 10164 10279
rect 10220 10223 10230 10279
rect 9782 10155 10230 10223
rect 9782 10099 9792 10155
rect 9848 10099 9916 10155
rect 9972 10099 10040 10155
rect 10096 10099 10164 10155
rect 10220 10099 10230 10155
rect 9782 10031 10230 10099
rect 9782 9975 9792 10031
rect 9848 9975 9916 10031
rect 9972 9975 10040 10031
rect 10096 9975 10164 10031
rect 10220 9975 10230 10031
rect 9782 9907 10230 9975
rect 9782 9851 9792 9907
rect 9848 9851 9916 9907
rect 9972 9851 10040 9907
rect 10096 9851 10164 9907
rect 10220 9851 10230 9907
rect 9782 9783 10230 9851
rect 9782 9727 9792 9783
rect 9848 9727 9916 9783
rect 9972 9727 10040 9783
rect 10096 9727 10164 9783
rect 10220 9727 10230 9783
rect 9782 9659 10230 9727
rect 9782 9603 9792 9659
rect 9848 9603 9916 9659
rect 9972 9603 10040 9659
rect 10096 9603 10164 9659
rect 10220 9603 10230 9659
rect 9782 9535 10230 9603
rect 9782 9479 9792 9535
rect 9848 9479 9916 9535
rect 9972 9479 10040 9535
rect 10096 9479 10164 9535
rect 10220 9479 10230 9535
rect 9782 9411 10230 9479
rect 9782 9355 9792 9411
rect 9848 9355 9916 9411
rect 9972 9355 10040 9411
rect 10096 9355 10164 9411
rect 10220 9355 10230 9411
rect 9782 9287 10230 9355
rect 9782 9231 9792 9287
rect 9848 9231 9916 9287
rect 9972 9231 10040 9287
rect 10096 9231 10164 9287
rect 10220 9231 10230 9287
rect 9782 9163 10230 9231
rect 9782 9107 9792 9163
rect 9848 9107 9916 9163
rect 9972 9107 10040 9163
rect 10096 9107 10164 9163
rect 10220 9107 10230 9163
rect 9782 9039 10230 9107
rect 9782 8983 9792 9039
rect 9848 8983 9916 9039
rect 9972 8983 10040 9039
rect 10096 8983 10164 9039
rect 10220 8983 10230 9039
rect 9782 8915 10230 8983
rect 9782 8859 9792 8915
rect 9848 8859 9916 8915
rect 9972 8859 10040 8915
rect 10096 8859 10164 8915
rect 10220 8859 10230 8915
rect 9782 8791 10230 8859
rect 9782 8735 9792 8791
rect 9848 8735 9916 8791
rect 9972 8735 10040 8791
rect 10096 8735 10164 8791
rect 10220 8735 10230 8791
rect 9782 8667 10230 8735
rect 9782 8611 9792 8667
rect 9848 8611 9916 8667
rect 9972 8611 10040 8667
rect 10096 8611 10164 8667
rect 10220 8611 10230 8667
rect 9782 8543 10230 8611
rect 9782 8487 9792 8543
rect 9848 8487 9916 8543
rect 9972 8487 10040 8543
rect 10096 8487 10164 8543
rect 10220 8487 10230 8543
rect 9782 8419 10230 8487
rect 9782 8363 9792 8419
rect 9848 8363 9916 8419
rect 9972 8363 10040 8419
rect 10096 8363 10164 8419
rect 10220 8363 10230 8419
rect 9782 8295 10230 8363
rect 9782 8239 9792 8295
rect 9848 8239 9916 8295
rect 9972 8239 10040 8295
rect 10096 8239 10164 8295
rect 10220 8239 10230 8295
rect 9782 8171 10230 8239
rect 9782 8115 9792 8171
rect 9848 8115 9916 8171
rect 9972 8115 10040 8171
rect 10096 8115 10164 8171
rect 10220 8115 10230 8171
rect 9782 8047 10230 8115
rect 9782 7991 9792 8047
rect 9848 7991 9916 8047
rect 9972 7991 10040 8047
rect 10096 7991 10164 8047
rect 10220 7991 10230 8047
rect 9782 7923 10230 7991
rect 9782 7867 9792 7923
rect 9848 7867 9916 7923
rect 9972 7867 10040 7923
rect 10096 7867 10164 7923
rect 10220 7867 10230 7923
rect 9782 7799 10230 7867
rect 9782 7743 9792 7799
rect 9848 7743 9916 7799
rect 9972 7743 10040 7799
rect 10096 7743 10164 7799
rect 10220 7743 10230 7799
rect 9782 7733 10230 7743
rect 12054 10651 12502 10661
rect 12054 10595 12064 10651
rect 12120 10595 12188 10651
rect 12244 10595 12312 10651
rect 12368 10595 12436 10651
rect 12492 10595 12502 10651
rect 12054 10527 12502 10595
rect 12054 10471 12064 10527
rect 12120 10471 12188 10527
rect 12244 10471 12312 10527
rect 12368 10471 12436 10527
rect 12492 10471 12502 10527
rect 12054 10403 12502 10471
rect 12054 10347 12064 10403
rect 12120 10347 12188 10403
rect 12244 10347 12312 10403
rect 12368 10347 12436 10403
rect 12492 10347 12502 10403
rect 12054 10279 12502 10347
rect 12054 10223 12064 10279
rect 12120 10223 12188 10279
rect 12244 10223 12312 10279
rect 12368 10223 12436 10279
rect 12492 10223 12502 10279
rect 12054 10155 12502 10223
rect 12054 10099 12064 10155
rect 12120 10099 12188 10155
rect 12244 10099 12312 10155
rect 12368 10099 12436 10155
rect 12492 10099 12502 10155
rect 12054 10031 12502 10099
rect 12054 9975 12064 10031
rect 12120 9975 12188 10031
rect 12244 9975 12312 10031
rect 12368 9975 12436 10031
rect 12492 9975 12502 10031
rect 12054 9907 12502 9975
rect 12054 9851 12064 9907
rect 12120 9851 12188 9907
rect 12244 9851 12312 9907
rect 12368 9851 12436 9907
rect 12492 9851 12502 9907
rect 12054 9783 12502 9851
rect 12054 9727 12064 9783
rect 12120 9727 12188 9783
rect 12244 9727 12312 9783
rect 12368 9727 12436 9783
rect 12492 9727 12502 9783
rect 12054 9659 12502 9727
rect 12054 9603 12064 9659
rect 12120 9603 12188 9659
rect 12244 9603 12312 9659
rect 12368 9603 12436 9659
rect 12492 9603 12502 9659
rect 12054 9535 12502 9603
rect 12054 9479 12064 9535
rect 12120 9479 12188 9535
rect 12244 9479 12312 9535
rect 12368 9479 12436 9535
rect 12492 9479 12502 9535
rect 12054 9411 12502 9479
rect 12054 9355 12064 9411
rect 12120 9355 12188 9411
rect 12244 9355 12312 9411
rect 12368 9355 12436 9411
rect 12492 9355 12502 9411
rect 12054 9287 12502 9355
rect 12054 9231 12064 9287
rect 12120 9231 12188 9287
rect 12244 9231 12312 9287
rect 12368 9231 12436 9287
rect 12492 9231 12502 9287
rect 12054 9163 12502 9231
rect 12054 9107 12064 9163
rect 12120 9107 12188 9163
rect 12244 9107 12312 9163
rect 12368 9107 12436 9163
rect 12492 9107 12502 9163
rect 12054 9039 12502 9107
rect 12054 8983 12064 9039
rect 12120 8983 12188 9039
rect 12244 8983 12312 9039
rect 12368 8983 12436 9039
rect 12492 8983 12502 9039
rect 12054 8915 12502 8983
rect 12054 8859 12064 8915
rect 12120 8859 12188 8915
rect 12244 8859 12312 8915
rect 12368 8859 12436 8915
rect 12492 8859 12502 8915
rect 12054 8791 12502 8859
rect 12054 8735 12064 8791
rect 12120 8735 12188 8791
rect 12244 8735 12312 8791
rect 12368 8735 12436 8791
rect 12492 8735 12502 8791
rect 12054 8667 12502 8735
rect 12054 8611 12064 8667
rect 12120 8611 12188 8667
rect 12244 8611 12312 8667
rect 12368 8611 12436 8667
rect 12492 8611 12502 8667
rect 12054 8543 12502 8611
rect 12054 8487 12064 8543
rect 12120 8487 12188 8543
rect 12244 8487 12312 8543
rect 12368 8487 12436 8543
rect 12492 8487 12502 8543
rect 12054 8419 12502 8487
rect 12054 8363 12064 8419
rect 12120 8363 12188 8419
rect 12244 8363 12312 8419
rect 12368 8363 12436 8419
rect 12492 8363 12502 8419
rect 12054 8295 12502 8363
rect 12054 8239 12064 8295
rect 12120 8239 12188 8295
rect 12244 8239 12312 8295
rect 12368 8239 12436 8295
rect 12492 8239 12502 8295
rect 12054 8171 12502 8239
rect 12054 8115 12064 8171
rect 12120 8115 12188 8171
rect 12244 8115 12312 8171
rect 12368 8115 12436 8171
rect 12492 8115 12502 8171
rect 12054 8047 12502 8115
rect 12054 7991 12064 8047
rect 12120 7991 12188 8047
rect 12244 7991 12312 8047
rect 12368 7991 12436 8047
rect 12492 7991 12502 8047
rect 12054 7923 12502 7991
rect 12054 7867 12064 7923
rect 12120 7867 12188 7923
rect 12244 7867 12312 7923
rect 12368 7867 12436 7923
rect 12492 7867 12502 7923
rect 12054 7799 12502 7867
rect 12054 7743 12064 7799
rect 12120 7743 12188 7799
rect 12244 7743 12312 7799
rect 12368 7743 12436 7799
rect 12492 7743 12502 7799
rect 12054 7733 12502 7743
rect 13190 10651 13638 10661
rect 13190 10595 13200 10651
rect 13256 10595 13324 10651
rect 13380 10595 13448 10651
rect 13504 10595 13572 10651
rect 13628 10595 13638 10651
rect 13190 10527 13638 10595
rect 13190 10471 13200 10527
rect 13256 10471 13324 10527
rect 13380 10471 13448 10527
rect 13504 10471 13572 10527
rect 13628 10471 13638 10527
rect 13190 10403 13638 10471
rect 13190 10347 13200 10403
rect 13256 10347 13324 10403
rect 13380 10347 13448 10403
rect 13504 10347 13572 10403
rect 13628 10347 13638 10403
rect 13190 10279 13638 10347
rect 13190 10223 13200 10279
rect 13256 10223 13324 10279
rect 13380 10223 13448 10279
rect 13504 10223 13572 10279
rect 13628 10223 13638 10279
rect 13190 10155 13638 10223
rect 13190 10099 13200 10155
rect 13256 10099 13324 10155
rect 13380 10099 13448 10155
rect 13504 10099 13572 10155
rect 13628 10099 13638 10155
rect 13190 10031 13638 10099
rect 13190 9975 13200 10031
rect 13256 9975 13324 10031
rect 13380 9975 13448 10031
rect 13504 9975 13572 10031
rect 13628 9975 13638 10031
rect 13190 9907 13638 9975
rect 13190 9851 13200 9907
rect 13256 9851 13324 9907
rect 13380 9851 13448 9907
rect 13504 9851 13572 9907
rect 13628 9851 13638 9907
rect 13190 9783 13638 9851
rect 13190 9727 13200 9783
rect 13256 9727 13324 9783
rect 13380 9727 13448 9783
rect 13504 9727 13572 9783
rect 13628 9727 13638 9783
rect 13190 9659 13638 9727
rect 13190 9603 13200 9659
rect 13256 9603 13324 9659
rect 13380 9603 13448 9659
rect 13504 9603 13572 9659
rect 13628 9603 13638 9659
rect 13190 9535 13638 9603
rect 13190 9479 13200 9535
rect 13256 9479 13324 9535
rect 13380 9479 13448 9535
rect 13504 9479 13572 9535
rect 13628 9479 13638 9535
rect 13190 9411 13638 9479
rect 13190 9355 13200 9411
rect 13256 9355 13324 9411
rect 13380 9355 13448 9411
rect 13504 9355 13572 9411
rect 13628 9355 13638 9411
rect 13190 9287 13638 9355
rect 13190 9231 13200 9287
rect 13256 9231 13324 9287
rect 13380 9231 13448 9287
rect 13504 9231 13572 9287
rect 13628 9231 13638 9287
rect 13190 9163 13638 9231
rect 13190 9107 13200 9163
rect 13256 9107 13324 9163
rect 13380 9107 13448 9163
rect 13504 9107 13572 9163
rect 13628 9107 13638 9163
rect 13190 9039 13638 9107
rect 13190 8983 13200 9039
rect 13256 8983 13324 9039
rect 13380 8983 13448 9039
rect 13504 8983 13572 9039
rect 13628 8983 13638 9039
rect 13190 8915 13638 8983
rect 13190 8859 13200 8915
rect 13256 8859 13324 8915
rect 13380 8859 13448 8915
rect 13504 8859 13572 8915
rect 13628 8859 13638 8915
rect 13190 8791 13638 8859
rect 13190 8735 13200 8791
rect 13256 8735 13324 8791
rect 13380 8735 13448 8791
rect 13504 8735 13572 8791
rect 13628 8735 13638 8791
rect 13190 8667 13638 8735
rect 13190 8611 13200 8667
rect 13256 8611 13324 8667
rect 13380 8611 13448 8667
rect 13504 8611 13572 8667
rect 13628 8611 13638 8667
rect 13190 8543 13638 8611
rect 13190 8487 13200 8543
rect 13256 8487 13324 8543
rect 13380 8487 13448 8543
rect 13504 8487 13572 8543
rect 13628 8487 13638 8543
rect 13190 8419 13638 8487
rect 13190 8363 13200 8419
rect 13256 8363 13324 8419
rect 13380 8363 13448 8419
rect 13504 8363 13572 8419
rect 13628 8363 13638 8419
rect 13190 8295 13638 8363
rect 13190 8239 13200 8295
rect 13256 8239 13324 8295
rect 13380 8239 13448 8295
rect 13504 8239 13572 8295
rect 13628 8239 13638 8295
rect 13190 8171 13638 8239
rect 13190 8115 13200 8171
rect 13256 8115 13324 8171
rect 13380 8115 13448 8171
rect 13504 8115 13572 8171
rect 13628 8115 13638 8171
rect 13190 8047 13638 8115
rect 13190 7991 13200 8047
rect 13256 7991 13324 8047
rect 13380 7991 13448 8047
rect 13504 7991 13572 8047
rect 13628 7991 13638 8047
rect 13190 7923 13638 7991
rect 13190 7867 13200 7923
rect 13256 7867 13324 7923
rect 13380 7867 13448 7923
rect 13504 7867 13572 7923
rect 13628 7867 13638 7923
rect 13190 7799 13638 7867
rect 13190 7743 13200 7799
rect 13256 7743 13324 7799
rect 13380 7743 13448 7799
rect 13504 7743 13572 7799
rect 13628 7743 13638 7799
rect 13190 7733 13638 7743
rect 1426 7451 1874 7461
rect 1426 7395 1436 7451
rect 1492 7395 1560 7451
rect 1616 7395 1684 7451
rect 1740 7395 1808 7451
rect 1864 7395 1874 7451
rect 1426 7327 1874 7395
rect 1426 7271 1436 7327
rect 1492 7271 1560 7327
rect 1616 7271 1684 7327
rect 1740 7271 1808 7327
rect 1864 7271 1874 7327
rect 1426 7203 1874 7271
rect 1426 7147 1436 7203
rect 1492 7147 1560 7203
rect 1616 7147 1684 7203
rect 1740 7147 1808 7203
rect 1864 7147 1874 7203
rect 1426 7079 1874 7147
rect 1426 7023 1436 7079
rect 1492 7023 1560 7079
rect 1616 7023 1684 7079
rect 1740 7023 1808 7079
rect 1864 7023 1874 7079
rect 1426 6955 1874 7023
rect 1426 6899 1436 6955
rect 1492 6899 1560 6955
rect 1616 6899 1684 6955
rect 1740 6899 1808 6955
rect 1864 6899 1874 6955
rect 1426 6831 1874 6899
rect 1426 6775 1436 6831
rect 1492 6775 1560 6831
rect 1616 6775 1684 6831
rect 1740 6775 1808 6831
rect 1864 6775 1874 6831
rect 1426 6707 1874 6775
rect 1426 6651 1436 6707
rect 1492 6651 1560 6707
rect 1616 6651 1684 6707
rect 1740 6651 1808 6707
rect 1864 6651 1874 6707
rect 1426 6583 1874 6651
rect 1426 6527 1436 6583
rect 1492 6527 1560 6583
rect 1616 6527 1684 6583
rect 1740 6527 1808 6583
rect 1864 6527 1874 6583
rect 1426 6459 1874 6527
rect 1426 6403 1436 6459
rect 1492 6403 1560 6459
rect 1616 6403 1684 6459
rect 1740 6403 1808 6459
rect 1864 6403 1874 6459
rect 1426 6335 1874 6403
rect 1426 6279 1436 6335
rect 1492 6279 1560 6335
rect 1616 6279 1684 6335
rect 1740 6279 1808 6335
rect 1864 6279 1874 6335
rect 1426 6211 1874 6279
rect 1426 6155 1436 6211
rect 1492 6155 1560 6211
rect 1616 6155 1684 6211
rect 1740 6155 1808 6211
rect 1864 6155 1874 6211
rect 1426 6087 1874 6155
rect 1426 6031 1436 6087
rect 1492 6031 1560 6087
rect 1616 6031 1684 6087
rect 1740 6031 1808 6087
rect 1864 6031 1874 6087
rect 1426 5963 1874 6031
rect 1426 5907 1436 5963
rect 1492 5907 1560 5963
rect 1616 5907 1684 5963
rect 1740 5907 1808 5963
rect 1864 5907 1874 5963
rect 1426 5839 1874 5907
rect 1426 5783 1436 5839
rect 1492 5783 1560 5839
rect 1616 5783 1684 5839
rect 1740 5783 1808 5839
rect 1864 5783 1874 5839
rect 1426 5715 1874 5783
rect 1426 5659 1436 5715
rect 1492 5659 1560 5715
rect 1616 5659 1684 5715
rect 1740 5659 1808 5715
rect 1864 5659 1874 5715
rect 1426 5591 1874 5659
rect 1426 5535 1436 5591
rect 1492 5535 1560 5591
rect 1616 5535 1684 5591
rect 1740 5535 1808 5591
rect 1864 5535 1874 5591
rect 1426 5467 1874 5535
rect 1426 5411 1436 5467
rect 1492 5411 1560 5467
rect 1616 5411 1684 5467
rect 1740 5411 1808 5467
rect 1864 5411 1874 5467
rect 1426 5343 1874 5411
rect 1426 5287 1436 5343
rect 1492 5287 1560 5343
rect 1616 5287 1684 5343
rect 1740 5287 1808 5343
rect 1864 5287 1874 5343
rect 1426 5219 1874 5287
rect 1426 5163 1436 5219
rect 1492 5163 1560 5219
rect 1616 5163 1684 5219
rect 1740 5163 1808 5219
rect 1864 5163 1874 5219
rect 1426 5095 1874 5163
rect 1426 5039 1436 5095
rect 1492 5039 1560 5095
rect 1616 5039 1684 5095
rect 1740 5039 1808 5095
rect 1864 5039 1874 5095
rect 1426 4971 1874 5039
rect 1426 4915 1436 4971
rect 1492 4915 1560 4971
rect 1616 4915 1684 4971
rect 1740 4915 1808 4971
rect 1864 4915 1874 4971
rect 1426 4847 1874 4915
rect 1426 4791 1436 4847
rect 1492 4791 1560 4847
rect 1616 4791 1684 4847
rect 1740 4791 1808 4847
rect 1864 4791 1874 4847
rect 1426 4723 1874 4791
rect 1426 4667 1436 4723
rect 1492 4667 1560 4723
rect 1616 4667 1684 4723
rect 1740 4667 1808 4723
rect 1864 4667 1874 4723
rect 1426 4599 1874 4667
rect 1426 4543 1436 4599
rect 1492 4543 1560 4599
rect 1616 4543 1684 4599
rect 1740 4543 1808 4599
rect 1864 4543 1874 4599
rect 1426 4533 1874 4543
rect 2562 7451 3010 7461
rect 2562 7395 2572 7451
rect 2628 7395 2696 7451
rect 2752 7395 2820 7451
rect 2876 7395 2944 7451
rect 3000 7395 3010 7451
rect 2562 7327 3010 7395
rect 2562 7271 2572 7327
rect 2628 7271 2696 7327
rect 2752 7271 2820 7327
rect 2876 7271 2944 7327
rect 3000 7271 3010 7327
rect 2562 7203 3010 7271
rect 2562 7147 2572 7203
rect 2628 7147 2696 7203
rect 2752 7147 2820 7203
rect 2876 7147 2944 7203
rect 3000 7147 3010 7203
rect 2562 7079 3010 7147
rect 2562 7023 2572 7079
rect 2628 7023 2696 7079
rect 2752 7023 2820 7079
rect 2876 7023 2944 7079
rect 3000 7023 3010 7079
rect 2562 6955 3010 7023
rect 2562 6899 2572 6955
rect 2628 6899 2696 6955
rect 2752 6899 2820 6955
rect 2876 6899 2944 6955
rect 3000 6899 3010 6955
rect 2562 6831 3010 6899
rect 2562 6775 2572 6831
rect 2628 6775 2696 6831
rect 2752 6775 2820 6831
rect 2876 6775 2944 6831
rect 3000 6775 3010 6831
rect 2562 6707 3010 6775
rect 2562 6651 2572 6707
rect 2628 6651 2696 6707
rect 2752 6651 2820 6707
rect 2876 6651 2944 6707
rect 3000 6651 3010 6707
rect 2562 6583 3010 6651
rect 2562 6527 2572 6583
rect 2628 6527 2696 6583
rect 2752 6527 2820 6583
rect 2876 6527 2944 6583
rect 3000 6527 3010 6583
rect 2562 6459 3010 6527
rect 2562 6403 2572 6459
rect 2628 6403 2696 6459
rect 2752 6403 2820 6459
rect 2876 6403 2944 6459
rect 3000 6403 3010 6459
rect 2562 6335 3010 6403
rect 2562 6279 2572 6335
rect 2628 6279 2696 6335
rect 2752 6279 2820 6335
rect 2876 6279 2944 6335
rect 3000 6279 3010 6335
rect 2562 6211 3010 6279
rect 2562 6155 2572 6211
rect 2628 6155 2696 6211
rect 2752 6155 2820 6211
rect 2876 6155 2944 6211
rect 3000 6155 3010 6211
rect 2562 6087 3010 6155
rect 2562 6031 2572 6087
rect 2628 6031 2696 6087
rect 2752 6031 2820 6087
rect 2876 6031 2944 6087
rect 3000 6031 3010 6087
rect 2562 5963 3010 6031
rect 2562 5907 2572 5963
rect 2628 5907 2696 5963
rect 2752 5907 2820 5963
rect 2876 5907 2944 5963
rect 3000 5907 3010 5963
rect 2562 5839 3010 5907
rect 2562 5783 2572 5839
rect 2628 5783 2696 5839
rect 2752 5783 2820 5839
rect 2876 5783 2944 5839
rect 3000 5783 3010 5839
rect 2562 5715 3010 5783
rect 2562 5659 2572 5715
rect 2628 5659 2696 5715
rect 2752 5659 2820 5715
rect 2876 5659 2944 5715
rect 3000 5659 3010 5715
rect 2562 5591 3010 5659
rect 2562 5535 2572 5591
rect 2628 5535 2696 5591
rect 2752 5535 2820 5591
rect 2876 5535 2944 5591
rect 3000 5535 3010 5591
rect 2562 5467 3010 5535
rect 2562 5411 2572 5467
rect 2628 5411 2696 5467
rect 2752 5411 2820 5467
rect 2876 5411 2944 5467
rect 3000 5411 3010 5467
rect 2562 5343 3010 5411
rect 2562 5287 2572 5343
rect 2628 5287 2696 5343
rect 2752 5287 2820 5343
rect 2876 5287 2944 5343
rect 3000 5287 3010 5343
rect 2562 5219 3010 5287
rect 2562 5163 2572 5219
rect 2628 5163 2696 5219
rect 2752 5163 2820 5219
rect 2876 5163 2944 5219
rect 3000 5163 3010 5219
rect 2562 5095 3010 5163
rect 2562 5039 2572 5095
rect 2628 5039 2696 5095
rect 2752 5039 2820 5095
rect 2876 5039 2944 5095
rect 3000 5039 3010 5095
rect 2562 4971 3010 5039
rect 2562 4915 2572 4971
rect 2628 4915 2696 4971
rect 2752 4915 2820 4971
rect 2876 4915 2944 4971
rect 3000 4915 3010 4971
rect 2562 4847 3010 4915
rect 2562 4791 2572 4847
rect 2628 4791 2696 4847
rect 2752 4791 2820 4847
rect 2876 4791 2944 4847
rect 3000 4791 3010 4847
rect 2562 4723 3010 4791
rect 2562 4667 2572 4723
rect 2628 4667 2696 4723
rect 2752 4667 2820 4723
rect 2876 4667 2944 4723
rect 3000 4667 3010 4723
rect 2562 4599 3010 4667
rect 2562 4543 2572 4599
rect 2628 4543 2696 4599
rect 2752 4543 2820 4599
rect 2876 4543 2944 4599
rect 3000 4543 3010 4599
rect 2562 4533 3010 4543
rect 4834 7451 5282 7461
rect 4834 7395 4844 7451
rect 4900 7395 4968 7451
rect 5024 7395 5092 7451
rect 5148 7395 5216 7451
rect 5272 7395 5282 7451
rect 4834 7327 5282 7395
rect 4834 7271 4844 7327
rect 4900 7271 4968 7327
rect 5024 7271 5092 7327
rect 5148 7271 5216 7327
rect 5272 7271 5282 7327
rect 4834 7203 5282 7271
rect 4834 7147 4844 7203
rect 4900 7147 4968 7203
rect 5024 7147 5092 7203
rect 5148 7147 5216 7203
rect 5272 7147 5282 7203
rect 4834 7079 5282 7147
rect 4834 7023 4844 7079
rect 4900 7023 4968 7079
rect 5024 7023 5092 7079
rect 5148 7023 5216 7079
rect 5272 7023 5282 7079
rect 4834 6955 5282 7023
rect 4834 6899 4844 6955
rect 4900 6899 4968 6955
rect 5024 6899 5092 6955
rect 5148 6899 5216 6955
rect 5272 6899 5282 6955
rect 4834 6831 5282 6899
rect 4834 6775 4844 6831
rect 4900 6775 4968 6831
rect 5024 6775 5092 6831
rect 5148 6775 5216 6831
rect 5272 6775 5282 6831
rect 4834 6707 5282 6775
rect 4834 6651 4844 6707
rect 4900 6651 4968 6707
rect 5024 6651 5092 6707
rect 5148 6651 5216 6707
rect 5272 6651 5282 6707
rect 4834 6583 5282 6651
rect 4834 6527 4844 6583
rect 4900 6527 4968 6583
rect 5024 6527 5092 6583
rect 5148 6527 5216 6583
rect 5272 6527 5282 6583
rect 4834 6459 5282 6527
rect 4834 6403 4844 6459
rect 4900 6403 4968 6459
rect 5024 6403 5092 6459
rect 5148 6403 5216 6459
rect 5272 6403 5282 6459
rect 4834 6335 5282 6403
rect 4834 6279 4844 6335
rect 4900 6279 4968 6335
rect 5024 6279 5092 6335
rect 5148 6279 5216 6335
rect 5272 6279 5282 6335
rect 4834 6211 5282 6279
rect 4834 6155 4844 6211
rect 4900 6155 4968 6211
rect 5024 6155 5092 6211
rect 5148 6155 5216 6211
rect 5272 6155 5282 6211
rect 4834 6087 5282 6155
rect 4834 6031 4844 6087
rect 4900 6031 4968 6087
rect 5024 6031 5092 6087
rect 5148 6031 5216 6087
rect 5272 6031 5282 6087
rect 4834 5963 5282 6031
rect 4834 5907 4844 5963
rect 4900 5907 4968 5963
rect 5024 5907 5092 5963
rect 5148 5907 5216 5963
rect 5272 5907 5282 5963
rect 4834 5839 5282 5907
rect 4834 5783 4844 5839
rect 4900 5783 4968 5839
rect 5024 5783 5092 5839
rect 5148 5783 5216 5839
rect 5272 5783 5282 5839
rect 4834 5715 5282 5783
rect 4834 5659 4844 5715
rect 4900 5659 4968 5715
rect 5024 5659 5092 5715
rect 5148 5659 5216 5715
rect 5272 5659 5282 5715
rect 4834 5591 5282 5659
rect 4834 5535 4844 5591
rect 4900 5535 4968 5591
rect 5024 5535 5092 5591
rect 5148 5535 5216 5591
rect 5272 5535 5282 5591
rect 4834 5467 5282 5535
rect 4834 5411 4844 5467
rect 4900 5411 4968 5467
rect 5024 5411 5092 5467
rect 5148 5411 5216 5467
rect 5272 5411 5282 5467
rect 4834 5343 5282 5411
rect 4834 5287 4844 5343
rect 4900 5287 4968 5343
rect 5024 5287 5092 5343
rect 5148 5287 5216 5343
rect 5272 5287 5282 5343
rect 4834 5219 5282 5287
rect 4834 5163 4844 5219
rect 4900 5163 4968 5219
rect 5024 5163 5092 5219
rect 5148 5163 5216 5219
rect 5272 5163 5282 5219
rect 4834 5095 5282 5163
rect 4834 5039 4844 5095
rect 4900 5039 4968 5095
rect 5024 5039 5092 5095
rect 5148 5039 5216 5095
rect 5272 5039 5282 5095
rect 4834 4971 5282 5039
rect 4834 4915 4844 4971
rect 4900 4915 4968 4971
rect 5024 4915 5092 4971
rect 5148 4915 5216 4971
rect 5272 4915 5282 4971
rect 4834 4847 5282 4915
rect 4834 4791 4844 4847
rect 4900 4791 4968 4847
rect 5024 4791 5092 4847
rect 5148 4791 5216 4847
rect 5272 4791 5282 4847
rect 4834 4723 5282 4791
rect 4834 4667 4844 4723
rect 4900 4667 4968 4723
rect 5024 4667 5092 4723
rect 5148 4667 5216 4723
rect 5272 4667 5282 4723
rect 4834 4599 5282 4667
rect 4834 4543 4844 4599
rect 4900 4543 4968 4599
rect 5024 4543 5092 4599
rect 5148 4543 5216 4599
rect 5272 4543 5282 4599
rect 4834 4533 5282 4543
rect 7127 7451 7451 7461
rect 7127 7395 7137 7451
rect 7193 7395 7261 7451
rect 7317 7395 7385 7451
rect 7441 7395 7451 7451
rect 7127 7327 7451 7395
rect 7127 7271 7137 7327
rect 7193 7271 7261 7327
rect 7317 7271 7385 7327
rect 7441 7271 7451 7327
rect 7127 7203 7451 7271
rect 7127 7147 7137 7203
rect 7193 7147 7261 7203
rect 7317 7147 7385 7203
rect 7441 7147 7451 7203
rect 7127 7079 7451 7147
rect 7127 7023 7137 7079
rect 7193 7023 7261 7079
rect 7317 7023 7385 7079
rect 7441 7023 7451 7079
rect 7127 6955 7451 7023
rect 7127 6899 7137 6955
rect 7193 6899 7261 6955
rect 7317 6899 7385 6955
rect 7441 6899 7451 6955
rect 7127 6831 7451 6899
rect 7127 6775 7137 6831
rect 7193 6775 7261 6831
rect 7317 6775 7385 6831
rect 7441 6775 7451 6831
rect 7127 6707 7451 6775
rect 7127 6651 7137 6707
rect 7193 6651 7261 6707
rect 7317 6651 7385 6707
rect 7441 6651 7451 6707
rect 7127 6583 7451 6651
rect 7127 6527 7137 6583
rect 7193 6527 7261 6583
rect 7317 6527 7385 6583
rect 7441 6527 7451 6583
rect 7127 6459 7451 6527
rect 7127 6403 7137 6459
rect 7193 6403 7261 6459
rect 7317 6403 7385 6459
rect 7441 6403 7451 6459
rect 7127 6335 7451 6403
rect 7127 6279 7137 6335
rect 7193 6279 7261 6335
rect 7317 6279 7385 6335
rect 7441 6279 7451 6335
rect 7127 6211 7451 6279
rect 7127 6155 7137 6211
rect 7193 6155 7261 6211
rect 7317 6155 7385 6211
rect 7441 6155 7451 6211
rect 7127 6087 7451 6155
rect 7127 6031 7137 6087
rect 7193 6031 7261 6087
rect 7317 6031 7385 6087
rect 7441 6031 7451 6087
rect 7127 5963 7451 6031
rect 7127 5907 7137 5963
rect 7193 5907 7261 5963
rect 7317 5907 7385 5963
rect 7441 5907 7451 5963
rect 7127 5839 7451 5907
rect 7127 5783 7137 5839
rect 7193 5783 7261 5839
rect 7317 5783 7385 5839
rect 7441 5783 7451 5839
rect 7127 5715 7451 5783
rect 7127 5659 7137 5715
rect 7193 5659 7261 5715
rect 7317 5659 7385 5715
rect 7441 5659 7451 5715
rect 7127 5591 7451 5659
rect 7127 5535 7137 5591
rect 7193 5535 7261 5591
rect 7317 5535 7385 5591
rect 7441 5535 7451 5591
rect 7127 5467 7451 5535
rect 7127 5411 7137 5467
rect 7193 5411 7261 5467
rect 7317 5411 7385 5467
rect 7441 5411 7451 5467
rect 7127 5343 7451 5411
rect 7127 5287 7137 5343
rect 7193 5287 7261 5343
rect 7317 5287 7385 5343
rect 7441 5287 7451 5343
rect 7127 5219 7451 5287
rect 7127 5163 7137 5219
rect 7193 5163 7261 5219
rect 7317 5163 7385 5219
rect 7441 5163 7451 5219
rect 7127 5095 7451 5163
rect 7127 5039 7137 5095
rect 7193 5039 7261 5095
rect 7317 5039 7385 5095
rect 7441 5039 7451 5095
rect 7127 4971 7451 5039
rect 7127 4915 7137 4971
rect 7193 4915 7261 4971
rect 7317 4915 7385 4971
rect 7441 4915 7451 4971
rect 7127 4847 7451 4915
rect 7127 4791 7137 4847
rect 7193 4791 7261 4847
rect 7317 4791 7385 4847
rect 7441 4791 7451 4847
rect 7127 4723 7451 4791
rect 7127 4667 7137 4723
rect 7193 4667 7261 4723
rect 7317 4667 7385 4723
rect 7441 4667 7451 4723
rect 7127 4599 7451 4667
rect 7127 4543 7137 4599
rect 7193 4543 7261 4599
rect 7317 4543 7385 4599
rect 7441 4543 7451 4599
rect 7127 4533 7451 4543
rect 7613 7451 7937 7461
rect 7613 7395 7623 7451
rect 7679 7395 7747 7451
rect 7803 7395 7871 7451
rect 7927 7395 7937 7451
rect 7613 7327 7937 7395
rect 7613 7271 7623 7327
rect 7679 7271 7747 7327
rect 7803 7271 7871 7327
rect 7927 7271 7937 7327
rect 7613 7203 7937 7271
rect 7613 7147 7623 7203
rect 7679 7147 7747 7203
rect 7803 7147 7871 7203
rect 7927 7147 7937 7203
rect 7613 7079 7937 7147
rect 7613 7023 7623 7079
rect 7679 7023 7747 7079
rect 7803 7023 7871 7079
rect 7927 7023 7937 7079
rect 7613 6955 7937 7023
rect 7613 6899 7623 6955
rect 7679 6899 7747 6955
rect 7803 6899 7871 6955
rect 7927 6899 7937 6955
rect 7613 6831 7937 6899
rect 7613 6775 7623 6831
rect 7679 6775 7747 6831
rect 7803 6775 7871 6831
rect 7927 6775 7937 6831
rect 7613 6707 7937 6775
rect 7613 6651 7623 6707
rect 7679 6651 7747 6707
rect 7803 6651 7871 6707
rect 7927 6651 7937 6707
rect 7613 6583 7937 6651
rect 7613 6527 7623 6583
rect 7679 6527 7747 6583
rect 7803 6527 7871 6583
rect 7927 6527 7937 6583
rect 7613 6459 7937 6527
rect 7613 6403 7623 6459
rect 7679 6403 7747 6459
rect 7803 6403 7871 6459
rect 7927 6403 7937 6459
rect 7613 6335 7937 6403
rect 7613 6279 7623 6335
rect 7679 6279 7747 6335
rect 7803 6279 7871 6335
rect 7927 6279 7937 6335
rect 7613 6211 7937 6279
rect 7613 6155 7623 6211
rect 7679 6155 7747 6211
rect 7803 6155 7871 6211
rect 7927 6155 7937 6211
rect 7613 6087 7937 6155
rect 7613 6031 7623 6087
rect 7679 6031 7747 6087
rect 7803 6031 7871 6087
rect 7927 6031 7937 6087
rect 7613 5963 7937 6031
rect 7613 5907 7623 5963
rect 7679 5907 7747 5963
rect 7803 5907 7871 5963
rect 7927 5907 7937 5963
rect 7613 5839 7937 5907
rect 7613 5783 7623 5839
rect 7679 5783 7747 5839
rect 7803 5783 7871 5839
rect 7927 5783 7937 5839
rect 7613 5715 7937 5783
rect 7613 5659 7623 5715
rect 7679 5659 7747 5715
rect 7803 5659 7871 5715
rect 7927 5659 7937 5715
rect 7613 5591 7937 5659
rect 7613 5535 7623 5591
rect 7679 5535 7747 5591
rect 7803 5535 7871 5591
rect 7927 5535 7937 5591
rect 7613 5467 7937 5535
rect 7613 5411 7623 5467
rect 7679 5411 7747 5467
rect 7803 5411 7871 5467
rect 7927 5411 7937 5467
rect 7613 5343 7937 5411
rect 7613 5287 7623 5343
rect 7679 5287 7747 5343
rect 7803 5287 7871 5343
rect 7927 5287 7937 5343
rect 7613 5219 7937 5287
rect 7613 5163 7623 5219
rect 7679 5163 7747 5219
rect 7803 5163 7871 5219
rect 7927 5163 7937 5219
rect 7613 5095 7937 5163
rect 7613 5039 7623 5095
rect 7679 5039 7747 5095
rect 7803 5039 7871 5095
rect 7927 5039 7937 5095
rect 7613 4971 7937 5039
rect 7613 4915 7623 4971
rect 7679 4915 7747 4971
rect 7803 4915 7871 4971
rect 7927 4915 7937 4971
rect 7613 4847 7937 4915
rect 7613 4791 7623 4847
rect 7679 4791 7747 4847
rect 7803 4791 7871 4847
rect 7927 4791 7937 4847
rect 7613 4723 7937 4791
rect 7613 4667 7623 4723
rect 7679 4667 7747 4723
rect 7803 4667 7871 4723
rect 7927 4667 7937 4723
rect 7613 4599 7937 4667
rect 7613 4543 7623 4599
rect 7679 4543 7747 4599
rect 7803 4543 7871 4599
rect 7927 4543 7937 4599
rect 7613 4533 7937 4543
rect 9782 7451 10230 7461
rect 9782 7395 9792 7451
rect 9848 7395 9916 7451
rect 9972 7395 10040 7451
rect 10096 7395 10164 7451
rect 10220 7395 10230 7451
rect 9782 7327 10230 7395
rect 9782 7271 9792 7327
rect 9848 7271 9916 7327
rect 9972 7271 10040 7327
rect 10096 7271 10164 7327
rect 10220 7271 10230 7327
rect 9782 7203 10230 7271
rect 9782 7147 9792 7203
rect 9848 7147 9916 7203
rect 9972 7147 10040 7203
rect 10096 7147 10164 7203
rect 10220 7147 10230 7203
rect 9782 7079 10230 7147
rect 9782 7023 9792 7079
rect 9848 7023 9916 7079
rect 9972 7023 10040 7079
rect 10096 7023 10164 7079
rect 10220 7023 10230 7079
rect 9782 6955 10230 7023
rect 9782 6899 9792 6955
rect 9848 6899 9916 6955
rect 9972 6899 10040 6955
rect 10096 6899 10164 6955
rect 10220 6899 10230 6955
rect 9782 6831 10230 6899
rect 9782 6775 9792 6831
rect 9848 6775 9916 6831
rect 9972 6775 10040 6831
rect 10096 6775 10164 6831
rect 10220 6775 10230 6831
rect 9782 6707 10230 6775
rect 9782 6651 9792 6707
rect 9848 6651 9916 6707
rect 9972 6651 10040 6707
rect 10096 6651 10164 6707
rect 10220 6651 10230 6707
rect 9782 6583 10230 6651
rect 9782 6527 9792 6583
rect 9848 6527 9916 6583
rect 9972 6527 10040 6583
rect 10096 6527 10164 6583
rect 10220 6527 10230 6583
rect 9782 6459 10230 6527
rect 9782 6403 9792 6459
rect 9848 6403 9916 6459
rect 9972 6403 10040 6459
rect 10096 6403 10164 6459
rect 10220 6403 10230 6459
rect 9782 6335 10230 6403
rect 9782 6279 9792 6335
rect 9848 6279 9916 6335
rect 9972 6279 10040 6335
rect 10096 6279 10164 6335
rect 10220 6279 10230 6335
rect 9782 6211 10230 6279
rect 9782 6155 9792 6211
rect 9848 6155 9916 6211
rect 9972 6155 10040 6211
rect 10096 6155 10164 6211
rect 10220 6155 10230 6211
rect 9782 6087 10230 6155
rect 9782 6031 9792 6087
rect 9848 6031 9916 6087
rect 9972 6031 10040 6087
rect 10096 6031 10164 6087
rect 10220 6031 10230 6087
rect 9782 5963 10230 6031
rect 9782 5907 9792 5963
rect 9848 5907 9916 5963
rect 9972 5907 10040 5963
rect 10096 5907 10164 5963
rect 10220 5907 10230 5963
rect 9782 5839 10230 5907
rect 9782 5783 9792 5839
rect 9848 5783 9916 5839
rect 9972 5783 10040 5839
rect 10096 5783 10164 5839
rect 10220 5783 10230 5839
rect 9782 5715 10230 5783
rect 9782 5659 9792 5715
rect 9848 5659 9916 5715
rect 9972 5659 10040 5715
rect 10096 5659 10164 5715
rect 10220 5659 10230 5715
rect 9782 5591 10230 5659
rect 9782 5535 9792 5591
rect 9848 5535 9916 5591
rect 9972 5535 10040 5591
rect 10096 5535 10164 5591
rect 10220 5535 10230 5591
rect 9782 5467 10230 5535
rect 9782 5411 9792 5467
rect 9848 5411 9916 5467
rect 9972 5411 10040 5467
rect 10096 5411 10164 5467
rect 10220 5411 10230 5467
rect 9782 5343 10230 5411
rect 9782 5287 9792 5343
rect 9848 5287 9916 5343
rect 9972 5287 10040 5343
rect 10096 5287 10164 5343
rect 10220 5287 10230 5343
rect 9782 5219 10230 5287
rect 9782 5163 9792 5219
rect 9848 5163 9916 5219
rect 9972 5163 10040 5219
rect 10096 5163 10164 5219
rect 10220 5163 10230 5219
rect 9782 5095 10230 5163
rect 9782 5039 9792 5095
rect 9848 5039 9916 5095
rect 9972 5039 10040 5095
rect 10096 5039 10164 5095
rect 10220 5039 10230 5095
rect 9782 4971 10230 5039
rect 9782 4915 9792 4971
rect 9848 4915 9916 4971
rect 9972 4915 10040 4971
rect 10096 4915 10164 4971
rect 10220 4915 10230 4971
rect 9782 4847 10230 4915
rect 9782 4791 9792 4847
rect 9848 4791 9916 4847
rect 9972 4791 10040 4847
rect 10096 4791 10164 4847
rect 10220 4791 10230 4847
rect 9782 4723 10230 4791
rect 9782 4667 9792 4723
rect 9848 4667 9916 4723
rect 9972 4667 10040 4723
rect 10096 4667 10164 4723
rect 10220 4667 10230 4723
rect 9782 4599 10230 4667
rect 9782 4543 9792 4599
rect 9848 4543 9916 4599
rect 9972 4543 10040 4599
rect 10096 4543 10164 4599
rect 10220 4543 10230 4599
rect 9782 4533 10230 4543
rect 12054 7451 12502 7461
rect 12054 7395 12064 7451
rect 12120 7395 12188 7451
rect 12244 7395 12312 7451
rect 12368 7395 12436 7451
rect 12492 7395 12502 7451
rect 12054 7327 12502 7395
rect 12054 7271 12064 7327
rect 12120 7271 12188 7327
rect 12244 7271 12312 7327
rect 12368 7271 12436 7327
rect 12492 7271 12502 7327
rect 12054 7203 12502 7271
rect 12054 7147 12064 7203
rect 12120 7147 12188 7203
rect 12244 7147 12312 7203
rect 12368 7147 12436 7203
rect 12492 7147 12502 7203
rect 12054 7079 12502 7147
rect 12054 7023 12064 7079
rect 12120 7023 12188 7079
rect 12244 7023 12312 7079
rect 12368 7023 12436 7079
rect 12492 7023 12502 7079
rect 12054 6955 12502 7023
rect 12054 6899 12064 6955
rect 12120 6899 12188 6955
rect 12244 6899 12312 6955
rect 12368 6899 12436 6955
rect 12492 6899 12502 6955
rect 12054 6831 12502 6899
rect 12054 6775 12064 6831
rect 12120 6775 12188 6831
rect 12244 6775 12312 6831
rect 12368 6775 12436 6831
rect 12492 6775 12502 6831
rect 12054 6707 12502 6775
rect 12054 6651 12064 6707
rect 12120 6651 12188 6707
rect 12244 6651 12312 6707
rect 12368 6651 12436 6707
rect 12492 6651 12502 6707
rect 12054 6583 12502 6651
rect 12054 6527 12064 6583
rect 12120 6527 12188 6583
rect 12244 6527 12312 6583
rect 12368 6527 12436 6583
rect 12492 6527 12502 6583
rect 12054 6459 12502 6527
rect 12054 6403 12064 6459
rect 12120 6403 12188 6459
rect 12244 6403 12312 6459
rect 12368 6403 12436 6459
rect 12492 6403 12502 6459
rect 12054 6335 12502 6403
rect 12054 6279 12064 6335
rect 12120 6279 12188 6335
rect 12244 6279 12312 6335
rect 12368 6279 12436 6335
rect 12492 6279 12502 6335
rect 12054 6211 12502 6279
rect 12054 6155 12064 6211
rect 12120 6155 12188 6211
rect 12244 6155 12312 6211
rect 12368 6155 12436 6211
rect 12492 6155 12502 6211
rect 12054 6087 12502 6155
rect 12054 6031 12064 6087
rect 12120 6031 12188 6087
rect 12244 6031 12312 6087
rect 12368 6031 12436 6087
rect 12492 6031 12502 6087
rect 12054 5963 12502 6031
rect 12054 5907 12064 5963
rect 12120 5907 12188 5963
rect 12244 5907 12312 5963
rect 12368 5907 12436 5963
rect 12492 5907 12502 5963
rect 12054 5839 12502 5907
rect 12054 5783 12064 5839
rect 12120 5783 12188 5839
rect 12244 5783 12312 5839
rect 12368 5783 12436 5839
rect 12492 5783 12502 5839
rect 12054 5715 12502 5783
rect 12054 5659 12064 5715
rect 12120 5659 12188 5715
rect 12244 5659 12312 5715
rect 12368 5659 12436 5715
rect 12492 5659 12502 5715
rect 12054 5591 12502 5659
rect 12054 5535 12064 5591
rect 12120 5535 12188 5591
rect 12244 5535 12312 5591
rect 12368 5535 12436 5591
rect 12492 5535 12502 5591
rect 12054 5467 12502 5535
rect 12054 5411 12064 5467
rect 12120 5411 12188 5467
rect 12244 5411 12312 5467
rect 12368 5411 12436 5467
rect 12492 5411 12502 5467
rect 12054 5343 12502 5411
rect 12054 5287 12064 5343
rect 12120 5287 12188 5343
rect 12244 5287 12312 5343
rect 12368 5287 12436 5343
rect 12492 5287 12502 5343
rect 12054 5219 12502 5287
rect 12054 5163 12064 5219
rect 12120 5163 12188 5219
rect 12244 5163 12312 5219
rect 12368 5163 12436 5219
rect 12492 5163 12502 5219
rect 12054 5095 12502 5163
rect 12054 5039 12064 5095
rect 12120 5039 12188 5095
rect 12244 5039 12312 5095
rect 12368 5039 12436 5095
rect 12492 5039 12502 5095
rect 12054 4971 12502 5039
rect 12054 4915 12064 4971
rect 12120 4915 12188 4971
rect 12244 4915 12312 4971
rect 12368 4915 12436 4971
rect 12492 4915 12502 4971
rect 12054 4847 12502 4915
rect 12054 4791 12064 4847
rect 12120 4791 12188 4847
rect 12244 4791 12312 4847
rect 12368 4791 12436 4847
rect 12492 4791 12502 4847
rect 12054 4723 12502 4791
rect 12054 4667 12064 4723
rect 12120 4667 12188 4723
rect 12244 4667 12312 4723
rect 12368 4667 12436 4723
rect 12492 4667 12502 4723
rect 12054 4599 12502 4667
rect 12054 4543 12064 4599
rect 12120 4543 12188 4599
rect 12244 4543 12312 4599
rect 12368 4543 12436 4599
rect 12492 4543 12502 4599
rect 12054 4533 12502 4543
rect 13190 7451 13638 7461
rect 13190 7395 13200 7451
rect 13256 7395 13324 7451
rect 13380 7395 13448 7451
rect 13504 7395 13572 7451
rect 13628 7395 13638 7451
rect 13190 7327 13638 7395
rect 13190 7271 13200 7327
rect 13256 7271 13324 7327
rect 13380 7271 13448 7327
rect 13504 7271 13572 7327
rect 13628 7271 13638 7327
rect 13190 7203 13638 7271
rect 13190 7147 13200 7203
rect 13256 7147 13324 7203
rect 13380 7147 13448 7203
rect 13504 7147 13572 7203
rect 13628 7147 13638 7203
rect 13190 7079 13638 7147
rect 13190 7023 13200 7079
rect 13256 7023 13324 7079
rect 13380 7023 13448 7079
rect 13504 7023 13572 7079
rect 13628 7023 13638 7079
rect 13190 6955 13638 7023
rect 13190 6899 13200 6955
rect 13256 6899 13324 6955
rect 13380 6899 13448 6955
rect 13504 6899 13572 6955
rect 13628 6899 13638 6955
rect 13190 6831 13638 6899
rect 13190 6775 13200 6831
rect 13256 6775 13324 6831
rect 13380 6775 13448 6831
rect 13504 6775 13572 6831
rect 13628 6775 13638 6831
rect 13190 6707 13638 6775
rect 13190 6651 13200 6707
rect 13256 6651 13324 6707
rect 13380 6651 13448 6707
rect 13504 6651 13572 6707
rect 13628 6651 13638 6707
rect 13190 6583 13638 6651
rect 13190 6527 13200 6583
rect 13256 6527 13324 6583
rect 13380 6527 13448 6583
rect 13504 6527 13572 6583
rect 13628 6527 13638 6583
rect 13190 6459 13638 6527
rect 13190 6403 13200 6459
rect 13256 6403 13324 6459
rect 13380 6403 13448 6459
rect 13504 6403 13572 6459
rect 13628 6403 13638 6459
rect 13190 6335 13638 6403
rect 13190 6279 13200 6335
rect 13256 6279 13324 6335
rect 13380 6279 13448 6335
rect 13504 6279 13572 6335
rect 13628 6279 13638 6335
rect 13190 6211 13638 6279
rect 13190 6155 13200 6211
rect 13256 6155 13324 6211
rect 13380 6155 13448 6211
rect 13504 6155 13572 6211
rect 13628 6155 13638 6211
rect 13190 6087 13638 6155
rect 13190 6031 13200 6087
rect 13256 6031 13324 6087
rect 13380 6031 13448 6087
rect 13504 6031 13572 6087
rect 13628 6031 13638 6087
rect 13190 5963 13638 6031
rect 13190 5907 13200 5963
rect 13256 5907 13324 5963
rect 13380 5907 13448 5963
rect 13504 5907 13572 5963
rect 13628 5907 13638 5963
rect 13190 5839 13638 5907
rect 13190 5783 13200 5839
rect 13256 5783 13324 5839
rect 13380 5783 13448 5839
rect 13504 5783 13572 5839
rect 13628 5783 13638 5839
rect 13190 5715 13638 5783
rect 13190 5659 13200 5715
rect 13256 5659 13324 5715
rect 13380 5659 13448 5715
rect 13504 5659 13572 5715
rect 13628 5659 13638 5715
rect 13190 5591 13638 5659
rect 13190 5535 13200 5591
rect 13256 5535 13324 5591
rect 13380 5535 13448 5591
rect 13504 5535 13572 5591
rect 13628 5535 13638 5591
rect 13190 5467 13638 5535
rect 13190 5411 13200 5467
rect 13256 5411 13324 5467
rect 13380 5411 13448 5467
rect 13504 5411 13572 5467
rect 13628 5411 13638 5467
rect 13190 5343 13638 5411
rect 13190 5287 13200 5343
rect 13256 5287 13324 5343
rect 13380 5287 13448 5343
rect 13504 5287 13572 5343
rect 13628 5287 13638 5343
rect 13190 5219 13638 5287
rect 13190 5163 13200 5219
rect 13256 5163 13324 5219
rect 13380 5163 13448 5219
rect 13504 5163 13572 5219
rect 13628 5163 13638 5219
rect 13190 5095 13638 5163
rect 13190 5039 13200 5095
rect 13256 5039 13324 5095
rect 13380 5039 13448 5095
rect 13504 5039 13572 5095
rect 13628 5039 13638 5095
rect 13190 4971 13638 5039
rect 13190 4915 13200 4971
rect 13256 4915 13324 4971
rect 13380 4915 13448 4971
rect 13504 4915 13572 4971
rect 13628 4915 13638 4971
rect 13190 4847 13638 4915
rect 13190 4791 13200 4847
rect 13256 4791 13324 4847
rect 13380 4791 13448 4847
rect 13504 4791 13572 4847
rect 13628 4791 13638 4847
rect 13190 4723 13638 4791
rect 13190 4667 13200 4723
rect 13256 4667 13324 4723
rect 13380 4667 13448 4723
rect 13504 4667 13572 4723
rect 13628 4667 13638 4723
rect 13190 4599 13638 4667
rect 13190 4543 13200 4599
rect 13256 4543 13324 4599
rect 13380 4543 13448 4599
rect 13504 4543 13572 4599
rect 13628 4543 13638 4599
rect 13190 4533 13638 4543
rect 1426 4251 1874 4261
rect 1426 4195 1436 4251
rect 1492 4195 1560 4251
rect 1616 4195 1684 4251
rect 1740 4195 1808 4251
rect 1864 4195 1874 4251
rect 1426 4127 1874 4195
rect 1426 4071 1436 4127
rect 1492 4071 1560 4127
rect 1616 4071 1684 4127
rect 1740 4071 1808 4127
rect 1864 4071 1874 4127
rect 1426 4003 1874 4071
rect 1426 3947 1436 4003
rect 1492 3947 1560 4003
rect 1616 3947 1684 4003
rect 1740 3947 1808 4003
rect 1864 3947 1874 4003
rect 1426 3879 1874 3947
rect 1426 3823 1436 3879
rect 1492 3823 1560 3879
rect 1616 3823 1684 3879
rect 1740 3823 1808 3879
rect 1864 3823 1874 3879
rect 1426 3755 1874 3823
rect 1426 3699 1436 3755
rect 1492 3699 1560 3755
rect 1616 3699 1684 3755
rect 1740 3699 1808 3755
rect 1864 3699 1874 3755
rect 1426 3631 1874 3699
rect 1426 3575 1436 3631
rect 1492 3575 1560 3631
rect 1616 3575 1684 3631
rect 1740 3575 1808 3631
rect 1864 3575 1874 3631
rect 1426 3507 1874 3575
rect 1426 3451 1436 3507
rect 1492 3451 1560 3507
rect 1616 3451 1684 3507
rect 1740 3451 1808 3507
rect 1864 3451 1874 3507
rect 1426 3383 1874 3451
rect 1426 3327 1436 3383
rect 1492 3327 1560 3383
rect 1616 3327 1684 3383
rect 1740 3327 1808 3383
rect 1864 3327 1874 3383
rect 1426 3259 1874 3327
rect 1426 3203 1436 3259
rect 1492 3203 1560 3259
rect 1616 3203 1684 3259
rect 1740 3203 1808 3259
rect 1864 3203 1874 3259
rect 1426 3135 1874 3203
rect 1426 3079 1436 3135
rect 1492 3079 1560 3135
rect 1616 3079 1684 3135
rect 1740 3079 1808 3135
rect 1864 3079 1874 3135
rect 1426 3011 1874 3079
rect 1426 2955 1436 3011
rect 1492 2955 1560 3011
rect 1616 2955 1684 3011
rect 1740 2955 1808 3011
rect 1864 2955 1874 3011
rect 1426 2887 1874 2955
rect 1426 2831 1436 2887
rect 1492 2831 1560 2887
rect 1616 2831 1684 2887
rect 1740 2831 1808 2887
rect 1864 2831 1874 2887
rect 1426 2763 1874 2831
rect 1426 2707 1436 2763
rect 1492 2707 1560 2763
rect 1616 2707 1684 2763
rect 1740 2707 1808 2763
rect 1864 2707 1874 2763
rect 1426 2639 1874 2707
rect 1426 2583 1436 2639
rect 1492 2583 1560 2639
rect 1616 2583 1684 2639
rect 1740 2583 1808 2639
rect 1864 2583 1874 2639
rect 1426 2515 1874 2583
rect 1426 2459 1436 2515
rect 1492 2459 1560 2515
rect 1616 2459 1684 2515
rect 1740 2459 1808 2515
rect 1864 2459 1874 2515
rect 1426 2391 1874 2459
rect 1426 2335 1436 2391
rect 1492 2335 1560 2391
rect 1616 2335 1684 2391
rect 1740 2335 1808 2391
rect 1864 2335 1874 2391
rect 1426 2267 1874 2335
rect 1426 2211 1436 2267
rect 1492 2211 1560 2267
rect 1616 2211 1684 2267
rect 1740 2211 1808 2267
rect 1864 2211 1874 2267
rect 1426 2143 1874 2211
rect 1426 2087 1436 2143
rect 1492 2087 1560 2143
rect 1616 2087 1684 2143
rect 1740 2087 1808 2143
rect 1864 2087 1874 2143
rect 1426 2019 1874 2087
rect 1426 1963 1436 2019
rect 1492 1963 1560 2019
rect 1616 1963 1684 2019
rect 1740 1963 1808 2019
rect 1864 1963 1874 2019
rect 1426 1895 1874 1963
rect 1426 1839 1436 1895
rect 1492 1839 1560 1895
rect 1616 1839 1684 1895
rect 1740 1839 1808 1895
rect 1864 1839 1874 1895
rect 1426 1771 1874 1839
rect 1426 1715 1436 1771
rect 1492 1715 1560 1771
rect 1616 1715 1684 1771
rect 1740 1715 1808 1771
rect 1864 1715 1874 1771
rect 1426 1647 1874 1715
rect 1426 1591 1436 1647
rect 1492 1591 1560 1647
rect 1616 1591 1684 1647
rect 1740 1591 1808 1647
rect 1864 1591 1874 1647
rect 1426 1523 1874 1591
rect 1426 1467 1436 1523
rect 1492 1467 1560 1523
rect 1616 1467 1684 1523
rect 1740 1467 1808 1523
rect 1864 1467 1874 1523
rect 1426 1399 1874 1467
rect 1426 1343 1436 1399
rect 1492 1343 1560 1399
rect 1616 1343 1684 1399
rect 1740 1343 1808 1399
rect 1864 1343 1874 1399
rect 1426 1333 1874 1343
rect 2562 4251 3010 4261
rect 2562 4195 2572 4251
rect 2628 4195 2696 4251
rect 2752 4195 2820 4251
rect 2876 4195 2944 4251
rect 3000 4195 3010 4251
rect 2562 4127 3010 4195
rect 2562 4071 2572 4127
rect 2628 4071 2696 4127
rect 2752 4071 2820 4127
rect 2876 4071 2944 4127
rect 3000 4071 3010 4127
rect 2562 4003 3010 4071
rect 2562 3947 2572 4003
rect 2628 3947 2696 4003
rect 2752 3947 2820 4003
rect 2876 3947 2944 4003
rect 3000 3947 3010 4003
rect 2562 3879 3010 3947
rect 2562 3823 2572 3879
rect 2628 3823 2696 3879
rect 2752 3823 2820 3879
rect 2876 3823 2944 3879
rect 3000 3823 3010 3879
rect 2562 3755 3010 3823
rect 2562 3699 2572 3755
rect 2628 3699 2696 3755
rect 2752 3699 2820 3755
rect 2876 3699 2944 3755
rect 3000 3699 3010 3755
rect 2562 3631 3010 3699
rect 2562 3575 2572 3631
rect 2628 3575 2696 3631
rect 2752 3575 2820 3631
rect 2876 3575 2944 3631
rect 3000 3575 3010 3631
rect 2562 3507 3010 3575
rect 2562 3451 2572 3507
rect 2628 3451 2696 3507
rect 2752 3451 2820 3507
rect 2876 3451 2944 3507
rect 3000 3451 3010 3507
rect 2562 3383 3010 3451
rect 2562 3327 2572 3383
rect 2628 3327 2696 3383
rect 2752 3327 2820 3383
rect 2876 3327 2944 3383
rect 3000 3327 3010 3383
rect 2562 3259 3010 3327
rect 2562 3203 2572 3259
rect 2628 3203 2696 3259
rect 2752 3203 2820 3259
rect 2876 3203 2944 3259
rect 3000 3203 3010 3259
rect 2562 3135 3010 3203
rect 2562 3079 2572 3135
rect 2628 3079 2696 3135
rect 2752 3079 2820 3135
rect 2876 3079 2944 3135
rect 3000 3079 3010 3135
rect 2562 3011 3010 3079
rect 2562 2955 2572 3011
rect 2628 2955 2696 3011
rect 2752 2955 2820 3011
rect 2876 2955 2944 3011
rect 3000 2955 3010 3011
rect 2562 2887 3010 2955
rect 2562 2831 2572 2887
rect 2628 2831 2696 2887
rect 2752 2831 2820 2887
rect 2876 2831 2944 2887
rect 3000 2831 3010 2887
rect 2562 2763 3010 2831
rect 2562 2707 2572 2763
rect 2628 2707 2696 2763
rect 2752 2707 2820 2763
rect 2876 2707 2944 2763
rect 3000 2707 3010 2763
rect 2562 2639 3010 2707
rect 2562 2583 2572 2639
rect 2628 2583 2696 2639
rect 2752 2583 2820 2639
rect 2876 2583 2944 2639
rect 3000 2583 3010 2639
rect 2562 2515 3010 2583
rect 2562 2459 2572 2515
rect 2628 2459 2696 2515
rect 2752 2459 2820 2515
rect 2876 2459 2944 2515
rect 3000 2459 3010 2515
rect 2562 2391 3010 2459
rect 2562 2335 2572 2391
rect 2628 2335 2696 2391
rect 2752 2335 2820 2391
rect 2876 2335 2944 2391
rect 3000 2335 3010 2391
rect 2562 2267 3010 2335
rect 2562 2211 2572 2267
rect 2628 2211 2696 2267
rect 2752 2211 2820 2267
rect 2876 2211 2944 2267
rect 3000 2211 3010 2267
rect 2562 2143 3010 2211
rect 2562 2087 2572 2143
rect 2628 2087 2696 2143
rect 2752 2087 2820 2143
rect 2876 2087 2944 2143
rect 3000 2087 3010 2143
rect 2562 2019 3010 2087
rect 2562 1963 2572 2019
rect 2628 1963 2696 2019
rect 2752 1963 2820 2019
rect 2876 1963 2944 2019
rect 3000 1963 3010 2019
rect 2562 1895 3010 1963
rect 2562 1839 2572 1895
rect 2628 1839 2696 1895
rect 2752 1839 2820 1895
rect 2876 1839 2944 1895
rect 3000 1839 3010 1895
rect 2562 1771 3010 1839
rect 2562 1715 2572 1771
rect 2628 1715 2696 1771
rect 2752 1715 2820 1771
rect 2876 1715 2944 1771
rect 3000 1715 3010 1771
rect 2562 1647 3010 1715
rect 2562 1591 2572 1647
rect 2628 1591 2696 1647
rect 2752 1591 2820 1647
rect 2876 1591 2944 1647
rect 3000 1591 3010 1647
rect 2562 1523 3010 1591
rect 2562 1467 2572 1523
rect 2628 1467 2696 1523
rect 2752 1467 2820 1523
rect 2876 1467 2944 1523
rect 3000 1467 3010 1523
rect 2562 1399 3010 1467
rect 2562 1343 2572 1399
rect 2628 1343 2696 1399
rect 2752 1343 2820 1399
rect 2876 1343 2944 1399
rect 3000 1343 3010 1399
rect 2562 1333 3010 1343
rect 4834 4251 5282 4261
rect 4834 4195 4844 4251
rect 4900 4195 4968 4251
rect 5024 4195 5092 4251
rect 5148 4195 5216 4251
rect 5272 4195 5282 4251
rect 4834 4127 5282 4195
rect 4834 4071 4844 4127
rect 4900 4071 4968 4127
rect 5024 4071 5092 4127
rect 5148 4071 5216 4127
rect 5272 4071 5282 4127
rect 4834 4003 5282 4071
rect 4834 3947 4844 4003
rect 4900 3947 4968 4003
rect 5024 3947 5092 4003
rect 5148 3947 5216 4003
rect 5272 3947 5282 4003
rect 4834 3879 5282 3947
rect 4834 3823 4844 3879
rect 4900 3823 4968 3879
rect 5024 3823 5092 3879
rect 5148 3823 5216 3879
rect 5272 3823 5282 3879
rect 4834 3755 5282 3823
rect 4834 3699 4844 3755
rect 4900 3699 4968 3755
rect 5024 3699 5092 3755
rect 5148 3699 5216 3755
rect 5272 3699 5282 3755
rect 4834 3631 5282 3699
rect 4834 3575 4844 3631
rect 4900 3575 4968 3631
rect 5024 3575 5092 3631
rect 5148 3575 5216 3631
rect 5272 3575 5282 3631
rect 4834 3507 5282 3575
rect 4834 3451 4844 3507
rect 4900 3451 4968 3507
rect 5024 3451 5092 3507
rect 5148 3451 5216 3507
rect 5272 3451 5282 3507
rect 4834 3383 5282 3451
rect 4834 3327 4844 3383
rect 4900 3327 4968 3383
rect 5024 3327 5092 3383
rect 5148 3327 5216 3383
rect 5272 3327 5282 3383
rect 4834 3259 5282 3327
rect 4834 3203 4844 3259
rect 4900 3203 4968 3259
rect 5024 3203 5092 3259
rect 5148 3203 5216 3259
rect 5272 3203 5282 3259
rect 4834 3135 5282 3203
rect 4834 3079 4844 3135
rect 4900 3079 4968 3135
rect 5024 3079 5092 3135
rect 5148 3079 5216 3135
rect 5272 3079 5282 3135
rect 4834 3011 5282 3079
rect 4834 2955 4844 3011
rect 4900 2955 4968 3011
rect 5024 2955 5092 3011
rect 5148 2955 5216 3011
rect 5272 2955 5282 3011
rect 4834 2887 5282 2955
rect 4834 2831 4844 2887
rect 4900 2831 4968 2887
rect 5024 2831 5092 2887
rect 5148 2831 5216 2887
rect 5272 2831 5282 2887
rect 4834 2763 5282 2831
rect 4834 2707 4844 2763
rect 4900 2707 4968 2763
rect 5024 2707 5092 2763
rect 5148 2707 5216 2763
rect 5272 2707 5282 2763
rect 4834 2639 5282 2707
rect 4834 2583 4844 2639
rect 4900 2583 4968 2639
rect 5024 2583 5092 2639
rect 5148 2583 5216 2639
rect 5272 2583 5282 2639
rect 4834 2515 5282 2583
rect 4834 2459 4844 2515
rect 4900 2459 4968 2515
rect 5024 2459 5092 2515
rect 5148 2459 5216 2515
rect 5272 2459 5282 2515
rect 4834 2391 5282 2459
rect 4834 2335 4844 2391
rect 4900 2335 4968 2391
rect 5024 2335 5092 2391
rect 5148 2335 5216 2391
rect 5272 2335 5282 2391
rect 4834 2267 5282 2335
rect 4834 2211 4844 2267
rect 4900 2211 4968 2267
rect 5024 2211 5092 2267
rect 5148 2211 5216 2267
rect 5272 2211 5282 2267
rect 4834 2143 5282 2211
rect 4834 2087 4844 2143
rect 4900 2087 4968 2143
rect 5024 2087 5092 2143
rect 5148 2087 5216 2143
rect 5272 2087 5282 2143
rect 4834 2019 5282 2087
rect 4834 1963 4844 2019
rect 4900 1963 4968 2019
rect 5024 1963 5092 2019
rect 5148 1963 5216 2019
rect 5272 1963 5282 2019
rect 4834 1895 5282 1963
rect 4834 1839 4844 1895
rect 4900 1839 4968 1895
rect 5024 1839 5092 1895
rect 5148 1839 5216 1895
rect 5272 1839 5282 1895
rect 4834 1771 5282 1839
rect 4834 1715 4844 1771
rect 4900 1715 4968 1771
rect 5024 1715 5092 1771
rect 5148 1715 5216 1771
rect 5272 1715 5282 1771
rect 4834 1647 5282 1715
rect 4834 1591 4844 1647
rect 4900 1591 4968 1647
rect 5024 1591 5092 1647
rect 5148 1591 5216 1647
rect 5272 1591 5282 1647
rect 4834 1523 5282 1591
rect 4834 1467 4844 1523
rect 4900 1467 4968 1523
rect 5024 1467 5092 1523
rect 5148 1467 5216 1523
rect 5272 1467 5282 1523
rect 4834 1399 5282 1467
rect 4834 1343 4844 1399
rect 4900 1343 4968 1399
rect 5024 1343 5092 1399
rect 5148 1343 5216 1399
rect 5272 1343 5282 1399
rect 4834 1333 5282 1343
rect 7127 4251 7451 4261
rect 7127 4195 7137 4251
rect 7193 4195 7261 4251
rect 7317 4195 7385 4251
rect 7441 4195 7451 4251
rect 7127 4127 7451 4195
rect 7127 4071 7137 4127
rect 7193 4071 7261 4127
rect 7317 4071 7385 4127
rect 7441 4071 7451 4127
rect 7127 4003 7451 4071
rect 7127 3947 7137 4003
rect 7193 3947 7261 4003
rect 7317 3947 7385 4003
rect 7441 3947 7451 4003
rect 7127 3879 7451 3947
rect 7127 3823 7137 3879
rect 7193 3823 7261 3879
rect 7317 3823 7385 3879
rect 7441 3823 7451 3879
rect 7127 3755 7451 3823
rect 7127 3699 7137 3755
rect 7193 3699 7261 3755
rect 7317 3699 7385 3755
rect 7441 3699 7451 3755
rect 7127 3631 7451 3699
rect 7127 3575 7137 3631
rect 7193 3575 7261 3631
rect 7317 3575 7385 3631
rect 7441 3575 7451 3631
rect 7127 3507 7451 3575
rect 7127 3451 7137 3507
rect 7193 3451 7261 3507
rect 7317 3451 7385 3507
rect 7441 3451 7451 3507
rect 7127 3383 7451 3451
rect 7127 3327 7137 3383
rect 7193 3327 7261 3383
rect 7317 3327 7385 3383
rect 7441 3327 7451 3383
rect 7127 3259 7451 3327
rect 7127 3203 7137 3259
rect 7193 3203 7261 3259
rect 7317 3203 7385 3259
rect 7441 3203 7451 3259
rect 7127 3135 7451 3203
rect 7127 3079 7137 3135
rect 7193 3079 7261 3135
rect 7317 3079 7385 3135
rect 7441 3079 7451 3135
rect 7127 3011 7451 3079
rect 7127 2955 7137 3011
rect 7193 2955 7261 3011
rect 7317 2955 7385 3011
rect 7441 2955 7451 3011
rect 7127 2887 7451 2955
rect 7127 2831 7137 2887
rect 7193 2831 7261 2887
rect 7317 2831 7385 2887
rect 7441 2831 7451 2887
rect 7127 2763 7451 2831
rect 7127 2707 7137 2763
rect 7193 2707 7261 2763
rect 7317 2707 7385 2763
rect 7441 2707 7451 2763
rect 7127 2639 7451 2707
rect 7127 2583 7137 2639
rect 7193 2583 7261 2639
rect 7317 2583 7385 2639
rect 7441 2583 7451 2639
rect 7127 2515 7451 2583
rect 7127 2459 7137 2515
rect 7193 2459 7261 2515
rect 7317 2459 7385 2515
rect 7441 2459 7451 2515
rect 7127 2391 7451 2459
rect 7127 2335 7137 2391
rect 7193 2335 7261 2391
rect 7317 2335 7385 2391
rect 7441 2335 7451 2391
rect 7127 2267 7451 2335
rect 7127 2211 7137 2267
rect 7193 2211 7261 2267
rect 7317 2211 7385 2267
rect 7441 2211 7451 2267
rect 7127 2143 7451 2211
rect 7127 2087 7137 2143
rect 7193 2087 7261 2143
rect 7317 2087 7385 2143
rect 7441 2087 7451 2143
rect 7127 2019 7451 2087
rect 7127 1963 7137 2019
rect 7193 1963 7261 2019
rect 7317 1963 7385 2019
rect 7441 1963 7451 2019
rect 7127 1895 7451 1963
rect 7127 1839 7137 1895
rect 7193 1839 7261 1895
rect 7317 1839 7385 1895
rect 7441 1839 7451 1895
rect 7127 1771 7451 1839
rect 7127 1715 7137 1771
rect 7193 1715 7261 1771
rect 7317 1715 7385 1771
rect 7441 1715 7451 1771
rect 7127 1647 7451 1715
rect 7127 1591 7137 1647
rect 7193 1591 7261 1647
rect 7317 1591 7385 1647
rect 7441 1591 7451 1647
rect 7127 1523 7451 1591
rect 7127 1467 7137 1523
rect 7193 1467 7261 1523
rect 7317 1467 7385 1523
rect 7441 1467 7451 1523
rect 7127 1399 7451 1467
rect 7127 1343 7137 1399
rect 7193 1343 7261 1399
rect 7317 1343 7385 1399
rect 7441 1343 7451 1399
rect 7127 1333 7451 1343
rect 7613 4251 7937 4261
rect 7613 4195 7623 4251
rect 7679 4195 7747 4251
rect 7803 4195 7871 4251
rect 7927 4195 7937 4251
rect 7613 4127 7937 4195
rect 7613 4071 7623 4127
rect 7679 4071 7747 4127
rect 7803 4071 7871 4127
rect 7927 4071 7937 4127
rect 7613 4003 7937 4071
rect 7613 3947 7623 4003
rect 7679 3947 7747 4003
rect 7803 3947 7871 4003
rect 7927 3947 7937 4003
rect 7613 3879 7937 3947
rect 7613 3823 7623 3879
rect 7679 3823 7747 3879
rect 7803 3823 7871 3879
rect 7927 3823 7937 3879
rect 7613 3755 7937 3823
rect 7613 3699 7623 3755
rect 7679 3699 7747 3755
rect 7803 3699 7871 3755
rect 7927 3699 7937 3755
rect 7613 3631 7937 3699
rect 7613 3575 7623 3631
rect 7679 3575 7747 3631
rect 7803 3575 7871 3631
rect 7927 3575 7937 3631
rect 7613 3507 7937 3575
rect 7613 3451 7623 3507
rect 7679 3451 7747 3507
rect 7803 3451 7871 3507
rect 7927 3451 7937 3507
rect 7613 3383 7937 3451
rect 7613 3327 7623 3383
rect 7679 3327 7747 3383
rect 7803 3327 7871 3383
rect 7927 3327 7937 3383
rect 7613 3259 7937 3327
rect 7613 3203 7623 3259
rect 7679 3203 7747 3259
rect 7803 3203 7871 3259
rect 7927 3203 7937 3259
rect 7613 3135 7937 3203
rect 7613 3079 7623 3135
rect 7679 3079 7747 3135
rect 7803 3079 7871 3135
rect 7927 3079 7937 3135
rect 7613 3011 7937 3079
rect 7613 2955 7623 3011
rect 7679 2955 7747 3011
rect 7803 2955 7871 3011
rect 7927 2955 7937 3011
rect 7613 2887 7937 2955
rect 7613 2831 7623 2887
rect 7679 2831 7747 2887
rect 7803 2831 7871 2887
rect 7927 2831 7937 2887
rect 7613 2763 7937 2831
rect 7613 2707 7623 2763
rect 7679 2707 7747 2763
rect 7803 2707 7871 2763
rect 7927 2707 7937 2763
rect 7613 2639 7937 2707
rect 7613 2583 7623 2639
rect 7679 2583 7747 2639
rect 7803 2583 7871 2639
rect 7927 2583 7937 2639
rect 7613 2515 7937 2583
rect 7613 2459 7623 2515
rect 7679 2459 7747 2515
rect 7803 2459 7871 2515
rect 7927 2459 7937 2515
rect 7613 2391 7937 2459
rect 7613 2335 7623 2391
rect 7679 2335 7747 2391
rect 7803 2335 7871 2391
rect 7927 2335 7937 2391
rect 7613 2267 7937 2335
rect 7613 2211 7623 2267
rect 7679 2211 7747 2267
rect 7803 2211 7871 2267
rect 7927 2211 7937 2267
rect 7613 2143 7937 2211
rect 7613 2087 7623 2143
rect 7679 2087 7747 2143
rect 7803 2087 7871 2143
rect 7927 2087 7937 2143
rect 7613 2019 7937 2087
rect 7613 1963 7623 2019
rect 7679 1963 7747 2019
rect 7803 1963 7871 2019
rect 7927 1963 7937 2019
rect 7613 1895 7937 1963
rect 7613 1839 7623 1895
rect 7679 1839 7747 1895
rect 7803 1839 7871 1895
rect 7927 1839 7937 1895
rect 7613 1771 7937 1839
rect 7613 1715 7623 1771
rect 7679 1715 7747 1771
rect 7803 1715 7871 1771
rect 7927 1715 7937 1771
rect 7613 1647 7937 1715
rect 7613 1591 7623 1647
rect 7679 1591 7747 1647
rect 7803 1591 7871 1647
rect 7927 1591 7937 1647
rect 7613 1523 7937 1591
rect 7613 1467 7623 1523
rect 7679 1467 7747 1523
rect 7803 1467 7871 1523
rect 7927 1467 7937 1523
rect 7613 1399 7937 1467
rect 7613 1343 7623 1399
rect 7679 1343 7747 1399
rect 7803 1343 7871 1399
rect 7927 1343 7937 1399
rect 7613 1333 7937 1343
rect 9782 4251 10230 4261
rect 9782 4195 9792 4251
rect 9848 4195 9916 4251
rect 9972 4195 10040 4251
rect 10096 4195 10164 4251
rect 10220 4195 10230 4251
rect 9782 4127 10230 4195
rect 9782 4071 9792 4127
rect 9848 4071 9916 4127
rect 9972 4071 10040 4127
rect 10096 4071 10164 4127
rect 10220 4071 10230 4127
rect 9782 4003 10230 4071
rect 9782 3947 9792 4003
rect 9848 3947 9916 4003
rect 9972 3947 10040 4003
rect 10096 3947 10164 4003
rect 10220 3947 10230 4003
rect 9782 3879 10230 3947
rect 9782 3823 9792 3879
rect 9848 3823 9916 3879
rect 9972 3823 10040 3879
rect 10096 3823 10164 3879
rect 10220 3823 10230 3879
rect 9782 3755 10230 3823
rect 9782 3699 9792 3755
rect 9848 3699 9916 3755
rect 9972 3699 10040 3755
rect 10096 3699 10164 3755
rect 10220 3699 10230 3755
rect 9782 3631 10230 3699
rect 9782 3575 9792 3631
rect 9848 3575 9916 3631
rect 9972 3575 10040 3631
rect 10096 3575 10164 3631
rect 10220 3575 10230 3631
rect 9782 3507 10230 3575
rect 9782 3451 9792 3507
rect 9848 3451 9916 3507
rect 9972 3451 10040 3507
rect 10096 3451 10164 3507
rect 10220 3451 10230 3507
rect 9782 3383 10230 3451
rect 9782 3327 9792 3383
rect 9848 3327 9916 3383
rect 9972 3327 10040 3383
rect 10096 3327 10164 3383
rect 10220 3327 10230 3383
rect 9782 3259 10230 3327
rect 9782 3203 9792 3259
rect 9848 3203 9916 3259
rect 9972 3203 10040 3259
rect 10096 3203 10164 3259
rect 10220 3203 10230 3259
rect 9782 3135 10230 3203
rect 9782 3079 9792 3135
rect 9848 3079 9916 3135
rect 9972 3079 10040 3135
rect 10096 3079 10164 3135
rect 10220 3079 10230 3135
rect 9782 3011 10230 3079
rect 9782 2955 9792 3011
rect 9848 2955 9916 3011
rect 9972 2955 10040 3011
rect 10096 2955 10164 3011
rect 10220 2955 10230 3011
rect 9782 2887 10230 2955
rect 9782 2831 9792 2887
rect 9848 2831 9916 2887
rect 9972 2831 10040 2887
rect 10096 2831 10164 2887
rect 10220 2831 10230 2887
rect 9782 2763 10230 2831
rect 9782 2707 9792 2763
rect 9848 2707 9916 2763
rect 9972 2707 10040 2763
rect 10096 2707 10164 2763
rect 10220 2707 10230 2763
rect 9782 2639 10230 2707
rect 9782 2583 9792 2639
rect 9848 2583 9916 2639
rect 9972 2583 10040 2639
rect 10096 2583 10164 2639
rect 10220 2583 10230 2639
rect 9782 2515 10230 2583
rect 9782 2459 9792 2515
rect 9848 2459 9916 2515
rect 9972 2459 10040 2515
rect 10096 2459 10164 2515
rect 10220 2459 10230 2515
rect 9782 2391 10230 2459
rect 9782 2335 9792 2391
rect 9848 2335 9916 2391
rect 9972 2335 10040 2391
rect 10096 2335 10164 2391
rect 10220 2335 10230 2391
rect 9782 2267 10230 2335
rect 9782 2211 9792 2267
rect 9848 2211 9916 2267
rect 9972 2211 10040 2267
rect 10096 2211 10164 2267
rect 10220 2211 10230 2267
rect 9782 2143 10230 2211
rect 9782 2087 9792 2143
rect 9848 2087 9916 2143
rect 9972 2087 10040 2143
rect 10096 2087 10164 2143
rect 10220 2087 10230 2143
rect 9782 2019 10230 2087
rect 9782 1963 9792 2019
rect 9848 1963 9916 2019
rect 9972 1963 10040 2019
rect 10096 1963 10164 2019
rect 10220 1963 10230 2019
rect 9782 1895 10230 1963
rect 9782 1839 9792 1895
rect 9848 1839 9916 1895
rect 9972 1839 10040 1895
rect 10096 1839 10164 1895
rect 10220 1839 10230 1895
rect 9782 1771 10230 1839
rect 9782 1715 9792 1771
rect 9848 1715 9916 1771
rect 9972 1715 10040 1771
rect 10096 1715 10164 1771
rect 10220 1715 10230 1771
rect 9782 1647 10230 1715
rect 9782 1591 9792 1647
rect 9848 1591 9916 1647
rect 9972 1591 10040 1647
rect 10096 1591 10164 1647
rect 10220 1591 10230 1647
rect 9782 1523 10230 1591
rect 9782 1467 9792 1523
rect 9848 1467 9916 1523
rect 9972 1467 10040 1523
rect 10096 1467 10164 1523
rect 10220 1467 10230 1523
rect 9782 1399 10230 1467
rect 9782 1343 9792 1399
rect 9848 1343 9916 1399
rect 9972 1343 10040 1399
rect 10096 1343 10164 1399
rect 10220 1343 10230 1399
rect 9782 1333 10230 1343
rect 12054 4251 12502 4261
rect 12054 4195 12064 4251
rect 12120 4195 12188 4251
rect 12244 4195 12312 4251
rect 12368 4195 12436 4251
rect 12492 4195 12502 4251
rect 12054 4127 12502 4195
rect 12054 4071 12064 4127
rect 12120 4071 12188 4127
rect 12244 4071 12312 4127
rect 12368 4071 12436 4127
rect 12492 4071 12502 4127
rect 12054 4003 12502 4071
rect 12054 3947 12064 4003
rect 12120 3947 12188 4003
rect 12244 3947 12312 4003
rect 12368 3947 12436 4003
rect 12492 3947 12502 4003
rect 12054 3879 12502 3947
rect 12054 3823 12064 3879
rect 12120 3823 12188 3879
rect 12244 3823 12312 3879
rect 12368 3823 12436 3879
rect 12492 3823 12502 3879
rect 12054 3755 12502 3823
rect 12054 3699 12064 3755
rect 12120 3699 12188 3755
rect 12244 3699 12312 3755
rect 12368 3699 12436 3755
rect 12492 3699 12502 3755
rect 12054 3631 12502 3699
rect 12054 3575 12064 3631
rect 12120 3575 12188 3631
rect 12244 3575 12312 3631
rect 12368 3575 12436 3631
rect 12492 3575 12502 3631
rect 12054 3507 12502 3575
rect 12054 3451 12064 3507
rect 12120 3451 12188 3507
rect 12244 3451 12312 3507
rect 12368 3451 12436 3507
rect 12492 3451 12502 3507
rect 12054 3383 12502 3451
rect 12054 3327 12064 3383
rect 12120 3327 12188 3383
rect 12244 3327 12312 3383
rect 12368 3327 12436 3383
rect 12492 3327 12502 3383
rect 12054 3259 12502 3327
rect 12054 3203 12064 3259
rect 12120 3203 12188 3259
rect 12244 3203 12312 3259
rect 12368 3203 12436 3259
rect 12492 3203 12502 3259
rect 12054 3135 12502 3203
rect 12054 3079 12064 3135
rect 12120 3079 12188 3135
rect 12244 3079 12312 3135
rect 12368 3079 12436 3135
rect 12492 3079 12502 3135
rect 12054 3011 12502 3079
rect 12054 2955 12064 3011
rect 12120 2955 12188 3011
rect 12244 2955 12312 3011
rect 12368 2955 12436 3011
rect 12492 2955 12502 3011
rect 12054 2887 12502 2955
rect 12054 2831 12064 2887
rect 12120 2831 12188 2887
rect 12244 2831 12312 2887
rect 12368 2831 12436 2887
rect 12492 2831 12502 2887
rect 12054 2763 12502 2831
rect 12054 2707 12064 2763
rect 12120 2707 12188 2763
rect 12244 2707 12312 2763
rect 12368 2707 12436 2763
rect 12492 2707 12502 2763
rect 12054 2639 12502 2707
rect 12054 2583 12064 2639
rect 12120 2583 12188 2639
rect 12244 2583 12312 2639
rect 12368 2583 12436 2639
rect 12492 2583 12502 2639
rect 12054 2515 12502 2583
rect 12054 2459 12064 2515
rect 12120 2459 12188 2515
rect 12244 2459 12312 2515
rect 12368 2459 12436 2515
rect 12492 2459 12502 2515
rect 12054 2391 12502 2459
rect 12054 2335 12064 2391
rect 12120 2335 12188 2391
rect 12244 2335 12312 2391
rect 12368 2335 12436 2391
rect 12492 2335 12502 2391
rect 12054 2267 12502 2335
rect 12054 2211 12064 2267
rect 12120 2211 12188 2267
rect 12244 2211 12312 2267
rect 12368 2211 12436 2267
rect 12492 2211 12502 2267
rect 12054 2143 12502 2211
rect 12054 2087 12064 2143
rect 12120 2087 12188 2143
rect 12244 2087 12312 2143
rect 12368 2087 12436 2143
rect 12492 2087 12502 2143
rect 12054 2019 12502 2087
rect 12054 1963 12064 2019
rect 12120 1963 12188 2019
rect 12244 1963 12312 2019
rect 12368 1963 12436 2019
rect 12492 1963 12502 2019
rect 12054 1895 12502 1963
rect 12054 1839 12064 1895
rect 12120 1839 12188 1895
rect 12244 1839 12312 1895
rect 12368 1839 12436 1895
rect 12492 1839 12502 1895
rect 12054 1771 12502 1839
rect 12054 1715 12064 1771
rect 12120 1715 12188 1771
rect 12244 1715 12312 1771
rect 12368 1715 12436 1771
rect 12492 1715 12502 1771
rect 12054 1647 12502 1715
rect 12054 1591 12064 1647
rect 12120 1591 12188 1647
rect 12244 1591 12312 1647
rect 12368 1591 12436 1647
rect 12492 1591 12502 1647
rect 12054 1523 12502 1591
rect 12054 1467 12064 1523
rect 12120 1467 12188 1523
rect 12244 1467 12312 1523
rect 12368 1467 12436 1523
rect 12492 1467 12502 1523
rect 12054 1399 12502 1467
rect 12054 1343 12064 1399
rect 12120 1343 12188 1399
rect 12244 1343 12312 1399
rect 12368 1343 12436 1399
rect 12492 1343 12502 1399
rect 12054 1333 12502 1343
rect 13190 4251 13638 4261
rect 13190 4195 13200 4251
rect 13256 4195 13324 4251
rect 13380 4195 13448 4251
rect 13504 4195 13572 4251
rect 13628 4195 13638 4251
rect 13190 4127 13638 4195
rect 13190 4071 13200 4127
rect 13256 4071 13324 4127
rect 13380 4071 13448 4127
rect 13504 4071 13572 4127
rect 13628 4071 13638 4127
rect 13190 4003 13638 4071
rect 13190 3947 13200 4003
rect 13256 3947 13324 4003
rect 13380 3947 13448 4003
rect 13504 3947 13572 4003
rect 13628 3947 13638 4003
rect 13190 3879 13638 3947
rect 13190 3823 13200 3879
rect 13256 3823 13324 3879
rect 13380 3823 13448 3879
rect 13504 3823 13572 3879
rect 13628 3823 13638 3879
rect 13190 3755 13638 3823
rect 13190 3699 13200 3755
rect 13256 3699 13324 3755
rect 13380 3699 13448 3755
rect 13504 3699 13572 3755
rect 13628 3699 13638 3755
rect 13190 3631 13638 3699
rect 13190 3575 13200 3631
rect 13256 3575 13324 3631
rect 13380 3575 13448 3631
rect 13504 3575 13572 3631
rect 13628 3575 13638 3631
rect 13190 3507 13638 3575
rect 13190 3451 13200 3507
rect 13256 3451 13324 3507
rect 13380 3451 13448 3507
rect 13504 3451 13572 3507
rect 13628 3451 13638 3507
rect 13190 3383 13638 3451
rect 13190 3327 13200 3383
rect 13256 3327 13324 3383
rect 13380 3327 13448 3383
rect 13504 3327 13572 3383
rect 13628 3327 13638 3383
rect 13190 3259 13638 3327
rect 13190 3203 13200 3259
rect 13256 3203 13324 3259
rect 13380 3203 13448 3259
rect 13504 3203 13572 3259
rect 13628 3203 13638 3259
rect 13190 3135 13638 3203
rect 13190 3079 13200 3135
rect 13256 3079 13324 3135
rect 13380 3079 13448 3135
rect 13504 3079 13572 3135
rect 13628 3079 13638 3135
rect 13190 3011 13638 3079
rect 13190 2955 13200 3011
rect 13256 2955 13324 3011
rect 13380 2955 13448 3011
rect 13504 2955 13572 3011
rect 13628 2955 13638 3011
rect 13190 2887 13638 2955
rect 13190 2831 13200 2887
rect 13256 2831 13324 2887
rect 13380 2831 13448 2887
rect 13504 2831 13572 2887
rect 13628 2831 13638 2887
rect 13190 2763 13638 2831
rect 13190 2707 13200 2763
rect 13256 2707 13324 2763
rect 13380 2707 13448 2763
rect 13504 2707 13572 2763
rect 13628 2707 13638 2763
rect 13190 2639 13638 2707
rect 13190 2583 13200 2639
rect 13256 2583 13324 2639
rect 13380 2583 13448 2639
rect 13504 2583 13572 2639
rect 13628 2583 13638 2639
rect 13190 2515 13638 2583
rect 13190 2459 13200 2515
rect 13256 2459 13324 2515
rect 13380 2459 13448 2515
rect 13504 2459 13572 2515
rect 13628 2459 13638 2515
rect 13190 2391 13638 2459
rect 13190 2335 13200 2391
rect 13256 2335 13324 2391
rect 13380 2335 13448 2391
rect 13504 2335 13572 2391
rect 13628 2335 13638 2391
rect 13190 2267 13638 2335
rect 13190 2211 13200 2267
rect 13256 2211 13324 2267
rect 13380 2211 13448 2267
rect 13504 2211 13572 2267
rect 13628 2211 13638 2267
rect 13190 2143 13638 2211
rect 13190 2087 13200 2143
rect 13256 2087 13324 2143
rect 13380 2087 13448 2143
rect 13504 2087 13572 2143
rect 13628 2087 13638 2143
rect 13190 2019 13638 2087
rect 13190 1963 13200 2019
rect 13256 1963 13324 2019
rect 13380 1963 13448 2019
rect 13504 1963 13572 2019
rect 13628 1963 13638 2019
rect 13190 1895 13638 1963
rect 13190 1839 13200 1895
rect 13256 1839 13324 1895
rect 13380 1839 13448 1895
rect 13504 1839 13572 1895
rect 13628 1839 13638 1895
rect 13190 1771 13638 1839
rect 13190 1715 13200 1771
rect 13256 1715 13324 1771
rect 13380 1715 13448 1771
rect 13504 1715 13572 1771
rect 13628 1715 13638 1771
rect 13190 1647 13638 1715
rect 13190 1591 13200 1647
rect 13256 1591 13324 1647
rect 13380 1591 13448 1647
rect 13504 1591 13572 1647
rect 13628 1591 13638 1647
rect 13190 1523 13638 1591
rect 13190 1467 13200 1523
rect 13256 1467 13324 1523
rect 13380 1467 13448 1523
rect 13504 1467 13572 1523
rect 13628 1467 13638 1523
rect 13190 1399 13638 1467
rect 13190 1343 13200 1399
rect 13256 1343 13324 1399
rect 13380 1343 13448 1399
rect 13504 1343 13572 1399
rect 13628 1343 13638 1399
rect 13190 1333 13638 1343
rect 13728 900 14236 10949
rect 14296 56922 14804 56975
rect 14296 56866 14336 56922
rect 14392 56866 14460 56922
rect 14516 56866 14584 56922
rect 14640 56866 14708 56922
rect 14764 56866 14804 56922
rect 14296 56798 14804 56866
rect 14296 56742 14336 56798
rect 14392 56742 14460 56798
rect 14516 56742 14584 56798
rect 14640 56742 14708 56798
rect 14764 56742 14804 56798
rect 14296 56711 14804 56742
rect 14296 56674 14352 56711
rect 14296 56618 14336 56674
rect 14404 56659 14460 56711
rect 14512 56674 14568 56711
rect 14620 56674 14804 56711
rect 14516 56659 14568 56674
rect 14392 56618 14460 56659
rect 14516 56618 14584 56659
rect 14640 56618 14708 56674
rect 14764 56618 14804 56674
rect 14296 56603 14804 56618
rect 14296 56551 14352 56603
rect 14404 56551 14460 56603
rect 14512 56551 14568 56603
rect 14620 56551 14804 56603
rect 14296 56550 14804 56551
rect 14296 56494 14336 56550
rect 14392 56495 14460 56550
rect 14516 56495 14584 56550
rect 14296 56443 14352 56494
rect 14404 56443 14460 56495
rect 14516 56494 14568 56495
rect 14640 56494 14708 56550
rect 14764 56494 14804 56550
rect 14512 56443 14568 56494
rect 14620 56443 14804 56494
rect 14296 56426 14804 56443
rect 14296 56370 14336 56426
rect 14392 56370 14460 56426
rect 14516 56370 14584 56426
rect 14640 56370 14708 56426
rect 14764 56370 14804 56426
rect 14296 56302 14804 56370
rect 14296 56246 14336 56302
rect 14392 56246 14460 56302
rect 14516 56246 14584 56302
rect 14640 56246 14708 56302
rect 14764 56246 14804 56302
rect 14296 56178 14804 56246
rect 14296 56122 14336 56178
rect 14392 56122 14460 56178
rect 14516 56122 14584 56178
rect 14640 56122 14708 56178
rect 14764 56122 14804 56178
rect 14296 56054 14804 56122
rect 14296 55998 14336 56054
rect 14392 55998 14460 56054
rect 14516 55998 14584 56054
rect 14640 55998 14708 56054
rect 14764 55998 14804 56054
rect 14296 55930 14804 55998
rect 14296 55874 14336 55930
rect 14392 55874 14460 55930
rect 14516 55874 14584 55930
rect 14640 55874 14708 55930
rect 14764 55874 14804 55930
rect 14296 55806 14804 55874
rect 14296 55750 14336 55806
rect 14392 55750 14460 55806
rect 14516 55750 14584 55806
rect 14640 55750 14708 55806
rect 14764 55750 14804 55806
rect 14296 53845 14804 55750
rect 14296 53789 14336 53845
rect 14392 53789 14460 53845
rect 14516 53789 14584 53845
rect 14640 53789 14708 53845
rect 14764 53789 14804 53845
rect 14296 53721 14804 53789
rect 14296 53665 14336 53721
rect 14392 53665 14460 53721
rect 14516 53665 14584 53721
rect 14640 53665 14708 53721
rect 14764 53665 14804 53721
rect 14296 53597 14804 53665
rect 14296 53541 14336 53597
rect 14392 53541 14460 53597
rect 14516 53541 14584 53597
rect 14640 53541 14708 53597
rect 14764 53541 14804 53597
rect 14296 53473 14804 53541
rect 14296 53417 14336 53473
rect 14392 53417 14460 53473
rect 14516 53417 14584 53473
rect 14640 53417 14708 53473
rect 14764 53417 14804 53473
rect 14296 53349 14804 53417
rect 14296 53293 14336 53349
rect 14392 53293 14460 53349
rect 14516 53293 14584 53349
rect 14640 53293 14708 53349
rect 14764 53293 14804 53349
rect 14296 53225 14804 53293
rect 14296 53169 14336 53225
rect 14392 53169 14460 53225
rect 14516 53169 14584 53225
rect 14640 53169 14708 53225
rect 14764 53169 14804 53225
rect 14296 53101 14804 53169
rect 14296 53045 14336 53101
rect 14392 53045 14460 53101
rect 14516 53045 14584 53101
rect 14640 53045 14708 53101
rect 14764 53045 14804 53101
rect 14296 53016 14804 53045
rect 14296 52977 14352 53016
rect 14296 52921 14336 52977
rect 14404 52964 14460 53016
rect 14512 52977 14568 53016
rect 14620 52977 14804 53016
rect 14516 52964 14568 52977
rect 14392 52921 14460 52964
rect 14516 52921 14584 52964
rect 14640 52921 14708 52977
rect 14764 52921 14804 52977
rect 14296 52908 14804 52921
rect 14296 52856 14352 52908
rect 14404 52856 14460 52908
rect 14512 52856 14568 52908
rect 14620 52856 14804 52908
rect 14296 52853 14804 52856
rect 14296 52797 14336 52853
rect 14392 52800 14460 52853
rect 14516 52800 14584 52853
rect 14296 52748 14352 52797
rect 14404 52748 14460 52800
rect 14516 52797 14568 52800
rect 14640 52797 14708 52853
rect 14764 52797 14804 52853
rect 14512 52748 14568 52797
rect 14620 52748 14804 52797
rect 14296 52729 14804 52748
rect 14296 52673 14336 52729
rect 14392 52692 14460 52729
rect 14516 52692 14584 52729
rect 14296 52640 14352 52673
rect 14404 52640 14460 52692
rect 14516 52673 14568 52692
rect 14640 52673 14708 52729
rect 14764 52673 14804 52729
rect 14512 52640 14568 52673
rect 14620 52640 14804 52673
rect 14296 52605 14804 52640
rect 14296 52549 14336 52605
rect 14392 52584 14460 52605
rect 14516 52584 14584 52605
rect 14296 52532 14352 52549
rect 14404 52532 14460 52584
rect 14516 52549 14568 52584
rect 14640 52549 14708 52605
rect 14764 52549 14804 52605
rect 14512 52532 14568 52549
rect 14620 52532 14804 52549
rect 14296 49068 14804 52532
rect 14942 52273 15032 52297
rect 14942 50921 14952 52273
rect 15008 50921 15032 52273
rect 14942 50897 15032 50921
rect 14296 49045 14352 49068
rect 14296 48989 14336 49045
rect 14404 49016 14460 49068
rect 14512 49045 14568 49068
rect 14620 49045 14804 49068
rect 14516 49016 14568 49045
rect 14392 48989 14460 49016
rect 14516 48989 14584 49016
rect 14640 48989 14708 49045
rect 14764 48989 14804 49045
rect 14296 48960 14804 48989
rect 14296 48921 14352 48960
rect 14296 48865 14336 48921
rect 14404 48908 14460 48960
rect 14512 48921 14568 48960
rect 14620 48921 14804 48960
rect 14516 48908 14568 48921
rect 14392 48865 14460 48908
rect 14516 48865 14584 48908
rect 14640 48865 14708 48921
rect 14764 48865 14804 48921
rect 14296 48852 14804 48865
rect 14296 48800 14352 48852
rect 14404 48800 14460 48852
rect 14512 48800 14568 48852
rect 14620 48800 14804 48852
rect 14296 48797 14804 48800
rect 14296 48741 14336 48797
rect 14392 48744 14460 48797
rect 14516 48744 14584 48797
rect 14296 48692 14352 48741
rect 14404 48692 14460 48744
rect 14516 48741 14568 48744
rect 14640 48741 14708 48797
rect 14764 48741 14804 48797
rect 14512 48692 14568 48741
rect 14620 48692 14804 48741
rect 14296 48673 14804 48692
rect 14296 48617 14336 48673
rect 14392 48636 14460 48673
rect 14516 48636 14584 48673
rect 14296 48584 14352 48617
rect 14404 48584 14460 48636
rect 14516 48617 14568 48636
rect 14640 48617 14708 48673
rect 14764 48617 14804 48673
rect 14512 48584 14568 48617
rect 14620 48584 14804 48617
rect 14296 48549 14804 48584
rect 14296 48493 14336 48549
rect 14392 48493 14460 48549
rect 14516 48493 14584 48549
rect 14640 48493 14708 48549
rect 14764 48493 14804 48549
rect 14296 48425 14804 48493
rect 14296 48369 14336 48425
rect 14392 48369 14460 48425
rect 14516 48369 14584 48425
rect 14640 48369 14708 48425
rect 14764 48369 14804 48425
rect 14296 48301 14804 48369
rect 14296 48245 14336 48301
rect 14392 48245 14460 48301
rect 14516 48245 14584 48301
rect 14640 48245 14708 48301
rect 14764 48245 14804 48301
rect 14296 48177 14804 48245
rect 14296 48121 14336 48177
rect 14392 48121 14460 48177
rect 14516 48121 14584 48177
rect 14640 48121 14708 48177
rect 14764 48121 14804 48177
rect 14296 48053 14804 48121
rect 14296 47997 14336 48053
rect 14392 47997 14460 48053
rect 14516 47997 14584 48053
rect 14640 47997 14708 48053
rect 14764 47997 14804 48053
rect 14296 47929 14804 47997
rect 14296 47873 14336 47929
rect 14392 47873 14460 47929
rect 14516 47873 14584 47929
rect 14640 47873 14708 47929
rect 14764 47873 14804 47929
rect 14296 47805 14804 47873
rect 14296 47749 14336 47805
rect 14392 47749 14460 47805
rect 14516 47749 14584 47805
rect 14640 47749 14708 47805
rect 14764 47749 14804 47805
rect 14296 45845 14804 47749
rect 14296 45789 14336 45845
rect 14392 45789 14460 45845
rect 14516 45789 14584 45845
rect 14640 45789 14708 45845
rect 14764 45789 14804 45845
rect 14296 45721 14804 45789
rect 14296 45665 14336 45721
rect 14392 45665 14460 45721
rect 14516 45665 14584 45721
rect 14640 45665 14708 45721
rect 14764 45665 14804 45721
rect 14296 45597 14804 45665
rect 14296 45541 14336 45597
rect 14392 45541 14460 45597
rect 14516 45541 14584 45597
rect 14640 45541 14708 45597
rect 14764 45541 14804 45597
rect 14296 45473 14804 45541
rect 14296 45417 14336 45473
rect 14392 45417 14460 45473
rect 14516 45417 14584 45473
rect 14640 45417 14708 45473
rect 14764 45417 14804 45473
rect 14296 45349 14804 45417
rect 14296 45293 14336 45349
rect 14392 45293 14460 45349
rect 14516 45293 14584 45349
rect 14640 45293 14708 45349
rect 14764 45293 14804 45349
rect 14296 45225 14804 45293
rect 14296 45169 14336 45225
rect 14392 45169 14460 45225
rect 14516 45169 14584 45225
rect 14640 45169 14708 45225
rect 14764 45169 14804 45225
rect 14296 45120 14804 45169
rect 14296 45101 14352 45120
rect 14296 45045 14336 45101
rect 14404 45068 14460 45120
rect 14512 45101 14568 45120
rect 14620 45101 14804 45120
rect 14516 45068 14568 45101
rect 14392 45045 14460 45068
rect 14516 45045 14584 45068
rect 14640 45045 14708 45101
rect 14764 45045 14804 45101
rect 14296 45012 14804 45045
rect 14296 44977 14352 45012
rect 14296 44921 14336 44977
rect 14404 44960 14460 45012
rect 14512 44977 14568 45012
rect 14620 44977 14804 45012
rect 14516 44960 14568 44977
rect 14392 44921 14460 44960
rect 14516 44921 14584 44960
rect 14640 44921 14708 44977
rect 14764 44921 14804 44977
rect 14296 44904 14804 44921
rect 14296 44853 14352 44904
rect 14296 44797 14336 44853
rect 14404 44852 14460 44904
rect 14512 44853 14568 44904
rect 14620 44853 14804 44904
rect 14516 44852 14568 44853
rect 14392 44797 14460 44852
rect 14516 44797 14584 44852
rect 14640 44797 14708 44853
rect 14764 44797 14804 44853
rect 14296 44796 14804 44797
rect 14296 44744 14352 44796
rect 14404 44744 14460 44796
rect 14512 44744 14568 44796
rect 14620 44744 14804 44796
rect 14296 44729 14804 44744
rect 14296 44673 14336 44729
rect 14392 44688 14460 44729
rect 14516 44688 14584 44729
rect 14296 44636 14352 44673
rect 14404 44636 14460 44688
rect 14516 44673 14568 44688
rect 14640 44673 14708 44729
rect 14764 44673 14804 44729
rect 14512 44636 14568 44673
rect 14620 44636 14804 44673
rect 14296 44605 14804 44636
rect 14296 44549 14336 44605
rect 14392 44549 14460 44605
rect 14516 44549 14584 44605
rect 14640 44549 14708 44605
rect 14764 44549 14804 44605
rect 14296 41172 14804 44549
rect 14296 41120 14352 41172
rect 14404 41120 14460 41172
rect 14512 41120 14568 41172
rect 14620 41120 14804 41172
rect 14296 41064 14804 41120
rect 14296 41012 14352 41064
rect 14404 41012 14460 41064
rect 14512 41012 14568 41064
rect 14620 41012 14804 41064
rect 14296 40956 14804 41012
rect 14296 40904 14352 40956
rect 14404 40904 14460 40956
rect 14512 40904 14568 40956
rect 14620 40904 14804 40956
rect 14296 40848 14804 40904
rect 14296 40796 14352 40848
rect 14404 40796 14460 40848
rect 14512 40796 14568 40848
rect 14620 40796 14804 40848
rect 14296 40740 14804 40796
rect 14296 40688 14352 40740
rect 14404 40688 14460 40740
rect 14512 40688 14568 40740
rect 14620 40688 14804 40740
rect 14296 37224 14804 40688
rect 14296 37172 14352 37224
rect 14404 37172 14460 37224
rect 14512 37172 14568 37224
rect 14620 37172 14804 37224
rect 14296 37116 14804 37172
rect 14296 37064 14352 37116
rect 14404 37064 14460 37116
rect 14512 37064 14568 37116
rect 14620 37064 14804 37116
rect 14296 37008 14804 37064
rect 14296 36956 14352 37008
rect 14404 36956 14460 37008
rect 14512 36956 14568 37008
rect 14620 36956 14804 37008
rect 14296 36900 14804 36956
rect 14296 36848 14352 36900
rect 14404 36848 14460 36900
rect 14512 36848 14568 36900
rect 14620 36848 14804 36900
rect 14296 36792 14804 36848
rect 14296 36740 14352 36792
rect 14404 36740 14460 36792
rect 14512 36740 14568 36792
rect 14620 36740 14804 36792
rect 14296 36251 14804 36740
rect 14942 37873 15032 37897
rect 14942 36521 14952 37873
rect 15008 36521 15032 37873
rect 14942 36497 15032 36521
rect 14296 36195 14336 36251
rect 14392 36195 14460 36251
rect 14516 36195 14584 36251
rect 14640 36195 14708 36251
rect 14764 36195 14804 36251
rect 14296 36127 14804 36195
rect 14296 36071 14336 36127
rect 14392 36071 14460 36127
rect 14516 36071 14584 36127
rect 14640 36071 14708 36127
rect 14764 36071 14804 36127
rect 14296 36003 14804 36071
rect 14296 35947 14336 36003
rect 14392 35947 14460 36003
rect 14516 35947 14584 36003
rect 14640 35947 14708 36003
rect 14764 35947 14804 36003
rect 14296 35879 14804 35947
rect 14296 35823 14336 35879
rect 14392 35823 14460 35879
rect 14516 35823 14584 35879
rect 14640 35823 14708 35879
rect 14764 35823 14804 35879
rect 14296 35755 14804 35823
rect 14296 35699 14336 35755
rect 14392 35699 14460 35755
rect 14516 35699 14584 35755
rect 14640 35699 14708 35755
rect 14764 35699 14804 35755
rect 14296 35631 14804 35699
rect 14296 35575 14336 35631
rect 14392 35575 14460 35631
rect 14516 35575 14584 35631
rect 14640 35575 14708 35631
rect 14764 35575 14804 35631
rect 14296 35507 14804 35575
rect 14296 35451 14336 35507
rect 14392 35451 14460 35507
rect 14516 35451 14584 35507
rect 14640 35451 14708 35507
rect 14764 35451 14804 35507
rect 14296 35383 14804 35451
rect 14296 35327 14336 35383
rect 14392 35327 14460 35383
rect 14516 35327 14584 35383
rect 14640 35327 14708 35383
rect 14764 35327 14804 35383
rect 14296 35259 14804 35327
rect 14296 35203 14336 35259
rect 14392 35203 14460 35259
rect 14516 35203 14584 35259
rect 14640 35203 14708 35259
rect 14764 35203 14804 35259
rect 14296 35135 14804 35203
rect 14296 35079 14336 35135
rect 14392 35079 14460 35135
rect 14516 35079 14584 35135
rect 14640 35079 14708 35135
rect 14764 35079 14804 35135
rect 14296 35011 14804 35079
rect 14296 34955 14336 35011
rect 14392 34955 14460 35011
rect 14516 34955 14584 35011
rect 14640 34955 14708 35011
rect 14764 34955 14804 35011
rect 14296 34887 14804 34955
rect 14296 34831 14336 34887
rect 14392 34831 14460 34887
rect 14516 34831 14584 34887
rect 14640 34831 14708 34887
rect 14764 34831 14804 34887
rect 14296 34763 14804 34831
rect 14296 34707 14336 34763
rect 14392 34707 14460 34763
rect 14516 34707 14584 34763
rect 14640 34707 14708 34763
rect 14764 34707 14804 34763
rect 14296 34639 14804 34707
rect 14296 34583 14336 34639
rect 14392 34583 14460 34639
rect 14516 34583 14584 34639
rect 14640 34583 14708 34639
rect 14764 34583 14804 34639
rect 14296 34515 14804 34583
rect 14296 34459 14336 34515
rect 14392 34459 14460 34515
rect 14516 34459 14584 34515
rect 14640 34459 14708 34515
rect 14764 34459 14804 34515
rect 14296 34391 14804 34459
rect 14296 34335 14336 34391
rect 14392 34335 14460 34391
rect 14516 34335 14584 34391
rect 14640 34335 14708 34391
rect 14764 34335 14804 34391
rect 14296 34267 14804 34335
rect 14296 34211 14336 34267
rect 14392 34211 14460 34267
rect 14516 34211 14584 34267
rect 14640 34211 14708 34267
rect 14764 34211 14804 34267
rect 14296 34143 14804 34211
rect 14296 34087 14336 34143
rect 14392 34087 14460 34143
rect 14516 34087 14584 34143
rect 14640 34087 14708 34143
rect 14764 34087 14804 34143
rect 14296 34019 14804 34087
rect 14296 33963 14336 34019
rect 14392 33963 14460 34019
rect 14516 33963 14584 34019
rect 14640 33963 14708 34019
rect 14764 33963 14804 34019
rect 14296 33895 14804 33963
rect 14296 33839 14336 33895
rect 14392 33839 14460 33895
rect 14516 33839 14584 33895
rect 14640 33839 14708 33895
rect 14764 33839 14804 33895
rect 14296 33771 14804 33839
rect 14296 33715 14336 33771
rect 14392 33715 14460 33771
rect 14516 33715 14584 33771
rect 14640 33715 14708 33771
rect 14764 33715 14804 33771
rect 14296 33647 14804 33715
rect 14296 33591 14336 33647
rect 14392 33591 14460 33647
rect 14516 33591 14584 33647
rect 14640 33591 14708 33647
rect 14764 33591 14804 33647
rect 14296 33523 14804 33591
rect 14296 33467 14336 33523
rect 14392 33467 14460 33523
rect 14516 33467 14584 33523
rect 14640 33467 14708 33523
rect 14764 33467 14804 33523
rect 14296 33399 14804 33467
rect 14296 33343 14336 33399
rect 14392 33343 14460 33399
rect 14516 33343 14584 33399
rect 14640 33343 14708 33399
rect 14764 33343 14804 33399
rect 14296 33276 14804 33343
rect 14296 33224 14352 33276
rect 14404 33224 14460 33276
rect 14512 33224 14568 33276
rect 14620 33224 14804 33276
rect 14296 33168 14804 33224
rect 14296 33116 14352 33168
rect 14404 33116 14460 33168
rect 14512 33116 14568 33168
rect 14620 33116 14804 33168
rect 14296 33060 14804 33116
rect 14296 33008 14352 33060
rect 14404 33008 14460 33060
rect 14512 33008 14568 33060
rect 14620 33008 14804 33060
rect 14296 32952 14804 33008
rect 14296 32900 14352 32952
rect 14404 32900 14460 32952
rect 14512 32900 14568 32952
rect 14620 32900 14804 32952
rect 14296 32844 14804 32900
rect 14296 32792 14352 32844
rect 14404 32792 14460 32844
rect 14512 32792 14568 32844
rect 14620 32792 14804 32844
rect 14296 29328 14804 32792
rect 14296 29276 14352 29328
rect 14404 29276 14460 29328
rect 14512 29276 14568 29328
rect 14620 29276 14804 29328
rect 14296 29220 14804 29276
rect 14296 29168 14352 29220
rect 14404 29168 14460 29220
rect 14512 29168 14568 29220
rect 14620 29168 14804 29220
rect 14296 29112 14804 29168
rect 14296 29060 14352 29112
rect 14404 29060 14460 29112
rect 14512 29060 14568 29112
rect 14620 29060 14804 29112
rect 14296 29004 14804 29060
rect 14296 28952 14352 29004
rect 14404 28952 14460 29004
rect 14512 28952 14568 29004
rect 14620 28952 14804 29004
rect 14296 28896 14804 28952
rect 14296 28844 14352 28896
rect 14404 28844 14460 28896
rect 14512 28844 14568 28896
rect 14620 28844 14804 28896
rect 14296 28245 14804 28844
rect 14296 28189 14336 28245
rect 14392 28189 14460 28245
rect 14516 28189 14584 28245
rect 14640 28189 14708 28245
rect 14764 28189 14804 28245
rect 14296 28121 14804 28189
rect 14296 28065 14336 28121
rect 14392 28065 14460 28121
rect 14516 28065 14584 28121
rect 14640 28065 14708 28121
rect 14764 28065 14804 28121
rect 14296 27997 14804 28065
rect 14296 27941 14336 27997
rect 14392 27941 14460 27997
rect 14516 27941 14584 27997
rect 14640 27941 14708 27997
rect 14764 27941 14804 27997
rect 14296 27873 14804 27941
rect 14296 27817 14336 27873
rect 14392 27817 14460 27873
rect 14516 27817 14584 27873
rect 14640 27817 14708 27873
rect 14764 27817 14804 27873
rect 14296 27749 14804 27817
rect 14296 27693 14336 27749
rect 14392 27693 14460 27749
rect 14516 27693 14584 27749
rect 14640 27693 14708 27749
rect 14764 27693 14804 27749
rect 14296 27625 14804 27693
rect 14296 27569 14336 27625
rect 14392 27569 14460 27625
rect 14516 27569 14584 27625
rect 14640 27569 14708 27625
rect 14764 27569 14804 27625
rect 14296 27501 14804 27569
rect 14296 27445 14336 27501
rect 14392 27445 14460 27501
rect 14516 27445 14584 27501
rect 14640 27445 14708 27501
rect 14764 27445 14804 27501
rect 14296 27377 14804 27445
rect 14296 27321 14336 27377
rect 14392 27321 14460 27377
rect 14516 27321 14584 27377
rect 14640 27321 14708 27377
rect 14764 27321 14804 27377
rect 14296 27253 14804 27321
rect 14296 27197 14336 27253
rect 14392 27197 14460 27253
rect 14516 27197 14584 27253
rect 14640 27197 14708 27253
rect 14764 27197 14804 27253
rect 14296 27129 14804 27197
rect 14296 27073 14336 27129
rect 14392 27073 14460 27129
rect 14516 27073 14584 27129
rect 14640 27073 14708 27129
rect 14764 27073 14804 27129
rect 14296 27005 14804 27073
rect 14296 26949 14336 27005
rect 14392 26949 14460 27005
rect 14516 26949 14584 27005
rect 14640 26949 14708 27005
rect 14764 26949 14804 27005
rect 14296 25380 14804 26949
rect 14296 25328 14352 25380
rect 14404 25328 14460 25380
rect 14512 25328 14568 25380
rect 14620 25328 14804 25380
rect 14296 25272 14804 25328
rect 14296 25220 14352 25272
rect 14404 25220 14460 25272
rect 14512 25220 14568 25272
rect 14620 25220 14804 25272
rect 14296 25164 14804 25220
rect 14296 25112 14352 25164
rect 14404 25112 14460 25164
rect 14512 25112 14568 25164
rect 14620 25112 14804 25164
rect 14296 25056 14804 25112
rect 14296 25004 14352 25056
rect 14404 25004 14460 25056
rect 14512 25004 14568 25056
rect 14620 25004 14804 25056
rect 14296 24948 14804 25004
rect 14296 24896 14352 24948
rect 14404 24896 14460 24948
rect 14512 24896 14568 24948
rect 14620 24896 14804 24948
rect 14296 21469 14804 24896
rect 14296 21417 14352 21469
rect 14404 21417 14460 21469
rect 14512 21417 14568 21469
rect 14620 21417 14804 21469
rect 14296 21361 14804 21417
rect 14296 21309 14352 21361
rect 14404 21309 14460 21361
rect 14512 21309 14568 21361
rect 14620 21309 14804 21361
rect 14296 21253 14804 21309
rect 14296 21201 14352 21253
rect 14404 21201 14460 21253
rect 14512 21201 14568 21253
rect 14620 21201 14804 21253
rect 14296 13845 14804 21201
rect 14296 13789 14336 13845
rect 14392 13789 14460 13845
rect 14516 13789 14584 13845
rect 14640 13789 14708 13845
rect 14764 13789 14804 13845
rect 14296 13721 14804 13789
rect 14296 13665 14336 13721
rect 14392 13665 14460 13721
rect 14516 13665 14584 13721
rect 14640 13665 14708 13721
rect 14764 13665 14804 13721
rect 14296 13597 14804 13665
rect 14296 13541 14336 13597
rect 14392 13541 14460 13597
rect 14516 13541 14584 13597
rect 14640 13541 14708 13597
rect 14764 13541 14804 13597
rect 14296 13473 14804 13541
rect 14296 13417 14336 13473
rect 14392 13417 14460 13473
rect 14516 13417 14584 13473
rect 14640 13417 14708 13473
rect 14764 13417 14804 13473
rect 14296 13349 14804 13417
rect 14296 13293 14336 13349
rect 14392 13293 14460 13349
rect 14516 13293 14584 13349
rect 14640 13293 14708 13349
rect 14764 13293 14804 13349
rect 14296 13225 14804 13293
rect 14296 13169 14336 13225
rect 14392 13169 14460 13225
rect 14516 13169 14584 13225
rect 14640 13169 14708 13225
rect 14764 13169 14804 13225
rect 14296 13101 14804 13169
rect 14296 13045 14336 13101
rect 14392 13045 14460 13101
rect 14516 13045 14584 13101
rect 14640 13045 14708 13101
rect 14764 13045 14804 13101
rect 14296 12977 14804 13045
rect 14296 12921 14336 12977
rect 14392 12921 14460 12977
rect 14516 12921 14584 12977
rect 14640 12921 14708 12977
rect 14764 12921 14804 12977
rect 14296 12853 14804 12921
rect 14296 12797 14336 12853
rect 14392 12797 14460 12853
rect 14516 12797 14584 12853
rect 14640 12797 14708 12853
rect 14764 12797 14804 12853
rect 14296 12729 14804 12797
rect 14296 12673 14336 12729
rect 14392 12673 14460 12729
rect 14516 12673 14584 12729
rect 14640 12673 14708 12729
rect 14764 12673 14804 12729
rect 14296 12605 14804 12673
rect 14296 12549 14336 12605
rect 14392 12549 14460 12605
rect 14516 12549 14584 12605
rect 14640 12549 14708 12605
rect 14764 12549 14804 12605
rect 14296 10651 14804 12549
rect 14296 10595 14336 10651
rect 14392 10595 14460 10651
rect 14516 10595 14584 10651
rect 14640 10595 14708 10651
rect 14764 10595 14804 10651
rect 14296 10527 14804 10595
rect 14296 10471 14336 10527
rect 14392 10471 14460 10527
rect 14516 10471 14584 10527
rect 14640 10471 14708 10527
rect 14764 10471 14804 10527
rect 14296 10403 14804 10471
rect 14296 10347 14336 10403
rect 14392 10347 14460 10403
rect 14516 10347 14584 10403
rect 14640 10347 14708 10403
rect 14764 10347 14804 10403
rect 14296 10279 14804 10347
rect 14296 10223 14336 10279
rect 14392 10223 14460 10279
rect 14516 10223 14584 10279
rect 14640 10223 14708 10279
rect 14764 10223 14804 10279
rect 14296 10155 14804 10223
rect 14296 10099 14336 10155
rect 14392 10099 14460 10155
rect 14516 10099 14584 10155
rect 14640 10099 14708 10155
rect 14764 10099 14804 10155
rect 14296 10031 14804 10099
rect 14296 9975 14336 10031
rect 14392 9975 14460 10031
rect 14516 9975 14584 10031
rect 14640 9975 14708 10031
rect 14764 9975 14804 10031
rect 14296 9907 14804 9975
rect 14296 9851 14336 9907
rect 14392 9851 14460 9907
rect 14516 9851 14584 9907
rect 14640 9851 14708 9907
rect 14764 9851 14804 9907
rect 14296 9783 14804 9851
rect 14296 9727 14336 9783
rect 14392 9727 14460 9783
rect 14516 9727 14584 9783
rect 14640 9727 14708 9783
rect 14764 9727 14804 9783
rect 14296 9659 14804 9727
rect 14296 9603 14336 9659
rect 14392 9603 14460 9659
rect 14516 9603 14584 9659
rect 14640 9603 14708 9659
rect 14764 9603 14804 9659
rect 14296 9535 14804 9603
rect 14296 9479 14336 9535
rect 14392 9479 14460 9535
rect 14516 9479 14584 9535
rect 14640 9479 14708 9535
rect 14764 9479 14804 9535
rect 14296 9411 14804 9479
rect 14296 9355 14336 9411
rect 14392 9355 14460 9411
rect 14516 9355 14584 9411
rect 14640 9355 14708 9411
rect 14764 9355 14804 9411
rect 14296 9287 14804 9355
rect 14296 9231 14336 9287
rect 14392 9231 14460 9287
rect 14516 9231 14584 9287
rect 14640 9231 14708 9287
rect 14764 9231 14804 9287
rect 14296 9163 14804 9231
rect 14296 9107 14336 9163
rect 14392 9107 14460 9163
rect 14516 9107 14584 9163
rect 14640 9107 14708 9163
rect 14764 9107 14804 9163
rect 14296 9039 14804 9107
rect 14296 8983 14336 9039
rect 14392 8983 14460 9039
rect 14516 8983 14584 9039
rect 14640 8983 14708 9039
rect 14764 8983 14804 9039
rect 14296 8915 14804 8983
rect 14296 8859 14336 8915
rect 14392 8859 14460 8915
rect 14516 8859 14584 8915
rect 14640 8859 14708 8915
rect 14764 8859 14804 8915
rect 14296 8791 14804 8859
rect 14296 8735 14336 8791
rect 14392 8735 14460 8791
rect 14516 8735 14584 8791
rect 14640 8735 14708 8791
rect 14764 8735 14804 8791
rect 14296 8667 14804 8735
rect 14296 8611 14336 8667
rect 14392 8611 14460 8667
rect 14516 8611 14584 8667
rect 14640 8611 14708 8667
rect 14764 8611 14804 8667
rect 14296 8543 14804 8611
rect 14296 8487 14336 8543
rect 14392 8487 14460 8543
rect 14516 8487 14584 8543
rect 14640 8487 14708 8543
rect 14764 8487 14804 8543
rect 14296 8419 14804 8487
rect 14296 8363 14336 8419
rect 14392 8363 14460 8419
rect 14516 8363 14584 8419
rect 14640 8363 14708 8419
rect 14764 8363 14804 8419
rect 14296 8295 14804 8363
rect 14296 8239 14336 8295
rect 14392 8239 14460 8295
rect 14516 8239 14584 8295
rect 14640 8239 14708 8295
rect 14764 8239 14804 8295
rect 14296 8171 14804 8239
rect 14296 8115 14336 8171
rect 14392 8115 14460 8171
rect 14516 8115 14584 8171
rect 14640 8115 14708 8171
rect 14764 8115 14804 8171
rect 14296 8047 14804 8115
rect 14296 7991 14336 8047
rect 14392 7991 14460 8047
rect 14516 7991 14584 8047
rect 14640 7991 14708 8047
rect 14764 7991 14804 8047
rect 14296 7923 14804 7991
rect 14296 7867 14336 7923
rect 14392 7867 14460 7923
rect 14516 7867 14584 7923
rect 14640 7867 14708 7923
rect 14764 7867 14804 7923
rect 14296 7799 14804 7867
rect 14296 7743 14336 7799
rect 14392 7743 14460 7799
rect 14516 7743 14584 7799
rect 14640 7743 14708 7799
rect 14764 7743 14804 7799
rect 14296 7451 14804 7743
rect 14296 7395 14336 7451
rect 14392 7395 14460 7451
rect 14516 7395 14584 7451
rect 14640 7395 14708 7451
rect 14764 7395 14804 7451
rect 14296 7327 14804 7395
rect 14296 7271 14336 7327
rect 14392 7271 14460 7327
rect 14516 7271 14584 7327
rect 14640 7271 14708 7327
rect 14764 7271 14804 7327
rect 14296 7203 14804 7271
rect 14296 7147 14336 7203
rect 14392 7147 14460 7203
rect 14516 7147 14584 7203
rect 14640 7147 14708 7203
rect 14764 7147 14804 7203
rect 14296 7079 14804 7147
rect 14296 7023 14336 7079
rect 14392 7023 14460 7079
rect 14516 7023 14584 7079
rect 14640 7023 14708 7079
rect 14764 7023 14804 7079
rect 14296 6955 14804 7023
rect 14296 6899 14336 6955
rect 14392 6899 14460 6955
rect 14516 6899 14584 6955
rect 14640 6899 14708 6955
rect 14764 6899 14804 6955
rect 14296 6831 14804 6899
rect 14296 6775 14336 6831
rect 14392 6775 14460 6831
rect 14516 6775 14584 6831
rect 14640 6775 14708 6831
rect 14764 6775 14804 6831
rect 14296 6707 14804 6775
rect 14296 6651 14336 6707
rect 14392 6651 14460 6707
rect 14516 6651 14584 6707
rect 14640 6651 14708 6707
rect 14764 6651 14804 6707
rect 14296 6583 14804 6651
rect 14296 6527 14336 6583
rect 14392 6527 14460 6583
rect 14516 6527 14584 6583
rect 14640 6527 14708 6583
rect 14764 6527 14804 6583
rect 14296 6459 14804 6527
rect 14296 6403 14336 6459
rect 14392 6403 14460 6459
rect 14516 6403 14584 6459
rect 14640 6403 14708 6459
rect 14764 6403 14804 6459
rect 14296 6335 14804 6403
rect 14296 6279 14336 6335
rect 14392 6279 14460 6335
rect 14516 6279 14584 6335
rect 14640 6279 14708 6335
rect 14764 6279 14804 6335
rect 14296 6211 14804 6279
rect 14296 6155 14336 6211
rect 14392 6155 14460 6211
rect 14516 6155 14584 6211
rect 14640 6155 14708 6211
rect 14764 6155 14804 6211
rect 14296 6087 14804 6155
rect 14296 6031 14336 6087
rect 14392 6031 14460 6087
rect 14516 6031 14584 6087
rect 14640 6031 14708 6087
rect 14764 6031 14804 6087
rect 14296 5963 14804 6031
rect 14296 5907 14336 5963
rect 14392 5907 14460 5963
rect 14516 5907 14584 5963
rect 14640 5907 14708 5963
rect 14764 5907 14804 5963
rect 14296 5839 14804 5907
rect 14296 5783 14336 5839
rect 14392 5783 14460 5839
rect 14516 5783 14584 5839
rect 14640 5783 14708 5839
rect 14764 5783 14804 5839
rect 14296 5715 14804 5783
rect 14296 5659 14336 5715
rect 14392 5659 14460 5715
rect 14516 5659 14584 5715
rect 14640 5659 14708 5715
rect 14764 5659 14804 5715
rect 14296 5591 14804 5659
rect 14296 5535 14336 5591
rect 14392 5535 14460 5591
rect 14516 5535 14584 5591
rect 14640 5535 14708 5591
rect 14764 5535 14804 5591
rect 14296 5467 14804 5535
rect 14296 5411 14336 5467
rect 14392 5411 14460 5467
rect 14516 5411 14584 5467
rect 14640 5411 14708 5467
rect 14764 5411 14804 5467
rect 14296 5343 14804 5411
rect 14296 5287 14336 5343
rect 14392 5287 14460 5343
rect 14516 5287 14584 5343
rect 14640 5287 14708 5343
rect 14764 5287 14804 5343
rect 14296 5219 14804 5287
rect 14296 5163 14336 5219
rect 14392 5163 14460 5219
rect 14516 5163 14584 5219
rect 14640 5163 14708 5219
rect 14764 5163 14804 5219
rect 14296 5095 14804 5163
rect 14296 5039 14336 5095
rect 14392 5039 14460 5095
rect 14516 5039 14584 5095
rect 14640 5039 14708 5095
rect 14764 5039 14804 5095
rect 14296 4971 14804 5039
rect 14296 4915 14336 4971
rect 14392 4915 14460 4971
rect 14516 4915 14584 4971
rect 14640 4915 14708 4971
rect 14764 4915 14804 4971
rect 14296 4847 14804 4915
rect 14296 4791 14336 4847
rect 14392 4791 14460 4847
rect 14516 4791 14584 4847
rect 14640 4791 14708 4847
rect 14764 4791 14804 4847
rect 14296 4723 14804 4791
rect 14296 4667 14336 4723
rect 14392 4667 14460 4723
rect 14516 4667 14584 4723
rect 14640 4667 14708 4723
rect 14764 4667 14804 4723
rect 14296 4599 14804 4667
rect 14296 4543 14336 4599
rect 14392 4543 14460 4599
rect 14516 4543 14584 4599
rect 14640 4543 14708 4599
rect 14764 4543 14804 4599
rect 14296 4251 14804 4543
rect 14296 4195 14336 4251
rect 14392 4195 14460 4251
rect 14516 4195 14584 4251
rect 14640 4195 14708 4251
rect 14764 4195 14804 4251
rect 14296 4127 14804 4195
rect 14296 4071 14336 4127
rect 14392 4071 14460 4127
rect 14516 4071 14584 4127
rect 14640 4071 14708 4127
rect 14764 4071 14804 4127
rect 14296 4003 14804 4071
rect 14296 3947 14336 4003
rect 14392 3947 14460 4003
rect 14516 3947 14584 4003
rect 14640 3947 14708 4003
rect 14764 3947 14804 4003
rect 14296 3879 14804 3947
rect 14296 3823 14336 3879
rect 14392 3823 14460 3879
rect 14516 3823 14584 3879
rect 14640 3823 14708 3879
rect 14764 3823 14804 3879
rect 14296 3755 14804 3823
rect 14296 3699 14336 3755
rect 14392 3699 14460 3755
rect 14516 3699 14584 3755
rect 14640 3699 14708 3755
rect 14764 3699 14804 3755
rect 14296 3631 14804 3699
rect 14296 3575 14336 3631
rect 14392 3575 14460 3631
rect 14516 3575 14584 3631
rect 14640 3575 14708 3631
rect 14764 3575 14804 3631
rect 14296 3507 14804 3575
rect 14296 3451 14336 3507
rect 14392 3451 14460 3507
rect 14516 3451 14584 3507
rect 14640 3451 14708 3507
rect 14764 3451 14804 3507
rect 14296 3383 14804 3451
rect 14296 3327 14336 3383
rect 14392 3327 14460 3383
rect 14516 3327 14584 3383
rect 14640 3327 14708 3383
rect 14764 3327 14804 3383
rect 14296 3259 14804 3327
rect 14296 3203 14336 3259
rect 14392 3203 14460 3259
rect 14516 3203 14584 3259
rect 14640 3203 14708 3259
rect 14764 3203 14804 3259
rect 14296 3135 14804 3203
rect 14296 3079 14336 3135
rect 14392 3079 14460 3135
rect 14516 3079 14584 3135
rect 14640 3079 14708 3135
rect 14764 3079 14804 3135
rect 14296 3011 14804 3079
rect 14296 2955 14336 3011
rect 14392 2955 14460 3011
rect 14516 2955 14584 3011
rect 14640 2955 14708 3011
rect 14764 2955 14804 3011
rect 14296 2887 14804 2955
rect 14296 2831 14336 2887
rect 14392 2831 14460 2887
rect 14516 2831 14584 2887
rect 14640 2831 14708 2887
rect 14764 2831 14804 2887
rect 14296 2763 14804 2831
rect 14296 2707 14336 2763
rect 14392 2707 14460 2763
rect 14516 2707 14584 2763
rect 14640 2707 14708 2763
rect 14764 2707 14804 2763
rect 14296 2639 14804 2707
rect 14296 2583 14336 2639
rect 14392 2583 14460 2639
rect 14516 2583 14584 2639
rect 14640 2583 14708 2639
rect 14764 2583 14804 2639
rect 14296 2515 14804 2583
rect 14296 2459 14336 2515
rect 14392 2459 14460 2515
rect 14516 2459 14584 2515
rect 14640 2459 14708 2515
rect 14764 2459 14804 2515
rect 14296 2391 14804 2459
rect 14296 2335 14336 2391
rect 14392 2335 14460 2391
rect 14516 2335 14584 2391
rect 14640 2335 14708 2391
rect 14764 2335 14804 2391
rect 14296 2267 14804 2335
rect 14296 2211 14336 2267
rect 14392 2211 14460 2267
rect 14516 2211 14584 2267
rect 14640 2211 14708 2267
rect 14764 2211 14804 2267
rect 14296 2143 14804 2211
rect 14296 2087 14336 2143
rect 14392 2087 14460 2143
rect 14516 2087 14584 2143
rect 14640 2087 14708 2143
rect 14764 2087 14804 2143
rect 14296 2019 14804 2087
rect 14296 1963 14336 2019
rect 14392 1963 14460 2019
rect 14516 1963 14584 2019
rect 14640 1963 14708 2019
rect 14764 1963 14804 2019
rect 14296 1895 14804 1963
rect 14296 1839 14336 1895
rect 14392 1839 14460 1895
rect 14516 1839 14584 1895
rect 14640 1839 14708 1895
rect 14764 1839 14804 1895
rect 14296 1771 14804 1839
rect 14296 1715 14336 1771
rect 14392 1715 14460 1771
rect 14516 1715 14584 1771
rect 14640 1715 14708 1771
rect 14764 1715 14804 1771
rect 14296 1647 14804 1715
rect 14296 1591 14336 1647
rect 14392 1591 14460 1647
rect 14516 1591 14584 1647
rect 14640 1591 14708 1647
rect 14764 1591 14804 1647
rect 14296 1523 14804 1591
rect 14296 1467 14336 1523
rect 14392 1467 14460 1523
rect 14516 1467 14584 1523
rect 14640 1467 14708 1523
rect 14764 1467 14804 1523
rect 14296 1399 14804 1467
rect 14296 1343 14336 1399
rect 14392 1343 14460 1399
rect 14516 1343 14584 1399
rect 14640 1343 14708 1399
rect 14764 1343 14804 1399
rect 14296 900 14804 1343
<< via2 >>
rect 300 56866 356 56922
rect 424 56866 480 56922
rect 548 56866 604 56922
rect 672 56866 728 56922
rect 300 56742 356 56798
rect 424 56742 480 56798
rect 548 56742 604 56798
rect 672 56742 728 56798
rect 300 56618 356 56674
rect 424 56659 444 56674
rect 444 56659 480 56674
rect 548 56659 552 56674
rect 552 56659 604 56674
rect 672 56659 712 56674
rect 712 56659 728 56674
rect 424 56618 480 56659
rect 548 56618 604 56659
rect 672 56618 728 56659
rect 300 56494 356 56550
rect 424 56495 480 56550
rect 548 56495 604 56550
rect 672 56495 728 56550
rect 424 56494 444 56495
rect 444 56494 480 56495
rect 548 56494 552 56495
rect 552 56494 604 56495
rect 672 56494 712 56495
rect 712 56494 728 56495
rect 300 56370 356 56426
rect 424 56370 480 56426
rect 548 56370 604 56426
rect 672 56370 728 56426
rect 1436 56866 1492 56922
rect 1560 56866 1616 56922
rect 1684 56866 1740 56922
rect 1808 56866 1864 56922
rect 1436 56742 1492 56798
rect 1560 56742 1616 56798
rect 1684 56742 1740 56798
rect 1808 56742 1864 56798
rect 1436 56659 1460 56674
rect 1460 56659 1492 56674
rect 1560 56659 1568 56674
rect 1568 56659 1616 56674
rect 1684 56659 1732 56674
rect 1732 56659 1740 56674
rect 1808 56659 1840 56674
rect 1840 56659 1864 56674
rect 1436 56618 1492 56659
rect 1560 56618 1616 56659
rect 1684 56618 1740 56659
rect 1808 56618 1864 56659
rect 1436 56495 1492 56550
rect 1560 56495 1616 56550
rect 1684 56495 1740 56550
rect 1808 56495 1864 56550
rect 1436 56494 1460 56495
rect 1460 56494 1492 56495
rect 1560 56494 1568 56495
rect 1568 56494 1616 56495
rect 1684 56494 1732 56495
rect 1732 56494 1740 56495
rect 1808 56494 1840 56495
rect 1840 56494 1864 56495
rect 1436 56370 1492 56426
rect 1560 56370 1616 56426
rect 1684 56370 1740 56426
rect 1808 56370 1864 56426
rect 300 56246 356 56302
rect 424 56246 480 56302
rect 548 56246 604 56302
rect 672 56246 728 56302
rect 300 56122 356 56178
rect 424 56122 480 56178
rect 548 56122 604 56178
rect 672 56122 728 56178
rect 300 55998 356 56054
rect 424 55998 480 56054
rect 548 55998 604 56054
rect 672 55998 728 56054
rect 300 55874 356 55930
rect 424 55874 480 55930
rect 548 55874 604 55930
rect 672 55874 728 55930
rect 300 55750 356 55806
rect 424 55750 480 55806
rect 548 55750 604 55806
rect 672 55750 728 55806
rect 1436 56246 1492 56302
rect 1560 56246 1616 56302
rect 1684 56246 1740 56302
rect 1808 56246 1864 56302
rect 1436 56122 1492 56178
rect 1560 56122 1616 56178
rect 1684 56122 1740 56178
rect 1808 56122 1864 56178
rect 1436 55998 1492 56054
rect 1560 55998 1616 56054
rect 1684 55998 1740 56054
rect 1808 55998 1864 56054
rect 1436 55874 1492 55930
rect 1560 55874 1616 55930
rect 1684 55874 1740 55930
rect 1808 55874 1864 55930
rect 1436 55750 1492 55806
rect 1560 55750 1616 55806
rect 1684 55750 1740 55806
rect 1808 55750 1864 55806
rect 868 55389 924 55445
rect 992 55404 1030 55445
rect 1030 55404 1048 55445
rect 1116 55404 1154 55445
rect 1154 55404 1172 55445
rect 1240 55404 1278 55445
rect 1278 55404 1296 55445
rect 992 55389 1048 55404
rect 1116 55389 1172 55404
rect 1240 55389 1296 55404
rect 868 55265 924 55321
rect 992 55280 1030 55321
rect 1030 55280 1048 55321
rect 1116 55280 1154 55321
rect 1154 55280 1172 55321
rect 1240 55280 1278 55321
rect 1278 55280 1296 55321
rect 992 55265 1048 55280
rect 1116 55265 1172 55280
rect 1240 55265 1296 55280
rect 868 55141 924 55197
rect 992 55156 1030 55197
rect 1030 55156 1048 55197
rect 1116 55156 1154 55197
rect 1154 55156 1172 55197
rect 1240 55156 1278 55197
rect 1278 55156 1296 55197
rect 992 55141 1048 55156
rect 1116 55141 1172 55156
rect 1240 55141 1296 55156
rect 868 55017 924 55073
rect 992 55032 1030 55073
rect 1030 55032 1048 55073
rect 1116 55032 1154 55073
rect 1154 55032 1172 55073
rect 1240 55032 1278 55073
rect 1278 55032 1296 55073
rect 992 55017 1048 55032
rect 1116 55017 1172 55032
rect 1240 55017 1296 55032
rect 868 54893 924 54949
rect 992 54908 1030 54949
rect 1030 54908 1048 54949
rect 1116 54908 1154 54949
rect 1154 54908 1172 54949
rect 1240 54908 1278 54949
rect 1278 54908 1296 54949
rect 992 54893 1048 54908
rect 1116 54893 1172 54908
rect 1240 54893 1296 54908
rect 868 54769 924 54825
rect 992 54784 1030 54825
rect 1030 54784 1048 54825
rect 1116 54784 1154 54825
rect 1154 54784 1172 54825
rect 1240 54784 1278 54825
rect 1278 54784 1296 54825
rect 992 54769 1048 54784
rect 1116 54769 1172 54784
rect 1240 54769 1296 54784
rect 868 54645 924 54701
rect 992 54660 1030 54701
rect 1030 54660 1048 54701
rect 1116 54660 1154 54701
rect 1154 54660 1172 54701
rect 1240 54660 1278 54701
rect 1278 54660 1296 54701
rect 992 54645 1048 54660
rect 1116 54645 1172 54660
rect 1240 54645 1296 54660
rect 868 54521 924 54577
rect 992 54536 1030 54577
rect 1030 54536 1048 54577
rect 1116 54536 1154 54577
rect 1154 54536 1172 54577
rect 1240 54536 1278 54577
rect 1278 54536 1296 54577
rect 992 54521 1048 54536
rect 1116 54521 1172 54536
rect 1240 54521 1296 54536
rect 868 54397 924 54453
rect 992 54412 1030 54453
rect 1030 54412 1048 54453
rect 1116 54412 1154 54453
rect 1154 54412 1172 54453
rect 1240 54412 1278 54453
rect 1278 54412 1296 54453
rect 992 54397 1048 54412
rect 1116 54397 1172 54412
rect 1240 54397 1296 54412
rect 868 54273 924 54329
rect 992 54288 1030 54329
rect 1030 54288 1048 54329
rect 1116 54288 1154 54329
rect 1154 54288 1172 54329
rect 1240 54288 1278 54329
rect 1278 54288 1296 54329
rect 992 54273 1048 54288
rect 1116 54273 1172 54288
rect 1240 54273 1296 54288
rect 868 54149 924 54205
rect 992 54164 1030 54205
rect 1030 54164 1048 54205
rect 1116 54164 1154 54205
rect 1154 54164 1172 54205
rect 1240 54164 1278 54205
rect 1278 54164 1296 54205
rect 992 54149 1048 54164
rect 1116 54149 1172 54164
rect 1240 54149 1296 54164
rect 300 53789 356 53845
rect 424 53789 480 53845
rect 548 53789 604 53845
rect 672 53789 728 53845
rect 300 53665 356 53721
rect 424 53665 480 53721
rect 548 53665 604 53721
rect 672 53665 728 53721
rect 300 53541 356 53597
rect 424 53541 480 53597
rect 548 53541 604 53597
rect 672 53541 728 53597
rect 300 53417 356 53473
rect 424 53417 480 53473
rect 548 53417 604 53473
rect 672 53417 728 53473
rect 300 53293 356 53349
rect 424 53293 480 53349
rect 548 53293 604 53349
rect 672 53293 728 53349
rect 300 53169 356 53225
rect 424 53169 480 53225
rect 548 53169 604 53225
rect 672 53169 728 53225
rect 1436 53789 1492 53845
rect 1560 53789 1616 53845
rect 1684 53789 1740 53845
rect 1808 53789 1864 53845
rect 1436 53665 1492 53721
rect 1560 53665 1616 53721
rect 1684 53665 1740 53721
rect 1808 53665 1864 53721
rect 1436 53541 1492 53597
rect 1560 53541 1616 53597
rect 1684 53541 1740 53597
rect 1808 53541 1864 53597
rect 1436 53417 1492 53473
rect 1560 53417 1616 53473
rect 1684 53417 1740 53473
rect 1808 53417 1864 53473
rect 1436 53293 1492 53349
rect 1560 53293 1616 53349
rect 1684 53293 1740 53349
rect 1808 53293 1864 53349
rect 1436 53169 1492 53225
rect 1560 53169 1616 53225
rect 1684 53169 1740 53225
rect 1808 53169 1864 53225
rect 300 53045 356 53101
rect 424 53045 480 53101
rect 548 53045 604 53101
rect 672 53045 728 53101
rect 300 52921 356 52977
rect 424 52964 444 52977
rect 444 52964 480 52977
rect 548 52964 552 52977
rect 552 52964 604 52977
rect 672 52964 712 52977
rect 712 52964 728 52977
rect 424 52921 480 52964
rect 548 52921 604 52964
rect 672 52921 728 52964
rect 300 52797 356 52853
rect 424 52800 480 52853
rect 548 52800 604 52853
rect 672 52800 728 52853
rect 424 52797 444 52800
rect 444 52797 480 52800
rect 548 52797 552 52800
rect 552 52797 604 52800
rect 672 52797 712 52800
rect 712 52797 728 52800
rect 300 52673 356 52729
rect 424 52692 480 52729
rect 548 52692 604 52729
rect 672 52692 728 52729
rect 424 52673 444 52692
rect 444 52673 480 52692
rect 548 52673 552 52692
rect 552 52673 604 52692
rect 672 52673 712 52692
rect 712 52673 728 52692
rect 300 52549 356 52605
rect 424 52584 480 52605
rect 548 52584 604 52605
rect 672 52584 728 52605
rect 424 52549 444 52584
rect 444 52549 480 52584
rect 548 52549 552 52584
rect 552 52549 604 52584
rect 672 52549 712 52584
rect 712 52549 728 52584
rect 56 52271 112 52273
rect 56 52219 58 52271
rect 58 52219 110 52271
rect 110 52219 112 52271
rect 56 52163 112 52219
rect 56 52111 58 52163
rect 58 52111 110 52163
rect 110 52111 112 52163
rect 56 52055 112 52111
rect 56 52003 58 52055
rect 58 52003 110 52055
rect 110 52003 112 52055
rect 56 51947 112 52003
rect 56 51895 58 51947
rect 58 51895 110 51947
rect 110 51895 112 51947
rect 56 51839 112 51895
rect 56 51787 58 51839
rect 58 51787 110 51839
rect 110 51787 112 51839
rect 56 51731 112 51787
rect 56 51679 58 51731
rect 58 51679 110 51731
rect 110 51679 112 51731
rect 56 51623 112 51679
rect 56 51571 58 51623
rect 58 51571 110 51623
rect 110 51571 112 51623
rect 56 51515 112 51571
rect 56 51463 58 51515
rect 58 51463 110 51515
rect 110 51463 112 51515
rect 56 51407 112 51463
rect 56 51355 58 51407
rect 58 51355 110 51407
rect 110 51355 112 51407
rect 56 51299 112 51355
rect 56 51247 58 51299
rect 58 51247 110 51299
rect 110 51247 112 51299
rect 56 51191 112 51247
rect 56 51139 58 51191
rect 58 51139 110 51191
rect 110 51139 112 51191
rect 56 51083 112 51139
rect 56 51031 58 51083
rect 58 51031 110 51083
rect 110 51031 112 51083
rect 56 50975 112 51031
rect 56 50923 58 50975
rect 58 50923 110 50975
rect 110 50923 112 50975
rect 56 50921 112 50923
rect 300 48989 356 49045
rect 424 49016 444 49045
rect 444 49016 480 49045
rect 548 49016 552 49045
rect 552 49016 604 49045
rect 672 49016 712 49045
rect 712 49016 728 49045
rect 424 48989 480 49016
rect 548 48989 604 49016
rect 672 48989 728 49016
rect 300 48865 356 48921
rect 424 48908 444 48921
rect 444 48908 480 48921
rect 548 48908 552 48921
rect 552 48908 604 48921
rect 672 48908 712 48921
rect 712 48908 728 48921
rect 424 48865 480 48908
rect 548 48865 604 48908
rect 672 48865 728 48908
rect 300 48741 356 48797
rect 424 48744 480 48797
rect 548 48744 604 48797
rect 672 48744 728 48797
rect 424 48741 444 48744
rect 444 48741 480 48744
rect 548 48741 552 48744
rect 552 48741 604 48744
rect 672 48741 712 48744
rect 712 48741 728 48744
rect 300 48617 356 48673
rect 424 48636 480 48673
rect 548 48636 604 48673
rect 672 48636 728 48673
rect 424 48617 444 48636
rect 444 48617 480 48636
rect 548 48617 552 48636
rect 552 48617 604 48636
rect 672 48617 712 48636
rect 712 48617 728 48636
rect 300 48493 356 48549
rect 424 48493 480 48549
rect 548 48493 604 48549
rect 672 48493 728 48549
rect 300 48369 356 48425
rect 424 48369 480 48425
rect 548 48369 604 48425
rect 672 48369 728 48425
rect 300 48245 356 48301
rect 424 48245 480 48301
rect 548 48245 604 48301
rect 672 48245 728 48301
rect 300 48121 356 48177
rect 424 48121 480 48177
rect 548 48121 604 48177
rect 672 48121 728 48177
rect 300 47997 356 48053
rect 424 47997 480 48053
rect 548 47997 604 48053
rect 672 47997 728 48053
rect 300 47873 356 47929
rect 424 47873 480 47929
rect 548 47873 604 47929
rect 672 47873 728 47929
rect 300 47749 356 47805
rect 424 47749 480 47805
rect 548 47749 604 47805
rect 672 47749 728 47805
rect 300 45789 356 45845
rect 424 45789 480 45845
rect 548 45789 604 45845
rect 672 45789 728 45845
rect 300 45665 356 45721
rect 424 45665 480 45721
rect 548 45665 604 45721
rect 672 45665 728 45721
rect 300 45541 356 45597
rect 424 45541 480 45597
rect 548 45541 604 45597
rect 672 45541 728 45597
rect 300 45417 356 45473
rect 424 45417 480 45473
rect 548 45417 604 45473
rect 672 45417 728 45473
rect 300 45293 356 45349
rect 424 45293 480 45349
rect 548 45293 604 45349
rect 672 45293 728 45349
rect 300 45169 356 45225
rect 424 45169 480 45225
rect 548 45169 604 45225
rect 672 45169 728 45225
rect 300 45045 356 45101
rect 424 45068 444 45101
rect 444 45068 480 45101
rect 548 45068 552 45101
rect 552 45068 604 45101
rect 672 45068 712 45101
rect 712 45068 728 45101
rect 424 45045 480 45068
rect 548 45045 604 45068
rect 672 45045 728 45068
rect 300 44921 356 44977
rect 424 44960 444 44977
rect 444 44960 480 44977
rect 548 44960 552 44977
rect 552 44960 604 44977
rect 672 44960 712 44977
rect 712 44960 728 44977
rect 424 44921 480 44960
rect 548 44921 604 44960
rect 672 44921 728 44960
rect 300 44797 356 44853
rect 424 44852 444 44853
rect 444 44852 480 44853
rect 548 44852 552 44853
rect 552 44852 604 44853
rect 672 44852 712 44853
rect 712 44852 728 44853
rect 424 44797 480 44852
rect 548 44797 604 44852
rect 672 44797 728 44852
rect 300 44673 356 44729
rect 424 44688 480 44729
rect 548 44688 604 44729
rect 672 44688 728 44729
rect 424 44673 444 44688
rect 444 44673 480 44688
rect 548 44673 552 44688
rect 552 44673 604 44688
rect 672 44673 712 44688
rect 712 44673 728 44688
rect 300 44549 356 44605
rect 424 44549 480 44605
rect 548 44549 604 44605
rect 672 44549 728 44605
rect 56 37871 112 37873
rect 56 37819 58 37871
rect 58 37819 110 37871
rect 110 37819 112 37871
rect 56 37763 112 37819
rect 56 37711 58 37763
rect 58 37711 110 37763
rect 110 37711 112 37763
rect 56 37655 112 37711
rect 56 37603 58 37655
rect 58 37603 110 37655
rect 110 37603 112 37655
rect 56 37547 112 37603
rect 56 37495 58 37547
rect 58 37495 110 37547
rect 110 37495 112 37547
rect 56 37439 112 37495
rect 56 37387 58 37439
rect 58 37387 110 37439
rect 110 37387 112 37439
rect 56 37331 112 37387
rect 56 37279 58 37331
rect 58 37279 110 37331
rect 110 37279 112 37331
rect 56 37223 112 37279
rect 56 37171 58 37223
rect 58 37171 110 37223
rect 110 37171 112 37223
rect 56 37115 112 37171
rect 56 37063 58 37115
rect 58 37063 110 37115
rect 110 37063 112 37115
rect 56 37007 112 37063
rect 56 36955 58 37007
rect 58 36955 110 37007
rect 110 36955 112 37007
rect 56 36899 112 36955
rect 56 36847 58 36899
rect 58 36847 110 36899
rect 110 36847 112 36899
rect 56 36791 112 36847
rect 56 36739 58 36791
rect 58 36739 110 36791
rect 110 36739 112 36791
rect 56 36683 112 36739
rect 56 36631 58 36683
rect 58 36631 110 36683
rect 110 36631 112 36683
rect 56 36575 112 36631
rect 56 36523 58 36575
rect 58 36523 110 36575
rect 110 36523 112 36575
rect 56 36521 112 36523
rect 838 50589 894 50645
rect 962 50589 1018 50645
rect 838 50465 894 50521
rect 962 50465 1018 50521
rect 838 50341 894 50397
rect 962 50341 1018 50397
rect 838 50217 894 50273
rect 962 50217 1018 50273
rect 838 50093 894 50149
rect 962 50093 1018 50149
rect 838 49969 894 50025
rect 962 49969 1018 50025
rect 838 49845 894 49901
rect 962 49845 1018 49901
rect 838 49721 894 49777
rect 962 49721 1018 49777
rect 838 49597 894 49653
rect 962 49597 1018 49653
rect 838 49473 894 49529
rect 962 49473 1018 49529
rect 838 49349 894 49405
rect 962 49349 1018 49405
rect 838 39389 894 39445
rect 962 39389 1018 39445
rect 838 39265 894 39321
rect 962 39265 1018 39321
rect 838 39141 894 39197
rect 962 39141 1018 39197
rect 838 39017 894 39073
rect 962 39017 1018 39073
rect 838 38893 894 38949
rect 962 38893 1018 38949
rect 838 38769 894 38825
rect 962 38769 1018 38825
rect 838 38645 894 38701
rect 962 38645 1018 38701
rect 838 38521 894 38577
rect 962 38521 1018 38577
rect 838 38397 894 38453
rect 962 38397 1018 38453
rect 838 38273 894 38329
rect 962 38273 1018 38329
rect 838 38149 894 38205
rect 962 38149 1018 38205
rect 1146 47436 1202 47445
rect 1146 47389 1148 47436
rect 1148 47389 1200 47436
rect 1200 47389 1202 47436
rect 1270 47436 1326 47445
rect 1270 47389 1272 47436
rect 1272 47389 1324 47436
rect 1324 47389 1326 47436
rect 1146 47312 1202 47321
rect 1146 47265 1148 47312
rect 1148 47265 1200 47312
rect 1200 47265 1202 47312
rect 1270 47312 1326 47321
rect 1270 47265 1272 47312
rect 1272 47265 1324 47312
rect 1324 47265 1326 47312
rect 1146 47188 1202 47197
rect 1146 47141 1148 47188
rect 1148 47141 1200 47188
rect 1200 47141 1202 47188
rect 1270 47188 1326 47197
rect 1270 47141 1272 47188
rect 1272 47141 1324 47188
rect 1324 47141 1326 47188
rect 1146 47064 1202 47073
rect 1146 47017 1148 47064
rect 1148 47017 1200 47064
rect 1200 47017 1202 47064
rect 1270 47064 1326 47073
rect 1270 47017 1272 47064
rect 1272 47017 1324 47064
rect 1324 47017 1326 47064
rect 1146 46940 1202 46949
rect 1146 46893 1148 46940
rect 1148 46893 1200 46940
rect 1200 46893 1202 46940
rect 1270 46940 1326 46949
rect 1270 46893 1272 46940
rect 1272 46893 1324 46940
rect 1324 46893 1326 46940
rect 1146 46816 1202 46825
rect 1146 46769 1148 46816
rect 1148 46769 1200 46816
rect 1200 46769 1202 46816
rect 1270 46816 1326 46825
rect 1270 46769 1272 46816
rect 1272 46769 1324 46816
rect 1324 46769 1326 46816
rect 1146 46692 1202 46701
rect 1146 46645 1148 46692
rect 1148 46645 1200 46692
rect 1200 46645 1202 46692
rect 1270 46692 1326 46701
rect 1270 46645 1272 46692
rect 1272 46645 1324 46692
rect 1324 46645 1326 46692
rect 1146 46568 1202 46577
rect 1146 46521 1148 46568
rect 1148 46521 1200 46568
rect 1200 46521 1202 46568
rect 1270 46568 1326 46577
rect 1270 46521 1272 46568
rect 1272 46521 1324 46568
rect 1324 46521 1326 46568
rect 1146 46444 1202 46453
rect 1146 46397 1148 46444
rect 1148 46397 1200 46444
rect 1200 46397 1202 46444
rect 1270 46444 1326 46453
rect 1270 46397 1272 46444
rect 1272 46397 1324 46444
rect 1324 46397 1326 46444
rect 1146 46320 1202 46329
rect 1146 46273 1148 46320
rect 1148 46273 1200 46320
rect 1200 46273 1202 46320
rect 1270 46320 1326 46329
rect 1270 46273 1272 46320
rect 1272 46273 1324 46320
rect 1324 46273 1326 46320
rect 1146 46196 1202 46205
rect 1146 46149 1148 46196
rect 1148 46149 1200 46196
rect 1200 46149 1202 46196
rect 1270 46196 1326 46205
rect 1270 46149 1272 46196
rect 1272 46149 1324 46196
rect 1324 46149 1326 46196
rect 1146 44232 1202 44245
rect 1146 44189 1148 44232
rect 1148 44189 1200 44232
rect 1200 44189 1202 44232
rect 1270 44232 1326 44245
rect 1270 44189 1272 44232
rect 1272 44189 1324 44232
rect 1324 44189 1326 44232
rect 1146 44108 1202 44121
rect 1146 44065 1148 44108
rect 1148 44065 1200 44108
rect 1200 44065 1202 44108
rect 1270 44108 1326 44121
rect 1270 44065 1272 44108
rect 1272 44065 1324 44108
rect 1324 44065 1326 44108
rect 1146 43984 1202 43997
rect 1146 43941 1148 43984
rect 1148 43941 1200 43984
rect 1200 43941 1202 43984
rect 1270 43984 1326 43997
rect 1270 43941 1272 43984
rect 1272 43941 1324 43984
rect 1324 43941 1326 43984
rect 1146 43860 1202 43873
rect 1146 43817 1148 43860
rect 1148 43817 1200 43860
rect 1200 43817 1202 43860
rect 1270 43860 1326 43873
rect 1270 43817 1272 43860
rect 1272 43817 1324 43860
rect 1324 43817 1326 43860
rect 1146 43736 1202 43749
rect 1146 43693 1148 43736
rect 1148 43693 1200 43736
rect 1200 43693 1202 43736
rect 1270 43736 1326 43749
rect 1270 43693 1272 43736
rect 1272 43693 1324 43736
rect 1324 43693 1326 43736
rect 1146 43612 1202 43625
rect 1146 43569 1148 43612
rect 1148 43569 1200 43612
rect 1200 43569 1202 43612
rect 1270 43612 1326 43625
rect 1270 43569 1272 43612
rect 1272 43569 1324 43612
rect 1324 43569 1326 43612
rect 1146 43488 1202 43501
rect 1146 43445 1148 43488
rect 1148 43445 1200 43488
rect 1200 43445 1202 43488
rect 1270 43488 1326 43501
rect 1270 43445 1272 43488
rect 1272 43445 1324 43488
rect 1324 43445 1326 43488
rect 1146 43364 1202 43377
rect 1146 43321 1148 43364
rect 1148 43321 1200 43364
rect 1200 43321 1202 43364
rect 1270 43364 1326 43377
rect 1270 43321 1272 43364
rect 1272 43321 1324 43364
rect 1324 43321 1326 43364
rect 1146 43240 1202 43253
rect 1146 43197 1148 43240
rect 1148 43197 1200 43240
rect 1200 43197 1202 43240
rect 1270 43240 1326 43253
rect 1270 43197 1272 43240
rect 1272 43197 1324 43240
rect 1324 43197 1326 43240
rect 1146 43116 1202 43129
rect 1146 43073 1148 43116
rect 1148 43073 1200 43116
rect 1200 43073 1202 43116
rect 1270 43116 1326 43129
rect 1270 43073 1272 43116
rect 1272 43073 1324 43116
rect 1324 43073 1326 43116
rect 1146 42992 1202 43005
rect 1146 42949 1148 42992
rect 1148 42949 1200 42992
rect 1200 42949 1202 42992
rect 1270 42992 1326 43005
rect 1270 42949 1272 42992
rect 1272 42949 1324 42992
rect 1324 42949 1326 42992
rect 1146 42620 1202 42645
rect 1146 42589 1148 42620
rect 1148 42589 1200 42620
rect 1200 42589 1202 42620
rect 1270 42620 1326 42645
rect 1270 42589 1272 42620
rect 1272 42589 1324 42620
rect 1324 42589 1326 42620
rect 1146 42496 1202 42521
rect 1146 42465 1148 42496
rect 1148 42465 1200 42496
rect 1200 42465 1202 42496
rect 1270 42496 1326 42521
rect 1270 42465 1272 42496
rect 1272 42465 1324 42496
rect 1324 42465 1326 42496
rect 1146 42372 1202 42397
rect 1146 42341 1148 42372
rect 1148 42341 1200 42372
rect 1200 42341 1202 42372
rect 1270 42372 1326 42397
rect 1270 42341 1272 42372
rect 1272 42341 1324 42372
rect 1324 42341 1326 42372
rect 1146 42248 1202 42273
rect 1146 42217 1148 42248
rect 1148 42217 1200 42248
rect 1200 42217 1202 42248
rect 1270 42248 1326 42273
rect 1270 42217 1272 42248
rect 1272 42217 1324 42248
rect 1324 42217 1326 42248
rect 1146 42124 1202 42149
rect 1146 42093 1148 42124
rect 1148 42093 1200 42124
rect 1200 42093 1202 42124
rect 1270 42124 1326 42149
rect 1270 42093 1272 42124
rect 1272 42093 1324 42124
rect 1324 42093 1326 42124
rect 1146 42000 1202 42025
rect 1146 41969 1148 42000
rect 1148 41969 1200 42000
rect 1200 41969 1202 42000
rect 1270 42000 1326 42025
rect 1270 41969 1272 42000
rect 1272 41969 1324 42000
rect 1324 41969 1326 42000
rect 1146 41876 1202 41901
rect 1146 41845 1148 41876
rect 1148 41845 1200 41876
rect 1200 41845 1202 41876
rect 1270 41876 1326 41901
rect 1270 41845 1272 41876
rect 1272 41845 1324 41876
rect 1324 41845 1326 41876
rect 1146 41752 1202 41777
rect 1146 41721 1148 41752
rect 1148 41721 1200 41752
rect 1200 41721 1202 41752
rect 1270 41752 1326 41777
rect 1270 41721 1272 41752
rect 1272 41721 1324 41752
rect 1324 41721 1326 41752
rect 1146 41628 1202 41653
rect 1146 41597 1148 41628
rect 1148 41597 1200 41628
rect 1200 41597 1202 41628
rect 1270 41628 1326 41653
rect 1270 41597 1272 41628
rect 1272 41597 1324 41628
rect 1324 41597 1326 41628
rect 1146 41504 1202 41529
rect 1146 41473 1148 41504
rect 1148 41473 1200 41504
rect 1200 41473 1202 41504
rect 1270 41504 1326 41529
rect 1270 41473 1272 41504
rect 1272 41473 1324 41504
rect 1324 41473 1326 41504
rect 1146 41380 1202 41405
rect 1146 41349 1148 41380
rect 1148 41349 1200 41380
rect 1200 41349 1202 41380
rect 1270 41380 1326 41405
rect 1270 41349 1272 41380
rect 1272 41349 1324 41380
rect 1324 41349 1326 41380
rect 1146 40989 1202 41045
rect 1270 40989 1326 41045
rect 1146 40865 1202 40921
rect 1270 40865 1326 40921
rect 1146 40741 1202 40797
rect 1270 40741 1326 40797
rect 1146 40617 1202 40673
rect 1270 40617 1326 40673
rect 1146 40532 1202 40549
rect 1146 40493 1148 40532
rect 1148 40493 1200 40532
rect 1200 40493 1202 40532
rect 1270 40532 1326 40549
rect 1270 40493 1272 40532
rect 1272 40493 1324 40532
rect 1324 40493 1326 40532
rect 1146 40408 1202 40425
rect 1146 40369 1148 40408
rect 1148 40369 1200 40408
rect 1200 40369 1202 40408
rect 1270 40408 1326 40425
rect 1270 40369 1272 40408
rect 1272 40369 1324 40408
rect 1324 40369 1326 40408
rect 1146 40284 1202 40301
rect 1146 40245 1148 40284
rect 1148 40245 1200 40284
rect 1200 40245 1202 40284
rect 1270 40284 1326 40301
rect 1270 40245 1272 40284
rect 1272 40245 1324 40284
rect 1324 40245 1326 40284
rect 1146 40160 1202 40177
rect 1146 40121 1148 40160
rect 1148 40121 1200 40160
rect 1200 40121 1202 40160
rect 1270 40160 1326 40177
rect 1270 40121 1272 40160
rect 1272 40121 1324 40160
rect 1324 40121 1326 40160
rect 1146 40036 1202 40053
rect 1146 39997 1148 40036
rect 1148 39997 1200 40036
rect 1200 39997 1202 40036
rect 1270 40036 1326 40053
rect 1270 39997 1272 40036
rect 1272 39997 1324 40036
rect 1324 39997 1326 40036
rect 1146 39912 1202 39929
rect 1146 39873 1148 39912
rect 1148 39873 1200 39912
rect 1200 39873 1202 39912
rect 1270 39912 1326 39929
rect 1270 39873 1272 39912
rect 1272 39873 1324 39912
rect 1324 39873 1326 39912
rect 1146 39788 1202 39805
rect 1146 39749 1148 39788
rect 1148 39749 1200 39788
rect 1200 39749 1202 39788
rect 1270 39788 1326 39805
rect 1270 39749 1272 39788
rect 1272 39749 1324 39788
rect 1324 39749 1326 39788
rect 300 36195 356 36251
rect 424 36195 480 36251
rect 548 36195 604 36251
rect 672 36195 728 36251
rect 300 36071 356 36127
rect 424 36071 480 36127
rect 548 36071 604 36127
rect 672 36071 728 36127
rect 300 35947 356 36003
rect 424 35947 480 36003
rect 548 35947 604 36003
rect 672 35947 728 36003
rect 300 35823 356 35879
rect 424 35823 480 35879
rect 548 35823 604 35879
rect 672 35823 728 35879
rect 300 35699 356 35755
rect 424 35699 480 35755
rect 548 35699 604 35755
rect 672 35699 728 35755
rect 300 35575 356 35631
rect 424 35575 480 35631
rect 548 35575 604 35631
rect 672 35575 728 35631
rect 300 35451 356 35507
rect 424 35451 480 35507
rect 548 35451 604 35507
rect 672 35451 728 35507
rect 300 35327 356 35383
rect 424 35327 480 35383
rect 548 35327 604 35383
rect 672 35327 728 35383
rect 300 35203 356 35259
rect 424 35203 480 35259
rect 548 35203 604 35259
rect 672 35203 728 35259
rect 300 35079 356 35135
rect 424 35079 480 35135
rect 548 35079 604 35135
rect 672 35079 728 35135
rect 300 34955 356 35011
rect 424 34955 480 35011
rect 548 34955 604 35011
rect 672 34955 728 35011
rect 300 34831 356 34887
rect 424 34831 480 34887
rect 548 34831 604 34887
rect 672 34831 728 34887
rect 300 34707 356 34763
rect 424 34707 480 34763
rect 548 34707 604 34763
rect 672 34707 728 34763
rect 300 34583 356 34639
rect 424 34583 480 34639
rect 548 34583 604 34639
rect 672 34583 728 34639
rect 300 34459 356 34515
rect 424 34459 480 34515
rect 548 34459 604 34515
rect 672 34459 728 34515
rect 300 34335 356 34391
rect 424 34335 480 34391
rect 548 34335 604 34391
rect 672 34335 728 34391
rect 300 34211 356 34267
rect 424 34211 480 34267
rect 548 34211 604 34267
rect 672 34211 728 34267
rect 300 34087 356 34143
rect 424 34087 480 34143
rect 548 34087 604 34143
rect 672 34087 728 34143
rect 300 33963 356 34019
rect 424 33963 480 34019
rect 548 33963 604 34019
rect 672 33963 728 34019
rect 300 33839 356 33895
rect 424 33839 480 33895
rect 548 33839 604 33895
rect 672 33839 728 33895
rect 300 33715 356 33771
rect 424 33715 480 33771
rect 548 33715 604 33771
rect 672 33715 728 33771
rect 300 33591 356 33647
rect 424 33591 480 33647
rect 548 33591 604 33647
rect 672 33591 728 33647
rect 300 33467 356 33523
rect 424 33467 480 33523
rect 548 33467 604 33523
rect 672 33467 728 33523
rect 300 33343 356 33399
rect 424 33343 480 33399
rect 548 33343 604 33399
rect 672 33343 728 33399
rect 868 32995 924 33051
rect 992 32995 1048 33051
rect 1116 32995 1172 33051
rect 1240 32995 1296 33051
rect 868 32871 924 32927
rect 992 32871 1048 32927
rect 1116 32871 1172 32927
rect 1240 32871 1296 32927
rect 868 32747 924 32803
rect 992 32747 1048 32803
rect 1116 32747 1172 32803
rect 1240 32747 1296 32803
rect 868 32623 924 32679
rect 992 32636 1048 32679
rect 1116 32636 1172 32679
rect 1240 32636 1296 32679
rect 992 32623 1030 32636
rect 1030 32623 1048 32636
rect 1116 32623 1154 32636
rect 1154 32623 1172 32636
rect 1240 32623 1278 32636
rect 1278 32623 1296 32636
rect 868 32499 924 32555
rect 992 32512 1048 32555
rect 1116 32512 1172 32555
rect 1240 32512 1296 32555
rect 992 32499 1030 32512
rect 1030 32499 1048 32512
rect 1116 32499 1154 32512
rect 1154 32499 1172 32512
rect 1240 32499 1278 32512
rect 1278 32499 1296 32512
rect 868 32375 924 32431
rect 992 32388 1048 32431
rect 1116 32388 1172 32431
rect 1240 32388 1296 32431
rect 992 32375 1030 32388
rect 1030 32375 1048 32388
rect 1116 32375 1154 32388
rect 1154 32375 1172 32388
rect 1240 32375 1278 32388
rect 1278 32375 1296 32388
rect 868 32251 924 32307
rect 992 32264 1048 32307
rect 1116 32264 1172 32307
rect 1240 32264 1296 32307
rect 992 32251 1030 32264
rect 1030 32251 1048 32264
rect 1116 32251 1154 32264
rect 1154 32251 1172 32264
rect 1240 32251 1278 32264
rect 1278 32251 1296 32264
rect 868 32127 924 32183
rect 992 32140 1048 32183
rect 1116 32140 1172 32183
rect 1240 32140 1296 32183
rect 992 32127 1030 32140
rect 1030 32127 1048 32140
rect 1116 32127 1154 32140
rect 1154 32127 1172 32140
rect 1240 32127 1278 32140
rect 1278 32127 1296 32140
rect 868 32003 924 32059
rect 992 32016 1048 32059
rect 1116 32016 1172 32059
rect 1240 32016 1296 32059
rect 992 32003 1030 32016
rect 1030 32003 1048 32016
rect 1116 32003 1154 32016
rect 1154 32003 1172 32016
rect 1240 32003 1278 32016
rect 1278 32003 1296 32016
rect 868 31879 924 31935
rect 992 31892 1048 31935
rect 1116 31892 1172 31935
rect 1240 31892 1296 31935
rect 992 31879 1030 31892
rect 1030 31879 1048 31892
rect 1116 31879 1154 31892
rect 1154 31879 1172 31892
rect 1240 31879 1278 31892
rect 1278 31879 1296 31892
rect 868 31755 924 31811
rect 992 31768 1048 31811
rect 1116 31768 1172 31811
rect 1240 31768 1296 31811
rect 992 31755 1030 31768
rect 1030 31755 1048 31768
rect 1116 31755 1154 31768
rect 1154 31755 1172 31768
rect 1240 31755 1278 31768
rect 1278 31755 1296 31768
rect 868 31631 924 31687
rect 992 31644 1048 31687
rect 1116 31644 1172 31687
rect 1240 31644 1296 31687
rect 992 31631 1030 31644
rect 1030 31631 1048 31644
rect 1116 31631 1154 31644
rect 1154 31631 1172 31644
rect 1240 31631 1278 31644
rect 1278 31631 1296 31644
rect 868 31507 924 31563
rect 992 31520 1048 31563
rect 1116 31520 1172 31563
rect 1240 31520 1296 31563
rect 992 31507 1030 31520
rect 1030 31507 1048 31520
rect 1116 31507 1154 31520
rect 1154 31507 1172 31520
rect 1240 31507 1278 31520
rect 1278 31507 1296 31520
rect 868 31383 924 31439
rect 992 31396 1048 31439
rect 1116 31396 1172 31439
rect 1240 31396 1296 31439
rect 992 31383 1030 31396
rect 1030 31383 1048 31396
rect 1116 31383 1154 31396
rect 1154 31383 1172 31396
rect 1240 31383 1278 31396
rect 1278 31383 1296 31396
rect 868 31259 924 31315
rect 992 31272 1048 31315
rect 1116 31272 1172 31315
rect 1240 31272 1296 31315
rect 992 31259 1030 31272
rect 1030 31259 1048 31272
rect 1116 31259 1154 31272
rect 1154 31259 1172 31272
rect 1240 31259 1278 31272
rect 1278 31259 1296 31272
rect 868 31135 924 31191
rect 992 31148 1048 31191
rect 1116 31148 1172 31191
rect 1240 31148 1296 31191
rect 992 31135 1030 31148
rect 1030 31135 1048 31148
rect 1116 31135 1154 31148
rect 1154 31135 1172 31148
rect 1240 31135 1278 31148
rect 1278 31135 1296 31148
rect 868 31011 924 31067
rect 992 31024 1048 31067
rect 1116 31024 1172 31067
rect 1240 31024 1296 31067
rect 992 31011 1030 31024
rect 1030 31011 1048 31024
rect 1116 31011 1154 31024
rect 1154 31011 1172 31024
rect 1240 31011 1278 31024
rect 1278 31011 1296 31024
rect 868 30887 924 30943
rect 992 30900 1048 30943
rect 1116 30900 1172 30943
rect 1240 30900 1296 30943
rect 992 30887 1030 30900
rect 1030 30887 1048 30900
rect 1116 30887 1154 30900
rect 1154 30887 1172 30900
rect 1240 30887 1278 30900
rect 1278 30887 1296 30900
rect 868 30763 924 30819
rect 992 30776 1048 30819
rect 1116 30776 1172 30819
rect 1240 30776 1296 30819
rect 992 30763 1030 30776
rect 1030 30763 1048 30776
rect 1116 30763 1154 30776
rect 1154 30763 1172 30776
rect 1240 30763 1278 30776
rect 1278 30763 1296 30776
rect 868 30639 924 30695
rect 992 30652 1048 30695
rect 1116 30652 1172 30695
rect 1240 30652 1296 30695
rect 992 30639 1030 30652
rect 1030 30639 1048 30652
rect 1116 30639 1154 30652
rect 1154 30639 1172 30652
rect 1240 30639 1278 30652
rect 1278 30639 1296 30652
rect 868 30515 924 30571
rect 992 30528 1048 30571
rect 1116 30528 1172 30571
rect 1240 30528 1296 30571
rect 992 30515 1030 30528
rect 1030 30515 1048 30528
rect 1116 30515 1154 30528
rect 1154 30515 1172 30528
rect 1240 30515 1278 30528
rect 1278 30515 1296 30528
rect 868 30391 924 30447
rect 992 30404 1048 30447
rect 1116 30404 1172 30447
rect 1240 30404 1296 30447
rect 992 30391 1030 30404
rect 1030 30391 1048 30404
rect 1116 30391 1154 30404
rect 1154 30391 1172 30404
rect 1240 30391 1278 30404
rect 1278 30391 1296 30404
rect 868 30267 924 30323
rect 992 30280 1048 30323
rect 1116 30280 1172 30323
rect 1240 30280 1296 30323
rect 992 30267 1030 30280
rect 1030 30267 1048 30280
rect 1116 30267 1154 30280
rect 1154 30267 1172 30280
rect 1240 30267 1278 30280
rect 1278 30267 1296 30280
rect 868 30143 924 30199
rect 992 30156 1048 30199
rect 1116 30156 1172 30199
rect 1240 30156 1296 30199
rect 992 30143 1030 30156
rect 1030 30143 1048 30156
rect 1116 30143 1154 30156
rect 1154 30143 1172 30156
rect 1240 30143 1278 30156
rect 1278 30143 1296 30156
rect 868 29789 924 29845
rect 992 29789 1048 29845
rect 1116 29789 1172 29845
rect 1240 29789 1296 29845
rect 868 29665 924 29721
rect 992 29665 1048 29721
rect 1116 29665 1172 29721
rect 1240 29665 1296 29721
rect 868 29541 924 29597
rect 992 29541 1048 29597
rect 1116 29541 1172 29597
rect 1240 29541 1296 29597
rect 868 29417 924 29473
rect 992 29417 1048 29473
rect 1116 29417 1172 29473
rect 1240 29417 1296 29473
rect 868 29293 924 29349
rect 992 29293 1048 29349
rect 1116 29293 1172 29349
rect 1240 29293 1296 29349
rect 868 29169 924 29225
rect 992 29169 1048 29225
rect 1116 29169 1172 29225
rect 1240 29169 1296 29225
rect 868 29045 924 29101
rect 992 29045 1048 29101
rect 1116 29045 1172 29101
rect 1240 29045 1296 29101
rect 868 28921 924 28977
rect 992 28921 1048 28977
rect 1116 28921 1172 28977
rect 1240 28921 1296 28977
rect 868 28797 924 28853
rect 992 28797 1048 28853
rect 1116 28797 1172 28853
rect 1240 28797 1296 28853
rect 868 28673 924 28729
rect 992 28688 1048 28729
rect 1116 28688 1172 28729
rect 1240 28688 1296 28729
rect 992 28673 1030 28688
rect 1030 28673 1048 28688
rect 1116 28673 1154 28688
rect 1154 28673 1172 28688
rect 1240 28673 1278 28688
rect 1278 28673 1296 28688
rect 868 28549 924 28605
rect 992 28564 1048 28605
rect 1116 28564 1172 28605
rect 1240 28564 1296 28605
rect 992 28549 1030 28564
rect 1030 28549 1048 28564
rect 1116 28549 1154 28564
rect 1154 28549 1172 28564
rect 1240 28549 1278 28564
rect 1278 28549 1296 28564
rect 300 28189 356 28245
rect 424 28189 480 28245
rect 548 28189 604 28245
rect 672 28189 728 28245
rect 300 28065 356 28121
rect 424 28065 480 28121
rect 548 28065 604 28121
rect 672 28065 728 28121
rect 300 27941 356 27997
rect 424 27941 480 27997
rect 548 27941 604 27997
rect 672 27941 728 27997
rect 300 27817 356 27873
rect 424 27817 480 27873
rect 548 27817 604 27873
rect 672 27817 728 27873
rect 300 27693 356 27749
rect 424 27693 480 27749
rect 548 27693 604 27749
rect 672 27693 728 27749
rect 300 27569 356 27625
rect 424 27569 480 27625
rect 548 27569 604 27625
rect 672 27569 728 27625
rect 300 27445 356 27501
rect 424 27445 480 27501
rect 548 27445 604 27501
rect 672 27445 728 27501
rect 300 27321 356 27377
rect 424 27321 480 27377
rect 548 27321 604 27377
rect 672 27321 728 27377
rect 300 27197 356 27253
rect 424 27197 480 27253
rect 548 27197 604 27253
rect 672 27197 728 27253
rect 300 27073 356 27129
rect 424 27073 480 27129
rect 548 27073 604 27129
rect 672 27073 728 27129
rect 300 26949 356 27005
rect 424 26949 480 27005
rect 548 26949 604 27005
rect 672 26949 728 27005
rect 868 26595 924 26651
rect 992 26595 1048 26651
rect 1116 26595 1172 26651
rect 1240 26595 1296 26651
rect 868 26471 924 26527
rect 992 26471 1048 26527
rect 1116 26471 1172 26527
rect 1240 26471 1296 26527
rect 868 26347 924 26403
rect 992 26347 1048 26403
rect 1116 26347 1172 26403
rect 1240 26347 1296 26403
rect 868 26223 924 26279
rect 992 26223 1048 26279
rect 1116 26223 1172 26279
rect 1240 26223 1296 26279
rect 868 26099 924 26155
rect 992 26099 1048 26155
rect 1116 26099 1172 26155
rect 1240 26099 1296 26155
rect 868 25975 924 26031
rect 992 25975 1048 26031
rect 1116 25975 1172 26031
rect 1240 25975 1296 26031
rect 868 25851 924 25907
rect 992 25851 1048 25907
rect 1116 25851 1172 25907
rect 1240 25851 1296 25907
rect 868 25727 924 25783
rect 992 25727 1048 25783
rect 1116 25727 1172 25783
rect 1240 25727 1296 25783
rect 868 25603 924 25659
rect 992 25603 1048 25659
rect 1116 25603 1172 25659
rect 1240 25603 1296 25659
rect 868 25479 924 25535
rect 992 25479 1048 25535
rect 1116 25479 1172 25535
rect 1240 25479 1296 25535
rect 868 25355 924 25411
rect 992 25355 1048 25411
rect 1116 25355 1172 25411
rect 1240 25355 1296 25411
rect 868 25231 924 25287
rect 992 25231 1048 25287
rect 1116 25231 1172 25287
rect 1240 25231 1296 25287
rect 868 25107 924 25163
rect 992 25107 1048 25163
rect 1116 25107 1172 25163
rect 1240 25107 1296 25163
rect 868 24983 924 25039
rect 992 24983 1048 25039
rect 1116 24983 1172 25039
rect 1240 24983 1296 25039
rect 868 24859 924 24915
rect 992 24859 1048 24915
rect 1116 24859 1172 24915
rect 1240 24859 1296 24915
rect 868 24735 924 24791
rect 992 24740 1048 24791
rect 1116 24740 1172 24791
rect 1240 24740 1296 24791
rect 992 24735 1030 24740
rect 1030 24735 1048 24740
rect 1116 24735 1154 24740
rect 1154 24735 1172 24740
rect 1240 24735 1278 24740
rect 1278 24735 1296 24740
rect 868 24611 924 24667
rect 992 24616 1048 24667
rect 1116 24616 1172 24667
rect 1240 24616 1296 24667
rect 992 24611 1030 24616
rect 1030 24611 1048 24616
rect 1116 24611 1154 24616
rect 1154 24611 1172 24616
rect 1240 24611 1278 24616
rect 1278 24611 1296 24616
rect 868 24487 924 24543
rect 992 24492 1048 24543
rect 1116 24492 1172 24543
rect 1240 24492 1296 24543
rect 992 24487 1030 24492
rect 1030 24487 1048 24492
rect 1116 24487 1154 24492
rect 1154 24487 1172 24492
rect 1240 24487 1278 24492
rect 1278 24487 1296 24492
rect 868 24363 924 24419
rect 992 24368 1048 24419
rect 1116 24368 1172 24419
rect 1240 24368 1296 24419
rect 992 24363 1030 24368
rect 1030 24363 1048 24368
rect 1116 24363 1154 24368
rect 1154 24363 1172 24368
rect 1240 24363 1278 24368
rect 1278 24363 1296 24368
rect 868 24239 924 24295
rect 992 24244 1048 24295
rect 1116 24244 1172 24295
rect 1240 24244 1296 24295
rect 992 24239 1030 24244
rect 1030 24239 1048 24244
rect 1116 24239 1154 24244
rect 1154 24239 1172 24244
rect 1240 24239 1278 24244
rect 1278 24239 1296 24244
rect 868 24115 924 24171
rect 992 24120 1048 24171
rect 1116 24120 1172 24171
rect 1240 24120 1296 24171
rect 992 24115 1030 24120
rect 1030 24115 1048 24120
rect 1116 24115 1154 24120
rect 1154 24115 1172 24120
rect 1240 24115 1278 24120
rect 1278 24115 1296 24120
rect 868 23991 924 24047
rect 992 23996 1048 24047
rect 1116 23996 1172 24047
rect 1240 23996 1296 24047
rect 992 23991 1030 23996
rect 1030 23991 1048 23996
rect 1116 23991 1154 23996
rect 1154 23991 1172 23996
rect 1240 23991 1278 23996
rect 1278 23991 1296 23996
rect 868 23867 924 23923
rect 992 23872 1048 23923
rect 1116 23872 1172 23923
rect 1240 23872 1296 23923
rect 992 23867 1030 23872
rect 1030 23867 1048 23872
rect 1116 23867 1154 23872
rect 1154 23867 1172 23872
rect 1240 23867 1278 23872
rect 1278 23867 1296 23872
rect 868 23743 924 23799
rect 992 23748 1048 23799
rect 1116 23748 1172 23799
rect 1240 23748 1296 23799
rect 992 23743 1030 23748
rect 1030 23743 1048 23748
rect 1116 23743 1154 23748
rect 1154 23743 1172 23748
rect 1240 23743 1278 23748
rect 1278 23743 1296 23748
rect 868 23395 924 23451
rect 992 23448 1030 23451
rect 1030 23448 1048 23451
rect 1116 23448 1154 23451
rect 1154 23448 1172 23451
rect 1240 23448 1278 23451
rect 1278 23448 1296 23451
rect 992 23395 1048 23448
rect 1116 23395 1172 23448
rect 1240 23395 1296 23448
rect 868 23271 924 23327
rect 992 23324 1030 23327
rect 1030 23324 1048 23327
rect 1116 23324 1154 23327
rect 1154 23324 1172 23327
rect 1240 23324 1278 23327
rect 1278 23324 1296 23327
rect 992 23271 1048 23324
rect 1116 23271 1172 23324
rect 1240 23271 1296 23324
rect 868 23147 924 23203
rect 992 23200 1030 23203
rect 1030 23200 1048 23203
rect 1116 23200 1154 23203
rect 1154 23200 1172 23203
rect 1240 23200 1278 23203
rect 1278 23200 1296 23203
rect 992 23147 1048 23200
rect 1116 23147 1172 23200
rect 1240 23147 1296 23200
rect 868 23023 924 23079
rect 992 23076 1030 23079
rect 1030 23076 1048 23079
rect 1116 23076 1154 23079
rect 1154 23076 1172 23079
rect 1240 23076 1278 23079
rect 1278 23076 1296 23079
rect 992 23023 1048 23076
rect 1116 23023 1172 23076
rect 1240 23023 1296 23076
rect 868 22899 924 22955
rect 992 22952 1030 22955
rect 1030 22952 1048 22955
rect 1116 22952 1154 22955
rect 1154 22952 1172 22955
rect 1240 22952 1278 22955
rect 1278 22952 1296 22955
rect 992 22899 1048 22952
rect 1116 22899 1172 22952
rect 1240 22899 1296 22952
rect 868 22775 924 22831
rect 992 22828 1030 22831
rect 1030 22828 1048 22831
rect 1116 22828 1154 22831
rect 1154 22828 1172 22831
rect 1240 22828 1278 22831
rect 1278 22828 1296 22831
rect 992 22775 1048 22828
rect 1116 22775 1172 22828
rect 1240 22775 1296 22828
rect 868 22651 924 22707
rect 992 22704 1030 22707
rect 1030 22704 1048 22707
rect 1116 22704 1154 22707
rect 1154 22704 1172 22707
rect 1240 22704 1278 22707
rect 1278 22704 1296 22707
rect 992 22651 1048 22704
rect 1116 22651 1172 22704
rect 1240 22651 1296 22704
rect 868 22527 924 22583
rect 992 22580 1030 22583
rect 1030 22580 1048 22583
rect 1116 22580 1154 22583
rect 1154 22580 1172 22583
rect 1240 22580 1278 22583
rect 1278 22580 1296 22583
rect 992 22527 1048 22580
rect 1116 22527 1172 22580
rect 1240 22527 1296 22580
rect 868 22403 924 22459
rect 992 22456 1030 22459
rect 1030 22456 1048 22459
rect 1116 22456 1154 22459
rect 1154 22456 1172 22459
rect 1240 22456 1278 22459
rect 1278 22456 1296 22459
rect 992 22403 1048 22456
rect 1116 22403 1172 22456
rect 1240 22403 1296 22456
rect 868 22279 924 22335
rect 992 22332 1030 22335
rect 1030 22332 1048 22335
rect 1116 22332 1154 22335
rect 1154 22332 1172 22335
rect 1240 22332 1278 22335
rect 1278 22332 1296 22335
rect 992 22279 1048 22332
rect 1116 22279 1172 22332
rect 1240 22279 1296 22332
rect 868 22155 924 22211
rect 992 22208 1030 22211
rect 1030 22208 1048 22211
rect 1116 22208 1154 22211
rect 1154 22208 1172 22211
rect 1240 22208 1278 22211
rect 1278 22208 1296 22211
rect 992 22155 1048 22208
rect 1116 22155 1172 22208
rect 1240 22155 1296 22208
rect 868 22031 924 22087
rect 992 22084 1030 22087
rect 1030 22084 1048 22087
rect 1116 22084 1154 22087
rect 1154 22084 1172 22087
rect 1240 22084 1278 22087
rect 1278 22084 1296 22087
rect 992 22031 1048 22084
rect 1116 22031 1172 22084
rect 1240 22031 1296 22084
rect 868 21907 924 21963
rect 992 21960 1030 21963
rect 1030 21960 1048 21963
rect 1116 21960 1154 21963
rect 1154 21960 1172 21963
rect 1240 21960 1278 21963
rect 1278 21960 1296 21963
rect 992 21907 1048 21960
rect 1116 21907 1172 21960
rect 1240 21907 1296 21960
rect 868 21783 924 21839
rect 992 21836 1030 21839
rect 1030 21836 1048 21839
rect 1116 21836 1154 21839
rect 1154 21836 1172 21839
rect 1240 21836 1278 21839
rect 1278 21836 1296 21839
rect 992 21783 1048 21836
rect 1116 21783 1172 21836
rect 1240 21783 1296 21836
rect 868 21659 924 21715
rect 992 21712 1030 21715
rect 1030 21712 1048 21715
rect 1116 21712 1154 21715
rect 1154 21712 1172 21715
rect 1240 21712 1278 21715
rect 1278 21712 1296 21715
rect 992 21659 1048 21712
rect 1116 21659 1172 21712
rect 1240 21659 1296 21712
rect 868 21535 924 21591
rect 992 21588 1030 21591
rect 1030 21588 1048 21591
rect 1116 21588 1154 21591
rect 1154 21588 1172 21591
rect 1240 21588 1278 21591
rect 1278 21588 1296 21591
rect 992 21535 1048 21588
rect 1116 21535 1172 21588
rect 1240 21535 1296 21588
rect 868 21411 924 21467
rect 992 21411 1048 21467
rect 1116 21411 1172 21467
rect 1240 21411 1296 21467
rect 868 21287 924 21343
rect 992 21287 1048 21343
rect 1116 21287 1172 21343
rect 1240 21287 1296 21343
rect 868 21163 924 21219
rect 992 21163 1048 21219
rect 1116 21163 1172 21219
rect 1240 21163 1296 21219
rect 868 21039 924 21095
rect 992 21039 1048 21095
rect 1116 21039 1172 21095
rect 1240 21039 1296 21095
rect 868 20915 924 20971
rect 992 20915 1048 20971
rect 1116 20915 1172 20971
rect 1240 20915 1296 20971
rect 868 20791 924 20847
rect 992 20791 1048 20847
rect 1116 20791 1172 20847
rect 1240 20791 1296 20847
rect 868 20667 924 20723
rect 992 20667 1048 20723
rect 1116 20667 1172 20723
rect 1240 20667 1296 20723
rect 868 20543 924 20599
rect 992 20543 1048 20599
rect 1116 20543 1172 20599
rect 1240 20543 1296 20599
rect 868 20195 924 20251
rect 992 20195 1048 20251
rect 1116 20195 1172 20251
rect 1240 20195 1296 20251
rect 868 20071 924 20127
rect 992 20071 1048 20127
rect 1116 20071 1172 20127
rect 1240 20071 1296 20127
rect 868 19947 924 20003
rect 992 19947 1048 20003
rect 1116 19947 1172 20003
rect 1240 19947 1296 20003
rect 868 19823 924 19879
rect 992 19823 1048 19879
rect 1116 19823 1172 19879
rect 1240 19823 1296 19879
rect 868 19699 924 19755
rect 992 19699 1048 19755
rect 1116 19699 1172 19755
rect 1240 19699 1296 19755
rect 868 19575 924 19631
rect 992 19575 1048 19631
rect 1116 19575 1172 19631
rect 1240 19575 1296 19631
rect 868 19451 924 19507
rect 992 19451 1048 19507
rect 1116 19451 1172 19507
rect 1240 19451 1296 19507
rect 868 19327 924 19383
rect 992 19327 1048 19383
rect 1116 19327 1172 19383
rect 1240 19327 1296 19383
rect 868 19203 924 19259
rect 992 19203 1048 19259
rect 1116 19203 1172 19259
rect 1240 19203 1296 19259
rect 868 19079 924 19135
rect 992 19079 1048 19135
rect 1116 19079 1172 19135
rect 1240 19079 1296 19135
rect 868 18955 924 19011
rect 992 18955 1048 19011
rect 1116 18955 1172 19011
rect 1240 18955 1296 19011
rect 868 18831 924 18887
rect 992 18831 1048 18887
rect 1116 18831 1172 18887
rect 1240 18831 1296 18887
rect 868 18707 924 18763
rect 992 18707 1048 18763
rect 1116 18707 1172 18763
rect 1240 18707 1296 18763
rect 868 18583 924 18639
rect 992 18583 1048 18639
rect 1116 18583 1172 18639
rect 1240 18583 1296 18639
rect 868 18459 924 18515
rect 992 18459 1048 18515
rect 1116 18459 1172 18515
rect 1240 18459 1296 18515
rect 868 18335 924 18391
rect 992 18335 1048 18391
rect 1116 18335 1172 18391
rect 1240 18335 1296 18391
rect 868 18211 924 18267
rect 992 18211 1048 18267
rect 1116 18211 1172 18267
rect 1240 18211 1296 18267
rect 868 18087 924 18143
rect 992 18087 1048 18143
rect 1116 18087 1172 18143
rect 1240 18087 1296 18143
rect 868 17963 924 18019
rect 992 17963 1048 18019
rect 1116 17963 1172 18019
rect 1240 17963 1296 18019
rect 868 17839 924 17895
rect 992 17839 1048 17895
rect 1116 17839 1172 17895
rect 1240 17839 1296 17895
rect 868 17715 924 17771
rect 992 17715 1048 17771
rect 1116 17715 1172 17771
rect 1240 17715 1296 17771
rect 868 17591 924 17647
rect 992 17591 1048 17647
rect 1116 17591 1172 17647
rect 1240 17591 1296 17647
rect 868 17467 924 17523
rect 992 17467 1048 17523
rect 1116 17467 1172 17523
rect 1240 17467 1296 17523
rect 868 17343 924 17399
rect 992 17343 1048 17399
rect 1116 17343 1172 17399
rect 1240 17343 1296 17399
rect 868 16995 924 17051
rect 992 16995 1048 17051
rect 1116 16995 1172 17051
rect 1240 16995 1296 17051
rect 868 16871 924 16927
rect 992 16871 1048 16927
rect 1116 16871 1172 16927
rect 1240 16871 1296 16927
rect 868 16747 924 16803
rect 992 16747 1048 16803
rect 1116 16747 1172 16803
rect 1240 16747 1296 16803
rect 868 16623 924 16679
rect 992 16623 1048 16679
rect 1116 16623 1172 16679
rect 1240 16623 1296 16679
rect 868 16499 924 16555
rect 992 16499 1048 16555
rect 1116 16499 1172 16555
rect 1240 16499 1296 16555
rect 868 16375 924 16431
rect 992 16375 1048 16431
rect 1116 16375 1172 16431
rect 1240 16375 1296 16431
rect 868 16251 924 16307
rect 992 16251 1048 16307
rect 1116 16251 1172 16307
rect 1240 16251 1296 16307
rect 868 16127 924 16183
rect 992 16127 1048 16183
rect 1116 16127 1172 16183
rect 1240 16127 1296 16183
rect 868 16003 924 16059
rect 992 16003 1048 16059
rect 1116 16003 1172 16059
rect 1240 16003 1296 16059
rect 868 15879 924 15935
rect 992 15879 1048 15935
rect 1116 15879 1172 15935
rect 1240 15879 1296 15935
rect 868 15755 924 15811
rect 992 15755 1048 15811
rect 1116 15755 1172 15811
rect 1240 15755 1296 15811
rect 1436 53048 1492 53101
rect 1436 53045 1438 53048
rect 1438 53045 1490 53048
rect 1490 53045 1492 53048
rect 1560 53048 1616 53101
rect 1560 53045 1562 53048
rect 1562 53045 1614 53048
rect 1614 53045 1616 53048
rect 1684 53048 1740 53101
rect 1684 53045 1686 53048
rect 1686 53045 1738 53048
rect 1738 53045 1740 53048
rect 1808 53048 1864 53101
rect 1808 53045 1810 53048
rect 1810 53045 1862 53048
rect 1862 53045 1864 53048
rect 1436 52924 1492 52977
rect 1436 52921 1438 52924
rect 1438 52921 1490 52924
rect 1490 52921 1492 52924
rect 1560 52924 1616 52977
rect 1560 52921 1562 52924
rect 1562 52921 1614 52924
rect 1614 52921 1616 52924
rect 1684 52924 1740 52977
rect 1684 52921 1686 52924
rect 1686 52921 1738 52924
rect 1738 52921 1740 52924
rect 1808 52924 1864 52977
rect 1808 52921 1810 52924
rect 1810 52921 1862 52924
rect 1862 52921 1864 52924
rect 1436 52800 1492 52853
rect 1436 52797 1438 52800
rect 1438 52797 1490 52800
rect 1490 52797 1492 52800
rect 1560 52800 1616 52853
rect 1560 52797 1562 52800
rect 1562 52797 1614 52800
rect 1614 52797 1616 52800
rect 1684 52800 1740 52853
rect 1684 52797 1686 52800
rect 1686 52797 1738 52800
rect 1738 52797 1740 52800
rect 1808 52800 1864 52853
rect 1808 52797 1810 52800
rect 1810 52797 1862 52800
rect 1862 52797 1864 52800
rect 1436 52676 1492 52729
rect 1436 52673 1438 52676
rect 1438 52673 1490 52676
rect 1490 52673 1492 52676
rect 1560 52676 1616 52729
rect 1560 52673 1562 52676
rect 1562 52673 1614 52676
rect 1614 52673 1616 52676
rect 1684 52676 1740 52729
rect 1684 52673 1686 52676
rect 1686 52673 1738 52676
rect 1738 52673 1740 52676
rect 1808 52676 1864 52729
rect 1808 52673 1810 52676
rect 1810 52673 1862 52676
rect 1862 52673 1864 52676
rect 1436 52552 1492 52605
rect 1436 52549 1438 52552
rect 1438 52549 1490 52552
rect 1490 52549 1492 52552
rect 1560 52552 1616 52605
rect 1560 52549 1562 52552
rect 1562 52549 1614 52552
rect 1614 52549 1616 52552
rect 1684 52552 1740 52605
rect 1684 52549 1686 52552
rect 1686 52549 1738 52552
rect 1738 52549 1740 52552
rect 1808 52552 1864 52605
rect 1808 52549 1810 52552
rect 1810 52549 1862 52552
rect 1862 52549 1864 52552
rect 1436 48989 1492 49045
rect 1560 48989 1616 49045
rect 1684 48989 1740 49045
rect 1808 48989 1864 49045
rect 1436 48865 1492 48921
rect 1560 48865 1616 48921
rect 1684 48865 1740 48921
rect 1808 48865 1864 48921
rect 1436 48741 1492 48797
rect 1560 48741 1616 48797
rect 1684 48741 1740 48797
rect 1808 48741 1864 48797
rect 1436 48617 1492 48673
rect 1560 48617 1616 48673
rect 1684 48617 1740 48673
rect 1808 48617 1864 48673
rect 1436 48493 1492 48549
rect 1560 48493 1616 48549
rect 1684 48493 1740 48549
rect 1808 48493 1864 48549
rect 1436 48369 1492 48425
rect 1560 48369 1616 48425
rect 1684 48369 1740 48425
rect 1808 48369 1864 48425
rect 1436 48245 1492 48301
rect 1560 48245 1616 48301
rect 1684 48245 1740 48301
rect 1808 48245 1864 48301
rect 1436 48121 1492 48177
rect 1560 48121 1616 48177
rect 1684 48121 1740 48177
rect 1808 48121 1864 48177
rect 1436 47997 1492 48053
rect 1560 47997 1616 48053
rect 1684 47997 1740 48053
rect 1808 47997 1864 48053
rect 1436 47873 1492 47929
rect 1560 47873 1616 47929
rect 1684 47873 1740 47929
rect 1808 47873 1864 47929
rect 1436 47749 1492 47805
rect 1560 47749 1616 47805
rect 1684 47749 1740 47805
rect 1808 47749 1864 47805
rect 1436 45789 1492 45845
rect 1560 45789 1616 45845
rect 1684 45789 1740 45845
rect 1808 45789 1864 45845
rect 1436 45665 1492 45721
rect 1560 45665 1616 45721
rect 1684 45665 1740 45721
rect 1808 45665 1864 45721
rect 1436 45541 1492 45597
rect 1560 45541 1616 45597
rect 1684 45541 1740 45597
rect 1808 45541 1864 45597
rect 1436 45417 1492 45473
rect 1560 45417 1616 45473
rect 1684 45417 1740 45473
rect 1808 45417 1864 45473
rect 1436 45293 1492 45349
rect 1560 45293 1616 45349
rect 1684 45293 1740 45349
rect 1808 45293 1864 45349
rect 1436 45169 1492 45225
rect 1560 45169 1616 45225
rect 1684 45169 1740 45225
rect 1808 45169 1864 45225
rect 1436 45100 1438 45101
rect 1438 45100 1490 45101
rect 1490 45100 1492 45101
rect 1436 45045 1492 45100
rect 1560 45100 1562 45101
rect 1562 45100 1614 45101
rect 1614 45100 1616 45101
rect 1560 45045 1616 45100
rect 1684 45100 1686 45101
rect 1686 45100 1738 45101
rect 1738 45100 1740 45101
rect 1684 45045 1740 45100
rect 1808 45100 1810 45101
rect 1810 45100 1862 45101
rect 1862 45100 1864 45101
rect 1808 45045 1864 45100
rect 1436 44976 1438 44977
rect 1438 44976 1490 44977
rect 1490 44976 1492 44977
rect 1436 44921 1492 44976
rect 1560 44976 1562 44977
rect 1562 44976 1614 44977
rect 1614 44976 1616 44977
rect 1560 44921 1616 44976
rect 1684 44976 1686 44977
rect 1686 44976 1738 44977
rect 1738 44976 1740 44977
rect 1684 44921 1740 44976
rect 1808 44976 1810 44977
rect 1810 44976 1862 44977
rect 1862 44976 1864 44977
rect 1808 44921 1864 44976
rect 1436 44852 1438 44853
rect 1438 44852 1490 44853
rect 1490 44852 1492 44853
rect 1436 44797 1492 44852
rect 1560 44852 1562 44853
rect 1562 44852 1614 44853
rect 1614 44852 1616 44853
rect 1560 44797 1616 44852
rect 1684 44852 1686 44853
rect 1686 44852 1738 44853
rect 1738 44852 1740 44853
rect 1684 44797 1740 44852
rect 1808 44852 1810 44853
rect 1810 44852 1862 44853
rect 1862 44852 1864 44853
rect 1808 44797 1864 44852
rect 1436 44728 1438 44729
rect 1438 44728 1490 44729
rect 1490 44728 1492 44729
rect 1436 44673 1492 44728
rect 1560 44728 1562 44729
rect 1562 44728 1614 44729
rect 1614 44728 1616 44729
rect 1560 44673 1616 44728
rect 1684 44728 1686 44729
rect 1686 44728 1738 44729
rect 1738 44728 1740 44729
rect 1684 44673 1740 44728
rect 1808 44728 1810 44729
rect 1810 44728 1862 44729
rect 1862 44728 1864 44729
rect 1808 44673 1864 44728
rect 1436 44604 1438 44605
rect 1438 44604 1490 44605
rect 1490 44604 1492 44605
rect 1436 44549 1492 44604
rect 1560 44604 1562 44605
rect 1562 44604 1614 44605
rect 1614 44604 1616 44605
rect 1560 44549 1616 44604
rect 1684 44604 1686 44605
rect 1686 44604 1738 44605
rect 1738 44604 1740 44605
rect 1684 44549 1740 44604
rect 1808 44604 1810 44605
rect 1810 44604 1862 44605
rect 1862 44604 1864 44605
rect 1808 44549 1864 44604
rect 1436 36195 1492 36251
rect 1560 36195 1616 36251
rect 1684 36195 1740 36251
rect 1808 36195 1864 36251
rect 1436 36071 1492 36127
rect 1560 36071 1616 36127
rect 1684 36071 1740 36127
rect 1808 36071 1864 36127
rect 1436 35947 1492 36003
rect 1560 35947 1616 36003
rect 1684 35947 1740 36003
rect 1808 35947 1864 36003
rect 1436 35823 1492 35879
rect 1560 35823 1616 35879
rect 1684 35823 1740 35879
rect 1808 35823 1864 35879
rect 1436 35699 1492 35755
rect 1560 35699 1616 35755
rect 1684 35699 1740 35755
rect 1808 35699 1864 35755
rect 1436 35575 1492 35631
rect 1560 35575 1616 35631
rect 1684 35575 1740 35631
rect 1808 35575 1864 35631
rect 1436 35451 1492 35507
rect 1560 35451 1616 35507
rect 1684 35451 1740 35507
rect 1808 35451 1864 35507
rect 1436 35327 1492 35383
rect 1560 35327 1616 35383
rect 1684 35327 1740 35383
rect 1808 35327 1864 35383
rect 1436 35203 1492 35259
rect 1560 35203 1616 35259
rect 1684 35203 1740 35259
rect 1808 35203 1864 35259
rect 1436 35079 1492 35135
rect 1560 35079 1616 35135
rect 1684 35079 1740 35135
rect 1808 35079 1864 35135
rect 1436 34955 1492 35011
rect 1560 34955 1616 35011
rect 1684 34955 1740 35011
rect 1808 34955 1864 35011
rect 1436 34831 1492 34887
rect 1560 34831 1616 34887
rect 1684 34831 1740 34887
rect 1808 34831 1864 34887
rect 1436 34707 1492 34763
rect 1560 34707 1616 34763
rect 1684 34707 1740 34763
rect 1808 34707 1864 34763
rect 1436 34583 1492 34639
rect 1560 34583 1616 34639
rect 1684 34583 1740 34639
rect 1808 34583 1864 34639
rect 1436 34459 1492 34515
rect 1560 34459 1616 34515
rect 1684 34459 1740 34515
rect 1808 34459 1864 34515
rect 1436 34335 1492 34391
rect 1560 34335 1616 34391
rect 1684 34335 1740 34391
rect 1808 34335 1864 34391
rect 1436 34211 1492 34267
rect 1560 34211 1616 34267
rect 1684 34211 1740 34267
rect 1808 34211 1864 34267
rect 1436 34087 1492 34143
rect 1560 34087 1616 34143
rect 1684 34087 1740 34143
rect 1808 34087 1864 34143
rect 1436 33963 1492 34019
rect 1560 33963 1616 34019
rect 1684 33963 1740 34019
rect 1808 33963 1864 34019
rect 1436 33839 1492 33895
rect 1560 33839 1616 33895
rect 1684 33839 1740 33895
rect 1808 33839 1864 33895
rect 1436 33715 1492 33771
rect 1560 33715 1616 33771
rect 1684 33715 1740 33771
rect 1808 33715 1864 33771
rect 1436 33591 1492 33647
rect 1560 33591 1616 33647
rect 1684 33591 1740 33647
rect 1808 33591 1864 33647
rect 1436 33467 1492 33523
rect 1560 33467 1616 33523
rect 1684 33467 1740 33523
rect 1808 33467 1864 33523
rect 1436 33343 1492 33399
rect 1560 33343 1616 33399
rect 1684 33343 1740 33399
rect 1808 33343 1864 33399
rect 1436 28189 1492 28245
rect 1560 28189 1616 28245
rect 1684 28189 1740 28245
rect 1808 28189 1864 28245
rect 1436 28065 1492 28121
rect 1560 28065 1616 28121
rect 1684 28065 1740 28121
rect 1808 28065 1864 28121
rect 1436 27941 1492 27997
rect 1560 27941 1616 27997
rect 1684 27941 1740 27997
rect 1808 27941 1864 27997
rect 1436 27817 1492 27873
rect 1560 27817 1616 27873
rect 1684 27817 1740 27873
rect 1808 27817 1864 27873
rect 1436 27693 1492 27749
rect 1560 27693 1616 27749
rect 1684 27693 1740 27749
rect 1808 27693 1864 27749
rect 1436 27569 1492 27625
rect 1560 27569 1616 27625
rect 1684 27569 1740 27625
rect 1808 27569 1864 27625
rect 1436 27445 1492 27501
rect 1560 27445 1616 27501
rect 1684 27445 1740 27501
rect 1808 27445 1864 27501
rect 1436 27321 1492 27377
rect 1560 27321 1616 27377
rect 1684 27321 1740 27377
rect 1808 27321 1864 27377
rect 1436 27197 1492 27253
rect 1560 27197 1616 27253
rect 1684 27197 1740 27253
rect 1808 27197 1864 27253
rect 1436 27073 1492 27129
rect 1560 27073 1616 27129
rect 1684 27073 1740 27129
rect 1808 27073 1864 27129
rect 1436 26949 1492 27005
rect 1560 26949 1616 27005
rect 1684 26949 1740 27005
rect 1808 26949 1864 27005
rect 2004 55389 2060 55445
rect 2128 55389 2184 55445
rect 2252 55389 2308 55445
rect 2376 55389 2432 55445
rect 2004 55265 2060 55321
rect 2128 55265 2184 55321
rect 2252 55265 2308 55321
rect 2376 55265 2432 55321
rect 2004 55141 2060 55197
rect 2128 55141 2184 55197
rect 2252 55141 2308 55197
rect 2376 55141 2432 55197
rect 2004 55017 2060 55073
rect 2128 55017 2184 55073
rect 2252 55017 2308 55073
rect 2376 55017 2432 55073
rect 2004 54893 2060 54949
rect 2128 54893 2184 54949
rect 2252 54893 2308 54949
rect 2376 54893 2432 54949
rect 2004 54769 2060 54825
rect 2128 54769 2184 54825
rect 2252 54769 2308 54825
rect 2376 54769 2432 54825
rect 2004 54645 2060 54701
rect 2128 54645 2184 54701
rect 2252 54645 2308 54701
rect 2376 54645 2432 54701
rect 2004 54521 2060 54577
rect 2128 54521 2184 54577
rect 2252 54521 2308 54577
rect 2376 54521 2432 54577
rect 2004 54397 2060 54453
rect 2128 54397 2184 54453
rect 2252 54397 2308 54453
rect 2376 54397 2432 54453
rect 2004 54273 2060 54329
rect 2128 54273 2184 54329
rect 2252 54273 2308 54329
rect 2376 54273 2432 54329
rect 2004 54149 2060 54205
rect 2128 54149 2184 54205
rect 2252 54149 2308 54205
rect 2376 54149 2432 54205
rect 2004 47389 2060 47445
rect 2128 47389 2184 47445
rect 2252 47389 2308 47445
rect 2376 47389 2432 47445
rect 2004 47265 2060 47321
rect 2128 47265 2184 47321
rect 2252 47265 2308 47321
rect 2376 47265 2432 47321
rect 2004 47141 2060 47197
rect 2128 47141 2184 47197
rect 2252 47141 2308 47197
rect 2376 47141 2432 47197
rect 2004 47017 2060 47073
rect 2128 47017 2184 47073
rect 2252 47017 2308 47073
rect 2376 47017 2432 47073
rect 2004 46893 2060 46949
rect 2128 46893 2184 46949
rect 2252 46893 2308 46949
rect 2376 46893 2432 46949
rect 2004 46769 2060 46825
rect 2128 46769 2184 46825
rect 2252 46769 2308 46825
rect 2376 46769 2432 46825
rect 2004 46645 2060 46701
rect 2128 46645 2184 46701
rect 2252 46645 2308 46701
rect 2376 46645 2432 46701
rect 2004 46521 2060 46577
rect 2128 46521 2184 46577
rect 2252 46521 2308 46577
rect 2376 46521 2432 46577
rect 2004 46397 2060 46453
rect 2128 46397 2184 46453
rect 2252 46397 2308 46453
rect 2376 46397 2432 46453
rect 2004 46273 2060 46329
rect 2128 46273 2184 46329
rect 2252 46273 2308 46329
rect 2376 46273 2432 46329
rect 2004 46149 2060 46205
rect 2128 46149 2184 46205
rect 2252 46149 2308 46205
rect 2376 46149 2432 46205
rect 2004 44189 2060 44245
rect 2128 44189 2184 44245
rect 2252 44189 2308 44245
rect 2376 44189 2432 44245
rect 2004 44065 2060 44121
rect 2128 44065 2184 44121
rect 2252 44065 2308 44121
rect 2376 44065 2432 44121
rect 2004 43941 2060 43997
rect 2128 43941 2184 43997
rect 2252 43941 2308 43997
rect 2376 43941 2432 43997
rect 2004 43817 2060 43873
rect 2128 43817 2184 43873
rect 2252 43817 2308 43873
rect 2376 43817 2432 43873
rect 2004 43693 2060 43749
rect 2128 43693 2184 43749
rect 2252 43693 2308 43749
rect 2376 43693 2432 43749
rect 2004 43569 2060 43625
rect 2128 43569 2184 43625
rect 2252 43569 2308 43625
rect 2376 43569 2432 43625
rect 2004 43445 2060 43501
rect 2128 43445 2184 43501
rect 2252 43445 2308 43501
rect 2376 43445 2432 43501
rect 2004 43321 2060 43377
rect 2128 43321 2184 43377
rect 2252 43321 2308 43377
rect 2376 43321 2432 43377
rect 2004 43197 2060 43253
rect 2128 43197 2184 43253
rect 2252 43197 2308 43253
rect 2376 43197 2432 43253
rect 2004 43073 2060 43129
rect 2128 43073 2184 43129
rect 2252 43073 2308 43129
rect 2376 43073 2432 43129
rect 2004 42949 2060 43005
rect 2128 42949 2184 43005
rect 2252 42949 2308 43005
rect 2376 42949 2432 43005
rect 2004 42589 2060 42645
rect 2128 42589 2184 42645
rect 2252 42589 2308 42645
rect 2376 42589 2432 42645
rect 2004 42465 2060 42521
rect 2128 42465 2184 42521
rect 2252 42465 2308 42521
rect 2376 42465 2432 42521
rect 2004 42341 2060 42397
rect 2128 42341 2184 42397
rect 2252 42341 2308 42397
rect 2376 42341 2432 42397
rect 2004 42217 2060 42273
rect 2128 42217 2184 42273
rect 2252 42217 2308 42273
rect 2376 42217 2432 42273
rect 2004 42093 2060 42149
rect 2128 42093 2184 42149
rect 2252 42093 2308 42149
rect 2376 42093 2432 42149
rect 2004 41969 2060 42025
rect 2128 41969 2184 42025
rect 2252 41969 2308 42025
rect 2376 41969 2432 42025
rect 2004 41845 2060 41901
rect 2128 41845 2184 41901
rect 2252 41845 2308 41901
rect 2376 41845 2432 41901
rect 2004 41721 2060 41777
rect 2128 41721 2184 41777
rect 2252 41721 2308 41777
rect 2376 41721 2432 41777
rect 2004 41597 2060 41653
rect 2128 41597 2184 41653
rect 2252 41597 2308 41653
rect 2376 41597 2432 41653
rect 2004 41473 2060 41529
rect 2128 41473 2184 41529
rect 2252 41473 2308 41529
rect 2376 41473 2432 41529
rect 2004 41349 2060 41405
rect 2128 41349 2184 41405
rect 2252 41349 2308 41405
rect 2376 41349 2432 41405
rect 2004 40989 2060 41045
rect 2128 40989 2184 41045
rect 2252 40989 2308 41045
rect 2376 40989 2432 41045
rect 2004 40865 2060 40921
rect 2128 40865 2184 40921
rect 2252 40865 2308 40921
rect 2376 40865 2432 40921
rect 2004 40741 2060 40797
rect 2128 40741 2184 40797
rect 2252 40741 2308 40797
rect 2376 40741 2432 40797
rect 2004 40617 2060 40673
rect 2128 40617 2184 40673
rect 2252 40617 2308 40673
rect 2376 40617 2432 40673
rect 2004 40493 2060 40549
rect 2128 40493 2184 40549
rect 2252 40493 2308 40549
rect 2376 40493 2432 40549
rect 2004 40369 2060 40425
rect 2128 40369 2184 40425
rect 2252 40369 2308 40425
rect 2376 40369 2432 40425
rect 2004 40245 2060 40301
rect 2128 40245 2184 40301
rect 2252 40245 2308 40301
rect 2376 40245 2432 40301
rect 2004 40121 2060 40177
rect 2128 40121 2184 40177
rect 2252 40121 2308 40177
rect 2376 40121 2432 40177
rect 2004 39997 2060 40053
rect 2128 39997 2184 40053
rect 2252 39997 2308 40053
rect 2376 39997 2432 40053
rect 2004 39873 2060 39929
rect 2128 39873 2184 39929
rect 2252 39873 2308 39929
rect 2376 39873 2432 39929
rect 2004 39749 2060 39805
rect 2128 39749 2184 39805
rect 2252 39749 2308 39805
rect 2376 39749 2432 39805
rect 2004 32995 2060 33051
rect 2128 32995 2184 33051
rect 2252 32995 2308 33051
rect 2376 32995 2432 33051
rect 2004 32871 2060 32927
rect 2128 32871 2184 32927
rect 2252 32871 2308 32927
rect 2376 32871 2432 32927
rect 2004 32747 2060 32803
rect 2128 32747 2184 32803
rect 2252 32747 2308 32803
rect 2376 32747 2432 32803
rect 2004 32623 2060 32679
rect 2128 32623 2184 32679
rect 2252 32623 2308 32679
rect 2376 32623 2432 32679
rect 2004 32499 2060 32555
rect 2128 32499 2184 32555
rect 2252 32499 2308 32555
rect 2376 32499 2432 32555
rect 2004 32375 2060 32431
rect 2128 32375 2184 32431
rect 2252 32375 2308 32431
rect 2376 32375 2432 32431
rect 2004 32251 2060 32307
rect 2128 32251 2184 32307
rect 2252 32251 2308 32307
rect 2376 32251 2432 32307
rect 2004 32127 2060 32183
rect 2128 32127 2184 32183
rect 2252 32127 2308 32183
rect 2376 32127 2432 32183
rect 2004 32003 2060 32059
rect 2128 32003 2184 32059
rect 2252 32003 2308 32059
rect 2376 32003 2432 32059
rect 2004 31879 2060 31935
rect 2128 31879 2184 31935
rect 2252 31879 2308 31935
rect 2376 31879 2432 31935
rect 2004 31755 2060 31811
rect 2128 31755 2184 31811
rect 2252 31755 2308 31811
rect 2376 31755 2432 31811
rect 2004 31631 2060 31687
rect 2128 31631 2184 31687
rect 2252 31631 2308 31687
rect 2376 31631 2432 31687
rect 2004 31507 2060 31563
rect 2128 31507 2184 31563
rect 2252 31507 2308 31563
rect 2376 31507 2432 31563
rect 2004 31383 2060 31439
rect 2128 31383 2184 31439
rect 2252 31383 2308 31439
rect 2376 31383 2432 31439
rect 2004 31259 2060 31315
rect 2128 31259 2184 31315
rect 2252 31259 2308 31315
rect 2376 31259 2432 31315
rect 2004 31135 2060 31191
rect 2128 31135 2184 31191
rect 2252 31135 2308 31191
rect 2376 31135 2432 31191
rect 2004 31011 2060 31067
rect 2128 31011 2184 31067
rect 2252 31011 2308 31067
rect 2376 31011 2432 31067
rect 2004 30887 2060 30943
rect 2128 30887 2184 30943
rect 2252 30887 2308 30943
rect 2376 30887 2432 30943
rect 2004 30763 2060 30819
rect 2128 30763 2184 30819
rect 2252 30763 2308 30819
rect 2376 30763 2432 30819
rect 2004 30639 2060 30695
rect 2128 30639 2184 30695
rect 2252 30639 2308 30695
rect 2376 30639 2432 30695
rect 2004 30515 2060 30571
rect 2128 30515 2184 30571
rect 2252 30515 2308 30571
rect 2376 30515 2432 30571
rect 2004 30391 2060 30447
rect 2128 30391 2184 30447
rect 2252 30391 2308 30447
rect 2376 30391 2432 30447
rect 2004 30267 2060 30323
rect 2128 30267 2184 30323
rect 2252 30267 2308 30323
rect 2376 30267 2432 30323
rect 2004 30143 2060 30199
rect 2128 30143 2184 30199
rect 2252 30143 2308 30199
rect 2376 30143 2432 30199
rect 2004 29789 2060 29845
rect 2128 29789 2184 29845
rect 2252 29789 2308 29845
rect 2376 29789 2432 29845
rect 2004 29665 2060 29721
rect 2128 29665 2184 29721
rect 2252 29665 2308 29721
rect 2376 29665 2432 29721
rect 2004 29541 2060 29597
rect 2128 29541 2184 29597
rect 2252 29541 2308 29597
rect 2376 29541 2432 29597
rect 2004 29417 2060 29473
rect 2128 29417 2184 29473
rect 2252 29417 2308 29473
rect 2376 29417 2432 29473
rect 2004 29293 2060 29349
rect 2128 29293 2184 29349
rect 2252 29293 2308 29349
rect 2376 29293 2432 29349
rect 2004 29169 2060 29225
rect 2128 29169 2184 29225
rect 2252 29169 2308 29225
rect 2376 29169 2432 29225
rect 2004 29045 2060 29101
rect 2128 29045 2184 29101
rect 2252 29045 2308 29101
rect 2376 29045 2432 29101
rect 2004 28921 2060 28977
rect 2128 28921 2184 28977
rect 2252 28921 2308 28977
rect 2376 28921 2432 28977
rect 2004 28797 2060 28853
rect 2128 28797 2184 28853
rect 2252 28797 2308 28853
rect 2376 28797 2432 28853
rect 2004 28673 2060 28729
rect 2128 28673 2184 28729
rect 2252 28673 2308 28729
rect 2376 28673 2432 28729
rect 2004 28549 2060 28605
rect 2128 28549 2184 28605
rect 2252 28549 2308 28605
rect 2376 28549 2432 28605
rect 2004 26595 2060 26651
rect 2128 26595 2184 26651
rect 2252 26595 2308 26651
rect 2376 26595 2432 26651
rect 2004 26471 2060 26527
rect 2128 26471 2184 26527
rect 2252 26471 2308 26527
rect 2376 26471 2432 26527
rect 2004 26347 2060 26403
rect 2128 26347 2184 26403
rect 2252 26347 2308 26403
rect 2376 26347 2432 26403
rect 2004 26223 2060 26279
rect 2128 26223 2184 26279
rect 2252 26223 2308 26279
rect 2376 26223 2432 26279
rect 2004 26099 2060 26155
rect 2128 26099 2184 26155
rect 2252 26099 2308 26155
rect 2376 26099 2432 26155
rect 2004 25975 2060 26031
rect 2128 25975 2184 26031
rect 2252 25975 2308 26031
rect 2376 25975 2432 26031
rect 2004 25851 2060 25907
rect 2128 25851 2184 25907
rect 2252 25851 2308 25907
rect 2376 25851 2432 25907
rect 2004 25727 2060 25783
rect 2128 25727 2184 25783
rect 2252 25727 2308 25783
rect 2376 25727 2432 25783
rect 2004 25603 2060 25659
rect 2128 25603 2184 25659
rect 2252 25603 2308 25659
rect 2376 25603 2432 25659
rect 2004 25479 2060 25535
rect 2128 25479 2184 25535
rect 2252 25479 2308 25535
rect 2376 25479 2432 25535
rect 2004 25355 2060 25411
rect 2128 25355 2184 25411
rect 2252 25355 2308 25411
rect 2376 25355 2432 25411
rect 2004 25231 2060 25287
rect 2128 25231 2184 25287
rect 2252 25231 2308 25287
rect 2376 25231 2432 25287
rect 2004 25107 2060 25163
rect 2128 25107 2184 25163
rect 2252 25107 2308 25163
rect 2376 25107 2432 25163
rect 2004 24983 2060 25039
rect 2128 24983 2184 25039
rect 2252 24983 2308 25039
rect 2376 24983 2432 25039
rect 2004 24859 2060 24915
rect 2128 24859 2184 24915
rect 2252 24859 2308 24915
rect 2376 24859 2432 24915
rect 2004 24735 2060 24791
rect 2128 24735 2184 24791
rect 2252 24735 2308 24791
rect 2376 24735 2432 24791
rect 2004 24611 2060 24667
rect 2128 24611 2184 24667
rect 2252 24611 2308 24667
rect 2376 24611 2432 24667
rect 2004 24487 2060 24543
rect 2128 24487 2184 24543
rect 2252 24487 2308 24543
rect 2376 24487 2432 24543
rect 2004 24363 2060 24419
rect 2128 24363 2184 24419
rect 2252 24363 2308 24419
rect 2376 24363 2432 24419
rect 2004 24239 2060 24295
rect 2128 24239 2184 24295
rect 2252 24239 2308 24295
rect 2376 24239 2432 24295
rect 2004 24115 2060 24171
rect 2128 24115 2184 24171
rect 2252 24115 2308 24171
rect 2376 24115 2432 24171
rect 2004 23991 2060 24047
rect 2128 23991 2184 24047
rect 2252 23991 2308 24047
rect 2376 23991 2432 24047
rect 2004 23867 2060 23923
rect 2128 23867 2184 23923
rect 2252 23867 2308 23923
rect 2376 23867 2432 23923
rect 2004 23743 2060 23799
rect 2128 23743 2184 23799
rect 2252 23743 2308 23799
rect 2376 23743 2432 23799
rect 2004 23395 2060 23451
rect 2128 23395 2184 23451
rect 2252 23395 2308 23451
rect 2376 23395 2432 23451
rect 2004 23271 2060 23327
rect 2128 23271 2184 23327
rect 2252 23271 2308 23327
rect 2376 23271 2432 23327
rect 2004 23147 2060 23203
rect 2128 23147 2184 23203
rect 2252 23147 2308 23203
rect 2376 23147 2432 23203
rect 2004 23023 2060 23079
rect 2128 23023 2184 23079
rect 2252 23023 2308 23079
rect 2376 23023 2432 23079
rect 2004 22899 2060 22955
rect 2128 22899 2184 22955
rect 2252 22899 2308 22955
rect 2376 22899 2432 22955
rect 2004 22775 2060 22831
rect 2128 22775 2184 22831
rect 2252 22775 2308 22831
rect 2376 22775 2432 22831
rect 2004 22651 2060 22707
rect 2128 22651 2184 22707
rect 2252 22651 2308 22707
rect 2376 22651 2432 22707
rect 2004 22527 2060 22583
rect 2128 22527 2184 22583
rect 2252 22527 2308 22583
rect 2376 22527 2432 22583
rect 2004 22403 2060 22459
rect 2128 22403 2184 22459
rect 2252 22403 2308 22459
rect 2376 22403 2432 22459
rect 2004 22279 2060 22335
rect 2128 22279 2184 22335
rect 2252 22279 2308 22335
rect 2376 22279 2432 22335
rect 2004 22155 2060 22211
rect 2128 22155 2184 22211
rect 2252 22155 2308 22211
rect 2376 22155 2432 22211
rect 2004 22031 2060 22087
rect 2128 22031 2184 22087
rect 2252 22031 2308 22087
rect 2376 22031 2432 22087
rect 2004 21907 2060 21963
rect 2128 21907 2184 21963
rect 2252 21907 2308 21963
rect 2376 21907 2432 21963
rect 2004 21783 2060 21839
rect 2128 21783 2184 21839
rect 2252 21783 2308 21839
rect 2376 21783 2432 21839
rect 2004 21659 2060 21715
rect 2128 21659 2184 21715
rect 2252 21659 2308 21715
rect 2376 21659 2432 21715
rect 2004 21535 2060 21591
rect 2128 21535 2184 21591
rect 2252 21535 2308 21591
rect 2376 21535 2432 21591
rect 2004 21411 2060 21467
rect 2128 21411 2184 21467
rect 2252 21411 2308 21467
rect 2376 21411 2432 21467
rect 2004 21287 2060 21343
rect 2128 21287 2184 21343
rect 2252 21287 2308 21343
rect 2376 21287 2432 21343
rect 2004 21163 2060 21219
rect 2128 21163 2184 21219
rect 2252 21163 2308 21219
rect 2376 21163 2432 21219
rect 2004 21039 2060 21095
rect 2128 21039 2184 21095
rect 2252 21039 2308 21095
rect 2376 21039 2432 21095
rect 2004 20915 2060 20971
rect 2128 20915 2184 20971
rect 2252 20915 2308 20971
rect 2376 20915 2432 20971
rect 2004 20791 2060 20847
rect 2128 20791 2184 20847
rect 2252 20791 2308 20847
rect 2376 20791 2432 20847
rect 2004 20667 2060 20723
rect 2128 20667 2184 20723
rect 2252 20667 2308 20723
rect 2376 20667 2432 20723
rect 2004 20543 2060 20599
rect 2128 20543 2184 20599
rect 2252 20543 2308 20599
rect 2376 20543 2432 20599
rect 2004 20195 2060 20251
rect 2128 20195 2184 20251
rect 2252 20195 2308 20251
rect 2376 20195 2432 20251
rect 2004 20071 2060 20127
rect 2128 20071 2184 20127
rect 2252 20071 2308 20127
rect 2376 20071 2432 20127
rect 2004 19947 2060 20003
rect 2128 19947 2184 20003
rect 2252 19947 2308 20003
rect 2376 19947 2432 20003
rect 2004 19823 2060 19879
rect 2128 19823 2184 19879
rect 2252 19823 2308 19879
rect 2376 19823 2432 19879
rect 2004 19699 2060 19755
rect 2128 19699 2184 19755
rect 2252 19699 2308 19755
rect 2376 19699 2432 19755
rect 2004 19575 2060 19631
rect 2128 19575 2184 19631
rect 2252 19575 2308 19631
rect 2376 19575 2432 19631
rect 2004 19451 2060 19507
rect 2128 19451 2184 19507
rect 2252 19451 2308 19507
rect 2376 19451 2432 19507
rect 2004 19327 2060 19383
rect 2128 19327 2184 19383
rect 2252 19327 2308 19383
rect 2376 19327 2432 19383
rect 2004 19203 2060 19259
rect 2128 19203 2184 19259
rect 2252 19203 2308 19259
rect 2376 19203 2432 19259
rect 2004 19079 2060 19135
rect 2128 19079 2184 19135
rect 2252 19079 2308 19135
rect 2376 19079 2432 19135
rect 2004 18955 2060 19011
rect 2128 18955 2184 19011
rect 2252 18955 2308 19011
rect 2376 18955 2432 19011
rect 2004 18831 2060 18887
rect 2128 18831 2184 18887
rect 2252 18831 2308 18887
rect 2376 18831 2432 18887
rect 2004 18707 2060 18763
rect 2128 18707 2184 18763
rect 2252 18707 2308 18763
rect 2376 18707 2432 18763
rect 2004 18583 2060 18639
rect 2128 18583 2184 18639
rect 2252 18583 2308 18639
rect 2376 18583 2432 18639
rect 2004 18459 2060 18515
rect 2128 18459 2184 18515
rect 2252 18459 2308 18515
rect 2376 18459 2432 18515
rect 2004 18335 2060 18391
rect 2128 18335 2184 18391
rect 2252 18335 2308 18391
rect 2376 18335 2432 18391
rect 2004 18211 2060 18267
rect 2128 18211 2184 18267
rect 2252 18211 2308 18267
rect 2376 18211 2432 18267
rect 2004 18087 2060 18143
rect 2128 18087 2184 18143
rect 2252 18087 2308 18143
rect 2376 18087 2432 18143
rect 2004 17963 2060 18019
rect 2128 17963 2184 18019
rect 2252 17963 2308 18019
rect 2376 17963 2432 18019
rect 2004 17839 2060 17895
rect 2128 17839 2184 17895
rect 2252 17839 2308 17895
rect 2376 17839 2432 17895
rect 2004 17715 2060 17771
rect 2128 17715 2184 17771
rect 2252 17715 2308 17771
rect 2376 17715 2432 17771
rect 2004 17591 2060 17647
rect 2128 17591 2184 17647
rect 2252 17591 2308 17647
rect 2376 17591 2432 17647
rect 2004 17467 2060 17523
rect 2128 17467 2184 17523
rect 2252 17467 2308 17523
rect 2376 17467 2432 17523
rect 2004 17343 2060 17399
rect 2128 17343 2184 17399
rect 2252 17343 2308 17399
rect 2376 17343 2432 17399
rect 2004 16995 2060 17051
rect 2128 16995 2184 17051
rect 2252 16995 2308 17051
rect 2376 16995 2432 17051
rect 2004 16871 2060 16927
rect 2128 16871 2184 16927
rect 2252 16871 2308 16927
rect 2376 16871 2432 16927
rect 2004 16747 2060 16803
rect 2128 16747 2184 16803
rect 2252 16747 2308 16803
rect 2376 16747 2432 16803
rect 2004 16623 2060 16679
rect 2128 16623 2184 16679
rect 2252 16623 2308 16679
rect 2376 16623 2432 16679
rect 2004 16499 2060 16555
rect 2128 16499 2184 16555
rect 2252 16499 2308 16555
rect 2376 16499 2432 16555
rect 2004 16375 2060 16431
rect 2128 16375 2184 16431
rect 2252 16375 2308 16431
rect 2376 16375 2432 16431
rect 2004 16251 2060 16307
rect 2128 16251 2184 16307
rect 2252 16251 2308 16307
rect 2376 16251 2432 16307
rect 2004 16127 2060 16183
rect 2128 16127 2184 16183
rect 2252 16127 2308 16183
rect 2376 16127 2432 16183
rect 2004 16003 2060 16059
rect 2128 16003 2184 16059
rect 2252 16003 2308 16059
rect 2376 16003 2432 16059
rect 2004 15879 2060 15935
rect 2128 15879 2184 15935
rect 2252 15879 2308 15935
rect 2376 15879 2432 15935
rect 868 15631 924 15687
rect 992 15631 1048 15687
rect 1116 15631 1172 15687
rect 1240 15631 1296 15687
rect 868 15507 924 15563
rect 992 15507 1048 15563
rect 1116 15507 1172 15563
rect 1240 15507 1296 15563
rect 868 15383 924 15439
rect 992 15383 1048 15439
rect 1116 15383 1172 15439
rect 1240 15383 1296 15439
rect 868 15259 924 15315
rect 992 15259 1048 15315
rect 1116 15259 1172 15315
rect 1240 15259 1296 15315
rect 868 15135 924 15191
rect 992 15135 1048 15191
rect 1116 15135 1172 15191
rect 1240 15135 1296 15191
rect 868 15011 924 15067
rect 992 15011 1048 15067
rect 1116 15011 1172 15067
rect 1240 15011 1296 15067
rect 868 14887 924 14943
rect 992 14887 1048 14943
rect 1116 14887 1172 14943
rect 1240 14887 1296 14943
rect 868 14763 924 14819
rect 992 14763 1048 14819
rect 1116 14763 1172 14819
rect 1240 14763 1296 14819
rect 868 14639 924 14695
rect 992 14639 1048 14695
rect 1116 14639 1172 14695
rect 1240 14639 1296 14695
rect 868 14515 924 14571
rect 992 14515 1048 14571
rect 1116 14515 1172 14571
rect 1240 14515 1296 14571
rect 868 14391 924 14447
rect 992 14391 1048 14447
rect 1116 14391 1172 14447
rect 1240 14391 1296 14447
rect 868 14267 924 14323
rect 992 14267 1048 14323
rect 1116 14267 1172 14323
rect 1240 14267 1296 14323
rect 868 14143 924 14199
rect 992 14143 1048 14199
rect 1116 14143 1172 14199
rect 1240 14143 1296 14199
rect 2004 15755 2060 15811
rect 2128 15755 2184 15811
rect 2252 15755 2308 15811
rect 2376 15755 2432 15811
rect 2572 56866 2628 56922
rect 2696 56866 2752 56922
rect 2820 56866 2876 56922
rect 2944 56866 3000 56922
rect 2572 56742 2628 56798
rect 2696 56742 2752 56798
rect 2820 56742 2876 56798
rect 2944 56742 3000 56798
rect 2572 56659 2596 56674
rect 2596 56659 2628 56674
rect 2696 56659 2704 56674
rect 2704 56659 2752 56674
rect 2820 56659 2868 56674
rect 2868 56659 2876 56674
rect 2944 56659 2976 56674
rect 2976 56659 3000 56674
rect 2572 56618 2628 56659
rect 2696 56618 2752 56659
rect 2820 56618 2876 56659
rect 2944 56618 3000 56659
rect 2572 56495 2628 56550
rect 2696 56495 2752 56550
rect 2820 56495 2876 56550
rect 2944 56495 3000 56550
rect 2572 56494 2596 56495
rect 2596 56494 2628 56495
rect 2696 56494 2704 56495
rect 2704 56494 2752 56495
rect 2820 56494 2868 56495
rect 2868 56494 2876 56495
rect 2944 56494 2976 56495
rect 2976 56494 3000 56495
rect 2572 56370 2628 56426
rect 2696 56370 2752 56426
rect 2820 56370 2876 56426
rect 2944 56370 3000 56426
rect 2572 56246 2628 56302
rect 2696 56246 2752 56302
rect 2820 56246 2876 56302
rect 2944 56246 3000 56302
rect 2572 56122 2628 56178
rect 2696 56122 2752 56178
rect 2820 56122 2876 56178
rect 2944 56122 3000 56178
rect 2572 55998 2628 56054
rect 2696 55998 2752 56054
rect 2820 55998 2876 56054
rect 2944 55998 3000 56054
rect 2572 55874 2628 55930
rect 2696 55874 2752 55930
rect 2820 55874 2876 55930
rect 2944 55874 3000 55930
rect 2572 55750 2628 55806
rect 2696 55750 2752 55806
rect 2820 55750 2876 55806
rect 2944 55750 3000 55806
rect 2572 53789 2628 53845
rect 2696 53789 2752 53845
rect 2820 53789 2876 53845
rect 2944 53789 3000 53845
rect 2572 53665 2628 53721
rect 2696 53665 2752 53721
rect 2820 53665 2876 53721
rect 2944 53665 3000 53721
rect 2572 53541 2628 53597
rect 2696 53541 2752 53597
rect 2820 53541 2876 53597
rect 2944 53541 3000 53597
rect 2572 53417 2628 53473
rect 2696 53417 2752 53473
rect 2820 53417 2876 53473
rect 2944 53417 3000 53473
rect 2572 53293 2628 53349
rect 2696 53293 2752 53349
rect 2820 53293 2876 53349
rect 2944 53293 3000 53349
rect 2572 53169 2628 53225
rect 2696 53169 2752 53225
rect 2820 53169 2876 53225
rect 2944 53169 3000 53225
rect 2572 53048 2628 53101
rect 2572 53045 2574 53048
rect 2574 53045 2626 53048
rect 2626 53045 2628 53048
rect 2696 53048 2752 53101
rect 2696 53045 2698 53048
rect 2698 53045 2750 53048
rect 2750 53045 2752 53048
rect 2820 53048 2876 53101
rect 2820 53045 2822 53048
rect 2822 53045 2874 53048
rect 2874 53045 2876 53048
rect 2944 53048 3000 53101
rect 2944 53045 2946 53048
rect 2946 53045 2998 53048
rect 2998 53045 3000 53048
rect 2572 52924 2628 52977
rect 2572 52921 2574 52924
rect 2574 52921 2626 52924
rect 2626 52921 2628 52924
rect 2696 52924 2752 52977
rect 2696 52921 2698 52924
rect 2698 52921 2750 52924
rect 2750 52921 2752 52924
rect 2820 52924 2876 52977
rect 2820 52921 2822 52924
rect 2822 52921 2874 52924
rect 2874 52921 2876 52924
rect 2944 52924 3000 52977
rect 2944 52921 2946 52924
rect 2946 52921 2998 52924
rect 2998 52921 3000 52924
rect 2572 52800 2628 52853
rect 2572 52797 2574 52800
rect 2574 52797 2626 52800
rect 2626 52797 2628 52800
rect 2696 52800 2752 52853
rect 2696 52797 2698 52800
rect 2698 52797 2750 52800
rect 2750 52797 2752 52800
rect 2820 52800 2876 52853
rect 2820 52797 2822 52800
rect 2822 52797 2874 52800
rect 2874 52797 2876 52800
rect 2944 52800 3000 52853
rect 2944 52797 2946 52800
rect 2946 52797 2998 52800
rect 2998 52797 3000 52800
rect 2572 52676 2628 52729
rect 2572 52673 2574 52676
rect 2574 52673 2626 52676
rect 2626 52673 2628 52676
rect 2696 52676 2752 52729
rect 2696 52673 2698 52676
rect 2698 52673 2750 52676
rect 2750 52673 2752 52676
rect 2820 52676 2876 52729
rect 2820 52673 2822 52676
rect 2822 52673 2874 52676
rect 2874 52673 2876 52676
rect 2944 52676 3000 52729
rect 2944 52673 2946 52676
rect 2946 52673 2998 52676
rect 2998 52673 3000 52676
rect 2572 52552 2628 52605
rect 2572 52549 2574 52552
rect 2574 52549 2626 52552
rect 2626 52549 2628 52552
rect 2696 52552 2752 52605
rect 2696 52549 2698 52552
rect 2698 52549 2750 52552
rect 2750 52549 2752 52552
rect 2820 52552 2876 52605
rect 2820 52549 2822 52552
rect 2822 52549 2874 52552
rect 2874 52549 2876 52552
rect 2944 52552 3000 52605
rect 2944 52549 2946 52552
rect 2946 52549 2998 52552
rect 2998 52549 3000 52552
rect 2572 48989 2628 49045
rect 2696 48989 2752 49045
rect 2820 48989 2876 49045
rect 2944 48989 3000 49045
rect 2572 48865 2628 48921
rect 2696 48865 2752 48921
rect 2820 48865 2876 48921
rect 2944 48865 3000 48921
rect 2572 48741 2628 48797
rect 2696 48741 2752 48797
rect 2820 48741 2876 48797
rect 2944 48741 3000 48797
rect 2572 48617 2628 48673
rect 2696 48617 2752 48673
rect 2820 48617 2876 48673
rect 2944 48617 3000 48673
rect 2572 48493 2628 48549
rect 2696 48493 2752 48549
rect 2820 48493 2876 48549
rect 2944 48493 3000 48549
rect 2572 48369 2628 48425
rect 2696 48369 2752 48425
rect 2820 48369 2876 48425
rect 2944 48369 3000 48425
rect 2572 48245 2628 48301
rect 2696 48245 2752 48301
rect 2820 48245 2876 48301
rect 2944 48245 3000 48301
rect 2572 48121 2628 48177
rect 2696 48121 2752 48177
rect 2820 48121 2876 48177
rect 2944 48121 3000 48177
rect 2572 47997 2628 48053
rect 2696 47997 2752 48053
rect 2820 47997 2876 48053
rect 2944 47997 3000 48053
rect 2572 47873 2628 47929
rect 2696 47873 2752 47929
rect 2820 47873 2876 47929
rect 2944 47873 3000 47929
rect 2572 47749 2628 47805
rect 2696 47749 2752 47805
rect 2820 47749 2876 47805
rect 2944 47749 3000 47805
rect 2572 45789 2628 45845
rect 2696 45789 2752 45845
rect 2820 45789 2876 45845
rect 2944 45789 3000 45845
rect 2572 45665 2628 45721
rect 2696 45665 2752 45721
rect 2820 45665 2876 45721
rect 2944 45665 3000 45721
rect 2572 45541 2628 45597
rect 2696 45541 2752 45597
rect 2820 45541 2876 45597
rect 2944 45541 3000 45597
rect 2572 45417 2628 45473
rect 2696 45417 2752 45473
rect 2820 45417 2876 45473
rect 2944 45417 3000 45473
rect 2572 45293 2628 45349
rect 2696 45293 2752 45349
rect 2820 45293 2876 45349
rect 2944 45293 3000 45349
rect 2572 45169 2628 45225
rect 2696 45169 2752 45225
rect 2820 45169 2876 45225
rect 2944 45169 3000 45225
rect 2572 45100 2574 45101
rect 2574 45100 2626 45101
rect 2626 45100 2628 45101
rect 2572 45045 2628 45100
rect 2696 45100 2698 45101
rect 2698 45100 2750 45101
rect 2750 45100 2752 45101
rect 2696 45045 2752 45100
rect 2820 45100 2822 45101
rect 2822 45100 2874 45101
rect 2874 45100 2876 45101
rect 2820 45045 2876 45100
rect 2944 45100 2946 45101
rect 2946 45100 2998 45101
rect 2998 45100 3000 45101
rect 2944 45045 3000 45100
rect 2572 44976 2574 44977
rect 2574 44976 2626 44977
rect 2626 44976 2628 44977
rect 2572 44921 2628 44976
rect 2696 44976 2698 44977
rect 2698 44976 2750 44977
rect 2750 44976 2752 44977
rect 2696 44921 2752 44976
rect 2820 44976 2822 44977
rect 2822 44976 2874 44977
rect 2874 44976 2876 44977
rect 2820 44921 2876 44976
rect 2944 44976 2946 44977
rect 2946 44976 2998 44977
rect 2998 44976 3000 44977
rect 2944 44921 3000 44976
rect 2572 44852 2574 44853
rect 2574 44852 2626 44853
rect 2626 44852 2628 44853
rect 2572 44797 2628 44852
rect 2696 44852 2698 44853
rect 2698 44852 2750 44853
rect 2750 44852 2752 44853
rect 2696 44797 2752 44852
rect 2820 44852 2822 44853
rect 2822 44852 2874 44853
rect 2874 44852 2876 44853
rect 2820 44797 2876 44852
rect 2944 44852 2946 44853
rect 2946 44852 2998 44853
rect 2998 44852 3000 44853
rect 2944 44797 3000 44852
rect 2572 44728 2574 44729
rect 2574 44728 2626 44729
rect 2626 44728 2628 44729
rect 2572 44673 2628 44728
rect 2696 44728 2698 44729
rect 2698 44728 2750 44729
rect 2750 44728 2752 44729
rect 2696 44673 2752 44728
rect 2820 44728 2822 44729
rect 2822 44728 2874 44729
rect 2874 44728 2876 44729
rect 2820 44673 2876 44728
rect 2944 44728 2946 44729
rect 2946 44728 2998 44729
rect 2998 44728 3000 44729
rect 2944 44673 3000 44728
rect 2572 44604 2574 44605
rect 2574 44604 2626 44605
rect 2626 44604 2628 44605
rect 2572 44549 2628 44604
rect 2696 44604 2698 44605
rect 2698 44604 2750 44605
rect 2750 44604 2752 44605
rect 2696 44549 2752 44604
rect 2820 44604 2822 44605
rect 2822 44604 2874 44605
rect 2874 44604 2876 44605
rect 2820 44549 2876 44604
rect 2944 44604 2946 44605
rect 2946 44604 2998 44605
rect 2998 44604 3000 44605
rect 2944 44549 3000 44604
rect 2572 36195 2628 36251
rect 2696 36195 2752 36251
rect 2820 36195 2876 36251
rect 2944 36195 3000 36251
rect 2572 36071 2628 36127
rect 2696 36071 2752 36127
rect 2820 36071 2876 36127
rect 2944 36071 3000 36127
rect 2572 35947 2628 36003
rect 2696 35947 2752 36003
rect 2820 35947 2876 36003
rect 2944 35947 3000 36003
rect 2572 35823 2628 35879
rect 2696 35823 2752 35879
rect 2820 35823 2876 35879
rect 2944 35823 3000 35879
rect 2572 35699 2628 35755
rect 2696 35699 2752 35755
rect 2820 35699 2876 35755
rect 2944 35699 3000 35755
rect 2572 35575 2628 35631
rect 2696 35575 2752 35631
rect 2820 35575 2876 35631
rect 2944 35575 3000 35631
rect 2572 35451 2628 35507
rect 2696 35451 2752 35507
rect 2820 35451 2876 35507
rect 2944 35451 3000 35507
rect 2572 35327 2628 35383
rect 2696 35327 2752 35383
rect 2820 35327 2876 35383
rect 2944 35327 3000 35383
rect 2572 35203 2628 35259
rect 2696 35203 2752 35259
rect 2820 35203 2876 35259
rect 2944 35203 3000 35259
rect 2572 35079 2628 35135
rect 2696 35079 2752 35135
rect 2820 35079 2876 35135
rect 2944 35079 3000 35135
rect 2572 34955 2628 35011
rect 2696 34955 2752 35011
rect 2820 34955 2876 35011
rect 2944 34955 3000 35011
rect 2572 34831 2628 34887
rect 2696 34831 2752 34887
rect 2820 34831 2876 34887
rect 2944 34831 3000 34887
rect 2572 34707 2628 34763
rect 2696 34707 2752 34763
rect 2820 34707 2876 34763
rect 2944 34707 3000 34763
rect 2572 34583 2628 34639
rect 2696 34583 2752 34639
rect 2820 34583 2876 34639
rect 2944 34583 3000 34639
rect 2572 34459 2628 34515
rect 2696 34459 2752 34515
rect 2820 34459 2876 34515
rect 2944 34459 3000 34515
rect 2572 34335 2628 34391
rect 2696 34335 2752 34391
rect 2820 34335 2876 34391
rect 2944 34335 3000 34391
rect 2572 34211 2628 34267
rect 2696 34211 2752 34267
rect 2820 34211 2876 34267
rect 2944 34211 3000 34267
rect 2572 34087 2628 34143
rect 2696 34087 2752 34143
rect 2820 34087 2876 34143
rect 2944 34087 3000 34143
rect 2572 33963 2628 34019
rect 2696 33963 2752 34019
rect 2820 33963 2876 34019
rect 2944 33963 3000 34019
rect 2572 33839 2628 33895
rect 2696 33839 2752 33895
rect 2820 33839 2876 33895
rect 2944 33839 3000 33895
rect 2572 33715 2628 33771
rect 2696 33715 2752 33771
rect 2820 33715 2876 33771
rect 2944 33715 3000 33771
rect 2572 33591 2628 33647
rect 2696 33591 2752 33647
rect 2820 33591 2876 33647
rect 2944 33591 3000 33647
rect 2572 33467 2628 33523
rect 2696 33467 2752 33523
rect 2820 33467 2876 33523
rect 2944 33467 3000 33523
rect 2572 33343 2628 33399
rect 2696 33343 2752 33399
rect 2820 33343 2876 33399
rect 2944 33343 3000 33399
rect 2572 28189 2628 28245
rect 2696 28189 2752 28245
rect 2820 28189 2876 28245
rect 2944 28189 3000 28245
rect 2572 28065 2628 28121
rect 2696 28065 2752 28121
rect 2820 28065 2876 28121
rect 2944 28065 3000 28121
rect 2572 27941 2628 27997
rect 2696 27941 2752 27997
rect 2820 27941 2876 27997
rect 2944 27941 3000 27997
rect 2572 27817 2628 27873
rect 2696 27817 2752 27873
rect 2820 27817 2876 27873
rect 2944 27817 3000 27873
rect 2572 27693 2628 27749
rect 2696 27693 2752 27749
rect 2820 27693 2876 27749
rect 2944 27693 3000 27749
rect 2572 27569 2628 27625
rect 2696 27569 2752 27625
rect 2820 27569 2876 27625
rect 2944 27569 3000 27625
rect 2572 27445 2628 27501
rect 2696 27445 2752 27501
rect 2820 27445 2876 27501
rect 2944 27445 3000 27501
rect 2572 27321 2628 27377
rect 2696 27321 2752 27377
rect 2820 27321 2876 27377
rect 2944 27321 3000 27377
rect 2572 27197 2628 27253
rect 2696 27197 2752 27253
rect 2820 27197 2876 27253
rect 2944 27197 3000 27253
rect 2572 27073 2628 27129
rect 2696 27073 2752 27129
rect 2820 27073 2876 27129
rect 2944 27073 3000 27129
rect 2572 26949 2628 27005
rect 2696 26949 2752 27005
rect 2820 26949 2876 27005
rect 2944 26949 3000 27005
rect 3708 55422 3764 55445
rect 3708 55389 3729 55422
rect 3729 55389 3764 55422
rect 3832 55389 3888 55445
rect 3956 55389 4012 55445
rect 4080 55389 4136 55445
rect 3708 55314 3764 55321
rect 3708 55265 3729 55314
rect 3729 55265 3764 55314
rect 3832 55265 3888 55321
rect 3956 55265 4012 55321
rect 4080 55265 4136 55321
rect 3708 55154 3729 55197
rect 3729 55154 3764 55197
rect 3708 55141 3764 55154
rect 3832 55141 3888 55197
rect 3956 55141 4012 55197
rect 4080 55141 4136 55197
rect 3708 55046 3729 55073
rect 3729 55046 3764 55073
rect 3708 55017 3764 55046
rect 3832 55017 3888 55073
rect 3956 55017 4012 55073
rect 4080 55017 4136 55073
rect 3708 54938 3729 54949
rect 3729 54938 3764 54949
rect 3708 54893 3764 54938
rect 3832 54893 3888 54949
rect 3956 54893 4012 54949
rect 4080 54893 4136 54949
rect 3708 54774 3764 54825
rect 3708 54769 3729 54774
rect 3729 54769 3764 54774
rect 3832 54769 3888 54825
rect 3956 54769 4012 54825
rect 4080 54769 4136 54825
rect 3708 54666 3764 54701
rect 3708 54645 3729 54666
rect 3729 54645 3764 54666
rect 3832 54645 3888 54701
rect 3956 54645 4012 54701
rect 4080 54645 4136 54701
rect 3708 54558 3764 54577
rect 3708 54521 3729 54558
rect 3729 54521 3764 54558
rect 3832 54521 3888 54577
rect 3956 54521 4012 54577
rect 4080 54521 4136 54577
rect 3708 54450 3764 54453
rect 3708 54398 3729 54450
rect 3729 54398 3764 54450
rect 3708 54397 3764 54398
rect 3832 54397 3888 54453
rect 3956 54397 4012 54453
rect 4080 54397 4136 54453
rect 3708 54290 3729 54329
rect 3729 54290 3764 54329
rect 3708 54273 3764 54290
rect 3832 54273 3888 54329
rect 3956 54273 4012 54329
rect 4080 54273 4136 54329
rect 3708 54182 3729 54205
rect 3729 54182 3764 54205
rect 3708 54149 3764 54182
rect 3832 54149 3888 54205
rect 3956 54149 4012 54205
rect 4080 54149 4136 54205
rect 3708 47418 3764 47445
rect 3708 47389 3729 47418
rect 3729 47389 3764 47418
rect 3832 47389 3888 47445
rect 3956 47389 4012 47445
rect 4080 47389 4136 47445
rect 3708 47310 3764 47321
rect 3708 47265 3729 47310
rect 3729 47265 3764 47310
rect 3832 47265 3888 47321
rect 3956 47265 4012 47321
rect 4080 47265 4136 47321
rect 3708 47150 3729 47197
rect 3729 47150 3764 47197
rect 3708 47141 3764 47150
rect 3832 47141 3888 47197
rect 3956 47141 4012 47197
rect 4080 47141 4136 47197
rect 3708 47042 3729 47073
rect 3729 47042 3764 47073
rect 3708 47017 3764 47042
rect 3832 47017 3888 47073
rect 3956 47017 4012 47073
rect 4080 47017 4136 47073
rect 3708 46934 3729 46949
rect 3729 46934 3764 46949
rect 3708 46893 3764 46934
rect 3832 46893 3888 46949
rect 3956 46893 4012 46949
rect 4080 46893 4136 46949
rect 3708 46770 3764 46825
rect 3708 46769 3729 46770
rect 3729 46769 3764 46770
rect 3832 46769 3888 46825
rect 3956 46769 4012 46825
rect 4080 46769 4136 46825
rect 3708 46662 3764 46701
rect 3708 46645 3729 46662
rect 3729 46645 3764 46662
rect 3832 46645 3888 46701
rect 3956 46645 4012 46701
rect 4080 46645 4136 46701
rect 3708 46554 3764 46577
rect 3708 46521 3729 46554
rect 3729 46521 3764 46554
rect 3832 46521 3888 46577
rect 3956 46521 4012 46577
rect 4080 46521 4136 46577
rect 3708 46446 3764 46453
rect 3708 46397 3729 46446
rect 3729 46397 3764 46446
rect 3832 46397 3888 46453
rect 3956 46397 4012 46453
rect 4080 46397 4136 46453
rect 3708 46286 3729 46329
rect 3729 46286 3764 46329
rect 3708 46273 3764 46286
rect 3832 46273 3888 46329
rect 3956 46273 4012 46329
rect 4080 46273 4136 46329
rect 3708 46178 3729 46205
rect 3729 46178 3764 46205
rect 3708 46149 3764 46178
rect 3832 46149 3888 46205
rect 3956 46149 4012 46205
rect 4080 46149 4136 46205
rect 3708 44226 3764 44245
rect 3708 44189 3729 44226
rect 3729 44189 3764 44226
rect 3832 44189 3888 44245
rect 3956 44189 4012 44245
rect 4080 44189 4136 44245
rect 3708 44118 3764 44121
rect 3708 44066 3729 44118
rect 3729 44066 3764 44118
rect 3708 44065 3764 44066
rect 3832 44065 3888 44121
rect 3956 44065 4012 44121
rect 4080 44065 4136 44121
rect 3708 43958 3729 43997
rect 3729 43958 3764 43997
rect 3708 43941 3764 43958
rect 3832 43941 3888 43997
rect 3956 43941 4012 43997
rect 4080 43941 4136 43997
rect 3708 43850 3729 43873
rect 3729 43850 3764 43873
rect 3708 43817 3764 43850
rect 3832 43817 3888 43873
rect 3956 43817 4012 43873
rect 4080 43817 4136 43873
rect 3708 43742 3729 43749
rect 3729 43742 3764 43749
rect 3708 43693 3764 43742
rect 3832 43693 3888 43749
rect 3956 43693 4012 43749
rect 4080 43693 4136 43749
rect 3708 43578 3764 43625
rect 3708 43569 3729 43578
rect 3729 43569 3764 43578
rect 3832 43569 3888 43625
rect 3956 43569 4012 43625
rect 4080 43569 4136 43625
rect 3708 43470 3764 43501
rect 3708 43445 3729 43470
rect 3729 43445 3764 43470
rect 3832 43445 3888 43501
rect 3956 43445 4012 43501
rect 4080 43445 4136 43501
rect 3708 43362 3764 43377
rect 3708 43321 3729 43362
rect 3729 43321 3764 43362
rect 3832 43321 3888 43377
rect 3956 43321 4012 43377
rect 4080 43321 4136 43377
rect 3708 43202 3729 43253
rect 3729 43202 3764 43253
rect 3708 43197 3764 43202
rect 3832 43197 3888 43253
rect 3956 43197 4012 43253
rect 4080 43197 4136 43253
rect 3708 43094 3729 43129
rect 3729 43094 3764 43129
rect 3708 43073 3764 43094
rect 3832 43073 3888 43129
rect 3956 43073 4012 43129
rect 4080 43073 4136 43129
rect 3708 42986 3729 43005
rect 3729 42986 3764 43005
rect 3708 42949 3764 42986
rect 3832 42949 3888 43005
rect 3956 42949 4012 43005
rect 4080 42949 4136 43005
rect 3708 42606 3764 42645
rect 3708 42589 3729 42606
rect 3729 42589 3764 42606
rect 3832 42589 3888 42645
rect 3956 42589 4012 42645
rect 4080 42589 4136 42645
rect 3708 42498 3764 42521
rect 3708 42465 3729 42498
rect 3729 42465 3764 42498
rect 3832 42465 3888 42521
rect 3956 42465 4012 42521
rect 4080 42465 4136 42521
rect 3708 42390 3764 42397
rect 3708 42341 3729 42390
rect 3729 42341 3764 42390
rect 3832 42341 3888 42397
rect 3956 42341 4012 42397
rect 4080 42341 4136 42397
rect 3708 42230 3729 42273
rect 3729 42230 3764 42273
rect 3708 42217 3764 42230
rect 3832 42217 3888 42273
rect 3956 42217 4012 42273
rect 4080 42217 4136 42273
rect 3708 42122 3729 42149
rect 3729 42122 3764 42149
rect 3708 42093 3764 42122
rect 3832 42093 3888 42149
rect 3956 42093 4012 42149
rect 4080 42093 4136 42149
rect 3708 42014 3729 42025
rect 3729 42014 3764 42025
rect 3708 41969 3764 42014
rect 3832 41969 3888 42025
rect 3956 41969 4012 42025
rect 4080 41969 4136 42025
rect 3708 41850 3764 41901
rect 3708 41845 3729 41850
rect 3729 41845 3764 41850
rect 3832 41845 3888 41901
rect 3956 41845 4012 41901
rect 4080 41845 4136 41901
rect 3708 41742 3764 41777
rect 3708 41721 3729 41742
rect 3729 41721 3764 41742
rect 3832 41721 3888 41777
rect 3956 41721 4012 41777
rect 4080 41721 4136 41777
rect 3708 41634 3764 41653
rect 3708 41597 3729 41634
rect 3729 41597 3764 41634
rect 3832 41597 3888 41653
rect 3956 41597 4012 41653
rect 4080 41597 4136 41653
rect 3708 41526 3764 41529
rect 3708 41474 3729 41526
rect 3729 41474 3764 41526
rect 3708 41473 3764 41474
rect 3832 41473 3888 41529
rect 3956 41473 4012 41529
rect 4080 41473 4136 41529
rect 3708 41366 3729 41405
rect 3729 41366 3764 41405
rect 3708 41349 3764 41366
rect 3832 41349 3888 41405
rect 3956 41349 4012 41405
rect 4080 41349 4136 41405
rect 3708 40989 3764 41045
rect 3832 40989 3888 41045
rect 3956 40989 4012 41045
rect 4080 40989 4136 41045
rect 3708 40865 3764 40921
rect 3832 40865 3888 40921
rect 3956 40865 4012 40921
rect 4080 40865 4136 40921
rect 3708 40741 3764 40797
rect 3832 40741 3888 40797
rect 3956 40741 4012 40797
rect 4080 40741 4136 40797
rect 3708 40617 3764 40673
rect 3832 40617 3888 40673
rect 3956 40617 4012 40673
rect 4080 40617 4136 40673
rect 3708 40494 3764 40549
rect 3708 40493 3729 40494
rect 3729 40493 3764 40494
rect 3832 40493 3888 40549
rect 3956 40493 4012 40549
rect 4080 40493 4136 40549
rect 3708 40386 3764 40425
rect 3708 40369 3729 40386
rect 3729 40369 3764 40386
rect 3832 40369 3888 40425
rect 3956 40369 4012 40425
rect 4080 40369 4136 40425
rect 3708 40278 3764 40301
rect 3708 40245 3729 40278
rect 3729 40245 3764 40278
rect 3832 40245 3888 40301
rect 3956 40245 4012 40301
rect 4080 40245 4136 40301
rect 3708 40170 3764 40177
rect 3708 40121 3729 40170
rect 3729 40121 3764 40170
rect 3832 40121 3888 40177
rect 3956 40121 4012 40177
rect 4080 40121 4136 40177
rect 3708 40010 3729 40053
rect 3729 40010 3764 40053
rect 3708 39997 3764 40010
rect 3832 39997 3888 40053
rect 3956 39997 4012 40053
rect 4080 39997 4136 40053
rect 3708 39902 3729 39929
rect 3729 39902 3764 39929
rect 3708 39873 3764 39902
rect 3832 39873 3888 39929
rect 3956 39873 4012 39929
rect 4080 39873 4136 39929
rect 3708 39794 3729 39805
rect 3729 39794 3764 39805
rect 3708 39749 3764 39794
rect 3832 39749 3888 39805
rect 3956 39749 4012 39805
rect 4080 39749 4136 39805
rect 3708 32995 3764 33051
rect 3832 32995 3888 33051
rect 3956 32995 4012 33051
rect 4080 32995 4136 33051
rect 3708 32871 3764 32927
rect 3832 32871 3888 32927
rect 3956 32871 4012 32927
rect 4080 32871 4136 32927
rect 3708 32747 3764 32803
rect 3832 32747 3888 32803
rect 3956 32747 4012 32803
rect 4080 32747 4136 32803
rect 3708 32623 3764 32679
rect 3832 32623 3888 32679
rect 3956 32623 4012 32679
rect 4080 32623 4136 32679
rect 3708 32546 3729 32555
rect 3729 32546 3764 32555
rect 3708 32499 3764 32546
rect 3832 32499 3888 32555
rect 3956 32499 4012 32555
rect 4080 32499 4136 32555
rect 3708 32382 3764 32431
rect 3708 32375 3729 32382
rect 3729 32375 3764 32382
rect 3832 32375 3888 32431
rect 3956 32375 4012 32431
rect 4080 32375 4136 32431
rect 3708 32274 3764 32307
rect 3708 32251 3729 32274
rect 3729 32251 3764 32274
rect 3832 32251 3888 32307
rect 3956 32251 4012 32307
rect 4080 32251 4136 32307
rect 3708 32166 3764 32183
rect 3708 32127 3729 32166
rect 3729 32127 3764 32166
rect 3832 32127 3888 32183
rect 3956 32127 4012 32183
rect 4080 32127 4136 32183
rect 3708 32058 3764 32059
rect 3708 32006 3729 32058
rect 3729 32006 3764 32058
rect 3708 32003 3764 32006
rect 3832 32003 3888 32059
rect 3956 32003 4012 32059
rect 4080 32003 4136 32059
rect 3708 31898 3729 31935
rect 3729 31898 3764 31935
rect 3708 31879 3764 31898
rect 3832 31879 3888 31935
rect 3956 31879 4012 31935
rect 4080 31879 4136 31935
rect 3708 31790 3729 31811
rect 3729 31790 3764 31811
rect 3708 31755 3764 31790
rect 3832 31755 3888 31811
rect 3956 31755 4012 31811
rect 4080 31755 4136 31811
rect 3708 31682 3729 31687
rect 3729 31682 3764 31687
rect 3708 31631 3764 31682
rect 3832 31631 3888 31687
rect 3956 31631 4012 31687
rect 4080 31631 4136 31687
rect 3708 31518 3764 31563
rect 3708 31507 3729 31518
rect 3729 31507 3764 31518
rect 3832 31507 3888 31563
rect 3956 31507 4012 31563
rect 4080 31507 4136 31563
rect 3708 31410 3764 31439
rect 3708 31383 3729 31410
rect 3729 31383 3764 31410
rect 3832 31383 3888 31439
rect 3956 31383 4012 31439
rect 4080 31383 4136 31439
rect 3708 31302 3764 31315
rect 3708 31259 3729 31302
rect 3729 31259 3764 31302
rect 3832 31259 3888 31315
rect 3956 31259 4012 31315
rect 4080 31259 4136 31315
rect 3708 31142 3729 31191
rect 3729 31142 3764 31191
rect 3708 31135 3764 31142
rect 3832 31135 3888 31191
rect 3956 31135 4012 31191
rect 4080 31135 4136 31191
rect 3708 31034 3729 31067
rect 3729 31034 3764 31067
rect 3708 31011 3764 31034
rect 3832 31011 3888 31067
rect 3956 31011 4012 31067
rect 4080 31011 4136 31067
rect 3708 30926 3729 30943
rect 3729 30926 3764 30943
rect 3708 30887 3764 30926
rect 3832 30887 3888 30943
rect 3956 30887 4012 30943
rect 4080 30887 4136 30943
rect 3708 30818 3729 30819
rect 3729 30818 3764 30819
rect 3708 30763 3764 30818
rect 3832 30763 3888 30819
rect 3956 30763 4012 30819
rect 4080 30763 4136 30819
rect 3708 30654 3764 30695
rect 3708 30639 3729 30654
rect 3729 30639 3764 30654
rect 3832 30639 3888 30695
rect 3956 30639 4012 30695
rect 4080 30639 4136 30695
rect 3708 30546 3764 30571
rect 3708 30515 3729 30546
rect 3729 30515 3764 30546
rect 3832 30515 3888 30571
rect 3956 30515 4012 30571
rect 4080 30515 4136 30571
rect 3708 30438 3764 30447
rect 3708 30391 3729 30438
rect 3729 30391 3764 30438
rect 3832 30391 3888 30447
rect 3956 30391 4012 30447
rect 4080 30391 4136 30447
rect 3708 30278 3729 30323
rect 3729 30278 3764 30323
rect 3708 30267 3764 30278
rect 3832 30267 3888 30323
rect 3956 30267 4012 30323
rect 4080 30267 4136 30323
rect 3708 30170 3729 30199
rect 3729 30170 3764 30199
rect 3708 30143 3764 30170
rect 3832 30143 3888 30199
rect 3956 30143 4012 30199
rect 4080 30143 4136 30199
rect 3708 29790 3764 29845
rect 3708 29789 3729 29790
rect 3729 29789 3764 29790
rect 3832 29789 3888 29845
rect 3956 29789 4012 29845
rect 4080 29789 4136 29845
rect 3708 29682 3764 29721
rect 3708 29665 3729 29682
rect 3729 29665 3764 29682
rect 3832 29665 3888 29721
rect 3956 29665 4012 29721
rect 4080 29665 4136 29721
rect 3708 29574 3764 29597
rect 3708 29541 3729 29574
rect 3729 29541 3764 29574
rect 3832 29541 3888 29597
rect 3956 29541 4012 29597
rect 4080 29541 4136 29597
rect 3708 29417 3764 29473
rect 3832 29417 3888 29473
rect 3956 29417 4012 29473
rect 4080 29417 4136 29473
rect 3708 29293 3764 29349
rect 3832 29293 3888 29349
rect 3956 29293 4012 29349
rect 4080 29293 4136 29349
rect 3708 29169 3764 29225
rect 3832 29169 3888 29225
rect 3956 29169 4012 29225
rect 4080 29169 4136 29225
rect 3708 29045 3764 29101
rect 3832 29045 3888 29101
rect 3956 29045 4012 29101
rect 4080 29045 4136 29101
rect 3708 28921 3764 28977
rect 3832 28921 3888 28977
rect 3956 28921 4012 28977
rect 4080 28921 4136 28977
rect 3708 28797 3764 28853
rect 3832 28797 3888 28853
rect 3956 28797 4012 28853
rect 4080 28797 4136 28853
rect 3708 28673 3764 28729
rect 3832 28673 3888 28729
rect 3956 28673 4012 28729
rect 4080 28673 4136 28729
rect 3708 28598 3729 28605
rect 3729 28598 3764 28605
rect 3708 28549 3764 28598
rect 3832 28549 3888 28605
rect 3956 28549 4012 28605
rect 4080 28549 4136 28605
rect 3708 26598 3764 26651
rect 3708 26595 3729 26598
rect 3729 26595 3764 26598
rect 3832 26595 3888 26651
rect 3956 26595 4012 26651
rect 4080 26595 4136 26651
rect 3708 26490 3764 26527
rect 3708 26471 3729 26490
rect 3729 26471 3764 26490
rect 3832 26471 3888 26527
rect 3956 26471 4012 26527
rect 4080 26471 4136 26527
rect 3708 26382 3764 26403
rect 3708 26347 3729 26382
rect 3729 26347 3764 26382
rect 3832 26347 3888 26403
rect 3956 26347 4012 26403
rect 4080 26347 4136 26403
rect 3708 26274 3764 26279
rect 3708 26223 3729 26274
rect 3729 26223 3764 26274
rect 3832 26223 3888 26279
rect 3956 26223 4012 26279
rect 4080 26223 4136 26279
rect 3708 26114 3729 26155
rect 3729 26114 3764 26155
rect 3708 26099 3764 26114
rect 3832 26099 3888 26155
rect 3956 26099 4012 26155
rect 4080 26099 4136 26155
rect 3708 26006 3729 26031
rect 3729 26006 3764 26031
rect 3708 25975 3764 26006
rect 3832 25975 3888 26031
rect 3956 25975 4012 26031
rect 4080 25975 4136 26031
rect 3708 25898 3729 25907
rect 3729 25898 3764 25907
rect 3708 25851 3764 25898
rect 3832 25851 3888 25907
rect 3956 25851 4012 25907
rect 4080 25851 4136 25907
rect 3708 25734 3764 25783
rect 3708 25727 3729 25734
rect 3729 25727 3764 25734
rect 3832 25727 3888 25783
rect 3956 25727 4012 25783
rect 4080 25727 4136 25783
rect 3708 25626 3764 25659
rect 3708 25603 3729 25626
rect 3729 25603 3764 25626
rect 3832 25603 3888 25659
rect 3956 25603 4012 25659
rect 4080 25603 4136 25659
rect 3708 25479 3764 25535
rect 3832 25479 3888 25535
rect 3956 25479 4012 25535
rect 4080 25479 4136 25535
rect 3708 25355 3764 25411
rect 3832 25355 3888 25411
rect 3956 25355 4012 25411
rect 4080 25355 4136 25411
rect 3708 25231 3764 25287
rect 3832 25231 3888 25287
rect 3956 25231 4012 25287
rect 4080 25231 4136 25287
rect 3708 25107 3764 25163
rect 3832 25107 3888 25163
rect 3956 25107 4012 25163
rect 4080 25107 4136 25163
rect 3708 24983 3764 25039
rect 3832 24983 3888 25039
rect 3956 24983 4012 25039
rect 4080 24983 4136 25039
rect 3708 24859 3764 24915
rect 3832 24859 3888 24915
rect 3956 24859 4012 24915
rect 4080 24859 4136 24915
rect 3708 24735 3764 24791
rect 3832 24735 3888 24791
rect 3956 24735 4012 24791
rect 4080 24735 4136 24791
rect 3708 24650 3729 24667
rect 3729 24650 3764 24667
rect 3708 24611 3764 24650
rect 3832 24611 3888 24667
rect 3956 24611 4012 24667
rect 4080 24611 4136 24667
rect 3708 24542 3729 24543
rect 3729 24542 3764 24543
rect 3708 24487 3764 24542
rect 3832 24487 3888 24543
rect 3956 24487 4012 24543
rect 4080 24487 4136 24543
rect 3708 24378 3764 24419
rect 3708 24363 3729 24378
rect 3729 24363 3764 24378
rect 3832 24363 3888 24419
rect 3956 24363 4012 24419
rect 4080 24363 4136 24419
rect 3708 24270 3764 24295
rect 3708 24239 3729 24270
rect 3729 24239 3764 24270
rect 3832 24239 3888 24295
rect 3956 24239 4012 24295
rect 4080 24239 4136 24295
rect 3708 24162 3764 24171
rect 3708 24115 3729 24162
rect 3729 24115 3764 24162
rect 3832 24115 3888 24171
rect 3956 24115 4012 24171
rect 4080 24115 4136 24171
rect 3708 24002 3729 24047
rect 3729 24002 3764 24047
rect 3708 23991 3764 24002
rect 3832 23991 3888 24047
rect 3956 23991 4012 24047
rect 4080 23991 4136 24047
rect 3708 23894 3729 23923
rect 3729 23894 3764 23923
rect 3708 23867 3764 23894
rect 3832 23867 3888 23923
rect 3956 23867 4012 23923
rect 4080 23867 4136 23923
rect 3708 23786 3729 23799
rect 3729 23786 3764 23799
rect 3708 23743 3764 23786
rect 3832 23743 3888 23799
rect 3956 23743 4012 23799
rect 4080 23743 4136 23799
rect 3708 23406 3764 23451
rect 3708 23395 3729 23406
rect 3729 23395 3764 23406
rect 3832 23395 3888 23451
rect 3956 23395 4012 23451
rect 4080 23395 4136 23451
rect 3708 23298 3764 23327
rect 3708 23271 3729 23298
rect 3729 23271 3764 23298
rect 3832 23271 3888 23327
rect 3956 23271 4012 23327
rect 4080 23271 4136 23327
rect 3708 23190 3764 23203
rect 3708 23147 3729 23190
rect 3729 23147 3764 23190
rect 3832 23147 3888 23203
rect 3956 23147 4012 23203
rect 4080 23147 4136 23203
rect 3708 23030 3729 23079
rect 3729 23030 3764 23079
rect 3708 23023 3764 23030
rect 3832 23023 3888 23079
rect 3956 23023 4012 23079
rect 4080 23023 4136 23079
rect 3708 22922 3729 22955
rect 3729 22922 3764 22955
rect 3708 22899 3764 22922
rect 3832 22899 3888 22955
rect 3956 22899 4012 22955
rect 4080 22899 4136 22955
rect 3708 22814 3729 22831
rect 3729 22814 3764 22831
rect 3708 22775 3764 22814
rect 3832 22775 3888 22831
rect 3956 22775 4012 22831
rect 4080 22775 4136 22831
rect 3708 22706 3729 22707
rect 3729 22706 3764 22707
rect 3708 22651 3764 22706
rect 3832 22651 3888 22707
rect 3956 22651 4012 22707
rect 4080 22651 4136 22707
rect 3708 22542 3764 22583
rect 3708 22527 3729 22542
rect 3729 22527 3764 22542
rect 3832 22527 3888 22583
rect 3956 22527 4012 22583
rect 4080 22527 4136 22583
rect 3708 22434 3764 22459
rect 3708 22403 3729 22434
rect 3729 22403 3764 22434
rect 3832 22403 3888 22459
rect 3956 22403 4012 22459
rect 4080 22403 4136 22459
rect 3708 22326 3764 22335
rect 3708 22279 3729 22326
rect 3729 22279 3764 22326
rect 3832 22279 3888 22335
rect 3956 22279 4012 22335
rect 4080 22279 4136 22335
rect 3708 22166 3729 22211
rect 3729 22166 3764 22211
rect 3708 22155 3764 22166
rect 3832 22155 3888 22211
rect 3956 22155 4012 22211
rect 4080 22155 4136 22211
rect 3708 22058 3729 22087
rect 3729 22058 3764 22087
rect 3708 22031 3764 22058
rect 3832 22031 3888 22087
rect 3956 22031 4012 22087
rect 4080 22031 4136 22087
rect 3708 21950 3729 21963
rect 3729 21950 3764 21963
rect 3708 21907 3764 21950
rect 3832 21907 3888 21963
rect 3956 21907 4012 21963
rect 4080 21907 4136 21963
rect 3708 21786 3764 21839
rect 3708 21783 3729 21786
rect 3729 21783 3764 21786
rect 3832 21783 3888 21839
rect 3956 21783 4012 21839
rect 4080 21783 4136 21839
rect 3708 21678 3764 21715
rect 3708 21659 3729 21678
rect 3729 21659 3764 21678
rect 3832 21659 3888 21715
rect 3956 21659 4012 21715
rect 4080 21659 4136 21715
rect 3708 21535 3764 21591
rect 3832 21535 3888 21591
rect 3956 21535 4012 21591
rect 4080 21535 4136 21591
rect 3708 21411 3764 21467
rect 3832 21411 3888 21467
rect 3956 21411 4012 21467
rect 4080 21411 4136 21467
rect 3708 21287 3764 21343
rect 3832 21287 3888 21343
rect 3956 21287 4012 21343
rect 4080 21287 4136 21343
rect 3708 21163 3764 21219
rect 3832 21163 3888 21219
rect 3956 21163 4012 21219
rect 4080 21163 4136 21219
rect 3708 21039 3764 21095
rect 3832 21039 3888 21095
rect 3956 21039 4012 21095
rect 4080 21039 4136 21095
rect 3708 20915 3764 20971
rect 3832 20915 3888 20971
rect 3956 20915 4012 20971
rect 4080 20915 4136 20971
rect 3708 20791 3764 20847
rect 3832 20791 3888 20847
rect 3956 20791 4012 20847
rect 4080 20791 4136 20847
rect 3708 20667 3764 20723
rect 3832 20667 3888 20723
rect 3956 20667 4012 20723
rect 4080 20667 4136 20723
rect 3708 20577 3764 20599
rect 3832 20577 3888 20599
rect 3956 20577 4012 20599
rect 4080 20577 4136 20599
rect 3708 20543 3732 20577
rect 3732 20543 3764 20577
rect 3832 20543 3840 20577
rect 3840 20543 3888 20577
rect 3956 20543 4004 20577
rect 4004 20543 4012 20577
rect 4080 20543 4112 20577
rect 4112 20543 4136 20577
rect 3708 20195 3764 20251
rect 3832 20195 3888 20251
rect 3956 20195 4012 20251
rect 4080 20195 4136 20251
rect 3708 20071 3764 20127
rect 3832 20071 3888 20127
rect 3956 20071 4012 20127
rect 4080 20071 4136 20127
rect 3708 19947 3764 20003
rect 3832 19947 3888 20003
rect 3956 19947 4012 20003
rect 4080 19947 4136 20003
rect 3708 19823 3764 19879
rect 3832 19823 3888 19879
rect 3956 19823 4012 19879
rect 4080 19823 4136 19879
rect 3708 19699 3764 19755
rect 3832 19699 3888 19755
rect 3956 19699 4012 19755
rect 4080 19699 4136 19755
rect 3708 19584 3764 19631
rect 3832 19584 3888 19631
rect 3956 19584 4012 19631
rect 4080 19584 4136 19631
rect 3708 19575 3732 19584
rect 3732 19575 3764 19584
rect 3832 19575 3840 19584
rect 3840 19575 3888 19584
rect 3956 19575 4004 19584
rect 4004 19575 4012 19584
rect 4080 19575 4112 19584
rect 4112 19575 4136 19584
rect 3708 19476 3764 19507
rect 3832 19476 3888 19507
rect 3956 19476 4012 19507
rect 4080 19476 4136 19507
rect 3708 19451 3732 19476
rect 3732 19451 3764 19476
rect 3832 19451 3840 19476
rect 3840 19451 3888 19476
rect 3956 19451 4004 19476
rect 4004 19451 4012 19476
rect 4080 19451 4112 19476
rect 4112 19451 4136 19476
rect 3708 19327 3764 19383
rect 3832 19327 3888 19383
rect 3956 19327 4012 19383
rect 4080 19327 4136 19383
rect 3708 19203 3764 19259
rect 3832 19203 3888 19259
rect 3956 19203 4012 19259
rect 4080 19203 4136 19259
rect 3708 19079 3764 19135
rect 3832 19079 3888 19135
rect 3956 19079 4012 19135
rect 4080 19079 4136 19135
rect 3708 18955 3764 19011
rect 3832 18955 3888 19011
rect 3956 18955 4012 19011
rect 4080 18955 4136 19011
rect 3708 18831 3764 18887
rect 3832 18831 3888 18887
rect 3956 18831 4012 18887
rect 4080 18831 4136 18887
rect 3708 18712 3764 18763
rect 3832 18712 3888 18763
rect 3956 18712 4012 18763
rect 4080 18712 4136 18763
rect 3708 18707 3732 18712
rect 3732 18707 3764 18712
rect 3832 18707 3840 18712
rect 3840 18707 3888 18712
rect 3956 18707 4004 18712
rect 4004 18707 4012 18712
rect 4080 18707 4112 18712
rect 4112 18707 4136 18712
rect 3708 18604 3764 18639
rect 3832 18604 3888 18639
rect 3956 18604 4012 18639
rect 4080 18604 4136 18639
rect 3708 18583 3732 18604
rect 3732 18583 3764 18604
rect 3832 18583 3840 18604
rect 3840 18583 3888 18604
rect 3956 18583 4004 18604
rect 4004 18583 4012 18604
rect 4080 18583 4112 18604
rect 4112 18583 4136 18604
rect 3708 18459 3764 18515
rect 3832 18459 3888 18515
rect 3956 18459 4012 18515
rect 4080 18459 4136 18515
rect 3708 18335 3764 18391
rect 3832 18335 3888 18391
rect 3956 18335 4012 18391
rect 4080 18335 4136 18391
rect 3708 18211 3764 18267
rect 3832 18211 3888 18267
rect 3956 18211 4012 18267
rect 4080 18211 4136 18267
rect 3708 18087 3764 18143
rect 3832 18087 3888 18143
rect 3956 18087 4012 18143
rect 4080 18087 4136 18143
rect 3708 17963 3764 18019
rect 3832 17963 3888 18019
rect 3956 17963 4012 18019
rect 4080 17963 4136 18019
rect 3708 17840 3764 17895
rect 3832 17840 3888 17895
rect 3956 17840 4012 17895
rect 4080 17840 4136 17895
rect 3708 17839 3732 17840
rect 3732 17839 3764 17840
rect 3832 17839 3840 17840
rect 3840 17839 3888 17840
rect 3956 17839 4004 17840
rect 4004 17839 4012 17840
rect 4080 17839 4112 17840
rect 4112 17839 4136 17840
rect 3708 17732 3764 17771
rect 3832 17732 3888 17771
rect 3956 17732 4012 17771
rect 4080 17732 4136 17771
rect 3708 17715 3732 17732
rect 3732 17715 3764 17732
rect 3832 17715 3840 17732
rect 3840 17715 3888 17732
rect 3956 17715 4004 17732
rect 4004 17715 4012 17732
rect 4080 17715 4112 17732
rect 4112 17715 4136 17732
rect 3708 17591 3764 17647
rect 3832 17591 3888 17647
rect 3956 17591 4012 17647
rect 4080 17591 4136 17647
rect 3708 17467 3764 17523
rect 3832 17467 3888 17523
rect 3956 17467 4012 17523
rect 4080 17467 4136 17523
rect 3708 17343 3764 17399
rect 3832 17343 3888 17399
rect 3956 17343 4012 17399
rect 4080 17343 4136 17399
rect 3708 16995 3764 17051
rect 3832 16995 3888 17051
rect 3956 16995 4012 17051
rect 4080 16995 4136 17051
rect 3708 16916 3732 16927
rect 3732 16916 3764 16927
rect 3832 16916 3840 16927
rect 3840 16916 3888 16927
rect 3956 16916 4004 16927
rect 4004 16916 4012 16927
rect 4080 16916 4112 16927
rect 4112 16916 4136 16927
rect 3708 16871 3764 16916
rect 3832 16871 3888 16916
rect 3956 16871 4012 16916
rect 4080 16871 4136 16916
rect 3708 16747 3764 16803
rect 3832 16747 3888 16803
rect 3956 16747 4012 16803
rect 4080 16747 4136 16803
rect 3708 16623 3764 16679
rect 3832 16623 3888 16679
rect 3956 16623 4012 16679
rect 4080 16623 4136 16679
rect 3708 16499 3764 16555
rect 3832 16499 3888 16555
rect 3956 16499 4012 16555
rect 4080 16499 4136 16555
rect 3708 16375 3764 16431
rect 3832 16375 3888 16431
rect 3956 16375 4012 16431
rect 4080 16375 4136 16431
rect 3708 16251 3764 16307
rect 3832 16251 3888 16307
rect 3956 16251 4012 16307
rect 4080 16251 4136 16307
rect 3708 16127 3764 16183
rect 3832 16127 3888 16183
rect 3956 16127 4012 16183
rect 4080 16127 4136 16183
rect 3708 16031 3732 16059
rect 3732 16031 3764 16059
rect 3832 16031 3840 16059
rect 3840 16031 3888 16059
rect 3956 16031 4004 16059
rect 4004 16031 4012 16059
rect 4080 16031 4112 16059
rect 4112 16031 4136 16059
rect 3708 16003 3764 16031
rect 3832 16003 3888 16031
rect 3956 16003 4012 16031
rect 4080 16003 4136 16031
rect 3708 15923 3732 15935
rect 3732 15923 3764 15935
rect 3832 15923 3840 15935
rect 3840 15923 3888 15935
rect 3956 15923 4004 15935
rect 4004 15923 4012 15935
rect 4080 15923 4112 15935
rect 4112 15923 4136 15935
rect 3708 15879 3764 15923
rect 3832 15879 3888 15923
rect 3956 15879 4012 15923
rect 4080 15879 4136 15923
rect 2004 15631 2060 15687
rect 2128 15631 2184 15687
rect 2252 15631 2308 15687
rect 2376 15631 2432 15687
rect 2004 15507 2060 15563
rect 2128 15507 2184 15563
rect 2252 15507 2308 15563
rect 2376 15507 2432 15563
rect 2004 15383 2060 15439
rect 2128 15383 2184 15439
rect 2252 15383 2308 15439
rect 2376 15383 2432 15439
rect 2004 15259 2060 15315
rect 2128 15259 2184 15315
rect 2252 15259 2308 15315
rect 2376 15259 2432 15315
rect 2004 15135 2060 15191
rect 2128 15135 2184 15191
rect 2252 15135 2308 15191
rect 2376 15135 2432 15191
rect 2004 15011 2060 15067
rect 2128 15011 2184 15067
rect 2252 15011 2308 15067
rect 2376 15011 2432 15067
rect 2004 14887 2060 14943
rect 2128 14887 2184 14943
rect 2252 14887 2308 14943
rect 2376 14887 2432 14943
rect 2004 14763 2060 14819
rect 2128 14763 2184 14819
rect 2252 14763 2308 14819
rect 2376 14763 2432 14819
rect 2004 14639 2060 14695
rect 2128 14639 2184 14695
rect 2252 14639 2308 14695
rect 2376 14639 2432 14695
rect 2004 14515 2060 14571
rect 2128 14515 2184 14571
rect 2252 14515 2308 14571
rect 2376 14515 2432 14571
rect 2004 14391 2060 14447
rect 2128 14391 2184 14447
rect 2252 14391 2308 14447
rect 2376 14391 2432 14447
rect 2004 14267 2060 14323
rect 2128 14267 2184 14323
rect 2252 14267 2308 14323
rect 2376 14267 2432 14323
rect 2004 14143 2060 14199
rect 2128 14143 2184 14199
rect 2252 14143 2308 14199
rect 2376 14143 2432 14199
rect 3708 15755 3764 15811
rect 3832 15755 3888 15811
rect 3956 15755 4012 15811
rect 4080 15755 4136 15811
rect 4844 56866 4900 56922
rect 4968 56866 5024 56922
rect 5092 56866 5148 56922
rect 5216 56866 5272 56922
rect 4844 56742 4900 56798
rect 4968 56742 5024 56798
rect 5092 56742 5148 56798
rect 5216 56742 5272 56798
rect 4844 56659 4868 56674
rect 4868 56659 4900 56674
rect 4968 56659 4976 56674
rect 4976 56659 5024 56674
rect 5092 56659 5140 56674
rect 5140 56659 5148 56674
rect 5216 56659 5248 56674
rect 5248 56659 5272 56674
rect 4844 56618 4900 56659
rect 4968 56618 5024 56659
rect 5092 56618 5148 56659
rect 5216 56618 5272 56659
rect 4844 56495 4900 56550
rect 4968 56495 5024 56550
rect 5092 56495 5148 56550
rect 5216 56495 5272 56550
rect 4844 56494 4868 56495
rect 4868 56494 4900 56495
rect 4968 56494 4976 56495
rect 4976 56494 5024 56495
rect 5092 56494 5140 56495
rect 5140 56494 5148 56495
rect 5216 56494 5248 56495
rect 5248 56494 5272 56495
rect 4844 56370 4900 56426
rect 4968 56370 5024 56426
rect 5092 56370 5148 56426
rect 5216 56370 5272 56426
rect 4844 56246 4900 56302
rect 4968 56246 5024 56302
rect 5092 56246 5148 56302
rect 5216 56246 5272 56302
rect 4844 56122 4900 56178
rect 4968 56122 5024 56178
rect 5092 56122 5148 56178
rect 5216 56122 5272 56178
rect 4844 55998 4900 56054
rect 4968 55998 5024 56054
rect 5092 55998 5148 56054
rect 5216 55998 5272 56054
rect 4844 55874 4900 55930
rect 4968 55874 5024 55930
rect 5092 55874 5148 55930
rect 5216 55874 5272 55930
rect 4844 55750 4900 55806
rect 4968 55750 5024 55806
rect 5092 55750 5148 55806
rect 5216 55750 5272 55806
rect 4844 53789 4900 53845
rect 4968 53789 5024 53845
rect 5092 53789 5148 53845
rect 5216 53789 5272 53845
rect 4844 53665 4900 53721
rect 4968 53665 5024 53721
rect 5092 53665 5148 53721
rect 5216 53665 5272 53721
rect 4844 53541 4900 53597
rect 4968 53541 5024 53597
rect 5092 53541 5148 53597
rect 5216 53541 5272 53597
rect 4844 53417 4900 53473
rect 4968 53417 5024 53473
rect 5092 53417 5148 53473
rect 5216 53417 5272 53473
rect 4844 53293 4900 53349
rect 4968 53293 5024 53349
rect 5092 53293 5148 53349
rect 5216 53293 5272 53349
rect 4844 53169 4900 53225
rect 4968 53169 5024 53225
rect 5092 53169 5148 53225
rect 5216 53169 5272 53225
rect 4844 53048 4900 53101
rect 4844 53045 4846 53048
rect 4846 53045 4898 53048
rect 4898 53045 4900 53048
rect 4968 53048 5024 53101
rect 4968 53045 4970 53048
rect 4970 53045 5022 53048
rect 5022 53045 5024 53048
rect 5092 53048 5148 53101
rect 5092 53045 5094 53048
rect 5094 53045 5146 53048
rect 5146 53045 5148 53048
rect 5216 53048 5272 53101
rect 5216 53045 5218 53048
rect 5218 53045 5270 53048
rect 5270 53045 5272 53048
rect 4844 52924 4900 52977
rect 4844 52921 4846 52924
rect 4846 52921 4898 52924
rect 4898 52921 4900 52924
rect 4968 52924 5024 52977
rect 4968 52921 4970 52924
rect 4970 52921 5022 52924
rect 5022 52921 5024 52924
rect 5092 52924 5148 52977
rect 5092 52921 5094 52924
rect 5094 52921 5146 52924
rect 5146 52921 5148 52924
rect 5216 52924 5272 52977
rect 5216 52921 5218 52924
rect 5218 52921 5270 52924
rect 5270 52921 5272 52924
rect 4844 52800 4900 52853
rect 4844 52797 4846 52800
rect 4846 52797 4898 52800
rect 4898 52797 4900 52800
rect 4968 52800 5024 52853
rect 4968 52797 4970 52800
rect 4970 52797 5022 52800
rect 5022 52797 5024 52800
rect 5092 52800 5148 52853
rect 5092 52797 5094 52800
rect 5094 52797 5146 52800
rect 5146 52797 5148 52800
rect 5216 52800 5272 52853
rect 5216 52797 5218 52800
rect 5218 52797 5270 52800
rect 5270 52797 5272 52800
rect 4844 52676 4900 52729
rect 4844 52673 4846 52676
rect 4846 52673 4898 52676
rect 4898 52673 4900 52676
rect 4968 52676 5024 52729
rect 4968 52673 4970 52676
rect 4970 52673 5022 52676
rect 5022 52673 5024 52676
rect 5092 52676 5148 52729
rect 5092 52673 5094 52676
rect 5094 52673 5146 52676
rect 5146 52673 5148 52676
rect 5216 52676 5272 52729
rect 5216 52673 5218 52676
rect 5218 52673 5270 52676
rect 5270 52673 5272 52676
rect 4844 52552 4900 52605
rect 4844 52549 4846 52552
rect 4846 52549 4898 52552
rect 4898 52549 4900 52552
rect 4968 52552 5024 52605
rect 4968 52549 4970 52552
rect 4970 52549 5022 52552
rect 5022 52549 5024 52552
rect 5092 52552 5148 52605
rect 5092 52549 5094 52552
rect 5094 52549 5146 52552
rect 5146 52549 5148 52552
rect 5216 52552 5272 52605
rect 5216 52549 5218 52552
rect 5218 52549 5270 52552
rect 5270 52549 5272 52552
rect 4844 48989 4900 49045
rect 4968 48989 5024 49045
rect 5092 48989 5148 49045
rect 5216 48989 5272 49045
rect 4844 48865 4900 48921
rect 4968 48865 5024 48921
rect 5092 48865 5148 48921
rect 5216 48865 5272 48921
rect 4844 48741 4900 48797
rect 4968 48741 5024 48797
rect 5092 48741 5148 48797
rect 5216 48741 5272 48797
rect 4844 48617 4900 48673
rect 4968 48617 5024 48673
rect 5092 48617 5148 48673
rect 5216 48617 5272 48673
rect 4844 48493 4900 48549
rect 4968 48493 5024 48549
rect 5092 48493 5148 48549
rect 5216 48493 5272 48549
rect 4844 48369 4900 48425
rect 4968 48369 5024 48425
rect 5092 48369 5148 48425
rect 5216 48369 5272 48425
rect 4844 48245 4900 48301
rect 4968 48245 5024 48301
rect 5092 48245 5148 48301
rect 5216 48245 5272 48301
rect 4844 48121 4900 48177
rect 4968 48121 5024 48177
rect 5092 48121 5148 48177
rect 5216 48121 5272 48177
rect 4844 47997 4900 48053
rect 4968 47997 5024 48053
rect 5092 47997 5148 48053
rect 5216 47997 5272 48053
rect 4844 47873 4900 47929
rect 4968 47873 5024 47929
rect 5092 47873 5148 47929
rect 5216 47873 5272 47929
rect 4844 47749 4900 47805
rect 4968 47749 5024 47805
rect 5092 47749 5148 47805
rect 5216 47749 5272 47805
rect 4844 45789 4900 45845
rect 4968 45789 5024 45845
rect 5092 45789 5148 45845
rect 5216 45789 5272 45845
rect 4844 45665 4900 45721
rect 4968 45665 5024 45721
rect 5092 45665 5148 45721
rect 5216 45665 5272 45721
rect 4844 45541 4900 45597
rect 4968 45541 5024 45597
rect 5092 45541 5148 45597
rect 5216 45541 5272 45597
rect 4844 45417 4900 45473
rect 4968 45417 5024 45473
rect 5092 45417 5148 45473
rect 5216 45417 5272 45473
rect 4844 45293 4900 45349
rect 4968 45293 5024 45349
rect 5092 45293 5148 45349
rect 5216 45293 5272 45349
rect 4844 45169 4900 45225
rect 4968 45169 5024 45225
rect 5092 45169 5148 45225
rect 5216 45169 5272 45225
rect 4844 45100 4846 45101
rect 4846 45100 4898 45101
rect 4898 45100 4900 45101
rect 4844 45045 4900 45100
rect 4968 45100 4970 45101
rect 4970 45100 5022 45101
rect 5022 45100 5024 45101
rect 4968 45045 5024 45100
rect 5092 45100 5094 45101
rect 5094 45100 5146 45101
rect 5146 45100 5148 45101
rect 5092 45045 5148 45100
rect 5216 45100 5218 45101
rect 5218 45100 5270 45101
rect 5270 45100 5272 45101
rect 5216 45045 5272 45100
rect 4844 44976 4846 44977
rect 4846 44976 4898 44977
rect 4898 44976 4900 44977
rect 4844 44921 4900 44976
rect 4968 44976 4970 44977
rect 4970 44976 5022 44977
rect 5022 44976 5024 44977
rect 4968 44921 5024 44976
rect 5092 44976 5094 44977
rect 5094 44976 5146 44977
rect 5146 44976 5148 44977
rect 5092 44921 5148 44976
rect 5216 44976 5218 44977
rect 5218 44976 5270 44977
rect 5270 44976 5272 44977
rect 5216 44921 5272 44976
rect 4844 44852 4846 44853
rect 4846 44852 4898 44853
rect 4898 44852 4900 44853
rect 4844 44797 4900 44852
rect 4968 44852 4970 44853
rect 4970 44852 5022 44853
rect 5022 44852 5024 44853
rect 4968 44797 5024 44852
rect 5092 44852 5094 44853
rect 5094 44852 5146 44853
rect 5146 44852 5148 44853
rect 5092 44797 5148 44852
rect 5216 44852 5218 44853
rect 5218 44852 5270 44853
rect 5270 44852 5272 44853
rect 5216 44797 5272 44852
rect 4844 44728 4846 44729
rect 4846 44728 4898 44729
rect 4898 44728 4900 44729
rect 4844 44673 4900 44728
rect 4968 44728 4970 44729
rect 4970 44728 5022 44729
rect 5022 44728 5024 44729
rect 4968 44673 5024 44728
rect 5092 44728 5094 44729
rect 5094 44728 5146 44729
rect 5146 44728 5148 44729
rect 5092 44673 5148 44728
rect 5216 44728 5218 44729
rect 5218 44728 5270 44729
rect 5270 44728 5272 44729
rect 5216 44673 5272 44728
rect 4844 44604 4846 44605
rect 4846 44604 4898 44605
rect 4898 44604 4900 44605
rect 4844 44549 4900 44604
rect 4968 44604 4970 44605
rect 4970 44604 5022 44605
rect 5022 44604 5024 44605
rect 4968 44549 5024 44604
rect 5092 44604 5094 44605
rect 5094 44604 5146 44605
rect 5146 44604 5148 44605
rect 5092 44549 5148 44604
rect 5216 44604 5218 44605
rect 5218 44604 5270 44605
rect 5270 44604 5272 44605
rect 5216 44549 5272 44604
rect 4844 36195 4900 36251
rect 4968 36195 5024 36251
rect 5092 36195 5148 36251
rect 5216 36195 5272 36251
rect 4844 36071 4900 36127
rect 4968 36071 5024 36127
rect 5092 36071 5148 36127
rect 5216 36071 5272 36127
rect 4844 35947 4900 36003
rect 4968 35947 5024 36003
rect 5092 35947 5148 36003
rect 5216 35947 5272 36003
rect 4844 35823 4900 35879
rect 4968 35823 5024 35879
rect 5092 35823 5148 35879
rect 5216 35823 5272 35879
rect 4844 35699 4900 35755
rect 4968 35699 5024 35755
rect 5092 35699 5148 35755
rect 5216 35699 5272 35755
rect 4844 35575 4900 35631
rect 4968 35575 5024 35631
rect 5092 35575 5148 35631
rect 5216 35575 5272 35631
rect 4844 35451 4900 35507
rect 4968 35451 5024 35507
rect 5092 35451 5148 35507
rect 5216 35451 5272 35507
rect 4844 35327 4900 35383
rect 4968 35327 5024 35383
rect 5092 35327 5148 35383
rect 5216 35327 5272 35383
rect 4844 35203 4900 35259
rect 4968 35203 5024 35259
rect 5092 35203 5148 35259
rect 5216 35203 5272 35259
rect 4844 35079 4900 35135
rect 4968 35079 5024 35135
rect 5092 35079 5148 35135
rect 5216 35079 5272 35135
rect 4844 34955 4900 35011
rect 4968 34955 5024 35011
rect 5092 34955 5148 35011
rect 5216 34955 5272 35011
rect 4844 34831 4900 34887
rect 4968 34831 5024 34887
rect 5092 34831 5148 34887
rect 5216 34831 5272 34887
rect 4844 34707 4900 34763
rect 4968 34707 5024 34763
rect 5092 34707 5148 34763
rect 5216 34707 5272 34763
rect 4844 34583 4900 34639
rect 4968 34583 5024 34639
rect 5092 34583 5148 34639
rect 5216 34583 5272 34639
rect 4844 34459 4900 34515
rect 4968 34459 5024 34515
rect 5092 34459 5148 34515
rect 5216 34459 5272 34515
rect 4844 34335 4900 34391
rect 4968 34335 5024 34391
rect 5092 34335 5148 34391
rect 5216 34335 5272 34391
rect 4844 34211 4900 34267
rect 4968 34211 5024 34267
rect 5092 34211 5148 34267
rect 5216 34211 5272 34267
rect 4844 34087 4900 34143
rect 4968 34087 5024 34143
rect 5092 34087 5148 34143
rect 5216 34087 5272 34143
rect 4844 33963 4900 34019
rect 4968 33963 5024 34019
rect 5092 33963 5148 34019
rect 5216 33963 5272 34019
rect 4844 33839 4900 33895
rect 4968 33839 5024 33895
rect 5092 33839 5148 33895
rect 5216 33839 5272 33895
rect 4844 33715 4900 33771
rect 4968 33715 5024 33771
rect 5092 33715 5148 33771
rect 5216 33715 5272 33771
rect 4844 33591 4900 33647
rect 4968 33591 5024 33647
rect 5092 33591 5148 33647
rect 5216 33591 5272 33647
rect 4844 33467 4900 33523
rect 4968 33467 5024 33523
rect 5092 33467 5148 33523
rect 5216 33467 5272 33523
rect 4844 33343 4900 33399
rect 4968 33343 5024 33399
rect 5092 33343 5148 33399
rect 5216 33343 5272 33399
rect 4844 28189 4900 28245
rect 4968 28189 5024 28245
rect 5092 28189 5148 28245
rect 5216 28189 5272 28245
rect 4844 28065 4900 28121
rect 4968 28065 5024 28121
rect 5092 28065 5148 28121
rect 5216 28065 5272 28121
rect 4844 27941 4900 27997
rect 4968 27941 5024 27997
rect 5092 27941 5148 27997
rect 5216 27941 5272 27997
rect 4844 27817 4900 27873
rect 4968 27817 5024 27873
rect 5092 27817 5148 27873
rect 5216 27817 5272 27873
rect 4844 27693 4900 27749
rect 4968 27693 5024 27749
rect 5092 27693 5148 27749
rect 5216 27693 5272 27749
rect 4844 27569 4900 27625
rect 4968 27569 5024 27625
rect 5092 27569 5148 27625
rect 5216 27569 5272 27625
rect 4844 27445 4900 27501
rect 4968 27445 5024 27501
rect 5092 27445 5148 27501
rect 5216 27445 5272 27501
rect 4844 27321 4900 27377
rect 4968 27321 5024 27377
rect 5092 27321 5148 27377
rect 5216 27321 5272 27377
rect 4844 27197 4900 27253
rect 4968 27197 5024 27253
rect 5092 27197 5148 27253
rect 5216 27197 5272 27253
rect 4844 27073 4900 27129
rect 4968 27073 5024 27129
rect 5092 27073 5148 27129
rect 5216 27073 5272 27129
rect 4844 26949 4900 27005
rect 4968 26949 5024 27005
rect 5092 26949 5148 27005
rect 5216 26949 5272 27005
rect 5980 55389 6036 55445
rect 6104 55389 6160 55445
rect 6228 55389 6284 55445
rect 6352 55422 6408 55445
rect 6352 55389 6387 55422
rect 6387 55389 6408 55422
rect 5980 55265 6036 55321
rect 6104 55265 6160 55321
rect 6228 55265 6284 55321
rect 6352 55314 6408 55321
rect 6352 55265 6387 55314
rect 6387 55265 6408 55314
rect 5980 55141 6036 55197
rect 6104 55141 6160 55197
rect 6228 55141 6284 55197
rect 6352 55154 6387 55197
rect 6387 55154 6408 55197
rect 6352 55141 6408 55154
rect 5980 55017 6036 55073
rect 6104 55017 6160 55073
rect 6228 55017 6284 55073
rect 6352 55046 6387 55073
rect 6387 55046 6408 55073
rect 6352 55017 6408 55046
rect 5980 54893 6036 54949
rect 6104 54893 6160 54949
rect 6228 54893 6284 54949
rect 6352 54938 6387 54949
rect 6387 54938 6408 54949
rect 6352 54893 6408 54938
rect 5980 54769 6036 54825
rect 6104 54769 6160 54825
rect 6228 54769 6284 54825
rect 6352 54774 6408 54825
rect 6352 54769 6387 54774
rect 6387 54769 6408 54774
rect 5980 54645 6036 54701
rect 6104 54645 6160 54701
rect 6228 54645 6284 54701
rect 6352 54666 6408 54701
rect 6352 54645 6387 54666
rect 6387 54645 6408 54666
rect 5980 54521 6036 54577
rect 6104 54521 6160 54577
rect 6228 54521 6284 54577
rect 6352 54558 6408 54577
rect 6352 54521 6387 54558
rect 6387 54521 6408 54558
rect 5980 54397 6036 54453
rect 6104 54397 6160 54453
rect 6228 54397 6284 54453
rect 6352 54450 6408 54453
rect 6352 54398 6387 54450
rect 6387 54398 6408 54450
rect 6352 54397 6408 54398
rect 5980 54273 6036 54329
rect 6104 54273 6160 54329
rect 6228 54273 6284 54329
rect 6352 54290 6387 54329
rect 6387 54290 6408 54329
rect 6352 54273 6408 54290
rect 5980 54149 6036 54205
rect 6104 54149 6160 54205
rect 6228 54149 6284 54205
rect 6352 54182 6387 54205
rect 6387 54182 6408 54205
rect 6352 54149 6408 54182
rect 5980 47389 6036 47445
rect 6104 47389 6160 47445
rect 6228 47389 6284 47445
rect 6352 47418 6408 47445
rect 6352 47389 6387 47418
rect 6387 47389 6408 47418
rect 5980 47265 6036 47321
rect 6104 47265 6160 47321
rect 6228 47265 6284 47321
rect 6352 47310 6408 47321
rect 6352 47265 6387 47310
rect 6387 47265 6408 47310
rect 5980 47141 6036 47197
rect 6104 47141 6160 47197
rect 6228 47141 6284 47197
rect 6352 47150 6387 47197
rect 6387 47150 6408 47197
rect 6352 47141 6408 47150
rect 5980 47017 6036 47073
rect 6104 47017 6160 47073
rect 6228 47017 6284 47073
rect 6352 47042 6387 47073
rect 6387 47042 6408 47073
rect 6352 47017 6408 47042
rect 5980 46893 6036 46949
rect 6104 46893 6160 46949
rect 6228 46893 6284 46949
rect 6352 46934 6387 46949
rect 6387 46934 6408 46949
rect 6352 46893 6408 46934
rect 5980 46769 6036 46825
rect 6104 46769 6160 46825
rect 6228 46769 6284 46825
rect 6352 46770 6408 46825
rect 6352 46769 6387 46770
rect 6387 46769 6408 46770
rect 5980 46645 6036 46701
rect 6104 46645 6160 46701
rect 6228 46645 6284 46701
rect 6352 46662 6408 46701
rect 6352 46645 6387 46662
rect 6387 46645 6408 46662
rect 5980 46521 6036 46577
rect 6104 46521 6160 46577
rect 6228 46521 6284 46577
rect 6352 46554 6408 46577
rect 6352 46521 6387 46554
rect 6387 46521 6408 46554
rect 5980 46397 6036 46453
rect 6104 46397 6160 46453
rect 6228 46397 6284 46453
rect 6352 46446 6408 46453
rect 6352 46397 6387 46446
rect 6387 46397 6408 46446
rect 5980 46273 6036 46329
rect 6104 46273 6160 46329
rect 6228 46273 6284 46329
rect 6352 46286 6387 46329
rect 6387 46286 6408 46329
rect 6352 46273 6408 46286
rect 5980 46149 6036 46205
rect 6104 46149 6160 46205
rect 6228 46149 6284 46205
rect 6352 46178 6387 46205
rect 6387 46178 6408 46205
rect 6352 46149 6408 46178
rect 5980 44189 6036 44245
rect 6104 44189 6160 44245
rect 6228 44189 6284 44245
rect 6352 44226 6408 44245
rect 6352 44189 6387 44226
rect 6387 44189 6408 44226
rect 5980 44065 6036 44121
rect 6104 44065 6160 44121
rect 6228 44065 6284 44121
rect 6352 44118 6408 44121
rect 6352 44066 6387 44118
rect 6387 44066 6408 44118
rect 6352 44065 6408 44066
rect 5980 43941 6036 43997
rect 6104 43941 6160 43997
rect 6228 43941 6284 43997
rect 6352 43958 6387 43997
rect 6387 43958 6408 43997
rect 6352 43941 6408 43958
rect 5980 43817 6036 43873
rect 6104 43817 6160 43873
rect 6228 43817 6284 43873
rect 6352 43850 6387 43873
rect 6387 43850 6408 43873
rect 6352 43817 6408 43850
rect 5980 43693 6036 43749
rect 6104 43693 6160 43749
rect 6228 43693 6284 43749
rect 6352 43742 6387 43749
rect 6387 43742 6408 43749
rect 6352 43693 6408 43742
rect 5980 43569 6036 43625
rect 6104 43569 6160 43625
rect 6228 43569 6284 43625
rect 6352 43578 6408 43625
rect 6352 43569 6387 43578
rect 6387 43569 6408 43578
rect 5980 43445 6036 43501
rect 6104 43445 6160 43501
rect 6228 43445 6284 43501
rect 6352 43470 6408 43501
rect 6352 43445 6387 43470
rect 6387 43445 6408 43470
rect 5980 43321 6036 43377
rect 6104 43321 6160 43377
rect 6228 43321 6284 43377
rect 6352 43362 6408 43377
rect 6352 43321 6387 43362
rect 6387 43321 6408 43362
rect 5980 43197 6036 43253
rect 6104 43197 6160 43253
rect 6228 43197 6284 43253
rect 6352 43202 6387 43253
rect 6387 43202 6408 43253
rect 6352 43197 6408 43202
rect 5980 43073 6036 43129
rect 6104 43073 6160 43129
rect 6228 43073 6284 43129
rect 6352 43094 6387 43129
rect 6387 43094 6408 43129
rect 6352 43073 6408 43094
rect 5980 42949 6036 43005
rect 6104 42949 6160 43005
rect 6228 42949 6284 43005
rect 6352 42986 6387 43005
rect 6387 42986 6408 43005
rect 6352 42949 6408 42986
rect 5980 42589 6036 42645
rect 6104 42589 6160 42645
rect 6228 42589 6284 42645
rect 6352 42606 6408 42645
rect 6352 42589 6387 42606
rect 6387 42589 6408 42606
rect 5980 42465 6036 42521
rect 6104 42465 6160 42521
rect 6228 42465 6284 42521
rect 6352 42498 6408 42521
rect 6352 42465 6387 42498
rect 6387 42465 6408 42498
rect 5980 42341 6036 42397
rect 6104 42341 6160 42397
rect 6228 42341 6284 42397
rect 6352 42390 6408 42397
rect 6352 42341 6387 42390
rect 6387 42341 6408 42390
rect 5980 42217 6036 42273
rect 6104 42217 6160 42273
rect 6228 42217 6284 42273
rect 6352 42230 6387 42273
rect 6387 42230 6408 42273
rect 6352 42217 6408 42230
rect 5980 42093 6036 42149
rect 6104 42093 6160 42149
rect 6228 42093 6284 42149
rect 6352 42122 6387 42149
rect 6387 42122 6408 42149
rect 6352 42093 6408 42122
rect 5980 41969 6036 42025
rect 6104 41969 6160 42025
rect 6228 41969 6284 42025
rect 6352 42014 6387 42025
rect 6387 42014 6408 42025
rect 6352 41969 6408 42014
rect 5980 41845 6036 41901
rect 6104 41845 6160 41901
rect 6228 41845 6284 41901
rect 6352 41850 6408 41901
rect 6352 41845 6387 41850
rect 6387 41845 6408 41850
rect 5980 41721 6036 41777
rect 6104 41721 6160 41777
rect 6228 41721 6284 41777
rect 6352 41742 6408 41777
rect 6352 41721 6387 41742
rect 6387 41721 6408 41742
rect 5980 41597 6036 41653
rect 6104 41597 6160 41653
rect 6228 41597 6284 41653
rect 6352 41634 6408 41653
rect 6352 41597 6387 41634
rect 6387 41597 6408 41634
rect 5980 41473 6036 41529
rect 6104 41473 6160 41529
rect 6228 41473 6284 41529
rect 6352 41526 6408 41529
rect 6352 41474 6387 41526
rect 6387 41474 6408 41526
rect 6352 41473 6408 41474
rect 5980 41349 6036 41405
rect 6104 41349 6160 41405
rect 6228 41349 6284 41405
rect 6352 41366 6387 41405
rect 6387 41366 6408 41405
rect 6352 41349 6408 41366
rect 5980 40989 6036 41045
rect 6104 40989 6160 41045
rect 6228 40989 6284 41045
rect 6352 40989 6408 41045
rect 5980 40865 6036 40921
rect 6104 40865 6160 40921
rect 6228 40865 6284 40921
rect 6352 40865 6408 40921
rect 5980 40741 6036 40797
rect 6104 40741 6160 40797
rect 6228 40741 6284 40797
rect 6352 40741 6408 40797
rect 5980 40617 6036 40673
rect 6104 40617 6160 40673
rect 6228 40617 6284 40673
rect 6352 40617 6408 40673
rect 5980 40493 6036 40549
rect 6104 40493 6160 40549
rect 6228 40493 6284 40549
rect 6352 40494 6408 40549
rect 6352 40493 6387 40494
rect 6387 40493 6408 40494
rect 5980 40369 6036 40425
rect 6104 40369 6160 40425
rect 6228 40369 6284 40425
rect 6352 40386 6408 40425
rect 6352 40369 6387 40386
rect 6387 40369 6408 40386
rect 5980 40245 6036 40301
rect 6104 40245 6160 40301
rect 6228 40245 6284 40301
rect 6352 40278 6408 40301
rect 6352 40245 6387 40278
rect 6387 40245 6408 40278
rect 5980 40121 6036 40177
rect 6104 40121 6160 40177
rect 6228 40121 6284 40177
rect 6352 40170 6408 40177
rect 6352 40121 6387 40170
rect 6387 40121 6408 40170
rect 5980 39997 6036 40053
rect 6104 39997 6160 40053
rect 6228 39997 6284 40053
rect 6352 40010 6387 40053
rect 6387 40010 6408 40053
rect 6352 39997 6408 40010
rect 5980 39873 6036 39929
rect 6104 39873 6160 39929
rect 6228 39873 6284 39929
rect 6352 39902 6387 39929
rect 6387 39902 6408 39929
rect 6352 39873 6408 39902
rect 5980 39749 6036 39805
rect 6104 39749 6160 39805
rect 6228 39749 6284 39805
rect 6352 39794 6387 39805
rect 6387 39794 6408 39805
rect 6352 39749 6408 39794
rect 5980 32995 6036 33051
rect 6104 32995 6160 33051
rect 6228 32995 6284 33051
rect 6352 32995 6408 33051
rect 5980 32871 6036 32927
rect 6104 32871 6160 32927
rect 6228 32871 6284 32927
rect 6352 32871 6408 32927
rect 5980 32747 6036 32803
rect 6104 32747 6160 32803
rect 6228 32747 6284 32803
rect 6352 32747 6408 32803
rect 5980 32623 6036 32679
rect 6104 32623 6160 32679
rect 6228 32623 6284 32679
rect 6352 32623 6408 32679
rect 5980 32499 6036 32555
rect 6104 32499 6160 32555
rect 6228 32499 6284 32555
rect 6352 32546 6387 32555
rect 6387 32546 6408 32555
rect 6352 32499 6408 32546
rect 5980 32375 6036 32431
rect 6104 32375 6160 32431
rect 6228 32375 6284 32431
rect 6352 32382 6408 32431
rect 6352 32375 6387 32382
rect 6387 32375 6408 32382
rect 5980 32251 6036 32307
rect 6104 32251 6160 32307
rect 6228 32251 6284 32307
rect 6352 32274 6408 32307
rect 6352 32251 6387 32274
rect 6387 32251 6408 32274
rect 5980 32127 6036 32183
rect 6104 32127 6160 32183
rect 6228 32127 6284 32183
rect 6352 32166 6408 32183
rect 6352 32127 6387 32166
rect 6387 32127 6408 32166
rect 5980 32003 6036 32059
rect 6104 32003 6160 32059
rect 6228 32003 6284 32059
rect 6352 32058 6408 32059
rect 6352 32006 6387 32058
rect 6387 32006 6408 32058
rect 6352 32003 6408 32006
rect 5980 31879 6036 31935
rect 6104 31879 6160 31935
rect 6228 31879 6284 31935
rect 6352 31898 6387 31935
rect 6387 31898 6408 31935
rect 6352 31879 6408 31898
rect 5980 31755 6036 31811
rect 6104 31755 6160 31811
rect 6228 31755 6284 31811
rect 6352 31790 6387 31811
rect 6387 31790 6408 31811
rect 6352 31755 6408 31790
rect 5980 31631 6036 31687
rect 6104 31631 6160 31687
rect 6228 31631 6284 31687
rect 6352 31682 6387 31687
rect 6387 31682 6408 31687
rect 6352 31631 6408 31682
rect 5980 31507 6036 31563
rect 6104 31507 6160 31563
rect 6228 31507 6284 31563
rect 6352 31518 6408 31563
rect 6352 31507 6387 31518
rect 6387 31507 6408 31518
rect 5980 31383 6036 31439
rect 6104 31383 6160 31439
rect 6228 31383 6284 31439
rect 6352 31410 6408 31439
rect 6352 31383 6387 31410
rect 6387 31383 6408 31410
rect 5980 31259 6036 31315
rect 6104 31259 6160 31315
rect 6228 31259 6284 31315
rect 6352 31302 6408 31315
rect 6352 31259 6387 31302
rect 6387 31259 6408 31302
rect 5980 31135 6036 31191
rect 6104 31135 6160 31191
rect 6228 31135 6284 31191
rect 6352 31142 6387 31191
rect 6387 31142 6408 31191
rect 6352 31135 6408 31142
rect 5980 31011 6036 31067
rect 6104 31011 6160 31067
rect 6228 31011 6284 31067
rect 6352 31034 6387 31067
rect 6387 31034 6408 31067
rect 6352 31011 6408 31034
rect 5980 30887 6036 30943
rect 6104 30887 6160 30943
rect 6228 30887 6284 30943
rect 6352 30926 6387 30943
rect 6387 30926 6408 30943
rect 6352 30887 6408 30926
rect 5980 30763 6036 30819
rect 6104 30763 6160 30819
rect 6228 30763 6284 30819
rect 6352 30818 6387 30819
rect 6387 30818 6408 30819
rect 6352 30763 6408 30818
rect 5980 30639 6036 30695
rect 6104 30639 6160 30695
rect 6228 30639 6284 30695
rect 6352 30654 6408 30695
rect 6352 30639 6387 30654
rect 6387 30639 6408 30654
rect 5980 30515 6036 30571
rect 6104 30515 6160 30571
rect 6228 30515 6284 30571
rect 6352 30546 6408 30571
rect 6352 30515 6387 30546
rect 6387 30515 6408 30546
rect 5980 30391 6036 30447
rect 6104 30391 6160 30447
rect 6228 30391 6284 30447
rect 6352 30438 6408 30447
rect 6352 30391 6387 30438
rect 6387 30391 6408 30438
rect 5980 30267 6036 30323
rect 6104 30267 6160 30323
rect 6228 30267 6284 30323
rect 6352 30278 6387 30323
rect 6387 30278 6408 30323
rect 6352 30267 6408 30278
rect 5980 30143 6036 30199
rect 6104 30143 6160 30199
rect 6228 30143 6284 30199
rect 6352 30170 6387 30199
rect 6387 30170 6408 30199
rect 6352 30143 6408 30170
rect 5980 29789 6036 29845
rect 6104 29789 6160 29845
rect 6228 29789 6284 29845
rect 6352 29790 6408 29845
rect 6352 29789 6387 29790
rect 6387 29789 6408 29790
rect 5980 29665 6036 29721
rect 6104 29665 6160 29721
rect 6228 29665 6284 29721
rect 6352 29682 6408 29721
rect 6352 29665 6387 29682
rect 6387 29665 6408 29682
rect 5980 29541 6036 29597
rect 6104 29541 6160 29597
rect 6228 29541 6284 29597
rect 6352 29574 6408 29597
rect 6352 29541 6387 29574
rect 6387 29541 6408 29574
rect 5980 29417 6036 29473
rect 6104 29417 6160 29473
rect 6228 29417 6284 29473
rect 6352 29417 6408 29473
rect 5980 29293 6036 29349
rect 6104 29293 6160 29349
rect 6228 29293 6284 29349
rect 6352 29293 6408 29349
rect 5980 29169 6036 29225
rect 6104 29169 6160 29225
rect 6228 29169 6284 29225
rect 6352 29169 6408 29225
rect 5980 29045 6036 29101
rect 6104 29045 6160 29101
rect 6228 29045 6284 29101
rect 6352 29045 6408 29101
rect 5980 28921 6036 28977
rect 6104 28921 6160 28977
rect 6228 28921 6284 28977
rect 6352 28921 6408 28977
rect 5980 28797 6036 28853
rect 6104 28797 6160 28853
rect 6228 28797 6284 28853
rect 6352 28797 6408 28853
rect 5980 28673 6036 28729
rect 6104 28673 6160 28729
rect 6228 28673 6284 28729
rect 6352 28673 6408 28729
rect 5980 28549 6036 28605
rect 6104 28549 6160 28605
rect 6228 28549 6284 28605
rect 6352 28598 6387 28605
rect 6387 28598 6408 28605
rect 6352 28549 6408 28598
rect 5980 26595 6036 26651
rect 6104 26595 6160 26651
rect 6228 26595 6284 26651
rect 6352 26598 6408 26651
rect 6352 26595 6387 26598
rect 6387 26595 6408 26598
rect 5980 26471 6036 26527
rect 6104 26471 6160 26527
rect 6228 26471 6284 26527
rect 6352 26490 6408 26527
rect 6352 26471 6387 26490
rect 6387 26471 6408 26490
rect 5980 26347 6036 26403
rect 6104 26347 6160 26403
rect 6228 26347 6284 26403
rect 6352 26382 6408 26403
rect 6352 26347 6387 26382
rect 6387 26347 6408 26382
rect 5980 26223 6036 26279
rect 6104 26223 6160 26279
rect 6228 26223 6284 26279
rect 6352 26274 6408 26279
rect 6352 26223 6387 26274
rect 6387 26223 6408 26274
rect 5980 26099 6036 26155
rect 6104 26099 6160 26155
rect 6228 26099 6284 26155
rect 6352 26114 6387 26155
rect 6387 26114 6408 26155
rect 6352 26099 6408 26114
rect 5980 25975 6036 26031
rect 6104 25975 6160 26031
rect 6228 25975 6284 26031
rect 6352 26006 6387 26031
rect 6387 26006 6408 26031
rect 6352 25975 6408 26006
rect 5980 25851 6036 25907
rect 6104 25851 6160 25907
rect 6228 25851 6284 25907
rect 6352 25898 6387 25907
rect 6387 25898 6408 25907
rect 6352 25851 6408 25898
rect 5980 25727 6036 25783
rect 6104 25727 6160 25783
rect 6228 25727 6284 25783
rect 6352 25734 6408 25783
rect 6352 25727 6387 25734
rect 6387 25727 6408 25734
rect 5980 25603 6036 25659
rect 6104 25603 6160 25659
rect 6228 25603 6284 25659
rect 6352 25626 6408 25659
rect 6352 25603 6387 25626
rect 6387 25603 6408 25626
rect 5980 25479 6036 25535
rect 6104 25479 6160 25535
rect 6228 25479 6284 25535
rect 6352 25479 6408 25535
rect 5980 25355 6036 25411
rect 6104 25355 6160 25411
rect 6228 25355 6284 25411
rect 6352 25355 6408 25411
rect 5980 25231 6036 25287
rect 6104 25231 6160 25287
rect 6228 25231 6284 25287
rect 6352 25231 6408 25287
rect 5980 25107 6036 25163
rect 6104 25107 6160 25163
rect 6228 25107 6284 25163
rect 6352 25107 6408 25163
rect 5980 24983 6036 25039
rect 6104 24983 6160 25039
rect 6228 24983 6284 25039
rect 6352 24983 6408 25039
rect 5980 24859 6036 24915
rect 6104 24859 6160 24915
rect 6228 24859 6284 24915
rect 6352 24859 6408 24915
rect 5980 24735 6036 24791
rect 6104 24735 6160 24791
rect 6228 24735 6284 24791
rect 6352 24735 6408 24791
rect 5980 24611 6036 24667
rect 6104 24611 6160 24667
rect 6228 24611 6284 24667
rect 6352 24650 6387 24667
rect 6387 24650 6408 24667
rect 6352 24611 6408 24650
rect 5980 24487 6036 24543
rect 6104 24487 6160 24543
rect 6228 24487 6284 24543
rect 6352 24542 6387 24543
rect 6387 24542 6408 24543
rect 6352 24487 6408 24542
rect 5980 24363 6036 24419
rect 6104 24363 6160 24419
rect 6228 24363 6284 24419
rect 6352 24378 6408 24419
rect 6352 24363 6387 24378
rect 6387 24363 6408 24378
rect 5980 24239 6036 24295
rect 6104 24239 6160 24295
rect 6228 24239 6284 24295
rect 6352 24270 6408 24295
rect 6352 24239 6387 24270
rect 6387 24239 6408 24270
rect 5980 24115 6036 24171
rect 6104 24115 6160 24171
rect 6228 24115 6284 24171
rect 6352 24162 6408 24171
rect 6352 24115 6387 24162
rect 6387 24115 6408 24162
rect 5980 23991 6036 24047
rect 6104 23991 6160 24047
rect 6228 23991 6284 24047
rect 6352 24002 6387 24047
rect 6387 24002 6408 24047
rect 6352 23991 6408 24002
rect 5980 23867 6036 23923
rect 6104 23867 6160 23923
rect 6228 23867 6284 23923
rect 6352 23894 6387 23923
rect 6387 23894 6408 23923
rect 6352 23867 6408 23894
rect 5980 23743 6036 23799
rect 6104 23743 6160 23799
rect 6228 23743 6284 23799
rect 6352 23786 6387 23799
rect 6387 23786 6408 23799
rect 6352 23743 6408 23786
rect 5980 23395 6036 23451
rect 6104 23395 6160 23451
rect 6228 23395 6284 23451
rect 6352 23406 6408 23451
rect 6352 23395 6387 23406
rect 6387 23395 6408 23406
rect 5980 23271 6036 23327
rect 6104 23271 6160 23327
rect 6228 23271 6284 23327
rect 6352 23298 6408 23327
rect 6352 23271 6387 23298
rect 6387 23271 6408 23298
rect 5980 23147 6036 23203
rect 6104 23147 6160 23203
rect 6228 23147 6284 23203
rect 6352 23190 6408 23203
rect 6352 23147 6387 23190
rect 6387 23147 6408 23190
rect 5980 23023 6036 23079
rect 6104 23023 6160 23079
rect 6228 23023 6284 23079
rect 6352 23030 6387 23079
rect 6387 23030 6408 23079
rect 6352 23023 6408 23030
rect 5980 22899 6036 22955
rect 6104 22899 6160 22955
rect 6228 22899 6284 22955
rect 6352 22922 6387 22955
rect 6387 22922 6408 22955
rect 6352 22899 6408 22922
rect 5980 22775 6036 22831
rect 6104 22775 6160 22831
rect 6228 22775 6284 22831
rect 6352 22814 6387 22831
rect 6387 22814 6408 22831
rect 6352 22775 6408 22814
rect 5980 22651 6036 22707
rect 6104 22651 6160 22707
rect 6228 22651 6284 22707
rect 6352 22706 6387 22707
rect 6387 22706 6408 22707
rect 6352 22651 6408 22706
rect 5980 22527 6036 22583
rect 6104 22527 6160 22583
rect 6228 22527 6284 22583
rect 6352 22542 6408 22583
rect 6352 22527 6387 22542
rect 6387 22527 6408 22542
rect 5980 22403 6036 22459
rect 6104 22403 6160 22459
rect 6228 22403 6284 22459
rect 6352 22434 6408 22459
rect 6352 22403 6387 22434
rect 6387 22403 6408 22434
rect 5980 22279 6036 22335
rect 6104 22279 6160 22335
rect 6228 22279 6284 22335
rect 6352 22326 6408 22335
rect 6352 22279 6387 22326
rect 6387 22279 6408 22326
rect 5980 22155 6036 22211
rect 6104 22155 6160 22211
rect 6228 22155 6284 22211
rect 6352 22166 6387 22211
rect 6387 22166 6408 22211
rect 6352 22155 6408 22166
rect 5980 22031 6036 22087
rect 6104 22031 6160 22087
rect 6228 22031 6284 22087
rect 6352 22058 6387 22087
rect 6387 22058 6408 22087
rect 6352 22031 6408 22058
rect 5980 21907 6036 21963
rect 6104 21907 6160 21963
rect 6228 21907 6284 21963
rect 6352 21950 6387 21963
rect 6387 21950 6408 21963
rect 6352 21907 6408 21950
rect 5980 21783 6036 21839
rect 6104 21783 6160 21839
rect 6228 21783 6284 21839
rect 6352 21786 6408 21839
rect 6352 21783 6387 21786
rect 6387 21783 6408 21786
rect 5980 21659 6036 21715
rect 6104 21659 6160 21715
rect 6228 21659 6284 21715
rect 6352 21678 6408 21715
rect 6352 21659 6387 21678
rect 6387 21659 6408 21678
rect 5980 21535 6036 21591
rect 6104 21535 6160 21591
rect 6228 21535 6284 21591
rect 6352 21535 6408 21591
rect 5980 21411 6036 21467
rect 6104 21411 6160 21467
rect 6228 21411 6284 21467
rect 6352 21411 6408 21467
rect 5980 21287 6036 21343
rect 6104 21287 6160 21343
rect 6228 21287 6284 21343
rect 6352 21287 6408 21343
rect 5980 21163 6036 21219
rect 6104 21163 6160 21219
rect 6228 21163 6284 21219
rect 6352 21163 6408 21219
rect 5980 21039 6036 21095
rect 6104 21039 6160 21095
rect 6228 21039 6284 21095
rect 6352 21039 6408 21095
rect 5980 20915 6036 20971
rect 6104 20915 6160 20971
rect 6228 20915 6284 20971
rect 6352 20915 6408 20971
rect 5980 20791 6036 20847
rect 6104 20791 6160 20847
rect 6228 20791 6284 20847
rect 6352 20791 6408 20847
rect 5980 20667 6036 20723
rect 6104 20667 6160 20723
rect 6228 20667 6284 20723
rect 6352 20667 6408 20723
rect 5980 20577 6036 20599
rect 6104 20577 6160 20599
rect 6228 20577 6284 20599
rect 6352 20577 6408 20599
rect 5980 20543 6004 20577
rect 6004 20543 6036 20577
rect 6104 20543 6112 20577
rect 6112 20543 6160 20577
rect 6228 20543 6276 20577
rect 6276 20543 6284 20577
rect 6352 20543 6384 20577
rect 6384 20543 6408 20577
rect 5980 20195 6036 20251
rect 6104 20195 6160 20251
rect 6228 20195 6284 20251
rect 6352 20195 6408 20251
rect 5980 20071 6036 20127
rect 6104 20071 6160 20127
rect 6228 20071 6284 20127
rect 6352 20071 6408 20127
rect 5980 19947 6036 20003
rect 6104 19947 6160 20003
rect 6228 19947 6284 20003
rect 6352 19947 6408 20003
rect 5980 19823 6036 19879
rect 6104 19823 6160 19879
rect 6228 19823 6284 19879
rect 6352 19823 6408 19879
rect 5980 19699 6036 19755
rect 6104 19699 6160 19755
rect 6228 19699 6284 19755
rect 6352 19699 6408 19755
rect 5980 19584 6036 19631
rect 6104 19584 6160 19631
rect 6228 19584 6284 19631
rect 6352 19584 6408 19631
rect 5980 19575 6004 19584
rect 6004 19575 6036 19584
rect 6104 19575 6112 19584
rect 6112 19575 6160 19584
rect 6228 19575 6276 19584
rect 6276 19575 6284 19584
rect 6352 19575 6384 19584
rect 6384 19575 6408 19584
rect 5980 19476 6036 19507
rect 6104 19476 6160 19507
rect 6228 19476 6284 19507
rect 6352 19476 6408 19507
rect 5980 19451 6004 19476
rect 6004 19451 6036 19476
rect 6104 19451 6112 19476
rect 6112 19451 6160 19476
rect 6228 19451 6276 19476
rect 6276 19451 6284 19476
rect 6352 19451 6384 19476
rect 6384 19451 6408 19476
rect 5980 19327 6036 19383
rect 6104 19327 6160 19383
rect 6228 19327 6284 19383
rect 6352 19327 6408 19383
rect 5980 19203 6036 19259
rect 6104 19203 6160 19259
rect 6228 19203 6284 19259
rect 6352 19203 6408 19259
rect 5980 19079 6036 19135
rect 6104 19079 6160 19135
rect 6228 19079 6284 19135
rect 6352 19079 6408 19135
rect 5980 18955 6036 19011
rect 6104 18955 6160 19011
rect 6228 18955 6284 19011
rect 6352 18955 6408 19011
rect 5980 18831 6036 18887
rect 6104 18831 6160 18887
rect 6228 18831 6284 18887
rect 6352 18831 6408 18887
rect 5980 18712 6036 18763
rect 6104 18712 6160 18763
rect 6228 18712 6284 18763
rect 6352 18712 6408 18763
rect 5980 18707 6004 18712
rect 6004 18707 6036 18712
rect 6104 18707 6112 18712
rect 6112 18707 6160 18712
rect 6228 18707 6276 18712
rect 6276 18707 6284 18712
rect 6352 18707 6384 18712
rect 6384 18707 6408 18712
rect 5980 18604 6036 18639
rect 6104 18604 6160 18639
rect 6228 18604 6284 18639
rect 6352 18604 6408 18639
rect 5980 18583 6004 18604
rect 6004 18583 6036 18604
rect 6104 18583 6112 18604
rect 6112 18583 6160 18604
rect 6228 18583 6276 18604
rect 6276 18583 6284 18604
rect 6352 18583 6384 18604
rect 6384 18583 6408 18604
rect 5980 18459 6036 18515
rect 6104 18459 6160 18515
rect 6228 18459 6284 18515
rect 6352 18459 6408 18515
rect 5980 18335 6036 18391
rect 6104 18335 6160 18391
rect 6228 18335 6284 18391
rect 6352 18335 6408 18391
rect 5980 18211 6036 18267
rect 6104 18211 6160 18267
rect 6228 18211 6284 18267
rect 6352 18211 6408 18267
rect 5980 18087 6036 18143
rect 6104 18087 6160 18143
rect 6228 18087 6284 18143
rect 6352 18087 6408 18143
rect 5980 17963 6036 18019
rect 6104 17963 6160 18019
rect 6228 17963 6284 18019
rect 6352 17963 6408 18019
rect 5980 17840 6036 17895
rect 6104 17840 6160 17895
rect 6228 17840 6284 17895
rect 6352 17840 6408 17895
rect 5980 17839 6004 17840
rect 6004 17839 6036 17840
rect 6104 17839 6112 17840
rect 6112 17839 6160 17840
rect 6228 17839 6276 17840
rect 6276 17839 6284 17840
rect 6352 17839 6384 17840
rect 6384 17839 6408 17840
rect 5980 17732 6036 17771
rect 6104 17732 6160 17771
rect 6228 17732 6284 17771
rect 6352 17732 6408 17771
rect 5980 17715 6004 17732
rect 6004 17715 6036 17732
rect 6104 17715 6112 17732
rect 6112 17715 6160 17732
rect 6228 17715 6276 17732
rect 6276 17715 6284 17732
rect 6352 17715 6384 17732
rect 6384 17715 6408 17732
rect 5980 17591 6036 17647
rect 6104 17591 6160 17647
rect 6228 17591 6284 17647
rect 6352 17591 6408 17647
rect 5980 17467 6036 17523
rect 6104 17467 6160 17523
rect 6228 17467 6284 17523
rect 6352 17467 6408 17523
rect 5980 17343 6036 17399
rect 6104 17343 6160 17399
rect 6228 17343 6284 17399
rect 6352 17343 6408 17399
rect 5980 16995 6036 17051
rect 6104 16995 6160 17051
rect 6228 16995 6284 17051
rect 6352 16995 6408 17051
rect 5980 16916 6004 16927
rect 6004 16916 6036 16927
rect 6104 16916 6112 16927
rect 6112 16916 6160 16927
rect 6228 16916 6276 16927
rect 6276 16916 6284 16927
rect 6352 16916 6384 16927
rect 6384 16916 6408 16927
rect 5980 16871 6036 16916
rect 6104 16871 6160 16916
rect 6228 16871 6284 16916
rect 6352 16871 6408 16916
rect 5980 16747 6036 16803
rect 6104 16747 6160 16803
rect 6228 16747 6284 16803
rect 6352 16747 6408 16803
rect 5980 16623 6036 16679
rect 6104 16623 6160 16679
rect 6228 16623 6284 16679
rect 6352 16623 6408 16679
rect 5980 16499 6036 16555
rect 6104 16499 6160 16555
rect 6228 16499 6284 16555
rect 6352 16499 6408 16555
rect 5980 16375 6036 16431
rect 6104 16375 6160 16431
rect 6228 16375 6284 16431
rect 6352 16375 6408 16431
rect 5980 16251 6036 16307
rect 6104 16251 6160 16307
rect 6228 16251 6284 16307
rect 6352 16251 6408 16307
rect 5980 16127 6036 16183
rect 6104 16127 6160 16183
rect 6228 16127 6284 16183
rect 6352 16127 6408 16183
rect 5980 16031 6004 16059
rect 6004 16031 6036 16059
rect 6104 16031 6112 16059
rect 6112 16031 6160 16059
rect 6228 16031 6276 16059
rect 6276 16031 6284 16059
rect 6352 16031 6384 16059
rect 6384 16031 6408 16059
rect 5980 16003 6036 16031
rect 6104 16003 6160 16031
rect 6228 16003 6284 16031
rect 6352 16003 6408 16031
rect 5980 15923 6004 15935
rect 6004 15923 6036 15935
rect 6104 15923 6112 15935
rect 6112 15923 6160 15935
rect 6228 15923 6276 15935
rect 6276 15923 6284 15935
rect 6352 15923 6384 15935
rect 6384 15923 6408 15935
rect 5980 15879 6036 15923
rect 6104 15879 6160 15923
rect 6228 15879 6284 15923
rect 6352 15879 6408 15923
rect 3708 15631 3764 15687
rect 3832 15631 3888 15687
rect 3956 15631 4012 15687
rect 4080 15631 4136 15687
rect 3708 15507 3764 15563
rect 3832 15507 3888 15563
rect 3956 15507 4012 15563
rect 4080 15507 4136 15563
rect 3708 15383 3764 15439
rect 3832 15383 3888 15439
rect 3956 15383 4012 15439
rect 4080 15383 4136 15439
rect 3708 15259 3764 15315
rect 3832 15259 3888 15315
rect 3956 15259 4012 15315
rect 4080 15259 4136 15315
rect 3708 15135 3764 15191
rect 3832 15135 3888 15191
rect 3956 15135 4012 15191
rect 4080 15135 4136 15191
rect 3708 15011 3764 15067
rect 3832 15011 3888 15067
rect 3956 15011 4012 15067
rect 4080 15011 4136 15067
rect 3708 14887 3764 14943
rect 3832 14887 3888 14943
rect 3956 14887 4012 14943
rect 4080 14887 4136 14943
rect 3708 14763 3764 14819
rect 3832 14763 3888 14819
rect 3956 14763 4012 14819
rect 4080 14763 4136 14819
rect 3708 14639 3764 14695
rect 3832 14639 3888 14695
rect 3956 14639 4012 14695
rect 4080 14639 4136 14695
rect 3708 14515 3764 14571
rect 3832 14515 3888 14571
rect 3956 14515 4012 14571
rect 4080 14515 4136 14571
rect 3708 14391 3764 14447
rect 3832 14391 3888 14447
rect 3956 14391 4012 14447
rect 4080 14391 4136 14447
rect 3708 14267 3764 14323
rect 3832 14267 3888 14323
rect 3956 14267 4012 14323
rect 4080 14267 4136 14323
rect 3708 14143 3764 14199
rect 3832 14143 3888 14199
rect 3956 14143 4012 14199
rect 4080 14143 4136 14199
rect 5980 15755 6036 15811
rect 6104 15755 6160 15811
rect 6228 15755 6284 15811
rect 6352 15755 6408 15811
rect 7137 56866 7193 56922
rect 7261 56866 7317 56922
rect 7385 56866 7441 56922
rect 7137 56742 7193 56798
rect 7261 56742 7317 56798
rect 7385 56742 7441 56798
rect 7137 56659 7153 56674
rect 7153 56659 7193 56674
rect 7137 56618 7193 56659
rect 7261 56618 7317 56674
rect 7385 56659 7425 56674
rect 7425 56659 7441 56674
rect 7385 56618 7441 56659
rect 7137 56495 7193 56550
rect 7137 56494 7153 56495
rect 7153 56494 7193 56495
rect 7261 56494 7317 56550
rect 7385 56495 7441 56550
rect 7385 56494 7425 56495
rect 7425 56494 7441 56495
rect 7137 56370 7193 56426
rect 7261 56370 7317 56426
rect 7385 56370 7441 56426
rect 7137 56246 7193 56302
rect 7261 56246 7317 56302
rect 7385 56246 7441 56302
rect 7137 56122 7193 56178
rect 7261 56122 7317 56178
rect 7385 56124 7441 56178
rect 7385 56122 7388 56124
rect 7388 56122 7440 56124
rect 7440 56122 7441 56124
rect 7137 55998 7193 56054
rect 7261 55998 7317 56054
rect 7385 56016 7441 56054
rect 7385 55998 7388 56016
rect 7388 55998 7440 56016
rect 7440 55998 7441 56016
rect 7137 55874 7193 55930
rect 7261 55874 7317 55930
rect 7385 55908 7441 55930
rect 7385 55874 7388 55908
rect 7388 55874 7440 55908
rect 7440 55874 7441 55908
rect 7137 55750 7193 55806
rect 7261 55750 7317 55806
rect 7385 55800 7441 55806
rect 7385 55750 7388 55800
rect 7388 55750 7440 55800
rect 7440 55750 7441 55800
rect 7137 53789 7193 53845
rect 7261 53789 7317 53845
rect 7385 53804 7388 53845
rect 7388 53804 7440 53845
rect 7440 53804 7441 53845
rect 7385 53789 7441 53804
rect 7137 53665 7193 53721
rect 7261 53665 7317 53721
rect 7385 53696 7388 53721
rect 7388 53696 7440 53721
rect 7440 53696 7441 53721
rect 7385 53665 7441 53696
rect 7137 53541 7193 53597
rect 7261 53541 7317 53597
rect 7385 53588 7388 53597
rect 7388 53588 7440 53597
rect 7440 53588 7441 53597
rect 7385 53541 7441 53588
rect 7137 53417 7193 53473
rect 7261 53417 7317 53473
rect 7385 53424 7441 53473
rect 7385 53417 7388 53424
rect 7388 53417 7440 53424
rect 7440 53417 7441 53424
rect 7137 53293 7193 53349
rect 7261 53293 7317 53349
rect 7385 53316 7441 53349
rect 7385 53293 7388 53316
rect 7388 53293 7440 53316
rect 7440 53293 7441 53316
rect 7137 53169 7193 53225
rect 7261 53169 7317 53225
rect 7385 53169 7441 53225
rect 7137 53048 7193 53101
rect 7137 53045 7139 53048
rect 7139 53045 7191 53048
rect 7191 53045 7193 53048
rect 7261 53048 7317 53101
rect 7261 53045 7263 53048
rect 7263 53045 7315 53048
rect 7315 53045 7317 53048
rect 7385 53048 7441 53101
rect 7385 53045 7387 53048
rect 7387 53045 7439 53048
rect 7439 53045 7441 53048
rect 7137 52924 7193 52977
rect 7137 52921 7139 52924
rect 7139 52921 7191 52924
rect 7191 52921 7193 52924
rect 7261 52924 7317 52977
rect 7261 52921 7263 52924
rect 7263 52921 7315 52924
rect 7315 52921 7317 52924
rect 7385 52924 7441 52977
rect 7385 52921 7387 52924
rect 7387 52921 7439 52924
rect 7439 52921 7441 52924
rect 7137 52800 7193 52853
rect 7137 52797 7139 52800
rect 7139 52797 7191 52800
rect 7191 52797 7193 52800
rect 7261 52800 7317 52853
rect 7261 52797 7263 52800
rect 7263 52797 7315 52800
rect 7315 52797 7317 52800
rect 7385 52800 7441 52853
rect 7385 52797 7387 52800
rect 7387 52797 7439 52800
rect 7439 52797 7441 52800
rect 7137 52676 7193 52729
rect 7137 52673 7139 52676
rect 7139 52673 7191 52676
rect 7191 52673 7193 52676
rect 7261 52676 7317 52729
rect 7261 52673 7263 52676
rect 7263 52673 7315 52676
rect 7315 52673 7317 52676
rect 7385 52676 7441 52729
rect 7385 52673 7387 52676
rect 7387 52673 7439 52676
rect 7439 52673 7441 52676
rect 7137 52552 7193 52605
rect 7137 52549 7139 52552
rect 7139 52549 7191 52552
rect 7191 52549 7193 52552
rect 7261 52552 7317 52605
rect 7261 52549 7263 52552
rect 7263 52549 7315 52552
rect 7315 52549 7317 52552
rect 7385 52552 7441 52605
rect 7385 52549 7387 52552
rect 7387 52549 7439 52552
rect 7439 52549 7441 52552
rect 7137 48989 7193 49045
rect 7261 48989 7317 49045
rect 7385 48989 7441 49045
rect 7137 48865 7193 48921
rect 7261 48865 7317 48921
rect 7385 48865 7441 48921
rect 7137 48741 7193 48797
rect 7261 48741 7317 48797
rect 7385 48741 7441 48797
rect 7137 48617 7193 48673
rect 7261 48617 7317 48673
rect 7385 48617 7441 48673
rect 7137 48493 7193 48549
rect 7261 48493 7317 48549
rect 7385 48493 7441 48549
rect 7137 48369 7193 48425
rect 7261 48369 7317 48425
rect 7385 48369 7441 48425
rect 7137 48245 7193 48301
rect 7261 48245 7317 48301
rect 7385 48284 7388 48301
rect 7388 48284 7440 48301
rect 7440 48284 7441 48301
rect 7385 48245 7441 48284
rect 7137 48121 7193 48177
rect 7261 48121 7317 48177
rect 7385 48176 7388 48177
rect 7388 48176 7440 48177
rect 7440 48176 7441 48177
rect 7385 48121 7441 48176
rect 7137 47997 7193 48053
rect 7261 47997 7317 48053
rect 7385 48012 7441 48053
rect 7385 47997 7388 48012
rect 7388 47997 7440 48012
rect 7440 47997 7441 48012
rect 7137 47873 7193 47929
rect 7261 47873 7317 47929
rect 7385 47904 7441 47929
rect 7385 47873 7388 47904
rect 7388 47873 7440 47904
rect 7440 47873 7441 47904
rect 7137 47749 7193 47805
rect 7261 47749 7317 47805
rect 7385 47796 7441 47805
rect 7385 47749 7388 47796
rect 7388 47749 7440 47796
rect 7440 47749 7441 47796
rect 7137 45789 7193 45845
rect 7261 45789 7317 45845
rect 7385 45800 7388 45845
rect 7388 45800 7440 45845
rect 7440 45800 7441 45845
rect 7385 45789 7441 45800
rect 7137 45665 7193 45721
rect 7261 45665 7317 45721
rect 7385 45692 7388 45721
rect 7388 45692 7440 45721
rect 7440 45692 7441 45721
rect 7385 45665 7441 45692
rect 7137 45541 7193 45597
rect 7261 45541 7317 45597
rect 7385 45584 7388 45597
rect 7388 45584 7440 45597
rect 7440 45584 7441 45597
rect 7385 45541 7441 45584
rect 7137 45417 7193 45473
rect 7261 45417 7317 45473
rect 7385 45420 7441 45473
rect 7385 45417 7388 45420
rect 7388 45417 7440 45420
rect 7440 45417 7441 45420
rect 7137 45293 7193 45349
rect 7261 45293 7317 45349
rect 7385 45293 7441 45349
rect 7137 45169 7193 45225
rect 7261 45169 7317 45225
rect 7385 45169 7441 45225
rect 7137 45100 7139 45101
rect 7139 45100 7191 45101
rect 7191 45100 7193 45101
rect 7137 45045 7193 45100
rect 7261 45100 7263 45101
rect 7263 45100 7315 45101
rect 7315 45100 7317 45101
rect 7261 45045 7317 45100
rect 7385 45100 7387 45101
rect 7387 45100 7439 45101
rect 7439 45100 7441 45101
rect 7385 45045 7441 45100
rect 7137 44976 7139 44977
rect 7139 44976 7191 44977
rect 7191 44976 7193 44977
rect 7137 44921 7193 44976
rect 7261 44976 7263 44977
rect 7263 44976 7315 44977
rect 7315 44976 7317 44977
rect 7261 44921 7317 44976
rect 7385 44976 7387 44977
rect 7387 44976 7439 44977
rect 7439 44976 7441 44977
rect 7385 44921 7441 44976
rect 7137 44852 7139 44853
rect 7139 44852 7191 44853
rect 7191 44852 7193 44853
rect 7137 44797 7193 44852
rect 7261 44852 7263 44853
rect 7263 44852 7315 44853
rect 7315 44852 7317 44853
rect 7261 44797 7317 44852
rect 7385 44852 7387 44853
rect 7387 44852 7439 44853
rect 7439 44852 7441 44853
rect 7385 44797 7441 44852
rect 7137 44728 7139 44729
rect 7139 44728 7191 44729
rect 7191 44728 7193 44729
rect 7137 44673 7193 44728
rect 7261 44728 7263 44729
rect 7263 44728 7315 44729
rect 7315 44728 7317 44729
rect 7261 44673 7317 44728
rect 7385 44728 7387 44729
rect 7387 44728 7439 44729
rect 7439 44728 7441 44729
rect 7385 44673 7441 44728
rect 7137 44604 7139 44605
rect 7139 44604 7191 44605
rect 7191 44604 7193 44605
rect 7137 44549 7193 44604
rect 7261 44604 7263 44605
rect 7263 44604 7315 44605
rect 7315 44604 7317 44605
rect 7261 44549 7317 44604
rect 7385 44604 7387 44605
rect 7387 44604 7439 44605
rect 7439 44604 7441 44605
rect 7385 44549 7441 44604
rect 7137 36195 7193 36251
rect 7261 36195 7317 36251
rect 7385 36224 7388 36251
rect 7388 36224 7440 36251
rect 7440 36224 7441 36251
rect 7385 36195 7441 36224
rect 7137 36071 7193 36127
rect 7261 36071 7317 36127
rect 7385 36116 7388 36127
rect 7388 36116 7440 36127
rect 7440 36116 7441 36127
rect 7385 36071 7441 36116
rect 7137 35947 7193 36003
rect 7261 35947 7317 36003
rect 7385 35952 7441 36003
rect 7385 35947 7388 35952
rect 7388 35947 7440 35952
rect 7440 35947 7441 35952
rect 7137 35823 7193 35879
rect 7261 35823 7317 35879
rect 7385 35844 7441 35879
rect 7385 35823 7388 35844
rect 7388 35823 7440 35844
rect 7440 35823 7441 35844
rect 7137 35699 7193 35755
rect 7261 35699 7317 35755
rect 7385 35736 7441 35755
rect 7385 35699 7388 35736
rect 7388 35699 7440 35736
rect 7440 35699 7441 35736
rect 7137 35575 7193 35631
rect 7261 35575 7317 35631
rect 7385 35628 7441 35631
rect 7385 35576 7388 35628
rect 7388 35576 7440 35628
rect 7440 35576 7441 35628
rect 7385 35575 7441 35576
rect 7137 35451 7193 35507
rect 7261 35451 7317 35507
rect 7385 35468 7388 35507
rect 7388 35468 7440 35507
rect 7440 35468 7441 35507
rect 7385 35451 7441 35468
rect 7137 35327 7193 35383
rect 7261 35327 7317 35383
rect 7385 35360 7388 35383
rect 7388 35360 7440 35383
rect 7440 35360 7441 35383
rect 7385 35327 7441 35360
rect 7137 35203 7193 35259
rect 7261 35203 7317 35259
rect 7385 35252 7388 35259
rect 7388 35252 7440 35259
rect 7440 35252 7441 35259
rect 7385 35203 7441 35252
rect 7137 35079 7193 35135
rect 7261 35079 7317 35135
rect 7385 35088 7441 35135
rect 7385 35079 7388 35088
rect 7388 35079 7440 35088
rect 7440 35079 7441 35088
rect 7137 34955 7193 35011
rect 7261 34955 7317 35011
rect 7385 34980 7441 35011
rect 7385 34955 7388 34980
rect 7388 34955 7440 34980
rect 7440 34955 7441 34980
rect 7137 34831 7193 34887
rect 7261 34831 7317 34887
rect 7385 34872 7441 34887
rect 7385 34831 7388 34872
rect 7388 34831 7440 34872
rect 7440 34831 7441 34872
rect 7137 34707 7193 34763
rect 7261 34707 7317 34763
rect 7385 34712 7388 34763
rect 7388 34712 7440 34763
rect 7440 34712 7441 34763
rect 7385 34707 7441 34712
rect 7137 34583 7193 34639
rect 7261 34583 7317 34639
rect 7385 34604 7388 34639
rect 7388 34604 7440 34639
rect 7440 34604 7441 34639
rect 7385 34583 7441 34604
rect 7137 34459 7193 34515
rect 7261 34459 7317 34515
rect 7385 34496 7388 34515
rect 7388 34496 7440 34515
rect 7440 34496 7441 34515
rect 7385 34459 7441 34496
rect 7137 34335 7193 34391
rect 7261 34335 7317 34391
rect 7385 34388 7388 34391
rect 7388 34388 7440 34391
rect 7440 34388 7441 34391
rect 7385 34335 7441 34388
rect 7137 34211 7193 34267
rect 7261 34211 7317 34267
rect 7385 34224 7441 34267
rect 7385 34211 7388 34224
rect 7388 34211 7440 34224
rect 7440 34211 7441 34224
rect 7137 34087 7193 34143
rect 7261 34087 7317 34143
rect 7385 34116 7441 34143
rect 7385 34087 7388 34116
rect 7388 34087 7440 34116
rect 7440 34087 7441 34116
rect 7137 33963 7193 34019
rect 7261 33963 7317 34019
rect 7385 34008 7441 34019
rect 7385 33963 7388 34008
rect 7388 33963 7440 34008
rect 7440 33963 7441 34008
rect 7137 33839 7193 33895
rect 7261 33839 7317 33895
rect 7385 33848 7388 33895
rect 7388 33848 7440 33895
rect 7440 33848 7441 33895
rect 7385 33839 7441 33848
rect 7137 33715 7193 33771
rect 7261 33715 7317 33771
rect 7385 33740 7388 33771
rect 7388 33740 7440 33771
rect 7440 33740 7441 33771
rect 7385 33715 7441 33740
rect 7137 33591 7193 33647
rect 7261 33591 7317 33647
rect 7385 33632 7388 33647
rect 7388 33632 7440 33647
rect 7440 33632 7441 33647
rect 7385 33591 7441 33632
rect 7137 33467 7193 33523
rect 7261 33467 7317 33523
rect 7385 33467 7441 33523
rect 7137 33343 7193 33399
rect 7261 33343 7317 33399
rect 7385 33343 7441 33399
rect 7137 28189 7193 28245
rect 7261 28189 7317 28245
rect 7385 28220 7388 28245
rect 7388 28220 7440 28245
rect 7440 28220 7441 28245
rect 7385 28189 7441 28220
rect 7137 28065 7193 28121
rect 7261 28065 7317 28121
rect 7385 28112 7388 28121
rect 7388 28112 7440 28121
rect 7440 28112 7441 28121
rect 7385 28065 7441 28112
rect 7137 27941 7193 27997
rect 7261 27941 7317 27997
rect 7385 27948 7441 27997
rect 7385 27941 7388 27948
rect 7388 27941 7440 27948
rect 7440 27941 7441 27948
rect 7137 27817 7193 27873
rect 7261 27817 7317 27873
rect 7385 27840 7441 27873
rect 7385 27817 7388 27840
rect 7388 27817 7440 27840
rect 7440 27817 7441 27840
rect 7137 27693 7193 27749
rect 7261 27693 7317 27749
rect 7385 27732 7441 27749
rect 7385 27693 7388 27732
rect 7388 27693 7440 27732
rect 7440 27693 7441 27732
rect 7137 27569 7193 27625
rect 7261 27569 7317 27625
rect 7385 27624 7441 27625
rect 7385 27572 7388 27624
rect 7388 27572 7440 27624
rect 7440 27572 7441 27624
rect 7385 27569 7441 27572
rect 7137 27445 7193 27501
rect 7261 27445 7317 27501
rect 7385 27464 7388 27501
rect 7388 27464 7440 27501
rect 7440 27464 7441 27501
rect 7385 27445 7441 27464
rect 7137 27321 7193 27377
rect 7261 27321 7317 27377
rect 7385 27356 7388 27377
rect 7388 27356 7440 27377
rect 7440 27356 7441 27377
rect 7385 27321 7441 27356
rect 7137 27197 7193 27253
rect 7261 27197 7317 27253
rect 7385 27248 7388 27253
rect 7388 27248 7440 27253
rect 7440 27248 7441 27253
rect 7385 27197 7441 27248
rect 7137 27073 7193 27129
rect 7261 27073 7317 27129
rect 7385 27084 7441 27129
rect 7385 27073 7388 27084
rect 7388 27073 7440 27084
rect 7440 27073 7441 27084
rect 7137 26949 7193 27005
rect 7261 26949 7317 27005
rect 7385 26976 7441 27005
rect 7385 26949 7388 26976
rect 7388 26949 7440 26976
rect 7440 26949 7441 26976
rect 7623 56866 7679 56922
rect 7747 56866 7803 56922
rect 7871 56866 7927 56922
rect 7623 56742 7679 56798
rect 7747 56742 7803 56798
rect 7871 56742 7927 56798
rect 7623 56659 7639 56674
rect 7639 56659 7679 56674
rect 7623 56618 7679 56659
rect 7747 56618 7803 56674
rect 7871 56659 7911 56674
rect 7911 56659 7927 56674
rect 7871 56618 7927 56659
rect 7623 56495 7679 56550
rect 7623 56494 7639 56495
rect 7639 56494 7679 56495
rect 7747 56494 7803 56550
rect 7871 56495 7927 56550
rect 7871 56494 7911 56495
rect 7911 56494 7927 56495
rect 7623 56370 7679 56426
rect 7747 56370 7803 56426
rect 7871 56370 7927 56426
rect 7623 56246 7679 56302
rect 7747 56246 7803 56302
rect 7871 56246 7927 56302
rect 7623 56124 7679 56178
rect 7623 56122 7624 56124
rect 7624 56122 7676 56124
rect 7676 56122 7679 56124
rect 7747 56122 7803 56178
rect 7871 56122 7927 56178
rect 7623 56016 7679 56054
rect 7623 55998 7624 56016
rect 7624 55998 7676 56016
rect 7676 55998 7679 56016
rect 7747 55998 7803 56054
rect 7871 55998 7927 56054
rect 7623 55908 7679 55930
rect 7623 55874 7624 55908
rect 7624 55874 7676 55908
rect 7676 55874 7679 55908
rect 7747 55874 7803 55930
rect 7871 55874 7927 55930
rect 7623 55800 7679 55806
rect 7623 55750 7624 55800
rect 7624 55750 7676 55800
rect 7676 55750 7679 55800
rect 7747 55750 7803 55806
rect 7871 55750 7927 55806
rect 7623 53804 7624 53845
rect 7624 53804 7676 53845
rect 7676 53804 7679 53845
rect 7623 53789 7679 53804
rect 7747 53789 7803 53845
rect 7871 53789 7927 53845
rect 7623 53696 7624 53721
rect 7624 53696 7676 53721
rect 7676 53696 7679 53721
rect 7623 53665 7679 53696
rect 7747 53665 7803 53721
rect 7871 53665 7927 53721
rect 7623 53588 7624 53597
rect 7624 53588 7676 53597
rect 7676 53588 7679 53597
rect 7623 53541 7679 53588
rect 7747 53541 7803 53597
rect 7871 53541 7927 53597
rect 7623 53424 7679 53473
rect 7623 53417 7624 53424
rect 7624 53417 7676 53424
rect 7676 53417 7679 53424
rect 7747 53417 7803 53473
rect 7871 53417 7927 53473
rect 7623 53316 7679 53349
rect 7623 53293 7624 53316
rect 7624 53293 7676 53316
rect 7676 53293 7679 53316
rect 7747 53293 7803 53349
rect 7871 53293 7927 53349
rect 7623 53169 7679 53225
rect 7747 53169 7803 53225
rect 7871 53169 7927 53225
rect 7623 53048 7679 53101
rect 7623 53045 7625 53048
rect 7625 53045 7677 53048
rect 7677 53045 7679 53048
rect 7747 53048 7803 53101
rect 7747 53045 7749 53048
rect 7749 53045 7801 53048
rect 7801 53045 7803 53048
rect 7871 53048 7927 53101
rect 7871 53045 7873 53048
rect 7873 53045 7925 53048
rect 7925 53045 7927 53048
rect 7623 52924 7679 52977
rect 7623 52921 7625 52924
rect 7625 52921 7677 52924
rect 7677 52921 7679 52924
rect 7747 52924 7803 52977
rect 7747 52921 7749 52924
rect 7749 52921 7801 52924
rect 7801 52921 7803 52924
rect 7871 52924 7927 52977
rect 7871 52921 7873 52924
rect 7873 52921 7925 52924
rect 7925 52921 7927 52924
rect 7623 52800 7679 52853
rect 7623 52797 7625 52800
rect 7625 52797 7677 52800
rect 7677 52797 7679 52800
rect 7747 52800 7803 52853
rect 7747 52797 7749 52800
rect 7749 52797 7801 52800
rect 7801 52797 7803 52800
rect 7871 52800 7927 52853
rect 7871 52797 7873 52800
rect 7873 52797 7925 52800
rect 7925 52797 7927 52800
rect 7623 52676 7679 52729
rect 7623 52673 7625 52676
rect 7625 52673 7677 52676
rect 7677 52673 7679 52676
rect 7747 52676 7803 52729
rect 7747 52673 7749 52676
rect 7749 52673 7801 52676
rect 7801 52673 7803 52676
rect 7871 52676 7927 52729
rect 7871 52673 7873 52676
rect 7873 52673 7925 52676
rect 7925 52673 7927 52676
rect 7623 52552 7679 52605
rect 7623 52549 7625 52552
rect 7625 52549 7677 52552
rect 7677 52549 7679 52552
rect 7747 52552 7803 52605
rect 7747 52549 7749 52552
rect 7749 52549 7801 52552
rect 7801 52549 7803 52552
rect 7871 52552 7927 52605
rect 7871 52549 7873 52552
rect 7873 52549 7925 52552
rect 7925 52549 7927 52552
rect 7623 48989 7679 49045
rect 7747 48989 7803 49045
rect 7871 48989 7927 49045
rect 7623 48865 7679 48921
rect 7747 48865 7803 48921
rect 7871 48865 7927 48921
rect 7623 48741 7679 48797
rect 7747 48741 7803 48797
rect 7871 48741 7927 48797
rect 7623 48617 7679 48673
rect 7747 48617 7803 48673
rect 7871 48617 7927 48673
rect 7623 48493 7679 48549
rect 7747 48493 7803 48549
rect 7871 48493 7927 48549
rect 7623 48369 7679 48425
rect 7747 48369 7803 48425
rect 7871 48369 7927 48425
rect 7623 48284 7624 48301
rect 7624 48284 7676 48301
rect 7676 48284 7679 48301
rect 7623 48245 7679 48284
rect 7747 48245 7803 48301
rect 7871 48245 7927 48301
rect 7623 48176 7624 48177
rect 7624 48176 7676 48177
rect 7676 48176 7679 48177
rect 7623 48121 7679 48176
rect 7747 48121 7803 48177
rect 7871 48121 7927 48177
rect 7623 48012 7679 48053
rect 7623 47997 7624 48012
rect 7624 47997 7676 48012
rect 7676 47997 7679 48012
rect 7747 47997 7803 48053
rect 7871 47997 7927 48053
rect 7623 47904 7679 47929
rect 7623 47873 7624 47904
rect 7624 47873 7676 47904
rect 7676 47873 7679 47904
rect 7747 47873 7803 47929
rect 7871 47873 7927 47929
rect 7623 47796 7679 47805
rect 7623 47749 7624 47796
rect 7624 47749 7676 47796
rect 7676 47749 7679 47796
rect 7747 47749 7803 47805
rect 7871 47749 7927 47805
rect 7623 45800 7624 45845
rect 7624 45800 7676 45845
rect 7676 45800 7679 45845
rect 7623 45789 7679 45800
rect 7747 45789 7803 45845
rect 7871 45789 7927 45845
rect 7623 45692 7624 45721
rect 7624 45692 7676 45721
rect 7676 45692 7679 45721
rect 7623 45665 7679 45692
rect 7747 45665 7803 45721
rect 7871 45665 7927 45721
rect 7623 45584 7624 45597
rect 7624 45584 7676 45597
rect 7676 45584 7679 45597
rect 7623 45541 7679 45584
rect 7747 45541 7803 45597
rect 7871 45541 7927 45597
rect 7623 45420 7679 45473
rect 7623 45417 7624 45420
rect 7624 45417 7676 45420
rect 7676 45417 7679 45420
rect 7747 45417 7803 45473
rect 7871 45417 7927 45473
rect 7623 45293 7679 45349
rect 7747 45293 7803 45349
rect 7871 45293 7927 45349
rect 7623 45169 7679 45225
rect 7747 45169 7803 45225
rect 7871 45169 7927 45225
rect 7623 45100 7625 45101
rect 7625 45100 7677 45101
rect 7677 45100 7679 45101
rect 7623 45045 7679 45100
rect 7747 45100 7749 45101
rect 7749 45100 7801 45101
rect 7801 45100 7803 45101
rect 7747 45045 7803 45100
rect 7871 45100 7873 45101
rect 7873 45100 7925 45101
rect 7925 45100 7927 45101
rect 7871 45045 7927 45100
rect 7623 44976 7625 44977
rect 7625 44976 7677 44977
rect 7677 44976 7679 44977
rect 7623 44921 7679 44976
rect 7747 44976 7749 44977
rect 7749 44976 7801 44977
rect 7801 44976 7803 44977
rect 7747 44921 7803 44976
rect 7871 44976 7873 44977
rect 7873 44976 7925 44977
rect 7925 44976 7927 44977
rect 7871 44921 7927 44976
rect 7623 44852 7625 44853
rect 7625 44852 7677 44853
rect 7677 44852 7679 44853
rect 7623 44797 7679 44852
rect 7747 44852 7749 44853
rect 7749 44852 7801 44853
rect 7801 44852 7803 44853
rect 7747 44797 7803 44852
rect 7871 44852 7873 44853
rect 7873 44852 7925 44853
rect 7925 44852 7927 44853
rect 7871 44797 7927 44852
rect 7623 44728 7625 44729
rect 7625 44728 7677 44729
rect 7677 44728 7679 44729
rect 7623 44673 7679 44728
rect 7747 44728 7749 44729
rect 7749 44728 7801 44729
rect 7801 44728 7803 44729
rect 7747 44673 7803 44728
rect 7871 44728 7873 44729
rect 7873 44728 7925 44729
rect 7925 44728 7927 44729
rect 7871 44673 7927 44728
rect 7623 44604 7625 44605
rect 7625 44604 7677 44605
rect 7677 44604 7679 44605
rect 7623 44549 7679 44604
rect 7747 44604 7749 44605
rect 7749 44604 7801 44605
rect 7801 44604 7803 44605
rect 7747 44549 7803 44604
rect 7871 44604 7873 44605
rect 7873 44604 7925 44605
rect 7925 44604 7927 44605
rect 7871 44549 7927 44604
rect 7623 36224 7624 36251
rect 7624 36224 7676 36251
rect 7676 36224 7679 36251
rect 7623 36195 7679 36224
rect 7747 36195 7803 36251
rect 7871 36195 7927 36251
rect 7623 36116 7624 36127
rect 7624 36116 7676 36127
rect 7676 36116 7679 36127
rect 7623 36071 7679 36116
rect 7747 36071 7803 36127
rect 7871 36071 7927 36127
rect 7623 35952 7679 36003
rect 7623 35947 7624 35952
rect 7624 35947 7676 35952
rect 7676 35947 7679 35952
rect 7747 35947 7803 36003
rect 7871 35947 7927 36003
rect 7623 35844 7679 35879
rect 7623 35823 7624 35844
rect 7624 35823 7676 35844
rect 7676 35823 7679 35844
rect 7747 35823 7803 35879
rect 7871 35823 7927 35879
rect 7623 35736 7679 35755
rect 7623 35699 7624 35736
rect 7624 35699 7676 35736
rect 7676 35699 7679 35736
rect 7747 35699 7803 35755
rect 7871 35699 7927 35755
rect 7623 35628 7679 35631
rect 7623 35576 7624 35628
rect 7624 35576 7676 35628
rect 7676 35576 7679 35628
rect 7623 35575 7679 35576
rect 7747 35575 7803 35631
rect 7871 35575 7927 35631
rect 7623 35468 7624 35507
rect 7624 35468 7676 35507
rect 7676 35468 7679 35507
rect 7623 35451 7679 35468
rect 7747 35451 7803 35507
rect 7871 35451 7927 35507
rect 7623 35360 7624 35383
rect 7624 35360 7676 35383
rect 7676 35360 7679 35383
rect 7623 35327 7679 35360
rect 7747 35327 7803 35383
rect 7871 35327 7927 35383
rect 7623 35252 7624 35259
rect 7624 35252 7676 35259
rect 7676 35252 7679 35259
rect 7623 35203 7679 35252
rect 7747 35203 7803 35259
rect 7871 35203 7927 35259
rect 7623 35088 7679 35135
rect 7623 35079 7624 35088
rect 7624 35079 7676 35088
rect 7676 35079 7679 35088
rect 7747 35079 7803 35135
rect 7871 35079 7927 35135
rect 7623 34980 7679 35011
rect 7623 34955 7624 34980
rect 7624 34955 7676 34980
rect 7676 34955 7679 34980
rect 7747 34955 7803 35011
rect 7871 34955 7927 35011
rect 7623 34872 7679 34887
rect 7623 34831 7624 34872
rect 7624 34831 7676 34872
rect 7676 34831 7679 34872
rect 7747 34831 7803 34887
rect 7871 34831 7927 34887
rect 7623 34712 7624 34763
rect 7624 34712 7676 34763
rect 7676 34712 7679 34763
rect 7623 34707 7679 34712
rect 7747 34707 7803 34763
rect 7871 34707 7927 34763
rect 7623 34604 7624 34639
rect 7624 34604 7676 34639
rect 7676 34604 7679 34639
rect 7623 34583 7679 34604
rect 7747 34583 7803 34639
rect 7871 34583 7927 34639
rect 7623 34496 7624 34515
rect 7624 34496 7676 34515
rect 7676 34496 7679 34515
rect 7623 34459 7679 34496
rect 7747 34459 7803 34515
rect 7871 34459 7927 34515
rect 7623 34388 7624 34391
rect 7624 34388 7676 34391
rect 7676 34388 7679 34391
rect 7623 34335 7679 34388
rect 7747 34335 7803 34391
rect 7871 34335 7927 34391
rect 7623 34224 7679 34267
rect 7623 34211 7624 34224
rect 7624 34211 7676 34224
rect 7676 34211 7679 34224
rect 7747 34211 7803 34267
rect 7871 34211 7927 34267
rect 7623 34116 7679 34143
rect 7623 34087 7624 34116
rect 7624 34087 7676 34116
rect 7676 34087 7679 34116
rect 7747 34087 7803 34143
rect 7871 34087 7927 34143
rect 7623 34008 7679 34019
rect 7623 33963 7624 34008
rect 7624 33963 7676 34008
rect 7676 33963 7679 34008
rect 7747 33963 7803 34019
rect 7871 33963 7927 34019
rect 7623 33848 7624 33895
rect 7624 33848 7676 33895
rect 7676 33848 7679 33895
rect 7623 33839 7679 33848
rect 7747 33839 7803 33895
rect 7871 33839 7927 33895
rect 7623 33740 7624 33771
rect 7624 33740 7676 33771
rect 7676 33740 7679 33771
rect 7623 33715 7679 33740
rect 7747 33715 7803 33771
rect 7871 33715 7927 33771
rect 7623 33632 7624 33647
rect 7624 33632 7676 33647
rect 7676 33632 7679 33647
rect 7623 33591 7679 33632
rect 7747 33591 7803 33647
rect 7871 33591 7927 33647
rect 7623 33467 7679 33523
rect 7747 33467 7803 33523
rect 7871 33467 7927 33523
rect 7623 33343 7679 33399
rect 7747 33343 7803 33399
rect 7871 33343 7927 33399
rect 7623 28220 7624 28245
rect 7624 28220 7676 28245
rect 7676 28220 7679 28245
rect 7623 28189 7679 28220
rect 7747 28189 7803 28245
rect 7871 28189 7927 28245
rect 7623 28112 7624 28121
rect 7624 28112 7676 28121
rect 7676 28112 7679 28121
rect 7623 28065 7679 28112
rect 7747 28065 7803 28121
rect 7871 28065 7927 28121
rect 7623 27948 7679 27997
rect 7623 27941 7624 27948
rect 7624 27941 7676 27948
rect 7676 27941 7679 27948
rect 7747 27941 7803 27997
rect 7871 27941 7927 27997
rect 7623 27840 7679 27873
rect 7623 27817 7624 27840
rect 7624 27817 7676 27840
rect 7676 27817 7679 27840
rect 7747 27817 7803 27873
rect 7871 27817 7927 27873
rect 7623 27732 7679 27749
rect 7623 27693 7624 27732
rect 7624 27693 7676 27732
rect 7676 27693 7679 27732
rect 7747 27693 7803 27749
rect 7871 27693 7927 27749
rect 7623 27624 7679 27625
rect 7623 27572 7624 27624
rect 7624 27572 7676 27624
rect 7676 27572 7679 27624
rect 7623 27569 7679 27572
rect 7747 27569 7803 27625
rect 7871 27569 7927 27625
rect 7623 27464 7624 27501
rect 7624 27464 7676 27501
rect 7676 27464 7679 27501
rect 7623 27445 7679 27464
rect 7747 27445 7803 27501
rect 7871 27445 7927 27501
rect 7623 27356 7624 27377
rect 7624 27356 7676 27377
rect 7676 27356 7679 27377
rect 7623 27321 7679 27356
rect 7747 27321 7803 27377
rect 7871 27321 7927 27377
rect 7623 27248 7624 27253
rect 7624 27248 7676 27253
rect 7676 27248 7679 27253
rect 7623 27197 7679 27248
rect 7747 27197 7803 27253
rect 7871 27197 7927 27253
rect 7623 27084 7679 27129
rect 7623 27073 7624 27084
rect 7624 27073 7676 27084
rect 7676 27073 7679 27084
rect 7747 27073 7803 27129
rect 7871 27073 7927 27129
rect 7623 26976 7679 27005
rect 7623 26949 7624 26976
rect 7624 26949 7676 26976
rect 7676 26949 7679 26976
rect 7747 26949 7803 27005
rect 7871 26949 7927 27005
rect 8656 55422 8712 55445
rect 8656 55389 8677 55422
rect 8677 55389 8712 55422
rect 8780 55389 8836 55445
rect 8904 55389 8960 55445
rect 9028 55389 9084 55445
rect 8656 55314 8712 55321
rect 8656 55265 8677 55314
rect 8677 55265 8712 55314
rect 8780 55265 8836 55321
rect 8904 55265 8960 55321
rect 9028 55265 9084 55321
rect 8656 55154 8677 55197
rect 8677 55154 8712 55197
rect 8656 55141 8712 55154
rect 8780 55141 8836 55197
rect 8904 55141 8960 55197
rect 9028 55141 9084 55197
rect 8656 55046 8677 55073
rect 8677 55046 8712 55073
rect 8656 55017 8712 55046
rect 8780 55017 8836 55073
rect 8904 55017 8960 55073
rect 9028 55017 9084 55073
rect 8656 54938 8677 54949
rect 8677 54938 8712 54949
rect 8656 54893 8712 54938
rect 8780 54893 8836 54949
rect 8904 54893 8960 54949
rect 9028 54893 9084 54949
rect 8656 54774 8712 54825
rect 8656 54769 8677 54774
rect 8677 54769 8712 54774
rect 8780 54769 8836 54825
rect 8904 54769 8960 54825
rect 9028 54769 9084 54825
rect 8656 54666 8712 54701
rect 8656 54645 8677 54666
rect 8677 54645 8712 54666
rect 8780 54645 8836 54701
rect 8904 54645 8960 54701
rect 9028 54645 9084 54701
rect 8656 54558 8712 54577
rect 8656 54521 8677 54558
rect 8677 54521 8712 54558
rect 8780 54521 8836 54577
rect 8904 54521 8960 54577
rect 9028 54521 9084 54577
rect 8656 54450 8712 54453
rect 8656 54398 8677 54450
rect 8677 54398 8712 54450
rect 8656 54397 8712 54398
rect 8780 54397 8836 54453
rect 8904 54397 8960 54453
rect 9028 54397 9084 54453
rect 8656 54290 8677 54329
rect 8677 54290 8712 54329
rect 8656 54273 8712 54290
rect 8780 54273 8836 54329
rect 8904 54273 8960 54329
rect 9028 54273 9084 54329
rect 8656 54182 8677 54205
rect 8677 54182 8712 54205
rect 8656 54149 8712 54182
rect 8780 54149 8836 54205
rect 8904 54149 8960 54205
rect 9028 54149 9084 54205
rect 8656 47418 8712 47445
rect 8656 47389 8677 47418
rect 8677 47389 8712 47418
rect 8780 47389 8836 47445
rect 8904 47389 8960 47445
rect 9028 47389 9084 47445
rect 8656 47310 8712 47321
rect 8656 47265 8677 47310
rect 8677 47265 8712 47310
rect 8780 47265 8836 47321
rect 8904 47265 8960 47321
rect 9028 47265 9084 47321
rect 8656 47150 8677 47197
rect 8677 47150 8712 47197
rect 8656 47141 8712 47150
rect 8780 47141 8836 47197
rect 8904 47141 8960 47197
rect 9028 47141 9084 47197
rect 8656 47042 8677 47073
rect 8677 47042 8712 47073
rect 8656 47017 8712 47042
rect 8780 47017 8836 47073
rect 8904 47017 8960 47073
rect 9028 47017 9084 47073
rect 8656 46934 8677 46949
rect 8677 46934 8712 46949
rect 8656 46893 8712 46934
rect 8780 46893 8836 46949
rect 8904 46893 8960 46949
rect 9028 46893 9084 46949
rect 8656 46770 8712 46825
rect 8656 46769 8677 46770
rect 8677 46769 8712 46770
rect 8780 46769 8836 46825
rect 8904 46769 8960 46825
rect 9028 46769 9084 46825
rect 8656 46662 8712 46701
rect 8656 46645 8677 46662
rect 8677 46645 8712 46662
rect 8780 46645 8836 46701
rect 8904 46645 8960 46701
rect 9028 46645 9084 46701
rect 8656 46554 8712 46577
rect 8656 46521 8677 46554
rect 8677 46521 8712 46554
rect 8780 46521 8836 46577
rect 8904 46521 8960 46577
rect 9028 46521 9084 46577
rect 8656 46446 8712 46453
rect 8656 46397 8677 46446
rect 8677 46397 8712 46446
rect 8780 46397 8836 46453
rect 8904 46397 8960 46453
rect 9028 46397 9084 46453
rect 8656 46286 8677 46329
rect 8677 46286 8712 46329
rect 8656 46273 8712 46286
rect 8780 46273 8836 46329
rect 8904 46273 8960 46329
rect 9028 46273 9084 46329
rect 8656 46178 8677 46205
rect 8677 46178 8712 46205
rect 8656 46149 8712 46178
rect 8780 46149 8836 46205
rect 8904 46149 8960 46205
rect 9028 46149 9084 46205
rect 8656 44226 8712 44245
rect 8656 44189 8677 44226
rect 8677 44189 8712 44226
rect 8780 44189 8836 44245
rect 8904 44189 8960 44245
rect 9028 44189 9084 44245
rect 8656 44118 8712 44121
rect 8656 44066 8677 44118
rect 8677 44066 8712 44118
rect 8656 44065 8712 44066
rect 8780 44065 8836 44121
rect 8904 44065 8960 44121
rect 9028 44065 9084 44121
rect 8656 43958 8677 43997
rect 8677 43958 8712 43997
rect 8656 43941 8712 43958
rect 8780 43941 8836 43997
rect 8904 43941 8960 43997
rect 9028 43941 9084 43997
rect 8656 43850 8677 43873
rect 8677 43850 8712 43873
rect 8656 43817 8712 43850
rect 8780 43817 8836 43873
rect 8904 43817 8960 43873
rect 9028 43817 9084 43873
rect 8656 43742 8677 43749
rect 8677 43742 8712 43749
rect 8656 43693 8712 43742
rect 8780 43693 8836 43749
rect 8904 43693 8960 43749
rect 9028 43693 9084 43749
rect 8656 43578 8712 43625
rect 8656 43569 8677 43578
rect 8677 43569 8712 43578
rect 8780 43569 8836 43625
rect 8904 43569 8960 43625
rect 9028 43569 9084 43625
rect 8656 43470 8712 43501
rect 8656 43445 8677 43470
rect 8677 43445 8712 43470
rect 8780 43445 8836 43501
rect 8904 43445 8960 43501
rect 9028 43445 9084 43501
rect 8656 43362 8712 43377
rect 8656 43321 8677 43362
rect 8677 43321 8712 43362
rect 8780 43321 8836 43377
rect 8904 43321 8960 43377
rect 9028 43321 9084 43377
rect 8656 43202 8677 43253
rect 8677 43202 8712 43253
rect 8656 43197 8712 43202
rect 8780 43197 8836 43253
rect 8904 43197 8960 43253
rect 9028 43197 9084 43253
rect 8656 43094 8677 43129
rect 8677 43094 8712 43129
rect 8656 43073 8712 43094
rect 8780 43073 8836 43129
rect 8904 43073 8960 43129
rect 9028 43073 9084 43129
rect 8656 42986 8677 43005
rect 8677 42986 8712 43005
rect 8656 42949 8712 42986
rect 8780 42949 8836 43005
rect 8904 42949 8960 43005
rect 9028 42949 9084 43005
rect 8656 42606 8712 42645
rect 8656 42589 8677 42606
rect 8677 42589 8712 42606
rect 8780 42589 8836 42645
rect 8904 42589 8960 42645
rect 9028 42589 9084 42645
rect 8656 42498 8712 42521
rect 8656 42465 8677 42498
rect 8677 42465 8712 42498
rect 8780 42465 8836 42521
rect 8904 42465 8960 42521
rect 9028 42465 9084 42521
rect 8656 42390 8712 42397
rect 8656 42341 8677 42390
rect 8677 42341 8712 42390
rect 8780 42341 8836 42397
rect 8904 42341 8960 42397
rect 9028 42341 9084 42397
rect 8656 42230 8677 42273
rect 8677 42230 8712 42273
rect 8656 42217 8712 42230
rect 8780 42217 8836 42273
rect 8904 42217 8960 42273
rect 9028 42217 9084 42273
rect 8656 42122 8677 42149
rect 8677 42122 8712 42149
rect 8656 42093 8712 42122
rect 8780 42093 8836 42149
rect 8904 42093 8960 42149
rect 9028 42093 9084 42149
rect 8656 42014 8677 42025
rect 8677 42014 8712 42025
rect 8656 41969 8712 42014
rect 8780 41969 8836 42025
rect 8904 41969 8960 42025
rect 9028 41969 9084 42025
rect 8656 41850 8712 41901
rect 8656 41845 8677 41850
rect 8677 41845 8712 41850
rect 8780 41845 8836 41901
rect 8904 41845 8960 41901
rect 9028 41845 9084 41901
rect 8656 41742 8712 41777
rect 8656 41721 8677 41742
rect 8677 41721 8712 41742
rect 8780 41721 8836 41777
rect 8904 41721 8960 41777
rect 9028 41721 9084 41777
rect 8656 41634 8712 41653
rect 8656 41597 8677 41634
rect 8677 41597 8712 41634
rect 8780 41597 8836 41653
rect 8904 41597 8960 41653
rect 9028 41597 9084 41653
rect 8656 41526 8712 41529
rect 8656 41474 8677 41526
rect 8677 41474 8712 41526
rect 8656 41473 8712 41474
rect 8780 41473 8836 41529
rect 8904 41473 8960 41529
rect 9028 41473 9084 41529
rect 8656 41366 8677 41405
rect 8677 41366 8712 41405
rect 8656 41349 8712 41366
rect 8780 41349 8836 41405
rect 8904 41349 8960 41405
rect 9028 41349 9084 41405
rect 8656 40989 8712 41045
rect 8780 40989 8836 41045
rect 8904 40989 8960 41045
rect 9028 40989 9084 41045
rect 8656 40865 8712 40921
rect 8780 40865 8836 40921
rect 8904 40865 8960 40921
rect 9028 40865 9084 40921
rect 8656 40741 8712 40797
rect 8780 40741 8836 40797
rect 8904 40741 8960 40797
rect 9028 40741 9084 40797
rect 8656 40617 8712 40673
rect 8780 40617 8836 40673
rect 8904 40617 8960 40673
rect 9028 40617 9084 40673
rect 8656 40494 8712 40549
rect 8656 40493 8677 40494
rect 8677 40493 8712 40494
rect 8780 40493 8836 40549
rect 8904 40493 8960 40549
rect 9028 40493 9084 40549
rect 8656 40386 8712 40425
rect 8656 40369 8677 40386
rect 8677 40369 8712 40386
rect 8780 40369 8836 40425
rect 8904 40369 8960 40425
rect 9028 40369 9084 40425
rect 8656 40278 8712 40301
rect 8656 40245 8677 40278
rect 8677 40245 8712 40278
rect 8780 40245 8836 40301
rect 8904 40245 8960 40301
rect 9028 40245 9084 40301
rect 8656 40170 8712 40177
rect 8656 40121 8677 40170
rect 8677 40121 8712 40170
rect 8780 40121 8836 40177
rect 8904 40121 8960 40177
rect 9028 40121 9084 40177
rect 8656 40010 8677 40053
rect 8677 40010 8712 40053
rect 8656 39997 8712 40010
rect 8780 39997 8836 40053
rect 8904 39997 8960 40053
rect 9028 39997 9084 40053
rect 8656 39902 8677 39929
rect 8677 39902 8712 39929
rect 8656 39873 8712 39902
rect 8780 39873 8836 39929
rect 8904 39873 8960 39929
rect 9028 39873 9084 39929
rect 8656 39794 8677 39805
rect 8677 39794 8712 39805
rect 8656 39749 8712 39794
rect 8780 39749 8836 39805
rect 8904 39749 8960 39805
rect 9028 39749 9084 39805
rect 8656 32995 8712 33051
rect 8780 32995 8836 33051
rect 8904 32995 8960 33051
rect 9028 32995 9084 33051
rect 8656 32871 8712 32927
rect 8780 32871 8836 32927
rect 8904 32871 8960 32927
rect 9028 32871 9084 32927
rect 8656 32747 8712 32803
rect 8780 32747 8836 32803
rect 8904 32747 8960 32803
rect 9028 32747 9084 32803
rect 8656 32623 8712 32679
rect 8780 32623 8836 32679
rect 8904 32623 8960 32679
rect 9028 32623 9084 32679
rect 8656 32546 8677 32555
rect 8677 32546 8712 32555
rect 8656 32499 8712 32546
rect 8780 32499 8836 32555
rect 8904 32499 8960 32555
rect 9028 32499 9084 32555
rect 8656 32382 8712 32431
rect 8656 32375 8677 32382
rect 8677 32375 8712 32382
rect 8780 32375 8836 32431
rect 8904 32375 8960 32431
rect 9028 32375 9084 32431
rect 8656 32274 8712 32307
rect 8656 32251 8677 32274
rect 8677 32251 8712 32274
rect 8780 32251 8836 32307
rect 8904 32251 8960 32307
rect 9028 32251 9084 32307
rect 8656 32166 8712 32183
rect 8656 32127 8677 32166
rect 8677 32127 8712 32166
rect 8780 32127 8836 32183
rect 8904 32127 8960 32183
rect 9028 32127 9084 32183
rect 8656 32058 8712 32059
rect 8656 32006 8677 32058
rect 8677 32006 8712 32058
rect 8656 32003 8712 32006
rect 8780 32003 8836 32059
rect 8904 32003 8960 32059
rect 9028 32003 9084 32059
rect 8656 31898 8677 31935
rect 8677 31898 8712 31935
rect 8656 31879 8712 31898
rect 8780 31879 8836 31935
rect 8904 31879 8960 31935
rect 9028 31879 9084 31935
rect 8656 31790 8677 31811
rect 8677 31790 8712 31811
rect 8656 31755 8712 31790
rect 8780 31755 8836 31811
rect 8904 31755 8960 31811
rect 9028 31755 9084 31811
rect 8656 31682 8677 31687
rect 8677 31682 8712 31687
rect 8656 31631 8712 31682
rect 8780 31631 8836 31687
rect 8904 31631 8960 31687
rect 9028 31631 9084 31687
rect 8656 31518 8712 31563
rect 8656 31507 8677 31518
rect 8677 31507 8712 31518
rect 8780 31507 8836 31563
rect 8904 31507 8960 31563
rect 9028 31507 9084 31563
rect 8656 31410 8712 31439
rect 8656 31383 8677 31410
rect 8677 31383 8712 31410
rect 8780 31383 8836 31439
rect 8904 31383 8960 31439
rect 9028 31383 9084 31439
rect 8656 31302 8712 31315
rect 8656 31259 8677 31302
rect 8677 31259 8712 31302
rect 8780 31259 8836 31315
rect 8904 31259 8960 31315
rect 9028 31259 9084 31315
rect 8656 31142 8677 31191
rect 8677 31142 8712 31191
rect 8656 31135 8712 31142
rect 8780 31135 8836 31191
rect 8904 31135 8960 31191
rect 9028 31135 9084 31191
rect 8656 31034 8677 31067
rect 8677 31034 8712 31067
rect 8656 31011 8712 31034
rect 8780 31011 8836 31067
rect 8904 31011 8960 31067
rect 9028 31011 9084 31067
rect 8656 30926 8677 30943
rect 8677 30926 8712 30943
rect 8656 30887 8712 30926
rect 8780 30887 8836 30943
rect 8904 30887 8960 30943
rect 9028 30887 9084 30943
rect 8656 30818 8677 30819
rect 8677 30818 8712 30819
rect 8656 30763 8712 30818
rect 8780 30763 8836 30819
rect 8904 30763 8960 30819
rect 9028 30763 9084 30819
rect 8656 30654 8712 30695
rect 8656 30639 8677 30654
rect 8677 30639 8712 30654
rect 8780 30639 8836 30695
rect 8904 30639 8960 30695
rect 9028 30639 9084 30695
rect 8656 30546 8712 30571
rect 8656 30515 8677 30546
rect 8677 30515 8712 30546
rect 8780 30515 8836 30571
rect 8904 30515 8960 30571
rect 9028 30515 9084 30571
rect 8656 30438 8712 30447
rect 8656 30391 8677 30438
rect 8677 30391 8712 30438
rect 8780 30391 8836 30447
rect 8904 30391 8960 30447
rect 9028 30391 9084 30447
rect 8656 30278 8677 30323
rect 8677 30278 8712 30323
rect 8656 30267 8712 30278
rect 8780 30267 8836 30323
rect 8904 30267 8960 30323
rect 9028 30267 9084 30323
rect 8656 30170 8677 30199
rect 8677 30170 8712 30199
rect 8656 30143 8712 30170
rect 8780 30143 8836 30199
rect 8904 30143 8960 30199
rect 9028 30143 9084 30199
rect 8656 29790 8712 29845
rect 8656 29789 8677 29790
rect 8677 29789 8712 29790
rect 8780 29789 8836 29845
rect 8904 29789 8960 29845
rect 9028 29789 9084 29845
rect 8656 29682 8712 29721
rect 8656 29665 8677 29682
rect 8677 29665 8712 29682
rect 8780 29665 8836 29721
rect 8904 29665 8960 29721
rect 9028 29665 9084 29721
rect 8656 29574 8712 29597
rect 8656 29541 8677 29574
rect 8677 29541 8712 29574
rect 8780 29541 8836 29597
rect 8904 29541 8960 29597
rect 9028 29541 9084 29597
rect 8656 29417 8712 29473
rect 8780 29417 8836 29473
rect 8904 29417 8960 29473
rect 9028 29417 9084 29473
rect 8656 29293 8712 29349
rect 8780 29293 8836 29349
rect 8904 29293 8960 29349
rect 9028 29293 9084 29349
rect 8656 29169 8712 29225
rect 8780 29169 8836 29225
rect 8904 29169 8960 29225
rect 9028 29169 9084 29225
rect 8656 29045 8712 29101
rect 8780 29045 8836 29101
rect 8904 29045 8960 29101
rect 9028 29045 9084 29101
rect 8656 28921 8712 28977
rect 8780 28921 8836 28977
rect 8904 28921 8960 28977
rect 9028 28921 9084 28977
rect 8656 28797 8712 28853
rect 8780 28797 8836 28853
rect 8904 28797 8960 28853
rect 9028 28797 9084 28853
rect 8656 28673 8712 28729
rect 8780 28673 8836 28729
rect 8904 28673 8960 28729
rect 9028 28673 9084 28729
rect 8656 28598 8677 28605
rect 8677 28598 8712 28605
rect 8656 28549 8712 28598
rect 8780 28549 8836 28605
rect 8904 28549 8960 28605
rect 9028 28549 9084 28605
rect 8656 26598 8712 26651
rect 8656 26595 8677 26598
rect 8677 26595 8712 26598
rect 8780 26595 8836 26651
rect 8904 26595 8960 26651
rect 9028 26595 9084 26651
rect 8656 26490 8712 26527
rect 8656 26471 8677 26490
rect 8677 26471 8712 26490
rect 8780 26471 8836 26527
rect 8904 26471 8960 26527
rect 9028 26471 9084 26527
rect 8656 26382 8712 26403
rect 8656 26347 8677 26382
rect 8677 26347 8712 26382
rect 8780 26347 8836 26403
rect 8904 26347 8960 26403
rect 9028 26347 9084 26403
rect 8656 26274 8712 26279
rect 8656 26223 8677 26274
rect 8677 26223 8712 26274
rect 8780 26223 8836 26279
rect 8904 26223 8960 26279
rect 9028 26223 9084 26279
rect 8656 26114 8677 26155
rect 8677 26114 8712 26155
rect 8656 26099 8712 26114
rect 8780 26099 8836 26155
rect 8904 26099 8960 26155
rect 9028 26099 9084 26155
rect 8656 26006 8677 26031
rect 8677 26006 8712 26031
rect 8656 25975 8712 26006
rect 8780 25975 8836 26031
rect 8904 25975 8960 26031
rect 9028 25975 9084 26031
rect 8656 25898 8677 25907
rect 8677 25898 8712 25907
rect 8656 25851 8712 25898
rect 8780 25851 8836 25907
rect 8904 25851 8960 25907
rect 9028 25851 9084 25907
rect 8656 25734 8712 25783
rect 8656 25727 8677 25734
rect 8677 25727 8712 25734
rect 8780 25727 8836 25783
rect 8904 25727 8960 25783
rect 9028 25727 9084 25783
rect 8656 25626 8712 25659
rect 8656 25603 8677 25626
rect 8677 25603 8712 25626
rect 8780 25603 8836 25659
rect 8904 25603 8960 25659
rect 9028 25603 9084 25659
rect 8656 25479 8712 25535
rect 8780 25479 8836 25535
rect 8904 25479 8960 25535
rect 9028 25479 9084 25535
rect 8656 25355 8712 25411
rect 8780 25355 8836 25411
rect 8904 25355 8960 25411
rect 9028 25355 9084 25411
rect 8656 25231 8712 25287
rect 8780 25231 8836 25287
rect 8904 25231 8960 25287
rect 9028 25231 9084 25287
rect 8656 25107 8712 25163
rect 8780 25107 8836 25163
rect 8904 25107 8960 25163
rect 9028 25107 9084 25163
rect 8656 24983 8712 25039
rect 8780 24983 8836 25039
rect 8904 24983 8960 25039
rect 9028 24983 9084 25039
rect 8656 24859 8712 24915
rect 8780 24859 8836 24915
rect 8904 24859 8960 24915
rect 9028 24859 9084 24915
rect 8656 24735 8712 24791
rect 8780 24735 8836 24791
rect 8904 24735 8960 24791
rect 9028 24735 9084 24791
rect 8656 24650 8677 24667
rect 8677 24650 8712 24667
rect 8656 24611 8712 24650
rect 8780 24611 8836 24667
rect 8904 24611 8960 24667
rect 9028 24611 9084 24667
rect 8656 24542 8677 24543
rect 8677 24542 8712 24543
rect 8656 24487 8712 24542
rect 8780 24487 8836 24543
rect 8904 24487 8960 24543
rect 9028 24487 9084 24543
rect 8656 24378 8712 24419
rect 8656 24363 8677 24378
rect 8677 24363 8712 24378
rect 8780 24363 8836 24419
rect 8904 24363 8960 24419
rect 9028 24363 9084 24419
rect 8656 24270 8712 24295
rect 8656 24239 8677 24270
rect 8677 24239 8712 24270
rect 8780 24239 8836 24295
rect 8904 24239 8960 24295
rect 9028 24239 9084 24295
rect 8656 24162 8712 24171
rect 8656 24115 8677 24162
rect 8677 24115 8712 24162
rect 8780 24115 8836 24171
rect 8904 24115 8960 24171
rect 9028 24115 9084 24171
rect 8656 24002 8677 24047
rect 8677 24002 8712 24047
rect 8656 23991 8712 24002
rect 8780 23991 8836 24047
rect 8904 23991 8960 24047
rect 9028 23991 9084 24047
rect 8656 23894 8677 23923
rect 8677 23894 8712 23923
rect 8656 23867 8712 23894
rect 8780 23867 8836 23923
rect 8904 23867 8960 23923
rect 9028 23867 9084 23923
rect 8656 23786 8677 23799
rect 8677 23786 8712 23799
rect 8656 23743 8712 23786
rect 8780 23743 8836 23799
rect 8904 23743 8960 23799
rect 9028 23743 9084 23799
rect 8656 23406 8712 23451
rect 8656 23395 8677 23406
rect 8677 23395 8712 23406
rect 8780 23395 8836 23451
rect 8904 23395 8960 23451
rect 9028 23395 9084 23451
rect 8656 23298 8712 23327
rect 8656 23271 8677 23298
rect 8677 23271 8712 23298
rect 8780 23271 8836 23327
rect 8904 23271 8960 23327
rect 9028 23271 9084 23327
rect 8656 23190 8712 23203
rect 8656 23147 8677 23190
rect 8677 23147 8712 23190
rect 8780 23147 8836 23203
rect 8904 23147 8960 23203
rect 9028 23147 9084 23203
rect 8656 23030 8677 23079
rect 8677 23030 8712 23079
rect 8656 23023 8712 23030
rect 8780 23023 8836 23079
rect 8904 23023 8960 23079
rect 9028 23023 9084 23079
rect 8656 22922 8677 22955
rect 8677 22922 8712 22955
rect 8656 22899 8712 22922
rect 8780 22899 8836 22955
rect 8904 22899 8960 22955
rect 9028 22899 9084 22955
rect 8656 22814 8677 22831
rect 8677 22814 8712 22831
rect 8656 22775 8712 22814
rect 8780 22775 8836 22831
rect 8904 22775 8960 22831
rect 9028 22775 9084 22831
rect 8656 22706 8677 22707
rect 8677 22706 8712 22707
rect 8656 22651 8712 22706
rect 8780 22651 8836 22707
rect 8904 22651 8960 22707
rect 9028 22651 9084 22707
rect 8656 22542 8712 22583
rect 8656 22527 8677 22542
rect 8677 22527 8712 22542
rect 8780 22527 8836 22583
rect 8904 22527 8960 22583
rect 9028 22527 9084 22583
rect 8656 22434 8712 22459
rect 8656 22403 8677 22434
rect 8677 22403 8712 22434
rect 8780 22403 8836 22459
rect 8904 22403 8960 22459
rect 9028 22403 9084 22459
rect 8656 22326 8712 22335
rect 8656 22279 8677 22326
rect 8677 22279 8712 22326
rect 8780 22279 8836 22335
rect 8904 22279 8960 22335
rect 9028 22279 9084 22335
rect 8656 22166 8677 22211
rect 8677 22166 8712 22211
rect 8656 22155 8712 22166
rect 8780 22155 8836 22211
rect 8904 22155 8960 22211
rect 9028 22155 9084 22211
rect 8656 22058 8677 22087
rect 8677 22058 8712 22087
rect 8656 22031 8712 22058
rect 8780 22031 8836 22087
rect 8904 22031 8960 22087
rect 9028 22031 9084 22087
rect 8656 21950 8677 21963
rect 8677 21950 8712 21963
rect 8656 21907 8712 21950
rect 8780 21907 8836 21963
rect 8904 21907 8960 21963
rect 9028 21907 9084 21963
rect 8656 21786 8712 21839
rect 8656 21783 8677 21786
rect 8677 21783 8712 21786
rect 8780 21783 8836 21839
rect 8904 21783 8960 21839
rect 9028 21783 9084 21839
rect 8656 21678 8712 21715
rect 8656 21659 8677 21678
rect 8677 21659 8712 21678
rect 8780 21659 8836 21715
rect 8904 21659 8960 21715
rect 9028 21659 9084 21715
rect 8656 21535 8712 21591
rect 8780 21535 8836 21591
rect 8904 21535 8960 21591
rect 9028 21535 9084 21591
rect 8656 21411 8712 21467
rect 8780 21411 8836 21467
rect 8904 21411 8960 21467
rect 9028 21411 9084 21467
rect 8656 21287 8712 21343
rect 8780 21287 8836 21343
rect 8904 21287 8960 21343
rect 9028 21287 9084 21343
rect 8656 21163 8712 21219
rect 8780 21163 8836 21219
rect 8904 21163 8960 21219
rect 9028 21163 9084 21219
rect 8656 21039 8712 21095
rect 8780 21039 8836 21095
rect 8904 21039 8960 21095
rect 9028 21039 9084 21095
rect 8656 20915 8712 20971
rect 8780 20915 8836 20971
rect 8904 20915 8960 20971
rect 9028 20915 9084 20971
rect 8656 20791 8712 20847
rect 8780 20791 8836 20847
rect 8904 20791 8960 20847
rect 9028 20791 9084 20847
rect 8656 20667 8712 20723
rect 8780 20667 8836 20723
rect 8904 20667 8960 20723
rect 9028 20667 9084 20723
rect 8656 20577 8712 20599
rect 8780 20577 8836 20599
rect 8904 20577 8960 20599
rect 9028 20577 9084 20599
rect 8656 20543 8680 20577
rect 8680 20543 8712 20577
rect 8780 20543 8788 20577
rect 8788 20543 8836 20577
rect 8904 20543 8952 20577
rect 8952 20543 8960 20577
rect 9028 20543 9060 20577
rect 9060 20543 9084 20577
rect 8656 20195 8712 20251
rect 8780 20195 8836 20251
rect 8904 20195 8960 20251
rect 9028 20195 9084 20251
rect 8656 20071 8712 20127
rect 8780 20071 8836 20127
rect 8904 20071 8960 20127
rect 9028 20071 9084 20127
rect 8656 19947 8712 20003
rect 8780 19947 8836 20003
rect 8904 19947 8960 20003
rect 9028 19947 9084 20003
rect 8656 19823 8712 19879
rect 8780 19823 8836 19879
rect 8904 19823 8960 19879
rect 9028 19823 9084 19879
rect 8656 19699 8712 19755
rect 8780 19699 8836 19755
rect 8904 19699 8960 19755
rect 9028 19699 9084 19755
rect 8656 19584 8712 19631
rect 8780 19584 8836 19631
rect 8904 19584 8960 19631
rect 9028 19584 9084 19631
rect 8656 19575 8680 19584
rect 8680 19575 8712 19584
rect 8780 19575 8788 19584
rect 8788 19575 8836 19584
rect 8904 19575 8952 19584
rect 8952 19575 8960 19584
rect 9028 19575 9060 19584
rect 9060 19575 9084 19584
rect 8656 19476 8712 19507
rect 8780 19476 8836 19507
rect 8904 19476 8960 19507
rect 9028 19476 9084 19507
rect 8656 19451 8680 19476
rect 8680 19451 8712 19476
rect 8780 19451 8788 19476
rect 8788 19451 8836 19476
rect 8904 19451 8952 19476
rect 8952 19451 8960 19476
rect 9028 19451 9060 19476
rect 9060 19451 9084 19476
rect 8656 19327 8712 19383
rect 8780 19327 8836 19383
rect 8904 19327 8960 19383
rect 9028 19327 9084 19383
rect 8656 19203 8712 19259
rect 8780 19203 8836 19259
rect 8904 19203 8960 19259
rect 9028 19203 9084 19259
rect 8656 19079 8712 19135
rect 8780 19079 8836 19135
rect 8904 19079 8960 19135
rect 9028 19079 9084 19135
rect 8656 18955 8712 19011
rect 8780 18955 8836 19011
rect 8904 18955 8960 19011
rect 9028 18955 9084 19011
rect 8656 18831 8712 18887
rect 8780 18831 8836 18887
rect 8904 18831 8960 18887
rect 9028 18831 9084 18887
rect 8656 18712 8712 18763
rect 8780 18712 8836 18763
rect 8904 18712 8960 18763
rect 9028 18712 9084 18763
rect 8656 18707 8680 18712
rect 8680 18707 8712 18712
rect 8780 18707 8788 18712
rect 8788 18707 8836 18712
rect 8904 18707 8952 18712
rect 8952 18707 8960 18712
rect 9028 18707 9060 18712
rect 9060 18707 9084 18712
rect 8656 18604 8712 18639
rect 8780 18604 8836 18639
rect 8904 18604 8960 18639
rect 9028 18604 9084 18639
rect 8656 18583 8680 18604
rect 8680 18583 8712 18604
rect 8780 18583 8788 18604
rect 8788 18583 8836 18604
rect 8904 18583 8952 18604
rect 8952 18583 8960 18604
rect 9028 18583 9060 18604
rect 9060 18583 9084 18604
rect 8656 18459 8712 18515
rect 8780 18459 8836 18515
rect 8904 18459 8960 18515
rect 9028 18459 9084 18515
rect 8656 18335 8712 18391
rect 8780 18335 8836 18391
rect 8904 18335 8960 18391
rect 9028 18335 9084 18391
rect 8656 18211 8712 18267
rect 8780 18211 8836 18267
rect 8904 18211 8960 18267
rect 9028 18211 9084 18267
rect 8656 18087 8712 18143
rect 8780 18087 8836 18143
rect 8904 18087 8960 18143
rect 9028 18087 9084 18143
rect 8656 17963 8712 18019
rect 8780 17963 8836 18019
rect 8904 17963 8960 18019
rect 9028 17963 9084 18019
rect 8656 17840 8712 17895
rect 8780 17840 8836 17895
rect 8904 17840 8960 17895
rect 9028 17840 9084 17895
rect 8656 17839 8680 17840
rect 8680 17839 8712 17840
rect 8780 17839 8788 17840
rect 8788 17839 8836 17840
rect 8904 17839 8952 17840
rect 8952 17839 8960 17840
rect 9028 17839 9060 17840
rect 9060 17839 9084 17840
rect 8656 17732 8712 17771
rect 8780 17732 8836 17771
rect 8904 17732 8960 17771
rect 9028 17732 9084 17771
rect 8656 17715 8680 17732
rect 8680 17715 8712 17732
rect 8780 17715 8788 17732
rect 8788 17715 8836 17732
rect 8904 17715 8952 17732
rect 8952 17715 8960 17732
rect 9028 17715 9060 17732
rect 9060 17715 9084 17732
rect 8656 17591 8712 17647
rect 8780 17591 8836 17647
rect 8904 17591 8960 17647
rect 9028 17591 9084 17647
rect 8656 17467 8712 17523
rect 8780 17467 8836 17523
rect 8904 17467 8960 17523
rect 9028 17467 9084 17523
rect 8656 17343 8712 17399
rect 8780 17343 8836 17399
rect 8904 17343 8960 17399
rect 9028 17343 9084 17399
rect 8656 16995 8712 17051
rect 8780 16995 8836 17051
rect 8904 16995 8960 17051
rect 9028 16995 9084 17051
rect 8656 16916 8680 16927
rect 8680 16916 8712 16927
rect 8780 16916 8788 16927
rect 8788 16916 8836 16927
rect 8904 16916 8952 16927
rect 8952 16916 8960 16927
rect 9028 16916 9060 16927
rect 9060 16916 9084 16927
rect 8656 16871 8712 16916
rect 8780 16871 8836 16916
rect 8904 16871 8960 16916
rect 9028 16871 9084 16916
rect 8656 16747 8712 16803
rect 8780 16747 8836 16803
rect 8904 16747 8960 16803
rect 9028 16747 9084 16803
rect 8656 16623 8712 16679
rect 8780 16623 8836 16679
rect 8904 16623 8960 16679
rect 9028 16623 9084 16679
rect 8656 16499 8712 16555
rect 8780 16499 8836 16555
rect 8904 16499 8960 16555
rect 9028 16499 9084 16555
rect 8656 16375 8712 16431
rect 8780 16375 8836 16431
rect 8904 16375 8960 16431
rect 9028 16375 9084 16431
rect 8656 16251 8712 16307
rect 8780 16251 8836 16307
rect 8904 16251 8960 16307
rect 9028 16251 9084 16307
rect 8656 16127 8712 16183
rect 8780 16127 8836 16183
rect 8904 16127 8960 16183
rect 9028 16127 9084 16183
rect 8656 16031 8680 16059
rect 8680 16031 8712 16059
rect 8780 16031 8788 16059
rect 8788 16031 8836 16059
rect 8904 16031 8952 16059
rect 8952 16031 8960 16059
rect 9028 16031 9060 16059
rect 9060 16031 9084 16059
rect 8656 16003 8712 16031
rect 8780 16003 8836 16031
rect 8904 16003 8960 16031
rect 9028 16003 9084 16031
rect 8656 15923 8680 15935
rect 8680 15923 8712 15935
rect 8780 15923 8788 15935
rect 8788 15923 8836 15935
rect 8904 15923 8952 15935
rect 8952 15923 8960 15935
rect 9028 15923 9060 15935
rect 9060 15923 9084 15935
rect 8656 15879 8712 15923
rect 8780 15879 8836 15923
rect 8904 15879 8960 15923
rect 9028 15879 9084 15923
rect 5980 15631 6036 15687
rect 6104 15631 6160 15687
rect 6228 15631 6284 15687
rect 6352 15631 6408 15687
rect 5980 15507 6036 15563
rect 6104 15507 6160 15563
rect 6228 15507 6284 15563
rect 6352 15507 6408 15563
rect 5980 15383 6036 15439
rect 6104 15383 6160 15439
rect 6228 15383 6284 15439
rect 6352 15383 6408 15439
rect 5980 15259 6036 15315
rect 6104 15259 6160 15315
rect 6228 15259 6284 15315
rect 6352 15259 6408 15315
rect 5980 15135 6036 15191
rect 6104 15135 6160 15191
rect 6228 15135 6284 15191
rect 6352 15135 6408 15191
rect 5980 15011 6036 15067
rect 6104 15011 6160 15067
rect 6228 15011 6284 15067
rect 6352 15011 6408 15067
rect 5980 14887 6036 14943
rect 6104 14887 6160 14943
rect 6228 14887 6284 14943
rect 6352 14887 6408 14943
rect 5980 14763 6036 14819
rect 6104 14763 6160 14819
rect 6228 14763 6284 14819
rect 6352 14763 6408 14819
rect 5980 14639 6036 14695
rect 6104 14639 6160 14695
rect 6228 14639 6284 14695
rect 6352 14639 6408 14695
rect 5980 14515 6036 14571
rect 6104 14515 6160 14571
rect 6228 14515 6284 14571
rect 6352 14515 6408 14571
rect 5980 14391 6036 14447
rect 6104 14391 6160 14447
rect 6228 14391 6284 14447
rect 6352 14391 6408 14447
rect 5980 14267 6036 14323
rect 6104 14267 6160 14323
rect 6228 14267 6284 14323
rect 6352 14267 6408 14323
rect 5980 14143 6036 14199
rect 6104 14143 6160 14199
rect 6228 14143 6284 14199
rect 6352 14143 6408 14199
rect 8656 15755 8712 15811
rect 8780 15755 8836 15811
rect 8904 15755 8960 15811
rect 9028 15755 9084 15811
rect 9792 56866 9848 56922
rect 9916 56866 9972 56922
rect 10040 56866 10096 56922
rect 10164 56866 10220 56922
rect 9792 56742 9848 56798
rect 9916 56742 9972 56798
rect 10040 56742 10096 56798
rect 10164 56742 10220 56798
rect 9792 56659 9816 56674
rect 9816 56659 9848 56674
rect 9916 56659 9924 56674
rect 9924 56659 9972 56674
rect 10040 56659 10088 56674
rect 10088 56659 10096 56674
rect 10164 56659 10196 56674
rect 10196 56659 10220 56674
rect 9792 56618 9848 56659
rect 9916 56618 9972 56659
rect 10040 56618 10096 56659
rect 10164 56618 10220 56659
rect 9792 56495 9848 56550
rect 9916 56495 9972 56550
rect 10040 56495 10096 56550
rect 10164 56495 10220 56550
rect 9792 56494 9816 56495
rect 9816 56494 9848 56495
rect 9916 56494 9924 56495
rect 9924 56494 9972 56495
rect 10040 56494 10088 56495
rect 10088 56494 10096 56495
rect 10164 56494 10196 56495
rect 10196 56494 10220 56495
rect 9792 56370 9848 56426
rect 9916 56370 9972 56426
rect 10040 56370 10096 56426
rect 10164 56370 10220 56426
rect 9792 56246 9848 56302
rect 9916 56246 9972 56302
rect 10040 56246 10096 56302
rect 10164 56246 10220 56302
rect 9792 56122 9848 56178
rect 9916 56122 9972 56178
rect 10040 56122 10096 56178
rect 10164 56122 10220 56178
rect 9792 55998 9848 56054
rect 9916 55998 9972 56054
rect 10040 55998 10096 56054
rect 10164 55998 10220 56054
rect 9792 55874 9848 55930
rect 9916 55874 9972 55930
rect 10040 55874 10096 55930
rect 10164 55874 10220 55930
rect 9792 55750 9848 55806
rect 9916 55750 9972 55806
rect 10040 55750 10096 55806
rect 10164 55750 10220 55806
rect 9792 53789 9848 53845
rect 9916 53789 9972 53845
rect 10040 53789 10096 53845
rect 10164 53789 10220 53845
rect 9792 53665 9848 53721
rect 9916 53665 9972 53721
rect 10040 53665 10096 53721
rect 10164 53665 10220 53721
rect 9792 53541 9848 53597
rect 9916 53541 9972 53597
rect 10040 53541 10096 53597
rect 10164 53541 10220 53597
rect 9792 53417 9848 53473
rect 9916 53417 9972 53473
rect 10040 53417 10096 53473
rect 10164 53417 10220 53473
rect 9792 53293 9848 53349
rect 9916 53293 9972 53349
rect 10040 53293 10096 53349
rect 10164 53293 10220 53349
rect 9792 53169 9848 53225
rect 9916 53169 9972 53225
rect 10040 53169 10096 53225
rect 10164 53169 10220 53225
rect 9792 53048 9848 53101
rect 9792 53045 9794 53048
rect 9794 53045 9846 53048
rect 9846 53045 9848 53048
rect 9916 53048 9972 53101
rect 9916 53045 9918 53048
rect 9918 53045 9970 53048
rect 9970 53045 9972 53048
rect 10040 53048 10096 53101
rect 10040 53045 10042 53048
rect 10042 53045 10094 53048
rect 10094 53045 10096 53048
rect 10164 53048 10220 53101
rect 10164 53045 10166 53048
rect 10166 53045 10218 53048
rect 10218 53045 10220 53048
rect 9792 52924 9848 52977
rect 9792 52921 9794 52924
rect 9794 52921 9846 52924
rect 9846 52921 9848 52924
rect 9916 52924 9972 52977
rect 9916 52921 9918 52924
rect 9918 52921 9970 52924
rect 9970 52921 9972 52924
rect 10040 52924 10096 52977
rect 10040 52921 10042 52924
rect 10042 52921 10094 52924
rect 10094 52921 10096 52924
rect 10164 52924 10220 52977
rect 10164 52921 10166 52924
rect 10166 52921 10218 52924
rect 10218 52921 10220 52924
rect 9792 52800 9848 52853
rect 9792 52797 9794 52800
rect 9794 52797 9846 52800
rect 9846 52797 9848 52800
rect 9916 52800 9972 52853
rect 9916 52797 9918 52800
rect 9918 52797 9970 52800
rect 9970 52797 9972 52800
rect 10040 52800 10096 52853
rect 10040 52797 10042 52800
rect 10042 52797 10094 52800
rect 10094 52797 10096 52800
rect 10164 52800 10220 52853
rect 10164 52797 10166 52800
rect 10166 52797 10218 52800
rect 10218 52797 10220 52800
rect 9792 52676 9848 52729
rect 9792 52673 9794 52676
rect 9794 52673 9846 52676
rect 9846 52673 9848 52676
rect 9916 52676 9972 52729
rect 9916 52673 9918 52676
rect 9918 52673 9970 52676
rect 9970 52673 9972 52676
rect 10040 52676 10096 52729
rect 10040 52673 10042 52676
rect 10042 52673 10094 52676
rect 10094 52673 10096 52676
rect 10164 52676 10220 52729
rect 10164 52673 10166 52676
rect 10166 52673 10218 52676
rect 10218 52673 10220 52676
rect 9792 52552 9848 52605
rect 9792 52549 9794 52552
rect 9794 52549 9846 52552
rect 9846 52549 9848 52552
rect 9916 52552 9972 52605
rect 9916 52549 9918 52552
rect 9918 52549 9970 52552
rect 9970 52549 9972 52552
rect 10040 52552 10096 52605
rect 10040 52549 10042 52552
rect 10042 52549 10094 52552
rect 10094 52549 10096 52552
rect 10164 52552 10220 52605
rect 10164 52549 10166 52552
rect 10166 52549 10218 52552
rect 10218 52549 10220 52552
rect 9792 48989 9848 49045
rect 9916 48989 9972 49045
rect 10040 48989 10096 49045
rect 10164 48989 10220 49045
rect 9792 48865 9848 48921
rect 9916 48865 9972 48921
rect 10040 48865 10096 48921
rect 10164 48865 10220 48921
rect 9792 48741 9848 48797
rect 9916 48741 9972 48797
rect 10040 48741 10096 48797
rect 10164 48741 10220 48797
rect 9792 48617 9848 48673
rect 9916 48617 9972 48673
rect 10040 48617 10096 48673
rect 10164 48617 10220 48673
rect 9792 48493 9848 48549
rect 9916 48493 9972 48549
rect 10040 48493 10096 48549
rect 10164 48493 10220 48549
rect 9792 48369 9848 48425
rect 9916 48369 9972 48425
rect 10040 48369 10096 48425
rect 10164 48369 10220 48425
rect 9792 48245 9848 48301
rect 9916 48245 9972 48301
rect 10040 48245 10096 48301
rect 10164 48245 10220 48301
rect 9792 48121 9848 48177
rect 9916 48121 9972 48177
rect 10040 48121 10096 48177
rect 10164 48121 10220 48177
rect 9792 47997 9848 48053
rect 9916 47997 9972 48053
rect 10040 47997 10096 48053
rect 10164 47997 10220 48053
rect 9792 47873 9848 47929
rect 9916 47873 9972 47929
rect 10040 47873 10096 47929
rect 10164 47873 10220 47929
rect 9792 47749 9848 47805
rect 9916 47749 9972 47805
rect 10040 47749 10096 47805
rect 10164 47749 10220 47805
rect 9792 45789 9848 45845
rect 9916 45789 9972 45845
rect 10040 45789 10096 45845
rect 10164 45789 10220 45845
rect 9792 45665 9848 45721
rect 9916 45665 9972 45721
rect 10040 45665 10096 45721
rect 10164 45665 10220 45721
rect 9792 45541 9848 45597
rect 9916 45541 9972 45597
rect 10040 45541 10096 45597
rect 10164 45541 10220 45597
rect 9792 45417 9848 45473
rect 9916 45417 9972 45473
rect 10040 45417 10096 45473
rect 10164 45417 10220 45473
rect 9792 45293 9848 45349
rect 9916 45293 9972 45349
rect 10040 45293 10096 45349
rect 10164 45293 10220 45349
rect 9792 45169 9848 45225
rect 9916 45169 9972 45225
rect 10040 45169 10096 45225
rect 10164 45169 10220 45225
rect 9792 45100 9794 45101
rect 9794 45100 9846 45101
rect 9846 45100 9848 45101
rect 9792 45045 9848 45100
rect 9916 45100 9918 45101
rect 9918 45100 9970 45101
rect 9970 45100 9972 45101
rect 9916 45045 9972 45100
rect 10040 45100 10042 45101
rect 10042 45100 10094 45101
rect 10094 45100 10096 45101
rect 10040 45045 10096 45100
rect 10164 45100 10166 45101
rect 10166 45100 10218 45101
rect 10218 45100 10220 45101
rect 10164 45045 10220 45100
rect 9792 44976 9794 44977
rect 9794 44976 9846 44977
rect 9846 44976 9848 44977
rect 9792 44921 9848 44976
rect 9916 44976 9918 44977
rect 9918 44976 9970 44977
rect 9970 44976 9972 44977
rect 9916 44921 9972 44976
rect 10040 44976 10042 44977
rect 10042 44976 10094 44977
rect 10094 44976 10096 44977
rect 10040 44921 10096 44976
rect 10164 44976 10166 44977
rect 10166 44976 10218 44977
rect 10218 44976 10220 44977
rect 10164 44921 10220 44976
rect 9792 44852 9794 44853
rect 9794 44852 9846 44853
rect 9846 44852 9848 44853
rect 9792 44797 9848 44852
rect 9916 44852 9918 44853
rect 9918 44852 9970 44853
rect 9970 44852 9972 44853
rect 9916 44797 9972 44852
rect 10040 44852 10042 44853
rect 10042 44852 10094 44853
rect 10094 44852 10096 44853
rect 10040 44797 10096 44852
rect 10164 44852 10166 44853
rect 10166 44852 10218 44853
rect 10218 44852 10220 44853
rect 10164 44797 10220 44852
rect 9792 44728 9794 44729
rect 9794 44728 9846 44729
rect 9846 44728 9848 44729
rect 9792 44673 9848 44728
rect 9916 44728 9918 44729
rect 9918 44728 9970 44729
rect 9970 44728 9972 44729
rect 9916 44673 9972 44728
rect 10040 44728 10042 44729
rect 10042 44728 10094 44729
rect 10094 44728 10096 44729
rect 10040 44673 10096 44728
rect 10164 44728 10166 44729
rect 10166 44728 10218 44729
rect 10218 44728 10220 44729
rect 10164 44673 10220 44728
rect 9792 44604 9794 44605
rect 9794 44604 9846 44605
rect 9846 44604 9848 44605
rect 9792 44549 9848 44604
rect 9916 44604 9918 44605
rect 9918 44604 9970 44605
rect 9970 44604 9972 44605
rect 9916 44549 9972 44604
rect 10040 44604 10042 44605
rect 10042 44604 10094 44605
rect 10094 44604 10096 44605
rect 10040 44549 10096 44604
rect 10164 44604 10166 44605
rect 10166 44604 10218 44605
rect 10218 44604 10220 44605
rect 10164 44549 10220 44604
rect 9792 36195 9848 36251
rect 9916 36195 9972 36251
rect 10040 36195 10096 36251
rect 10164 36195 10220 36251
rect 9792 36071 9848 36127
rect 9916 36071 9972 36127
rect 10040 36071 10096 36127
rect 10164 36071 10220 36127
rect 9792 35947 9848 36003
rect 9916 35947 9972 36003
rect 10040 35947 10096 36003
rect 10164 35947 10220 36003
rect 9792 35823 9848 35879
rect 9916 35823 9972 35879
rect 10040 35823 10096 35879
rect 10164 35823 10220 35879
rect 9792 35699 9848 35755
rect 9916 35699 9972 35755
rect 10040 35699 10096 35755
rect 10164 35699 10220 35755
rect 9792 35575 9848 35631
rect 9916 35575 9972 35631
rect 10040 35575 10096 35631
rect 10164 35575 10220 35631
rect 9792 35451 9848 35507
rect 9916 35451 9972 35507
rect 10040 35451 10096 35507
rect 10164 35451 10220 35507
rect 9792 35327 9848 35383
rect 9916 35327 9972 35383
rect 10040 35327 10096 35383
rect 10164 35327 10220 35383
rect 9792 35203 9848 35259
rect 9916 35203 9972 35259
rect 10040 35203 10096 35259
rect 10164 35203 10220 35259
rect 9792 35079 9848 35135
rect 9916 35079 9972 35135
rect 10040 35079 10096 35135
rect 10164 35079 10220 35135
rect 9792 34955 9848 35011
rect 9916 34955 9972 35011
rect 10040 34955 10096 35011
rect 10164 34955 10220 35011
rect 9792 34831 9848 34887
rect 9916 34831 9972 34887
rect 10040 34831 10096 34887
rect 10164 34831 10220 34887
rect 9792 34707 9848 34763
rect 9916 34707 9972 34763
rect 10040 34707 10096 34763
rect 10164 34707 10220 34763
rect 9792 34583 9848 34639
rect 9916 34583 9972 34639
rect 10040 34583 10096 34639
rect 10164 34583 10220 34639
rect 9792 34459 9848 34515
rect 9916 34459 9972 34515
rect 10040 34459 10096 34515
rect 10164 34459 10220 34515
rect 9792 34335 9848 34391
rect 9916 34335 9972 34391
rect 10040 34335 10096 34391
rect 10164 34335 10220 34391
rect 9792 34211 9848 34267
rect 9916 34211 9972 34267
rect 10040 34211 10096 34267
rect 10164 34211 10220 34267
rect 9792 34087 9848 34143
rect 9916 34087 9972 34143
rect 10040 34087 10096 34143
rect 10164 34087 10220 34143
rect 9792 33963 9848 34019
rect 9916 33963 9972 34019
rect 10040 33963 10096 34019
rect 10164 33963 10220 34019
rect 9792 33839 9848 33895
rect 9916 33839 9972 33895
rect 10040 33839 10096 33895
rect 10164 33839 10220 33895
rect 9792 33715 9848 33771
rect 9916 33715 9972 33771
rect 10040 33715 10096 33771
rect 10164 33715 10220 33771
rect 9792 33591 9848 33647
rect 9916 33591 9972 33647
rect 10040 33591 10096 33647
rect 10164 33591 10220 33647
rect 9792 33467 9848 33523
rect 9916 33467 9972 33523
rect 10040 33467 10096 33523
rect 10164 33467 10220 33523
rect 9792 33343 9848 33399
rect 9916 33343 9972 33399
rect 10040 33343 10096 33399
rect 10164 33343 10220 33399
rect 9792 28189 9848 28245
rect 9916 28189 9972 28245
rect 10040 28189 10096 28245
rect 10164 28189 10220 28245
rect 9792 28065 9848 28121
rect 9916 28065 9972 28121
rect 10040 28065 10096 28121
rect 10164 28065 10220 28121
rect 9792 27941 9848 27997
rect 9916 27941 9972 27997
rect 10040 27941 10096 27997
rect 10164 27941 10220 27997
rect 9792 27817 9848 27873
rect 9916 27817 9972 27873
rect 10040 27817 10096 27873
rect 10164 27817 10220 27873
rect 9792 27693 9848 27749
rect 9916 27693 9972 27749
rect 10040 27693 10096 27749
rect 10164 27693 10220 27749
rect 9792 27569 9848 27625
rect 9916 27569 9972 27625
rect 10040 27569 10096 27625
rect 10164 27569 10220 27625
rect 9792 27445 9848 27501
rect 9916 27445 9972 27501
rect 10040 27445 10096 27501
rect 10164 27445 10220 27501
rect 9792 27321 9848 27377
rect 9916 27321 9972 27377
rect 10040 27321 10096 27377
rect 10164 27321 10220 27377
rect 9792 27197 9848 27253
rect 9916 27197 9972 27253
rect 10040 27197 10096 27253
rect 10164 27197 10220 27253
rect 9792 27073 9848 27129
rect 9916 27073 9972 27129
rect 10040 27073 10096 27129
rect 10164 27073 10220 27129
rect 9792 26949 9848 27005
rect 9916 26949 9972 27005
rect 10040 26949 10096 27005
rect 10164 26949 10220 27005
rect 10928 55389 10984 55445
rect 11052 55389 11108 55445
rect 11176 55389 11232 55445
rect 11300 55422 11356 55445
rect 11300 55389 11335 55422
rect 11335 55389 11356 55422
rect 10928 55265 10984 55321
rect 11052 55265 11108 55321
rect 11176 55265 11232 55321
rect 11300 55314 11356 55321
rect 11300 55265 11335 55314
rect 11335 55265 11356 55314
rect 10928 55141 10984 55197
rect 11052 55141 11108 55197
rect 11176 55141 11232 55197
rect 11300 55154 11335 55197
rect 11335 55154 11356 55197
rect 11300 55141 11356 55154
rect 10928 55017 10984 55073
rect 11052 55017 11108 55073
rect 11176 55017 11232 55073
rect 11300 55046 11335 55073
rect 11335 55046 11356 55073
rect 11300 55017 11356 55046
rect 10928 54893 10984 54949
rect 11052 54893 11108 54949
rect 11176 54893 11232 54949
rect 11300 54938 11335 54949
rect 11335 54938 11356 54949
rect 11300 54893 11356 54938
rect 10928 54769 10984 54825
rect 11052 54769 11108 54825
rect 11176 54769 11232 54825
rect 11300 54774 11356 54825
rect 11300 54769 11335 54774
rect 11335 54769 11356 54774
rect 10928 54645 10984 54701
rect 11052 54645 11108 54701
rect 11176 54645 11232 54701
rect 11300 54666 11356 54701
rect 11300 54645 11335 54666
rect 11335 54645 11356 54666
rect 10928 54521 10984 54577
rect 11052 54521 11108 54577
rect 11176 54521 11232 54577
rect 11300 54558 11356 54577
rect 11300 54521 11335 54558
rect 11335 54521 11356 54558
rect 10928 54397 10984 54453
rect 11052 54397 11108 54453
rect 11176 54397 11232 54453
rect 11300 54450 11356 54453
rect 11300 54398 11335 54450
rect 11335 54398 11356 54450
rect 11300 54397 11356 54398
rect 10928 54273 10984 54329
rect 11052 54273 11108 54329
rect 11176 54273 11232 54329
rect 11300 54290 11335 54329
rect 11335 54290 11356 54329
rect 11300 54273 11356 54290
rect 10928 54149 10984 54205
rect 11052 54149 11108 54205
rect 11176 54149 11232 54205
rect 11300 54182 11335 54205
rect 11335 54182 11356 54205
rect 11300 54149 11356 54182
rect 10928 47389 10984 47445
rect 11052 47389 11108 47445
rect 11176 47389 11232 47445
rect 11300 47418 11356 47445
rect 11300 47389 11335 47418
rect 11335 47389 11356 47418
rect 10928 47265 10984 47321
rect 11052 47265 11108 47321
rect 11176 47265 11232 47321
rect 11300 47310 11356 47321
rect 11300 47265 11335 47310
rect 11335 47265 11356 47310
rect 10928 47141 10984 47197
rect 11052 47141 11108 47197
rect 11176 47141 11232 47197
rect 11300 47150 11335 47197
rect 11335 47150 11356 47197
rect 11300 47141 11356 47150
rect 10928 47017 10984 47073
rect 11052 47017 11108 47073
rect 11176 47017 11232 47073
rect 11300 47042 11335 47073
rect 11335 47042 11356 47073
rect 11300 47017 11356 47042
rect 10928 46893 10984 46949
rect 11052 46893 11108 46949
rect 11176 46893 11232 46949
rect 11300 46934 11335 46949
rect 11335 46934 11356 46949
rect 11300 46893 11356 46934
rect 10928 46769 10984 46825
rect 11052 46769 11108 46825
rect 11176 46769 11232 46825
rect 11300 46770 11356 46825
rect 11300 46769 11335 46770
rect 11335 46769 11356 46770
rect 10928 46645 10984 46701
rect 11052 46645 11108 46701
rect 11176 46645 11232 46701
rect 11300 46662 11356 46701
rect 11300 46645 11335 46662
rect 11335 46645 11356 46662
rect 10928 46521 10984 46577
rect 11052 46521 11108 46577
rect 11176 46521 11232 46577
rect 11300 46554 11356 46577
rect 11300 46521 11335 46554
rect 11335 46521 11356 46554
rect 10928 46397 10984 46453
rect 11052 46397 11108 46453
rect 11176 46397 11232 46453
rect 11300 46446 11356 46453
rect 11300 46397 11335 46446
rect 11335 46397 11356 46446
rect 10928 46273 10984 46329
rect 11052 46273 11108 46329
rect 11176 46273 11232 46329
rect 11300 46286 11335 46329
rect 11335 46286 11356 46329
rect 11300 46273 11356 46286
rect 10928 46149 10984 46205
rect 11052 46149 11108 46205
rect 11176 46149 11232 46205
rect 11300 46178 11335 46205
rect 11335 46178 11356 46205
rect 11300 46149 11356 46178
rect 10928 44189 10984 44245
rect 11052 44189 11108 44245
rect 11176 44189 11232 44245
rect 11300 44226 11356 44245
rect 11300 44189 11335 44226
rect 11335 44189 11356 44226
rect 10928 44065 10984 44121
rect 11052 44065 11108 44121
rect 11176 44065 11232 44121
rect 11300 44118 11356 44121
rect 11300 44066 11335 44118
rect 11335 44066 11356 44118
rect 11300 44065 11356 44066
rect 10928 43941 10984 43997
rect 11052 43941 11108 43997
rect 11176 43941 11232 43997
rect 11300 43958 11335 43997
rect 11335 43958 11356 43997
rect 11300 43941 11356 43958
rect 10928 43817 10984 43873
rect 11052 43817 11108 43873
rect 11176 43817 11232 43873
rect 11300 43850 11335 43873
rect 11335 43850 11356 43873
rect 11300 43817 11356 43850
rect 10928 43693 10984 43749
rect 11052 43693 11108 43749
rect 11176 43693 11232 43749
rect 11300 43742 11335 43749
rect 11335 43742 11356 43749
rect 11300 43693 11356 43742
rect 10928 43569 10984 43625
rect 11052 43569 11108 43625
rect 11176 43569 11232 43625
rect 11300 43578 11356 43625
rect 11300 43569 11335 43578
rect 11335 43569 11356 43578
rect 10928 43445 10984 43501
rect 11052 43445 11108 43501
rect 11176 43445 11232 43501
rect 11300 43470 11356 43501
rect 11300 43445 11335 43470
rect 11335 43445 11356 43470
rect 10928 43321 10984 43377
rect 11052 43321 11108 43377
rect 11176 43321 11232 43377
rect 11300 43362 11356 43377
rect 11300 43321 11335 43362
rect 11335 43321 11356 43362
rect 10928 43197 10984 43253
rect 11052 43197 11108 43253
rect 11176 43197 11232 43253
rect 11300 43202 11335 43253
rect 11335 43202 11356 43253
rect 11300 43197 11356 43202
rect 10928 43073 10984 43129
rect 11052 43073 11108 43129
rect 11176 43073 11232 43129
rect 11300 43094 11335 43129
rect 11335 43094 11356 43129
rect 11300 43073 11356 43094
rect 10928 42949 10984 43005
rect 11052 42949 11108 43005
rect 11176 42949 11232 43005
rect 11300 42986 11335 43005
rect 11335 42986 11356 43005
rect 11300 42949 11356 42986
rect 10928 42589 10984 42645
rect 11052 42589 11108 42645
rect 11176 42589 11232 42645
rect 11300 42606 11356 42645
rect 11300 42589 11335 42606
rect 11335 42589 11356 42606
rect 10928 42465 10984 42521
rect 11052 42465 11108 42521
rect 11176 42465 11232 42521
rect 11300 42498 11356 42521
rect 11300 42465 11335 42498
rect 11335 42465 11356 42498
rect 10928 42341 10984 42397
rect 11052 42341 11108 42397
rect 11176 42341 11232 42397
rect 11300 42390 11356 42397
rect 11300 42341 11335 42390
rect 11335 42341 11356 42390
rect 10928 42217 10984 42273
rect 11052 42217 11108 42273
rect 11176 42217 11232 42273
rect 11300 42230 11335 42273
rect 11335 42230 11356 42273
rect 11300 42217 11356 42230
rect 10928 42093 10984 42149
rect 11052 42093 11108 42149
rect 11176 42093 11232 42149
rect 11300 42122 11335 42149
rect 11335 42122 11356 42149
rect 11300 42093 11356 42122
rect 10928 41969 10984 42025
rect 11052 41969 11108 42025
rect 11176 41969 11232 42025
rect 11300 42014 11335 42025
rect 11335 42014 11356 42025
rect 11300 41969 11356 42014
rect 10928 41845 10984 41901
rect 11052 41845 11108 41901
rect 11176 41845 11232 41901
rect 11300 41850 11356 41901
rect 11300 41845 11335 41850
rect 11335 41845 11356 41850
rect 10928 41721 10984 41777
rect 11052 41721 11108 41777
rect 11176 41721 11232 41777
rect 11300 41742 11356 41777
rect 11300 41721 11335 41742
rect 11335 41721 11356 41742
rect 10928 41597 10984 41653
rect 11052 41597 11108 41653
rect 11176 41597 11232 41653
rect 11300 41634 11356 41653
rect 11300 41597 11335 41634
rect 11335 41597 11356 41634
rect 10928 41473 10984 41529
rect 11052 41473 11108 41529
rect 11176 41473 11232 41529
rect 11300 41526 11356 41529
rect 11300 41474 11335 41526
rect 11335 41474 11356 41526
rect 11300 41473 11356 41474
rect 10928 41349 10984 41405
rect 11052 41349 11108 41405
rect 11176 41349 11232 41405
rect 11300 41366 11335 41405
rect 11335 41366 11356 41405
rect 11300 41349 11356 41366
rect 10928 40989 10984 41045
rect 11052 40989 11108 41045
rect 11176 40989 11232 41045
rect 11300 40989 11356 41045
rect 10928 40865 10984 40921
rect 11052 40865 11108 40921
rect 11176 40865 11232 40921
rect 11300 40865 11356 40921
rect 10928 40741 10984 40797
rect 11052 40741 11108 40797
rect 11176 40741 11232 40797
rect 11300 40741 11356 40797
rect 10928 40617 10984 40673
rect 11052 40617 11108 40673
rect 11176 40617 11232 40673
rect 11300 40617 11356 40673
rect 10928 40493 10984 40549
rect 11052 40493 11108 40549
rect 11176 40493 11232 40549
rect 11300 40494 11356 40549
rect 11300 40493 11335 40494
rect 11335 40493 11356 40494
rect 10928 40369 10984 40425
rect 11052 40369 11108 40425
rect 11176 40369 11232 40425
rect 11300 40386 11356 40425
rect 11300 40369 11335 40386
rect 11335 40369 11356 40386
rect 10928 40245 10984 40301
rect 11052 40245 11108 40301
rect 11176 40245 11232 40301
rect 11300 40278 11356 40301
rect 11300 40245 11335 40278
rect 11335 40245 11356 40278
rect 10928 40121 10984 40177
rect 11052 40121 11108 40177
rect 11176 40121 11232 40177
rect 11300 40170 11356 40177
rect 11300 40121 11335 40170
rect 11335 40121 11356 40170
rect 10928 39997 10984 40053
rect 11052 39997 11108 40053
rect 11176 39997 11232 40053
rect 11300 40010 11335 40053
rect 11335 40010 11356 40053
rect 11300 39997 11356 40010
rect 10928 39873 10984 39929
rect 11052 39873 11108 39929
rect 11176 39873 11232 39929
rect 11300 39902 11335 39929
rect 11335 39902 11356 39929
rect 11300 39873 11356 39902
rect 10928 39749 10984 39805
rect 11052 39749 11108 39805
rect 11176 39749 11232 39805
rect 11300 39794 11335 39805
rect 11335 39794 11356 39805
rect 11300 39749 11356 39794
rect 10928 32995 10984 33051
rect 11052 32995 11108 33051
rect 11176 32995 11232 33051
rect 11300 32995 11356 33051
rect 10928 32871 10984 32927
rect 11052 32871 11108 32927
rect 11176 32871 11232 32927
rect 11300 32871 11356 32927
rect 10928 32747 10984 32803
rect 11052 32747 11108 32803
rect 11176 32747 11232 32803
rect 11300 32747 11356 32803
rect 10928 32623 10984 32679
rect 11052 32623 11108 32679
rect 11176 32623 11232 32679
rect 11300 32623 11356 32679
rect 10928 32499 10984 32555
rect 11052 32499 11108 32555
rect 11176 32499 11232 32555
rect 11300 32546 11335 32555
rect 11335 32546 11356 32555
rect 11300 32499 11356 32546
rect 10928 32375 10984 32431
rect 11052 32375 11108 32431
rect 11176 32375 11232 32431
rect 11300 32382 11356 32431
rect 11300 32375 11335 32382
rect 11335 32375 11356 32382
rect 10928 32251 10984 32307
rect 11052 32251 11108 32307
rect 11176 32251 11232 32307
rect 11300 32274 11356 32307
rect 11300 32251 11335 32274
rect 11335 32251 11356 32274
rect 10928 32127 10984 32183
rect 11052 32127 11108 32183
rect 11176 32127 11232 32183
rect 11300 32166 11356 32183
rect 11300 32127 11335 32166
rect 11335 32127 11356 32166
rect 10928 32003 10984 32059
rect 11052 32003 11108 32059
rect 11176 32003 11232 32059
rect 11300 32058 11356 32059
rect 11300 32006 11335 32058
rect 11335 32006 11356 32058
rect 11300 32003 11356 32006
rect 10928 31879 10984 31935
rect 11052 31879 11108 31935
rect 11176 31879 11232 31935
rect 11300 31898 11335 31935
rect 11335 31898 11356 31935
rect 11300 31879 11356 31898
rect 10928 31755 10984 31811
rect 11052 31755 11108 31811
rect 11176 31755 11232 31811
rect 11300 31790 11335 31811
rect 11335 31790 11356 31811
rect 11300 31755 11356 31790
rect 10928 31631 10984 31687
rect 11052 31631 11108 31687
rect 11176 31631 11232 31687
rect 11300 31682 11335 31687
rect 11335 31682 11356 31687
rect 11300 31631 11356 31682
rect 10928 31507 10984 31563
rect 11052 31507 11108 31563
rect 11176 31507 11232 31563
rect 11300 31518 11356 31563
rect 11300 31507 11335 31518
rect 11335 31507 11356 31518
rect 10928 31383 10984 31439
rect 11052 31383 11108 31439
rect 11176 31383 11232 31439
rect 11300 31410 11356 31439
rect 11300 31383 11335 31410
rect 11335 31383 11356 31410
rect 10928 31259 10984 31315
rect 11052 31259 11108 31315
rect 11176 31259 11232 31315
rect 11300 31302 11356 31315
rect 11300 31259 11335 31302
rect 11335 31259 11356 31302
rect 10928 31135 10984 31191
rect 11052 31135 11108 31191
rect 11176 31135 11232 31191
rect 11300 31142 11335 31191
rect 11335 31142 11356 31191
rect 11300 31135 11356 31142
rect 10928 31011 10984 31067
rect 11052 31011 11108 31067
rect 11176 31011 11232 31067
rect 11300 31034 11335 31067
rect 11335 31034 11356 31067
rect 11300 31011 11356 31034
rect 10928 30887 10984 30943
rect 11052 30887 11108 30943
rect 11176 30887 11232 30943
rect 11300 30926 11335 30943
rect 11335 30926 11356 30943
rect 11300 30887 11356 30926
rect 10928 30763 10984 30819
rect 11052 30763 11108 30819
rect 11176 30763 11232 30819
rect 11300 30818 11335 30819
rect 11335 30818 11356 30819
rect 11300 30763 11356 30818
rect 10928 30639 10984 30695
rect 11052 30639 11108 30695
rect 11176 30639 11232 30695
rect 11300 30654 11356 30695
rect 11300 30639 11335 30654
rect 11335 30639 11356 30654
rect 10928 30515 10984 30571
rect 11052 30515 11108 30571
rect 11176 30515 11232 30571
rect 11300 30546 11356 30571
rect 11300 30515 11335 30546
rect 11335 30515 11356 30546
rect 10928 30391 10984 30447
rect 11052 30391 11108 30447
rect 11176 30391 11232 30447
rect 11300 30438 11356 30447
rect 11300 30391 11335 30438
rect 11335 30391 11356 30438
rect 10928 30267 10984 30323
rect 11052 30267 11108 30323
rect 11176 30267 11232 30323
rect 11300 30278 11335 30323
rect 11335 30278 11356 30323
rect 11300 30267 11356 30278
rect 10928 30143 10984 30199
rect 11052 30143 11108 30199
rect 11176 30143 11232 30199
rect 11300 30170 11335 30199
rect 11335 30170 11356 30199
rect 11300 30143 11356 30170
rect 10928 29789 10984 29845
rect 11052 29789 11108 29845
rect 11176 29789 11232 29845
rect 11300 29790 11356 29845
rect 11300 29789 11335 29790
rect 11335 29789 11356 29790
rect 10928 29665 10984 29721
rect 11052 29665 11108 29721
rect 11176 29665 11232 29721
rect 11300 29682 11356 29721
rect 11300 29665 11335 29682
rect 11335 29665 11356 29682
rect 10928 29541 10984 29597
rect 11052 29541 11108 29597
rect 11176 29541 11232 29597
rect 11300 29574 11356 29597
rect 11300 29541 11335 29574
rect 11335 29541 11356 29574
rect 10928 29417 10984 29473
rect 11052 29417 11108 29473
rect 11176 29417 11232 29473
rect 11300 29417 11356 29473
rect 10928 29293 10984 29349
rect 11052 29293 11108 29349
rect 11176 29293 11232 29349
rect 11300 29293 11356 29349
rect 10928 29169 10984 29225
rect 11052 29169 11108 29225
rect 11176 29169 11232 29225
rect 11300 29169 11356 29225
rect 10928 29045 10984 29101
rect 11052 29045 11108 29101
rect 11176 29045 11232 29101
rect 11300 29045 11356 29101
rect 10928 28921 10984 28977
rect 11052 28921 11108 28977
rect 11176 28921 11232 28977
rect 11300 28921 11356 28977
rect 10928 28797 10984 28853
rect 11052 28797 11108 28853
rect 11176 28797 11232 28853
rect 11300 28797 11356 28853
rect 10928 28673 10984 28729
rect 11052 28673 11108 28729
rect 11176 28673 11232 28729
rect 11300 28673 11356 28729
rect 10928 28549 10984 28605
rect 11052 28549 11108 28605
rect 11176 28549 11232 28605
rect 11300 28598 11335 28605
rect 11335 28598 11356 28605
rect 11300 28549 11356 28598
rect 10928 26595 10984 26651
rect 11052 26595 11108 26651
rect 11176 26595 11232 26651
rect 11300 26598 11356 26651
rect 11300 26595 11335 26598
rect 11335 26595 11356 26598
rect 10928 26471 10984 26527
rect 11052 26471 11108 26527
rect 11176 26471 11232 26527
rect 11300 26490 11356 26527
rect 11300 26471 11335 26490
rect 11335 26471 11356 26490
rect 10928 26347 10984 26403
rect 11052 26347 11108 26403
rect 11176 26347 11232 26403
rect 11300 26382 11356 26403
rect 11300 26347 11335 26382
rect 11335 26347 11356 26382
rect 10928 26223 10984 26279
rect 11052 26223 11108 26279
rect 11176 26223 11232 26279
rect 11300 26274 11356 26279
rect 11300 26223 11335 26274
rect 11335 26223 11356 26274
rect 10928 26099 10984 26155
rect 11052 26099 11108 26155
rect 11176 26099 11232 26155
rect 11300 26114 11335 26155
rect 11335 26114 11356 26155
rect 11300 26099 11356 26114
rect 10928 25975 10984 26031
rect 11052 25975 11108 26031
rect 11176 25975 11232 26031
rect 11300 26006 11335 26031
rect 11335 26006 11356 26031
rect 11300 25975 11356 26006
rect 10928 25851 10984 25907
rect 11052 25851 11108 25907
rect 11176 25851 11232 25907
rect 11300 25898 11335 25907
rect 11335 25898 11356 25907
rect 11300 25851 11356 25898
rect 10928 25727 10984 25783
rect 11052 25727 11108 25783
rect 11176 25727 11232 25783
rect 11300 25734 11356 25783
rect 11300 25727 11335 25734
rect 11335 25727 11356 25734
rect 10928 25603 10984 25659
rect 11052 25603 11108 25659
rect 11176 25603 11232 25659
rect 11300 25626 11356 25659
rect 11300 25603 11335 25626
rect 11335 25603 11356 25626
rect 10928 25479 10984 25535
rect 11052 25479 11108 25535
rect 11176 25479 11232 25535
rect 11300 25479 11356 25535
rect 10928 25355 10984 25411
rect 11052 25355 11108 25411
rect 11176 25355 11232 25411
rect 11300 25355 11356 25411
rect 10928 25231 10984 25287
rect 11052 25231 11108 25287
rect 11176 25231 11232 25287
rect 11300 25231 11356 25287
rect 10928 25107 10984 25163
rect 11052 25107 11108 25163
rect 11176 25107 11232 25163
rect 11300 25107 11356 25163
rect 10928 24983 10984 25039
rect 11052 24983 11108 25039
rect 11176 24983 11232 25039
rect 11300 24983 11356 25039
rect 10928 24859 10984 24915
rect 11052 24859 11108 24915
rect 11176 24859 11232 24915
rect 11300 24859 11356 24915
rect 10928 24735 10984 24791
rect 11052 24735 11108 24791
rect 11176 24735 11232 24791
rect 11300 24735 11356 24791
rect 10928 24611 10984 24667
rect 11052 24611 11108 24667
rect 11176 24611 11232 24667
rect 11300 24650 11335 24667
rect 11335 24650 11356 24667
rect 11300 24611 11356 24650
rect 10928 24487 10984 24543
rect 11052 24487 11108 24543
rect 11176 24487 11232 24543
rect 11300 24542 11335 24543
rect 11335 24542 11356 24543
rect 11300 24487 11356 24542
rect 10928 24363 10984 24419
rect 11052 24363 11108 24419
rect 11176 24363 11232 24419
rect 11300 24378 11356 24419
rect 11300 24363 11335 24378
rect 11335 24363 11356 24378
rect 10928 24239 10984 24295
rect 11052 24239 11108 24295
rect 11176 24239 11232 24295
rect 11300 24270 11356 24295
rect 11300 24239 11335 24270
rect 11335 24239 11356 24270
rect 10928 24115 10984 24171
rect 11052 24115 11108 24171
rect 11176 24115 11232 24171
rect 11300 24162 11356 24171
rect 11300 24115 11335 24162
rect 11335 24115 11356 24162
rect 10928 23991 10984 24047
rect 11052 23991 11108 24047
rect 11176 23991 11232 24047
rect 11300 24002 11335 24047
rect 11335 24002 11356 24047
rect 11300 23991 11356 24002
rect 10928 23867 10984 23923
rect 11052 23867 11108 23923
rect 11176 23867 11232 23923
rect 11300 23894 11335 23923
rect 11335 23894 11356 23923
rect 11300 23867 11356 23894
rect 10928 23743 10984 23799
rect 11052 23743 11108 23799
rect 11176 23743 11232 23799
rect 11300 23786 11335 23799
rect 11335 23786 11356 23799
rect 11300 23743 11356 23786
rect 10928 23395 10984 23451
rect 11052 23395 11108 23451
rect 11176 23395 11232 23451
rect 11300 23406 11356 23451
rect 11300 23395 11335 23406
rect 11335 23395 11356 23406
rect 10928 23271 10984 23327
rect 11052 23271 11108 23327
rect 11176 23271 11232 23327
rect 11300 23298 11356 23327
rect 11300 23271 11335 23298
rect 11335 23271 11356 23298
rect 10928 23147 10984 23203
rect 11052 23147 11108 23203
rect 11176 23147 11232 23203
rect 11300 23190 11356 23203
rect 11300 23147 11335 23190
rect 11335 23147 11356 23190
rect 10928 23023 10984 23079
rect 11052 23023 11108 23079
rect 11176 23023 11232 23079
rect 11300 23030 11335 23079
rect 11335 23030 11356 23079
rect 11300 23023 11356 23030
rect 10928 22899 10984 22955
rect 11052 22899 11108 22955
rect 11176 22899 11232 22955
rect 11300 22922 11335 22955
rect 11335 22922 11356 22955
rect 11300 22899 11356 22922
rect 10928 22775 10984 22831
rect 11052 22775 11108 22831
rect 11176 22775 11232 22831
rect 11300 22814 11335 22831
rect 11335 22814 11356 22831
rect 11300 22775 11356 22814
rect 10928 22651 10984 22707
rect 11052 22651 11108 22707
rect 11176 22651 11232 22707
rect 11300 22706 11335 22707
rect 11335 22706 11356 22707
rect 11300 22651 11356 22706
rect 10928 22527 10984 22583
rect 11052 22527 11108 22583
rect 11176 22527 11232 22583
rect 11300 22542 11356 22583
rect 11300 22527 11335 22542
rect 11335 22527 11356 22542
rect 10928 22403 10984 22459
rect 11052 22403 11108 22459
rect 11176 22403 11232 22459
rect 11300 22434 11356 22459
rect 11300 22403 11335 22434
rect 11335 22403 11356 22434
rect 10928 22279 10984 22335
rect 11052 22279 11108 22335
rect 11176 22279 11232 22335
rect 11300 22326 11356 22335
rect 11300 22279 11335 22326
rect 11335 22279 11356 22326
rect 10928 22155 10984 22211
rect 11052 22155 11108 22211
rect 11176 22155 11232 22211
rect 11300 22166 11335 22211
rect 11335 22166 11356 22211
rect 11300 22155 11356 22166
rect 10928 22031 10984 22087
rect 11052 22031 11108 22087
rect 11176 22031 11232 22087
rect 11300 22058 11335 22087
rect 11335 22058 11356 22087
rect 11300 22031 11356 22058
rect 10928 21907 10984 21963
rect 11052 21907 11108 21963
rect 11176 21907 11232 21963
rect 11300 21950 11335 21963
rect 11335 21950 11356 21963
rect 11300 21907 11356 21950
rect 10928 21783 10984 21839
rect 11052 21783 11108 21839
rect 11176 21783 11232 21839
rect 11300 21786 11356 21839
rect 11300 21783 11335 21786
rect 11335 21783 11356 21786
rect 10928 21659 10984 21715
rect 11052 21659 11108 21715
rect 11176 21659 11232 21715
rect 11300 21678 11356 21715
rect 11300 21659 11335 21678
rect 11335 21659 11356 21678
rect 10928 21535 10984 21591
rect 11052 21535 11108 21591
rect 11176 21535 11232 21591
rect 11300 21535 11356 21591
rect 10928 21411 10984 21467
rect 11052 21411 11108 21467
rect 11176 21411 11232 21467
rect 11300 21411 11356 21467
rect 10928 21287 10984 21343
rect 11052 21287 11108 21343
rect 11176 21287 11232 21343
rect 11300 21287 11356 21343
rect 10928 21163 10984 21219
rect 11052 21163 11108 21219
rect 11176 21163 11232 21219
rect 11300 21163 11356 21219
rect 10928 21039 10984 21095
rect 11052 21039 11108 21095
rect 11176 21039 11232 21095
rect 11300 21039 11356 21095
rect 10928 20915 10984 20971
rect 11052 20915 11108 20971
rect 11176 20915 11232 20971
rect 11300 20915 11356 20971
rect 10928 20791 10984 20847
rect 11052 20791 11108 20847
rect 11176 20791 11232 20847
rect 11300 20791 11356 20847
rect 10928 20667 10984 20723
rect 11052 20667 11108 20723
rect 11176 20667 11232 20723
rect 11300 20667 11356 20723
rect 10928 20577 10984 20599
rect 11052 20577 11108 20599
rect 11176 20577 11232 20599
rect 11300 20577 11356 20599
rect 10928 20543 10952 20577
rect 10952 20543 10984 20577
rect 11052 20543 11060 20577
rect 11060 20543 11108 20577
rect 11176 20543 11224 20577
rect 11224 20543 11232 20577
rect 11300 20543 11332 20577
rect 11332 20543 11356 20577
rect 10928 20195 10984 20251
rect 11052 20195 11108 20251
rect 11176 20195 11232 20251
rect 11300 20195 11356 20251
rect 10928 20071 10984 20127
rect 11052 20071 11108 20127
rect 11176 20071 11232 20127
rect 11300 20071 11356 20127
rect 10928 19947 10984 20003
rect 11052 19947 11108 20003
rect 11176 19947 11232 20003
rect 11300 19947 11356 20003
rect 10928 19823 10984 19879
rect 11052 19823 11108 19879
rect 11176 19823 11232 19879
rect 11300 19823 11356 19879
rect 10928 19699 10984 19755
rect 11052 19699 11108 19755
rect 11176 19699 11232 19755
rect 11300 19699 11356 19755
rect 10928 19584 10984 19631
rect 11052 19584 11108 19631
rect 11176 19584 11232 19631
rect 11300 19584 11356 19631
rect 10928 19575 10952 19584
rect 10952 19575 10984 19584
rect 11052 19575 11060 19584
rect 11060 19575 11108 19584
rect 11176 19575 11224 19584
rect 11224 19575 11232 19584
rect 11300 19575 11332 19584
rect 11332 19575 11356 19584
rect 10928 19476 10984 19507
rect 11052 19476 11108 19507
rect 11176 19476 11232 19507
rect 11300 19476 11356 19507
rect 10928 19451 10952 19476
rect 10952 19451 10984 19476
rect 11052 19451 11060 19476
rect 11060 19451 11108 19476
rect 11176 19451 11224 19476
rect 11224 19451 11232 19476
rect 11300 19451 11332 19476
rect 11332 19451 11356 19476
rect 10928 19327 10984 19383
rect 11052 19327 11108 19383
rect 11176 19327 11232 19383
rect 11300 19327 11356 19383
rect 10928 19203 10984 19259
rect 11052 19203 11108 19259
rect 11176 19203 11232 19259
rect 11300 19203 11356 19259
rect 10928 19079 10984 19135
rect 11052 19079 11108 19135
rect 11176 19079 11232 19135
rect 11300 19079 11356 19135
rect 10928 18955 10984 19011
rect 11052 18955 11108 19011
rect 11176 18955 11232 19011
rect 11300 18955 11356 19011
rect 10928 18831 10984 18887
rect 11052 18831 11108 18887
rect 11176 18831 11232 18887
rect 11300 18831 11356 18887
rect 10928 18712 10984 18763
rect 11052 18712 11108 18763
rect 11176 18712 11232 18763
rect 11300 18712 11356 18763
rect 10928 18707 10952 18712
rect 10952 18707 10984 18712
rect 11052 18707 11060 18712
rect 11060 18707 11108 18712
rect 11176 18707 11224 18712
rect 11224 18707 11232 18712
rect 11300 18707 11332 18712
rect 11332 18707 11356 18712
rect 10928 18604 10984 18639
rect 11052 18604 11108 18639
rect 11176 18604 11232 18639
rect 11300 18604 11356 18639
rect 10928 18583 10952 18604
rect 10952 18583 10984 18604
rect 11052 18583 11060 18604
rect 11060 18583 11108 18604
rect 11176 18583 11224 18604
rect 11224 18583 11232 18604
rect 11300 18583 11332 18604
rect 11332 18583 11356 18604
rect 10928 18459 10984 18515
rect 11052 18459 11108 18515
rect 11176 18459 11232 18515
rect 11300 18459 11356 18515
rect 10928 18335 10984 18391
rect 11052 18335 11108 18391
rect 11176 18335 11232 18391
rect 11300 18335 11356 18391
rect 10928 18211 10984 18267
rect 11052 18211 11108 18267
rect 11176 18211 11232 18267
rect 11300 18211 11356 18267
rect 10928 18087 10984 18143
rect 11052 18087 11108 18143
rect 11176 18087 11232 18143
rect 11300 18087 11356 18143
rect 10928 17963 10984 18019
rect 11052 17963 11108 18019
rect 11176 17963 11232 18019
rect 11300 17963 11356 18019
rect 10928 17840 10984 17895
rect 11052 17840 11108 17895
rect 11176 17840 11232 17895
rect 11300 17840 11356 17895
rect 10928 17839 10952 17840
rect 10952 17839 10984 17840
rect 11052 17839 11060 17840
rect 11060 17839 11108 17840
rect 11176 17839 11224 17840
rect 11224 17839 11232 17840
rect 11300 17839 11332 17840
rect 11332 17839 11356 17840
rect 10928 17732 10984 17771
rect 11052 17732 11108 17771
rect 11176 17732 11232 17771
rect 11300 17732 11356 17771
rect 10928 17715 10952 17732
rect 10952 17715 10984 17732
rect 11052 17715 11060 17732
rect 11060 17715 11108 17732
rect 11176 17715 11224 17732
rect 11224 17715 11232 17732
rect 11300 17715 11332 17732
rect 11332 17715 11356 17732
rect 10928 17591 10984 17647
rect 11052 17591 11108 17647
rect 11176 17591 11232 17647
rect 11300 17591 11356 17647
rect 10928 17467 10984 17523
rect 11052 17467 11108 17523
rect 11176 17467 11232 17523
rect 11300 17467 11356 17523
rect 10928 17343 10984 17399
rect 11052 17343 11108 17399
rect 11176 17343 11232 17399
rect 11300 17343 11356 17399
rect 10928 16995 10984 17051
rect 11052 16995 11108 17051
rect 11176 16995 11232 17051
rect 11300 16995 11356 17051
rect 10928 16916 10952 16927
rect 10952 16916 10984 16927
rect 11052 16916 11060 16927
rect 11060 16916 11108 16927
rect 11176 16916 11224 16927
rect 11224 16916 11232 16927
rect 11300 16916 11332 16927
rect 11332 16916 11356 16927
rect 10928 16871 10984 16916
rect 11052 16871 11108 16916
rect 11176 16871 11232 16916
rect 11300 16871 11356 16916
rect 10928 16747 10984 16803
rect 11052 16747 11108 16803
rect 11176 16747 11232 16803
rect 11300 16747 11356 16803
rect 10928 16623 10984 16679
rect 11052 16623 11108 16679
rect 11176 16623 11232 16679
rect 11300 16623 11356 16679
rect 10928 16499 10984 16555
rect 11052 16499 11108 16555
rect 11176 16499 11232 16555
rect 11300 16499 11356 16555
rect 10928 16375 10984 16431
rect 11052 16375 11108 16431
rect 11176 16375 11232 16431
rect 11300 16375 11356 16431
rect 10928 16251 10984 16307
rect 11052 16251 11108 16307
rect 11176 16251 11232 16307
rect 11300 16251 11356 16307
rect 10928 16127 10984 16183
rect 11052 16127 11108 16183
rect 11176 16127 11232 16183
rect 11300 16127 11356 16183
rect 10928 16031 10952 16059
rect 10952 16031 10984 16059
rect 11052 16031 11060 16059
rect 11060 16031 11108 16059
rect 11176 16031 11224 16059
rect 11224 16031 11232 16059
rect 11300 16031 11332 16059
rect 11332 16031 11356 16059
rect 10928 16003 10984 16031
rect 11052 16003 11108 16031
rect 11176 16003 11232 16031
rect 11300 16003 11356 16031
rect 10928 15923 10952 15935
rect 10952 15923 10984 15935
rect 11052 15923 11060 15935
rect 11060 15923 11108 15935
rect 11176 15923 11224 15935
rect 11224 15923 11232 15935
rect 11300 15923 11332 15935
rect 11332 15923 11356 15935
rect 10928 15879 10984 15923
rect 11052 15879 11108 15923
rect 11176 15879 11232 15923
rect 11300 15879 11356 15923
rect 8656 15631 8712 15687
rect 8780 15631 8836 15687
rect 8904 15631 8960 15687
rect 9028 15631 9084 15687
rect 8656 15507 8712 15563
rect 8780 15507 8836 15563
rect 8904 15507 8960 15563
rect 9028 15507 9084 15563
rect 8656 15383 8712 15439
rect 8780 15383 8836 15439
rect 8904 15383 8960 15439
rect 9028 15383 9084 15439
rect 8656 15259 8712 15315
rect 8780 15259 8836 15315
rect 8904 15259 8960 15315
rect 9028 15259 9084 15315
rect 8656 15135 8712 15191
rect 8780 15135 8836 15191
rect 8904 15135 8960 15191
rect 9028 15135 9084 15191
rect 8656 15011 8712 15067
rect 8780 15011 8836 15067
rect 8904 15011 8960 15067
rect 9028 15011 9084 15067
rect 8656 14887 8712 14943
rect 8780 14887 8836 14943
rect 8904 14887 8960 14943
rect 9028 14887 9084 14943
rect 8656 14763 8712 14819
rect 8780 14763 8836 14819
rect 8904 14763 8960 14819
rect 9028 14763 9084 14819
rect 8656 14639 8712 14695
rect 8780 14639 8836 14695
rect 8904 14639 8960 14695
rect 9028 14639 9084 14695
rect 8656 14515 8712 14571
rect 8780 14515 8836 14571
rect 8904 14515 8960 14571
rect 9028 14515 9084 14571
rect 8656 14391 8712 14447
rect 8780 14391 8836 14447
rect 8904 14391 8960 14447
rect 9028 14391 9084 14447
rect 8656 14267 8712 14323
rect 8780 14267 8836 14323
rect 8904 14267 8960 14323
rect 9028 14267 9084 14323
rect 8656 14143 8712 14199
rect 8780 14143 8836 14199
rect 8904 14143 8960 14199
rect 9028 14143 9084 14199
rect 10928 15755 10984 15811
rect 11052 15755 11108 15811
rect 11176 15755 11232 15811
rect 11300 15755 11356 15811
rect 12064 56866 12120 56922
rect 12188 56866 12244 56922
rect 12312 56866 12368 56922
rect 12436 56866 12492 56922
rect 12064 56742 12120 56798
rect 12188 56742 12244 56798
rect 12312 56742 12368 56798
rect 12436 56742 12492 56798
rect 12064 56659 12088 56674
rect 12088 56659 12120 56674
rect 12188 56659 12196 56674
rect 12196 56659 12244 56674
rect 12312 56659 12360 56674
rect 12360 56659 12368 56674
rect 12436 56659 12468 56674
rect 12468 56659 12492 56674
rect 12064 56618 12120 56659
rect 12188 56618 12244 56659
rect 12312 56618 12368 56659
rect 12436 56618 12492 56659
rect 12064 56495 12120 56550
rect 12188 56495 12244 56550
rect 12312 56495 12368 56550
rect 12436 56495 12492 56550
rect 12064 56494 12088 56495
rect 12088 56494 12120 56495
rect 12188 56494 12196 56495
rect 12196 56494 12244 56495
rect 12312 56494 12360 56495
rect 12360 56494 12368 56495
rect 12436 56494 12468 56495
rect 12468 56494 12492 56495
rect 12064 56370 12120 56426
rect 12188 56370 12244 56426
rect 12312 56370 12368 56426
rect 12436 56370 12492 56426
rect 12064 56246 12120 56302
rect 12188 56246 12244 56302
rect 12312 56246 12368 56302
rect 12436 56246 12492 56302
rect 12064 56122 12120 56178
rect 12188 56122 12244 56178
rect 12312 56122 12368 56178
rect 12436 56122 12492 56178
rect 12064 55998 12120 56054
rect 12188 55998 12244 56054
rect 12312 55998 12368 56054
rect 12436 55998 12492 56054
rect 12064 55874 12120 55930
rect 12188 55874 12244 55930
rect 12312 55874 12368 55930
rect 12436 55874 12492 55930
rect 12064 55750 12120 55806
rect 12188 55750 12244 55806
rect 12312 55750 12368 55806
rect 12436 55750 12492 55806
rect 12064 53789 12120 53845
rect 12188 53789 12244 53845
rect 12312 53789 12368 53845
rect 12436 53789 12492 53845
rect 12064 53665 12120 53721
rect 12188 53665 12244 53721
rect 12312 53665 12368 53721
rect 12436 53665 12492 53721
rect 12064 53541 12120 53597
rect 12188 53541 12244 53597
rect 12312 53541 12368 53597
rect 12436 53541 12492 53597
rect 12064 53417 12120 53473
rect 12188 53417 12244 53473
rect 12312 53417 12368 53473
rect 12436 53417 12492 53473
rect 12064 53293 12120 53349
rect 12188 53293 12244 53349
rect 12312 53293 12368 53349
rect 12436 53293 12492 53349
rect 12064 53169 12120 53225
rect 12188 53169 12244 53225
rect 12312 53169 12368 53225
rect 12436 53169 12492 53225
rect 12064 53048 12120 53101
rect 12064 53045 12066 53048
rect 12066 53045 12118 53048
rect 12118 53045 12120 53048
rect 12188 53048 12244 53101
rect 12188 53045 12190 53048
rect 12190 53045 12242 53048
rect 12242 53045 12244 53048
rect 12312 53048 12368 53101
rect 12312 53045 12314 53048
rect 12314 53045 12366 53048
rect 12366 53045 12368 53048
rect 12436 53048 12492 53101
rect 12436 53045 12438 53048
rect 12438 53045 12490 53048
rect 12490 53045 12492 53048
rect 12064 52924 12120 52977
rect 12064 52921 12066 52924
rect 12066 52921 12118 52924
rect 12118 52921 12120 52924
rect 12188 52924 12244 52977
rect 12188 52921 12190 52924
rect 12190 52921 12242 52924
rect 12242 52921 12244 52924
rect 12312 52924 12368 52977
rect 12312 52921 12314 52924
rect 12314 52921 12366 52924
rect 12366 52921 12368 52924
rect 12436 52924 12492 52977
rect 12436 52921 12438 52924
rect 12438 52921 12490 52924
rect 12490 52921 12492 52924
rect 12064 52800 12120 52853
rect 12064 52797 12066 52800
rect 12066 52797 12118 52800
rect 12118 52797 12120 52800
rect 12188 52800 12244 52853
rect 12188 52797 12190 52800
rect 12190 52797 12242 52800
rect 12242 52797 12244 52800
rect 12312 52800 12368 52853
rect 12312 52797 12314 52800
rect 12314 52797 12366 52800
rect 12366 52797 12368 52800
rect 12436 52800 12492 52853
rect 12436 52797 12438 52800
rect 12438 52797 12490 52800
rect 12490 52797 12492 52800
rect 12064 52676 12120 52729
rect 12064 52673 12066 52676
rect 12066 52673 12118 52676
rect 12118 52673 12120 52676
rect 12188 52676 12244 52729
rect 12188 52673 12190 52676
rect 12190 52673 12242 52676
rect 12242 52673 12244 52676
rect 12312 52676 12368 52729
rect 12312 52673 12314 52676
rect 12314 52673 12366 52676
rect 12366 52673 12368 52676
rect 12436 52676 12492 52729
rect 12436 52673 12438 52676
rect 12438 52673 12490 52676
rect 12490 52673 12492 52676
rect 12064 52552 12120 52605
rect 12064 52549 12066 52552
rect 12066 52549 12118 52552
rect 12118 52549 12120 52552
rect 12188 52552 12244 52605
rect 12188 52549 12190 52552
rect 12190 52549 12242 52552
rect 12242 52549 12244 52552
rect 12312 52552 12368 52605
rect 12312 52549 12314 52552
rect 12314 52549 12366 52552
rect 12366 52549 12368 52552
rect 12436 52552 12492 52605
rect 12436 52549 12438 52552
rect 12438 52549 12490 52552
rect 12490 52549 12492 52552
rect 12064 48989 12120 49045
rect 12188 48989 12244 49045
rect 12312 48989 12368 49045
rect 12436 48989 12492 49045
rect 12064 48865 12120 48921
rect 12188 48865 12244 48921
rect 12312 48865 12368 48921
rect 12436 48865 12492 48921
rect 12064 48741 12120 48797
rect 12188 48741 12244 48797
rect 12312 48741 12368 48797
rect 12436 48741 12492 48797
rect 12064 48617 12120 48673
rect 12188 48617 12244 48673
rect 12312 48617 12368 48673
rect 12436 48617 12492 48673
rect 12064 48493 12120 48549
rect 12188 48493 12244 48549
rect 12312 48493 12368 48549
rect 12436 48493 12492 48549
rect 12064 48369 12120 48425
rect 12188 48369 12244 48425
rect 12312 48369 12368 48425
rect 12436 48369 12492 48425
rect 12064 48245 12120 48301
rect 12188 48245 12244 48301
rect 12312 48245 12368 48301
rect 12436 48245 12492 48301
rect 12064 48121 12120 48177
rect 12188 48121 12244 48177
rect 12312 48121 12368 48177
rect 12436 48121 12492 48177
rect 12064 47997 12120 48053
rect 12188 47997 12244 48053
rect 12312 47997 12368 48053
rect 12436 47997 12492 48053
rect 12064 47873 12120 47929
rect 12188 47873 12244 47929
rect 12312 47873 12368 47929
rect 12436 47873 12492 47929
rect 12064 47749 12120 47805
rect 12188 47749 12244 47805
rect 12312 47749 12368 47805
rect 12436 47749 12492 47805
rect 12064 45789 12120 45845
rect 12188 45789 12244 45845
rect 12312 45789 12368 45845
rect 12436 45789 12492 45845
rect 12064 45665 12120 45721
rect 12188 45665 12244 45721
rect 12312 45665 12368 45721
rect 12436 45665 12492 45721
rect 12064 45541 12120 45597
rect 12188 45541 12244 45597
rect 12312 45541 12368 45597
rect 12436 45541 12492 45597
rect 12064 45417 12120 45473
rect 12188 45417 12244 45473
rect 12312 45417 12368 45473
rect 12436 45417 12492 45473
rect 12064 45293 12120 45349
rect 12188 45293 12244 45349
rect 12312 45293 12368 45349
rect 12436 45293 12492 45349
rect 12064 45169 12120 45225
rect 12188 45169 12244 45225
rect 12312 45169 12368 45225
rect 12436 45169 12492 45225
rect 12064 45100 12066 45101
rect 12066 45100 12118 45101
rect 12118 45100 12120 45101
rect 12064 45045 12120 45100
rect 12188 45100 12190 45101
rect 12190 45100 12242 45101
rect 12242 45100 12244 45101
rect 12188 45045 12244 45100
rect 12312 45100 12314 45101
rect 12314 45100 12366 45101
rect 12366 45100 12368 45101
rect 12312 45045 12368 45100
rect 12436 45100 12438 45101
rect 12438 45100 12490 45101
rect 12490 45100 12492 45101
rect 12436 45045 12492 45100
rect 12064 44976 12066 44977
rect 12066 44976 12118 44977
rect 12118 44976 12120 44977
rect 12064 44921 12120 44976
rect 12188 44976 12190 44977
rect 12190 44976 12242 44977
rect 12242 44976 12244 44977
rect 12188 44921 12244 44976
rect 12312 44976 12314 44977
rect 12314 44976 12366 44977
rect 12366 44976 12368 44977
rect 12312 44921 12368 44976
rect 12436 44976 12438 44977
rect 12438 44976 12490 44977
rect 12490 44976 12492 44977
rect 12436 44921 12492 44976
rect 12064 44852 12066 44853
rect 12066 44852 12118 44853
rect 12118 44852 12120 44853
rect 12064 44797 12120 44852
rect 12188 44852 12190 44853
rect 12190 44852 12242 44853
rect 12242 44852 12244 44853
rect 12188 44797 12244 44852
rect 12312 44852 12314 44853
rect 12314 44852 12366 44853
rect 12366 44852 12368 44853
rect 12312 44797 12368 44852
rect 12436 44852 12438 44853
rect 12438 44852 12490 44853
rect 12490 44852 12492 44853
rect 12436 44797 12492 44852
rect 12064 44728 12066 44729
rect 12066 44728 12118 44729
rect 12118 44728 12120 44729
rect 12064 44673 12120 44728
rect 12188 44728 12190 44729
rect 12190 44728 12242 44729
rect 12242 44728 12244 44729
rect 12188 44673 12244 44728
rect 12312 44728 12314 44729
rect 12314 44728 12366 44729
rect 12366 44728 12368 44729
rect 12312 44673 12368 44728
rect 12436 44728 12438 44729
rect 12438 44728 12490 44729
rect 12490 44728 12492 44729
rect 12436 44673 12492 44728
rect 12064 44604 12066 44605
rect 12066 44604 12118 44605
rect 12118 44604 12120 44605
rect 12064 44549 12120 44604
rect 12188 44604 12190 44605
rect 12190 44604 12242 44605
rect 12242 44604 12244 44605
rect 12188 44549 12244 44604
rect 12312 44604 12314 44605
rect 12314 44604 12366 44605
rect 12366 44604 12368 44605
rect 12312 44549 12368 44604
rect 12436 44604 12438 44605
rect 12438 44604 12490 44605
rect 12490 44604 12492 44605
rect 12436 44549 12492 44604
rect 12064 36195 12120 36251
rect 12188 36195 12244 36251
rect 12312 36195 12368 36251
rect 12436 36195 12492 36251
rect 12064 36071 12120 36127
rect 12188 36071 12244 36127
rect 12312 36071 12368 36127
rect 12436 36071 12492 36127
rect 12064 35947 12120 36003
rect 12188 35947 12244 36003
rect 12312 35947 12368 36003
rect 12436 35947 12492 36003
rect 12064 35823 12120 35879
rect 12188 35823 12244 35879
rect 12312 35823 12368 35879
rect 12436 35823 12492 35879
rect 12064 35699 12120 35755
rect 12188 35699 12244 35755
rect 12312 35699 12368 35755
rect 12436 35699 12492 35755
rect 12064 35575 12120 35631
rect 12188 35575 12244 35631
rect 12312 35575 12368 35631
rect 12436 35575 12492 35631
rect 12064 35451 12120 35507
rect 12188 35451 12244 35507
rect 12312 35451 12368 35507
rect 12436 35451 12492 35507
rect 12064 35327 12120 35383
rect 12188 35327 12244 35383
rect 12312 35327 12368 35383
rect 12436 35327 12492 35383
rect 12064 35203 12120 35259
rect 12188 35203 12244 35259
rect 12312 35203 12368 35259
rect 12436 35203 12492 35259
rect 12064 35079 12120 35135
rect 12188 35079 12244 35135
rect 12312 35079 12368 35135
rect 12436 35079 12492 35135
rect 12064 34955 12120 35011
rect 12188 34955 12244 35011
rect 12312 34955 12368 35011
rect 12436 34955 12492 35011
rect 12064 34831 12120 34887
rect 12188 34831 12244 34887
rect 12312 34831 12368 34887
rect 12436 34831 12492 34887
rect 12064 34707 12120 34763
rect 12188 34707 12244 34763
rect 12312 34707 12368 34763
rect 12436 34707 12492 34763
rect 12064 34583 12120 34639
rect 12188 34583 12244 34639
rect 12312 34583 12368 34639
rect 12436 34583 12492 34639
rect 12064 34459 12120 34515
rect 12188 34459 12244 34515
rect 12312 34459 12368 34515
rect 12436 34459 12492 34515
rect 12064 34335 12120 34391
rect 12188 34335 12244 34391
rect 12312 34335 12368 34391
rect 12436 34335 12492 34391
rect 12064 34211 12120 34267
rect 12188 34211 12244 34267
rect 12312 34211 12368 34267
rect 12436 34211 12492 34267
rect 12064 34087 12120 34143
rect 12188 34087 12244 34143
rect 12312 34087 12368 34143
rect 12436 34087 12492 34143
rect 12064 33963 12120 34019
rect 12188 33963 12244 34019
rect 12312 33963 12368 34019
rect 12436 33963 12492 34019
rect 12064 33839 12120 33895
rect 12188 33839 12244 33895
rect 12312 33839 12368 33895
rect 12436 33839 12492 33895
rect 12064 33715 12120 33771
rect 12188 33715 12244 33771
rect 12312 33715 12368 33771
rect 12436 33715 12492 33771
rect 12064 33591 12120 33647
rect 12188 33591 12244 33647
rect 12312 33591 12368 33647
rect 12436 33591 12492 33647
rect 12064 33467 12120 33523
rect 12188 33467 12244 33523
rect 12312 33467 12368 33523
rect 12436 33467 12492 33523
rect 12064 33343 12120 33399
rect 12188 33343 12244 33399
rect 12312 33343 12368 33399
rect 12436 33343 12492 33399
rect 12064 28189 12120 28245
rect 12188 28189 12244 28245
rect 12312 28189 12368 28245
rect 12436 28189 12492 28245
rect 12064 28065 12120 28121
rect 12188 28065 12244 28121
rect 12312 28065 12368 28121
rect 12436 28065 12492 28121
rect 12064 27941 12120 27997
rect 12188 27941 12244 27997
rect 12312 27941 12368 27997
rect 12436 27941 12492 27997
rect 12064 27817 12120 27873
rect 12188 27817 12244 27873
rect 12312 27817 12368 27873
rect 12436 27817 12492 27873
rect 12064 27693 12120 27749
rect 12188 27693 12244 27749
rect 12312 27693 12368 27749
rect 12436 27693 12492 27749
rect 12064 27569 12120 27625
rect 12188 27569 12244 27625
rect 12312 27569 12368 27625
rect 12436 27569 12492 27625
rect 12064 27445 12120 27501
rect 12188 27445 12244 27501
rect 12312 27445 12368 27501
rect 12436 27445 12492 27501
rect 12064 27321 12120 27377
rect 12188 27321 12244 27377
rect 12312 27321 12368 27377
rect 12436 27321 12492 27377
rect 12064 27197 12120 27253
rect 12188 27197 12244 27253
rect 12312 27197 12368 27253
rect 12436 27197 12492 27253
rect 12064 27073 12120 27129
rect 12188 27073 12244 27129
rect 12312 27073 12368 27129
rect 12436 27073 12492 27129
rect 12064 26949 12120 27005
rect 12188 26949 12244 27005
rect 12312 26949 12368 27005
rect 12436 26949 12492 27005
rect 12632 55389 12688 55445
rect 12756 55389 12812 55445
rect 12880 55389 12936 55445
rect 13004 55389 13060 55445
rect 12632 55265 12688 55321
rect 12756 55265 12812 55321
rect 12880 55265 12936 55321
rect 13004 55265 13060 55321
rect 12632 55141 12688 55197
rect 12756 55141 12812 55197
rect 12880 55141 12936 55197
rect 13004 55141 13060 55197
rect 12632 55017 12688 55073
rect 12756 55017 12812 55073
rect 12880 55017 12936 55073
rect 13004 55017 13060 55073
rect 12632 54893 12688 54949
rect 12756 54893 12812 54949
rect 12880 54893 12936 54949
rect 13004 54893 13060 54949
rect 12632 54769 12688 54825
rect 12756 54769 12812 54825
rect 12880 54769 12936 54825
rect 13004 54769 13060 54825
rect 12632 54645 12688 54701
rect 12756 54645 12812 54701
rect 12880 54645 12936 54701
rect 13004 54645 13060 54701
rect 12632 54521 12688 54577
rect 12756 54521 12812 54577
rect 12880 54521 12936 54577
rect 13004 54521 13060 54577
rect 12632 54397 12688 54453
rect 12756 54397 12812 54453
rect 12880 54397 12936 54453
rect 13004 54397 13060 54453
rect 12632 54273 12688 54329
rect 12756 54273 12812 54329
rect 12880 54273 12936 54329
rect 13004 54273 13060 54329
rect 12632 54149 12688 54205
rect 12756 54149 12812 54205
rect 12880 54149 12936 54205
rect 13004 54149 13060 54205
rect 13200 56866 13256 56922
rect 13324 56866 13380 56922
rect 13448 56866 13504 56922
rect 13572 56866 13628 56922
rect 13200 56742 13256 56798
rect 13324 56742 13380 56798
rect 13448 56742 13504 56798
rect 13572 56742 13628 56798
rect 13200 56659 13224 56674
rect 13224 56659 13256 56674
rect 13324 56659 13332 56674
rect 13332 56659 13380 56674
rect 13448 56659 13496 56674
rect 13496 56659 13504 56674
rect 13572 56659 13604 56674
rect 13604 56659 13628 56674
rect 13200 56618 13256 56659
rect 13324 56618 13380 56659
rect 13448 56618 13504 56659
rect 13572 56618 13628 56659
rect 13200 56495 13256 56550
rect 13324 56495 13380 56550
rect 13448 56495 13504 56550
rect 13572 56495 13628 56550
rect 13200 56494 13224 56495
rect 13224 56494 13256 56495
rect 13324 56494 13332 56495
rect 13332 56494 13380 56495
rect 13448 56494 13496 56495
rect 13496 56494 13504 56495
rect 13572 56494 13604 56495
rect 13604 56494 13628 56495
rect 13200 56370 13256 56426
rect 13324 56370 13380 56426
rect 13448 56370 13504 56426
rect 13572 56370 13628 56426
rect 13200 56246 13256 56302
rect 13324 56246 13380 56302
rect 13448 56246 13504 56302
rect 13572 56246 13628 56302
rect 13200 56122 13256 56178
rect 13324 56122 13380 56178
rect 13448 56122 13504 56178
rect 13572 56122 13628 56178
rect 13200 55998 13256 56054
rect 13324 55998 13380 56054
rect 13448 55998 13504 56054
rect 13572 55998 13628 56054
rect 13200 55874 13256 55930
rect 13324 55874 13380 55930
rect 13448 55874 13504 55930
rect 13572 55874 13628 55930
rect 13200 55750 13256 55806
rect 13324 55750 13380 55806
rect 13448 55750 13504 55806
rect 13572 55750 13628 55806
rect 13200 53789 13256 53845
rect 13324 53789 13380 53845
rect 13448 53789 13504 53845
rect 13572 53789 13628 53845
rect 13200 53665 13256 53721
rect 13324 53665 13380 53721
rect 13448 53665 13504 53721
rect 13572 53665 13628 53721
rect 13200 53541 13256 53597
rect 13324 53541 13380 53597
rect 13448 53541 13504 53597
rect 13572 53541 13628 53597
rect 13200 53417 13256 53473
rect 13324 53417 13380 53473
rect 13448 53417 13504 53473
rect 13572 53417 13628 53473
rect 13200 53293 13256 53349
rect 13324 53293 13380 53349
rect 13448 53293 13504 53349
rect 13572 53293 13628 53349
rect 13200 53169 13256 53225
rect 13324 53169 13380 53225
rect 13448 53169 13504 53225
rect 13572 53169 13628 53225
rect 13200 53048 13256 53101
rect 13200 53045 13202 53048
rect 13202 53045 13254 53048
rect 13254 53045 13256 53048
rect 13324 53048 13380 53101
rect 13324 53045 13326 53048
rect 13326 53045 13378 53048
rect 13378 53045 13380 53048
rect 13448 53048 13504 53101
rect 13448 53045 13450 53048
rect 13450 53045 13502 53048
rect 13502 53045 13504 53048
rect 13572 53048 13628 53101
rect 13572 53045 13574 53048
rect 13574 53045 13626 53048
rect 13626 53045 13628 53048
rect 13200 52924 13256 52977
rect 13200 52921 13202 52924
rect 13202 52921 13254 52924
rect 13254 52921 13256 52924
rect 13324 52924 13380 52977
rect 13324 52921 13326 52924
rect 13326 52921 13378 52924
rect 13378 52921 13380 52924
rect 13448 52924 13504 52977
rect 13448 52921 13450 52924
rect 13450 52921 13502 52924
rect 13502 52921 13504 52924
rect 13572 52924 13628 52977
rect 13572 52921 13574 52924
rect 13574 52921 13626 52924
rect 13626 52921 13628 52924
rect 13200 52800 13256 52853
rect 13200 52797 13202 52800
rect 13202 52797 13254 52800
rect 13254 52797 13256 52800
rect 13324 52800 13380 52853
rect 13324 52797 13326 52800
rect 13326 52797 13378 52800
rect 13378 52797 13380 52800
rect 13448 52800 13504 52853
rect 13448 52797 13450 52800
rect 13450 52797 13502 52800
rect 13502 52797 13504 52800
rect 13572 52800 13628 52853
rect 13572 52797 13574 52800
rect 13574 52797 13626 52800
rect 13626 52797 13628 52800
rect 13200 52676 13256 52729
rect 13200 52673 13202 52676
rect 13202 52673 13254 52676
rect 13254 52673 13256 52676
rect 13324 52676 13380 52729
rect 13324 52673 13326 52676
rect 13326 52673 13378 52676
rect 13378 52673 13380 52676
rect 13448 52676 13504 52729
rect 13448 52673 13450 52676
rect 13450 52673 13502 52676
rect 13502 52673 13504 52676
rect 13572 52676 13628 52729
rect 13572 52673 13574 52676
rect 13574 52673 13626 52676
rect 13626 52673 13628 52676
rect 13200 52552 13256 52605
rect 13200 52549 13202 52552
rect 13202 52549 13254 52552
rect 13254 52549 13256 52552
rect 13324 52552 13380 52605
rect 13324 52549 13326 52552
rect 13326 52549 13378 52552
rect 13378 52549 13380 52552
rect 13448 52552 13504 52605
rect 13448 52549 13450 52552
rect 13450 52549 13502 52552
rect 13502 52549 13504 52552
rect 13572 52552 13628 52605
rect 13572 52549 13574 52552
rect 13574 52549 13626 52552
rect 13626 52549 13628 52552
rect 12632 47389 12688 47445
rect 12756 47389 12812 47445
rect 12880 47389 12936 47445
rect 13004 47389 13060 47445
rect 12632 47265 12688 47321
rect 12756 47265 12812 47321
rect 12880 47265 12936 47321
rect 13004 47265 13060 47321
rect 12632 47141 12688 47197
rect 12756 47141 12812 47197
rect 12880 47141 12936 47197
rect 13004 47141 13060 47197
rect 12632 47017 12688 47073
rect 12756 47017 12812 47073
rect 12880 47017 12936 47073
rect 13004 47017 13060 47073
rect 12632 46893 12688 46949
rect 12756 46893 12812 46949
rect 12880 46893 12936 46949
rect 13004 46893 13060 46949
rect 12632 46769 12688 46825
rect 12756 46769 12812 46825
rect 12880 46769 12936 46825
rect 13004 46769 13060 46825
rect 12632 46645 12688 46701
rect 12756 46645 12812 46701
rect 12880 46645 12936 46701
rect 13004 46645 13060 46701
rect 12632 46521 12688 46577
rect 12756 46521 12812 46577
rect 12880 46521 12936 46577
rect 13004 46521 13060 46577
rect 12632 46397 12688 46453
rect 12756 46397 12812 46453
rect 12880 46397 12936 46453
rect 13004 46397 13060 46453
rect 12632 46273 12688 46329
rect 12756 46273 12812 46329
rect 12880 46273 12936 46329
rect 13004 46273 13060 46329
rect 12632 46149 12688 46205
rect 12756 46149 12812 46205
rect 12880 46149 12936 46205
rect 13004 46149 13060 46205
rect 12632 44189 12688 44245
rect 12756 44189 12812 44245
rect 12880 44189 12936 44245
rect 13004 44189 13060 44245
rect 12632 44065 12688 44121
rect 12756 44065 12812 44121
rect 12880 44065 12936 44121
rect 13004 44065 13060 44121
rect 12632 43941 12688 43997
rect 12756 43941 12812 43997
rect 12880 43941 12936 43997
rect 13004 43941 13060 43997
rect 12632 43817 12688 43873
rect 12756 43817 12812 43873
rect 12880 43817 12936 43873
rect 13004 43817 13060 43873
rect 12632 43693 12688 43749
rect 12756 43693 12812 43749
rect 12880 43693 12936 43749
rect 13004 43693 13060 43749
rect 12632 43569 12688 43625
rect 12756 43569 12812 43625
rect 12880 43569 12936 43625
rect 13004 43569 13060 43625
rect 12632 43445 12688 43501
rect 12756 43445 12812 43501
rect 12880 43445 12936 43501
rect 13004 43445 13060 43501
rect 12632 43321 12688 43377
rect 12756 43321 12812 43377
rect 12880 43321 12936 43377
rect 13004 43321 13060 43377
rect 12632 43197 12688 43253
rect 12756 43197 12812 43253
rect 12880 43197 12936 43253
rect 13004 43197 13060 43253
rect 12632 43073 12688 43129
rect 12756 43073 12812 43129
rect 12880 43073 12936 43129
rect 13004 43073 13060 43129
rect 12632 42949 12688 43005
rect 12756 42949 12812 43005
rect 12880 42949 12936 43005
rect 13004 42949 13060 43005
rect 12632 42589 12688 42645
rect 12756 42589 12812 42645
rect 12880 42589 12936 42645
rect 13004 42589 13060 42645
rect 12632 42465 12688 42521
rect 12756 42465 12812 42521
rect 12880 42465 12936 42521
rect 13004 42465 13060 42521
rect 12632 42341 12688 42397
rect 12756 42341 12812 42397
rect 12880 42341 12936 42397
rect 13004 42341 13060 42397
rect 12632 42217 12688 42273
rect 12756 42217 12812 42273
rect 12880 42217 12936 42273
rect 13004 42217 13060 42273
rect 12632 42093 12688 42149
rect 12756 42093 12812 42149
rect 12880 42093 12936 42149
rect 13004 42093 13060 42149
rect 12632 41969 12688 42025
rect 12756 41969 12812 42025
rect 12880 41969 12936 42025
rect 13004 41969 13060 42025
rect 12632 41845 12688 41901
rect 12756 41845 12812 41901
rect 12880 41845 12936 41901
rect 13004 41845 13060 41901
rect 12632 41721 12688 41777
rect 12756 41721 12812 41777
rect 12880 41721 12936 41777
rect 13004 41721 13060 41777
rect 12632 41597 12688 41653
rect 12756 41597 12812 41653
rect 12880 41597 12936 41653
rect 13004 41597 13060 41653
rect 12632 41473 12688 41529
rect 12756 41473 12812 41529
rect 12880 41473 12936 41529
rect 13004 41473 13060 41529
rect 12632 41349 12688 41405
rect 12756 41349 12812 41405
rect 12880 41349 12936 41405
rect 13004 41349 13060 41405
rect 12632 40989 12688 41045
rect 12756 40989 12812 41045
rect 12880 40989 12936 41045
rect 13004 40989 13060 41045
rect 12632 40865 12688 40921
rect 12756 40865 12812 40921
rect 12880 40865 12936 40921
rect 13004 40865 13060 40921
rect 12632 40741 12688 40797
rect 12756 40741 12812 40797
rect 12880 40741 12936 40797
rect 13004 40741 13060 40797
rect 12632 40617 12688 40673
rect 12756 40617 12812 40673
rect 12880 40617 12936 40673
rect 13004 40617 13060 40673
rect 12632 40493 12688 40549
rect 12756 40493 12812 40549
rect 12880 40493 12936 40549
rect 13004 40493 13060 40549
rect 12632 40369 12688 40425
rect 12756 40369 12812 40425
rect 12880 40369 12936 40425
rect 13004 40369 13060 40425
rect 12632 40245 12688 40301
rect 12756 40245 12812 40301
rect 12880 40245 12936 40301
rect 13004 40245 13060 40301
rect 12632 40121 12688 40177
rect 12756 40121 12812 40177
rect 12880 40121 12936 40177
rect 13004 40121 13060 40177
rect 12632 39997 12688 40053
rect 12756 39997 12812 40053
rect 12880 39997 12936 40053
rect 13004 39997 13060 40053
rect 12632 39873 12688 39929
rect 12756 39873 12812 39929
rect 12880 39873 12936 39929
rect 13004 39873 13060 39929
rect 12632 39749 12688 39805
rect 12756 39749 12812 39805
rect 12880 39749 12936 39805
rect 13004 39749 13060 39805
rect 13170 52189 13226 52245
rect 13294 52189 13350 52245
rect 13170 52065 13226 52121
rect 13294 52065 13350 52121
rect 13170 51941 13226 51997
rect 13294 51941 13350 51997
rect 13170 51817 13226 51873
rect 13294 51817 13350 51873
rect 13170 51693 13226 51749
rect 13294 51693 13350 51749
rect 13170 51569 13226 51625
rect 13294 51569 13350 51625
rect 13170 51445 13226 51501
rect 13294 51445 13350 51501
rect 13170 51321 13226 51377
rect 13294 51321 13350 51377
rect 13170 51197 13226 51253
rect 13294 51197 13350 51253
rect 13170 51073 13226 51129
rect 13294 51073 13350 51129
rect 13170 50949 13226 51005
rect 13294 50949 13350 51005
rect 13170 37789 13226 37845
rect 13294 37789 13350 37845
rect 13170 37665 13226 37721
rect 13294 37665 13350 37721
rect 13170 37541 13226 37597
rect 13294 37541 13350 37597
rect 13170 37417 13226 37473
rect 13294 37417 13350 37473
rect 13170 37293 13226 37349
rect 13294 37293 13350 37349
rect 13170 37169 13226 37225
rect 13294 37169 13350 37225
rect 13170 37045 13226 37101
rect 13294 37045 13350 37101
rect 13170 36921 13226 36977
rect 13294 36921 13350 36977
rect 13170 36797 13226 36853
rect 13294 36797 13350 36853
rect 13170 36673 13226 36729
rect 13294 36673 13350 36729
rect 13170 36549 13226 36605
rect 13294 36549 13350 36605
rect 13478 48989 13534 49045
rect 13602 48989 13658 49045
rect 13478 48865 13534 48921
rect 13602 48865 13658 48921
rect 13478 48741 13534 48797
rect 13602 48741 13658 48797
rect 13478 48617 13534 48673
rect 13602 48617 13658 48673
rect 13478 48493 13534 48549
rect 13602 48493 13658 48549
rect 13478 48369 13534 48425
rect 13602 48369 13658 48425
rect 13478 48245 13534 48301
rect 13602 48245 13658 48301
rect 13478 48121 13534 48177
rect 13602 48121 13658 48177
rect 13478 47997 13534 48053
rect 13602 47997 13658 48053
rect 13478 47873 13534 47929
rect 13602 47873 13658 47929
rect 13478 47749 13534 47805
rect 13602 47749 13658 47805
rect 13478 45789 13534 45845
rect 13602 45789 13658 45845
rect 13478 45665 13534 45721
rect 13602 45665 13658 45721
rect 13478 45541 13534 45597
rect 13602 45541 13658 45597
rect 13478 45417 13534 45473
rect 13602 45417 13658 45473
rect 13478 45293 13534 45349
rect 13602 45293 13658 45349
rect 13478 45169 13534 45225
rect 13602 45169 13658 45225
rect 13478 45100 13480 45101
rect 13480 45100 13532 45101
rect 13532 45100 13534 45101
rect 13478 45045 13534 45100
rect 13602 45100 13604 45101
rect 13604 45100 13656 45101
rect 13656 45100 13658 45101
rect 13602 45045 13658 45100
rect 13478 44976 13480 44977
rect 13480 44976 13532 44977
rect 13532 44976 13534 44977
rect 13478 44921 13534 44976
rect 13602 44976 13604 44977
rect 13604 44976 13656 44977
rect 13656 44976 13658 44977
rect 13602 44921 13658 44976
rect 13478 44852 13480 44853
rect 13480 44852 13532 44853
rect 13532 44852 13534 44853
rect 13478 44797 13534 44852
rect 13602 44852 13604 44853
rect 13604 44852 13656 44853
rect 13656 44852 13658 44853
rect 13602 44797 13658 44852
rect 13478 44728 13480 44729
rect 13480 44728 13532 44729
rect 13532 44728 13534 44729
rect 13478 44673 13534 44728
rect 13602 44728 13604 44729
rect 13604 44728 13656 44729
rect 13656 44728 13658 44729
rect 13602 44673 13658 44728
rect 13478 44604 13480 44605
rect 13480 44604 13532 44605
rect 13532 44604 13534 44605
rect 13478 44549 13534 44604
rect 13602 44604 13604 44605
rect 13604 44604 13656 44605
rect 13656 44604 13658 44605
rect 13602 44549 13658 44604
rect 12632 32995 12688 33051
rect 12756 32995 12812 33051
rect 12880 32995 12936 33051
rect 13004 32995 13060 33051
rect 12632 32871 12688 32927
rect 12756 32871 12812 32927
rect 12880 32871 12936 32927
rect 13004 32871 13060 32927
rect 12632 32747 12688 32803
rect 12756 32747 12812 32803
rect 12880 32747 12936 32803
rect 13004 32747 13060 32803
rect 12632 32623 12688 32679
rect 12756 32623 12812 32679
rect 12880 32623 12936 32679
rect 13004 32623 13060 32679
rect 12632 32499 12688 32555
rect 12756 32499 12812 32555
rect 12880 32499 12936 32555
rect 13004 32499 13060 32555
rect 12632 32375 12688 32431
rect 12756 32375 12812 32431
rect 12880 32375 12936 32431
rect 13004 32375 13060 32431
rect 12632 32251 12688 32307
rect 12756 32251 12812 32307
rect 12880 32251 12936 32307
rect 13004 32251 13060 32307
rect 12632 32127 12688 32183
rect 12756 32127 12812 32183
rect 12880 32127 12936 32183
rect 13004 32127 13060 32183
rect 12632 32003 12688 32059
rect 12756 32003 12812 32059
rect 12880 32003 12936 32059
rect 13004 32003 13060 32059
rect 12632 31879 12688 31935
rect 12756 31879 12812 31935
rect 12880 31879 12936 31935
rect 13004 31879 13060 31935
rect 12632 31755 12688 31811
rect 12756 31755 12812 31811
rect 12880 31755 12936 31811
rect 13004 31755 13060 31811
rect 12632 31631 12688 31687
rect 12756 31631 12812 31687
rect 12880 31631 12936 31687
rect 13004 31631 13060 31687
rect 12632 31507 12688 31563
rect 12756 31507 12812 31563
rect 12880 31507 12936 31563
rect 13004 31507 13060 31563
rect 12632 31383 12688 31439
rect 12756 31383 12812 31439
rect 12880 31383 12936 31439
rect 13004 31383 13060 31439
rect 12632 31259 12688 31315
rect 12756 31259 12812 31315
rect 12880 31259 12936 31315
rect 13004 31259 13060 31315
rect 12632 31135 12688 31191
rect 12756 31135 12812 31191
rect 12880 31135 12936 31191
rect 13004 31135 13060 31191
rect 12632 31011 12688 31067
rect 12756 31011 12812 31067
rect 12880 31011 12936 31067
rect 13004 31011 13060 31067
rect 12632 30887 12688 30943
rect 12756 30887 12812 30943
rect 12880 30887 12936 30943
rect 13004 30887 13060 30943
rect 12632 30763 12688 30819
rect 12756 30763 12812 30819
rect 12880 30763 12936 30819
rect 13004 30763 13060 30819
rect 12632 30639 12688 30695
rect 12756 30639 12812 30695
rect 12880 30639 12936 30695
rect 13004 30639 13060 30695
rect 12632 30515 12688 30571
rect 12756 30515 12812 30571
rect 12880 30515 12936 30571
rect 13004 30515 13060 30571
rect 12632 30391 12688 30447
rect 12756 30391 12812 30447
rect 12880 30391 12936 30447
rect 13004 30391 13060 30447
rect 12632 30267 12688 30323
rect 12756 30267 12812 30323
rect 12880 30267 12936 30323
rect 13004 30267 13060 30323
rect 12632 30143 12688 30199
rect 12756 30143 12812 30199
rect 12880 30143 12936 30199
rect 13004 30143 13060 30199
rect 12632 29789 12688 29845
rect 12756 29789 12812 29845
rect 12880 29789 12936 29845
rect 13004 29789 13060 29845
rect 12632 29665 12688 29721
rect 12756 29665 12812 29721
rect 12880 29665 12936 29721
rect 13004 29665 13060 29721
rect 12632 29541 12688 29597
rect 12756 29541 12812 29597
rect 12880 29541 12936 29597
rect 13004 29541 13060 29597
rect 12632 29417 12688 29473
rect 12756 29417 12812 29473
rect 12880 29417 12936 29473
rect 13004 29417 13060 29473
rect 12632 29293 12688 29349
rect 12756 29293 12812 29349
rect 12880 29293 12936 29349
rect 13004 29293 13060 29349
rect 12632 29169 12688 29225
rect 12756 29169 12812 29225
rect 12880 29169 12936 29225
rect 13004 29169 13060 29225
rect 12632 29045 12688 29101
rect 12756 29045 12812 29101
rect 12880 29045 12936 29101
rect 13004 29045 13060 29101
rect 12632 28921 12688 28977
rect 12756 28921 12812 28977
rect 12880 28921 12936 28977
rect 13004 28921 13060 28977
rect 12632 28797 12688 28853
rect 12756 28797 12812 28853
rect 12880 28797 12936 28853
rect 13004 28797 13060 28853
rect 12632 28673 12688 28729
rect 12756 28673 12812 28729
rect 12880 28673 12936 28729
rect 13004 28673 13060 28729
rect 12632 28549 12688 28605
rect 12756 28549 12812 28605
rect 12880 28549 12936 28605
rect 13004 28549 13060 28605
rect 12632 26595 12688 26651
rect 12756 26595 12812 26651
rect 12880 26595 12936 26651
rect 13004 26595 13060 26651
rect 12632 26471 12688 26527
rect 12756 26471 12812 26527
rect 12880 26471 12936 26527
rect 13004 26471 13060 26527
rect 12632 26347 12688 26403
rect 12756 26347 12812 26403
rect 12880 26347 12936 26403
rect 13004 26347 13060 26403
rect 12632 26223 12688 26279
rect 12756 26223 12812 26279
rect 12880 26223 12936 26279
rect 13004 26223 13060 26279
rect 12632 26099 12688 26155
rect 12756 26099 12812 26155
rect 12880 26099 12936 26155
rect 13004 26099 13060 26155
rect 12632 25975 12688 26031
rect 12756 25975 12812 26031
rect 12880 25975 12936 26031
rect 13004 25975 13060 26031
rect 12632 25851 12688 25907
rect 12756 25851 12812 25907
rect 12880 25851 12936 25907
rect 13004 25851 13060 25907
rect 12632 25727 12688 25783
rect 12756 25727 12812 25783
rect 12880 25727 12936 25783
rect 13004 25727 13060 25783
rect 12632 25603 12688 25659
rect 12756 25603 12812 25659
rect 12880 25603 12936 25659
rect 13004 25603 13060 25659
rect 12632 25479 12688 25535
rect 12756 25479 12812 25535
rect 12880 25479 12936 25535
rect 13004 25479 13060 25535
rect 12632 25355 12688 25411
rect 12756 25355 12812 25411
rect 12880 25355 12936 25411
rect 13004 25355 13060 25411
rect 12632 25231 12688 25287
rect 12756 25231 12812 25287
rect 12880 25231 12936 25287
rect 13004 25231 13060 25287
rect 12632 25107 12688 25163
rect 12756 25107 12812 25163
rect 12880 25107 12936 25163
rect 13004 25107 13060 25163
rect 12632 24983 12688 25039
rect 12756 24983 12812 25039
rect 12880 24983 12936 25039
rect 13004 24983 13060 25039
rect 12632 24859 12688 24915
rect 12756 24859 12812 24915
rect 12880 24859 12936 24915
rect 13004 24859 13060 24915
rect 12632 24735 12688 24791
rect 12756 24735 12812 24791
rect 12880 24735 12936 24791
rect 13004 24735 13060 24791
rect 12632 24611 12688 24667
rect 12756 24611 12812 24667
rect 12880 24611 12936 24667
rect 13004 24611 13060 24667
rect 12632 24487 12688 24543
rect 12756 24487 12812 24543
rect 12880 24487 12936 24543
rect 13004 24487 13060 24543
rect 12632 24363 12688 24419
rect 12756 24363 12812 24419
rect 12880 24363 12936 24419
rect 13004 24363 13060 24419
rect 12632 24239 12688 24295
rect 12756 24239 12812 24295
rect 12880 24239 12936 24295
rect 13004 24239 13060 24295
rect 12632 24115 12688 24171
rect 12756 24115 12812 24171
rect 12880 24115 12936 24171
rect 13004 24115 13060 24171
rect 12632 23991 12688 24047
rect 12756 23991 12812 24047
rect 12880 23991 12936 24047
rect 13004 23991 13060 24047
rect 12632 23867 12688 23923
rect 12756 23867 12812 23923
rect 12880 23867 12936 23923
rect 13004 23867 13060 23923
rect 12632 23743 12688 23799
rect 12756 23743 12812 23799
rect 12880 23743 12936 23799
rect 13004 23743 13060 23799
rect 12632 23395 12688 23451
rect 12756 23395 12812 23451
rect 12880 23395 12936 23451
rect 13004 23395 13060 23451
rect 12632 23271 12688 23327
rect 12756 23271 12812 23327
rect 12880 23271 12936 23327
rect 13004 23271 13060 23327
rect 12632 23147 12688 23203
rect 12756 23147 12812 23203
rect 12880 23147 12936 23203
rect 13004 23147 13060 23203
rect 12632 23023 12688 23079
rect 12756 23023 12812 23079
rect 12880 23023 12936 23079
rect 13004 23023 13060 23079
rect 12632 22899 12688 22955
rect 12756 22899 12812 22955
rect 12880 22899 12936 22955
rect 13004 22899 13060 22955
rect 12632 22775 12688 22831
rect 12756 22775 12812 22831
rect 12880 22775 12936 22831
rect 13004 22775 13060 22831
rect 12632 22651 12688 22707
rect 12756 22651 12812 22707
rect 12880 22651 12936 22707
rect 13004 22651 13060 22707
rect 12632 22527 12688 22583
rect 12756 22527 12812 22583
rect 12880 22527 12936 22583
rect 13004 22527 13060 22583
rect 12632 22403 12688 22459
rect 12756 22403 12812 22459
rect 12880 22403 12936 22459
rect 13004 22403 13060 22459
rect 12632 22279 12688 22335
rect 12756 22279 12812 22335
rect 12880 22279 12936 22335
rect 13004 22279 13060 22335
rect 12632 22155 12688 22211
rect 12756 22155 12812 22211
rect 12880 22155 12936 22211
rect 13004 22155 13060 22211
rect 12632 22031 12688 22087
rect 12756 22031 12812 22087
rect 12880 22031 12936 22087
rect 13004 22031 13060 22087
rect 12632 21907 12688 21963
rect 12756 21907 12812 21963
rect 12880 21907 12936 21963
rect 13004 21907 13060 21963
rect 12632 21783 12688 21839
rect 12756 21783 12812 21839
rect 12880 21783 12936 21839
rect 13004 21783 13060 21839
rect 12632 21659 12688 21715
rect 12756 21659 12812 21715
rect 12880 21659 12936 21715
rect 13004 21659 13060 21715
rect 12632 21535 12688 21591
rect 12756 21535 12812 21591
rect 12880 21535 12936 21591
rect 13004 21535 13060 21591
rect 12632 21411 12688 21467
rect 12756 21411 12812 21467
rect 12880 21411 12936 21467
rect 13004 21411 13060 21467
rect 12632 21287 12688 21343
rect 12756 21287 12812 21343
rect 12880 21287 12936 21343
rect 13004 21287 13060 21343
rect 12632 21163 12688 21219
rect 12756 21163 12812 21219
rect 12880 21163 12936 21219
rect 13004 21163 13060 21219
rect 12632 21039 12688 21095
rect 12756 21039 12812 21095
rect 12880 21039 12936 21095
rect 13004 21039 13060 21095
rect 12632 20915 12688 20971
rect 12756 20915 12812 20971
rect 12880 20915 12936 20971
rect 13004 20915 13060 20971
rect 12632 20791 12688 20847
rect 12756 20791 12812 20847
rect 12880 20791 12936 20847
rect 13004 20791 13060 20847
rect 12632 20667 12688 20723
rect 12756 20667 12812 20723
rect 12880 20667 12936 20723
rect 13004 20667 13060 20723
rect 12632 20543 12688 20599
rect 12756 20543 12812 20599
rect 12880 20543 12936 20599
rect 13004 20543 13060 20599
rect 12632 20195 12688 20251
rect 12756 20195 12812 20251
rect 12880 20195 12936 20251
rect 13004 20195 13060 20251
rect 12632 20071 12688 20127
rect 12756 20071 12812 20127
rect 12880 20071 12936 20127
rect 13004 20071 13060 20127
rect 12632 19947 12688 20003
rect 12756 19947 12812 20003
rect 12880 19947 12936 20003
rect 13004 19947 13060 20003
rect 12632 19823 12688 19879
rect 12756 19823 12812 19879
rect 12880 19823 12936 19879
rect 13004 19823 13060 19879
rect 12632 19699 12688 19755
rect 12756 19699 12812 19755
rect 12880 19699 12936 19755
rect 13004 19699 13060 19755
rect 12632 19575 12688 19631
rect 12756 19575 12812 19631
rect 12880 19575 12936 19631
rect 13004 19575 13060 19631
rect 12632 19451 12688 19507
rect 12756 19451 12812 19507
rect 12880 19451 12936 19507
rect 13004 19451 13060 19507
rect 12632 19327 12688 19383
rect 12756 19327 12812 19383
rect 12880 19327 12936 19383
rect 13004 19327 13060 19383
rect 12632 19203 12688 19259
rect 12756 19203 12812 19259
rect 12880 19203 12936 19259
rect 13004 19203 13060 19259
rect 12632 19079 12688 19135
rect 12756 19079 12812 19135
rect 12880 19079 12936 19135
rect 13004 19079 13060 19135
rect 12632 18955 12688 19011
rect 12756 18955 12812 19011
rect 12880 18955 12936 19011
rect 13004 18955 13060 19011
rect 12632 18831 12688 18887
rect 12756 18831 12812 18887
rect 12880 18831 12936 18887
rect 13004 18831 13060 18887
rect 12632 18707 12688 18763
rect 12756 18707 12812 18763
rect 12880 18707 12936 18763
rect 13004 18707 13060 18763
rect 12632 18583 12688 18639
rect 12756 18583 12812 18639
rect 12880 18583 12936 18639
rect 13004 18583 13060 18639
rect 12632 18459 12688 18515
rect 12756 18459 12812 18515
rect 12880 18459 12936 18515
rect 13004 18459 13060 18515
rect 12632 18335 12688 18391
rect 12756 18335 12812 18391
rect 12880 18335 12936 18391
rect 13004 18335 13060 18391
rect 12632 18211 12688 18267
rect 12756 18211 12812 18267
rect 12880 18211 12936 18267
rect 13004 18211 13060 18267
rect 12632 18087 12688 18143
rect 12756 18087 12812 18143
rect 12880 18087 12936 18143
rect 13004 18087 13060 18143
rect 12632 17963 12688 18019
rect 12756 17963 12812 18019
rect 12880 17963 12936 18019
rect 13004 17963 13060 18019
rect 12632 17839 12688 17895
rect 12756 17839 12812 17895
rect 12880 17839 12936 17895
rect 13004 17839 13060 17895
rect 12632 17715 12688 17771
rect 12756 17715 12812 17771
rect 12880 17715 12936 17771
rect 13004 17715 13060 17771
rect 12632 17591 12688 17647
rect 12756 17591 12812 17647
rect 12880 17591 12936 17647
rect 13004 17591 13060 17647
rect 12632 17467 12688 17523
rect 12756 17467 12812 17523
rect 12880 17467 12936 17523
rect 13004 17467 13060 17523
rect 12632 17343 12688 17399
rect 12756 17343 12812 17399
rect 12880 17343 12936 17399
rect 13004 17343 13060 17399
rect 12632 16995 12688 17051
rect 12756 16995 12812 17051
rect 12880 16995 12936 17051
rect 13004 16995 13060 17051
rect 12632 16871 12688 16927
rect 12756 16871 12812 16927
rect 12880 16871 12936 16927
rect 13004 16871 13060 16927
rect 12632 16747 12688 16803
rect 12756 16747 12812 16803
rect 12880 16747 12936 16803
rect 13004 16747 13060 16803
rect 12632 16623 12688 16679
rect 12756 16623 12812 16679
rect 12880 16623 12936 16679
rect 13004 16623 13060 16679
rect 12632 16499 12688 16555
rect 12756 16499 12812 16555
rect 12880 16499 12936 16555
rect 13004 16499 13060 16555
rect 12632 16375 12688 16431
rect 12756 16375 12812 16431
rect 12880 16375 12936 16431
rect 13004 16375 13060 16431
rect 12632 16251 12688 16307
rect 12756 16251 12812 16307
rect 12880 16251 12936 16307
rect 13004 16251 13060 16307
rect 12632 16127 12688 16183
rect 12756 16127 12812 16183
rect 12880 16127 12936 16183
rect 13004 16127 13060 16183
rect 12632 16003 12688 16059
rect 12756 16003 12812 16059
rect 12880 16003 12936 16059
rect 13004 16003 13060 16059
rect 12632 15879 12688 15935
rect 12756 15879 12812 15935
rect 12880 15879 12936 15935
rect 13004 15879 13060 15935
rect 10928 15631 10984 15687
rect 11052 15631 11108 15687
rect 11176 15631 11232 15687
rect 11300 15631 11356 15687
rect 10928 15507 10984 15563
rect 11052 15507 11108 15563
rect 11176 15507 11232 15563
rect 11300 15507 11356 15563
rect 10928 15383 10984 15439
rect 11052 15383 11108 15439
rect 11176 15383 11232 15439
rect 11300 15383 11356 15439
rect 10928 15259 10984 15315
rect 11052 15259 11108 15315
rect 11176 15259 11232 15315
rect 11300 15259 11356 15315
rect 10928 15135 10984 15191
rect 11052 15135 11108 15191
rect 11176 15135 11232 15191
rect 11300 15135 11356 15191
rect 10928 15011 10984 15067
rect 11052 15011 11108 15067
rect 11176 15011 11232 15067
rect 11300 15011 11356 15067
rect 10928 14887 10984 14943
rect 11052 14887 11108 14943
rect 11176 14887 11232 14943
rect 11300 14887 11356 14943
rect 10928 14763 10984 14819
rect 11052 14763 11108 14819
rect 11176 14763 11232 14819
rect 11300 14763 11356 14819
rect 10928 14639 10984 14695
rect 11052 14639 11108 14695
rect 11176 14639 11232 14695
rect 11300 14639 11356 14695
rect 10928 14515 10984 14571
rect 11052 14515 11108 14571
rect 11176 14515 11232 14571
rect 11300 14515 11356 14571
rect 10928 14391 10984 14447
rect 11052 14391 11108 14447
rect 11176 14391 11232 14447
rect 11300 14391 11356 14447
rect 10928 14267 10984 14323
rect 11052 14267 11108 14323
rect 11176 14267 11232 14323
rect 11300 14267 11356 14323
rect 10928 14143 10984 14199
rect 11052 14143 11108 14199
rect 11176 14143 11232 14199
rect 11300 14143 11356 14199
rect 12632 15755 12688 15811
rect 12756 15755 12812 15811
rect 12880 15755 12936 15811
rect 13004 15755 13060 15811
rect 13200 36195 13256 36251
rect 13324 36195 13380 36251
rect 13448 36195 13504 36251
rect 13572 36195 13628 36251
rect 13200 36071 13256 36127
rect 13324 36071 13380 36127
rect 13448 36071 13504 36127
rect 13572 36071 13628 36127
rect 13200 35947 13256 36003
rect 13324 35947 13380 36003
rect 13448 35947 13504 36003
rect 13572 35947 13628 36003
rect 13200 35823 13256 35879
rect 13324 35823 13380 35879
rect 13448 35823 13504 35879
rect 13572 35823 13628 35879
rect 13200 35699 13256 35755
rect 13324 35699 13380 35755
rect 13448 35699 13504 35755
rect 13572 35699 13628 35755
rect 13200 35575 13256 35631
rect 13324 35575 13380 35631
rect 13448 35575 13504 35631
rect 13572 35575 13628 35631
rect 13200 35451 13256 35507
rect 13324 35451 13380 35507
rect 13448 35451 13504 35507
rect 13572 35451 13628 35507
rect 13200 35327 13256 35383
rect 13324 35327 13380 35383
rect 13448 35327 13504 35383
rect 13572 35327 13628 35383
rect 13200 35203 13256 35259
rect 13324 35203 13380 35259
rect 13448 35203 13504 35259
rect 13572 35203 13628 35259
rect 13200 35079 13256 35135
rect 13324 35079 13380 35135
rect 13448 35079 13504 35135
rect 13572 35079 13628 35135
rect 13200 34955 13256 35011
rect 13324 34955 13380 35011
rect 13448 34955 13504 35011
rect 13572 34955 13628 35011
rect 13200 34831 13256 34887
rect 13324 34831 13380 34887
rect 13448 34831 13504 34887
rect 13572 34831 13628 34887
rect 13200 34707 13256 34763
rect 13324 34707 13380 34763
rect 13448 34707 13504 34763
rect 13572 34707 13628 34763
rect 13200 34583 13256 34639
rect 13324 34583 13380 34639
rect 13448 34583 13504 34639
rect 13572 34583 13628 34639
rect 13200 34459 13256 34515
rect 13324 34459 13380 34515
rect 13448 34459 13504 34515
rect 13572 34459 13628 34515
rect 13200 34335 13256 34391
rect 13324 34335 13380 34391
rect 13448 34335 13504 34391
rect 13572 34335 13628 34391
rect 13200 34211 13256 34267
rect 13324 34211 13380 34267
rect 13448 34211 13504 34267
rect 13572 34211 13628 34267
rect 13200 34087 13256 34143
rect 13324 34087 13380 34143
rect 13448 34087 13504 34143
rect 13572 34087 13628 34143
rect 13200 33963 13256 34019
rect 13324 33963 13380 34019
rect 13448 33963 13504 34019
rect 13572 33963 13628 34019
rect 13200 33839 13256 33895
rect 13324 33839 13380 33895
rect 13448 33839 13504 33895
rect 13572 33839 13628 33895
rect 13200 33715 13256 33771
rect 13324 33715 13380 33771
rect 13448 33715 13504 33771
rect 13572 33715 13628 33771
rect 13200 33591 13256 33647
rect 13324 33591 13380 33647
rect 13448 33591 13504 33647
rect 13572 33591 13628 33647
rect 13200 33467 13256 33523
rect 13324 33467 13380 33523
rect 13448 33467 13504 33523
rect 13572 33467 13628 33523
rect 13200 33343 13256 33399
rect 13324 33343 13380 33399
rect 13448 33343 13504 33399
rect 13572 33343 13628 33399
rect 13200 28189 13256 28245
rect 13324 28189 13380 28245
rect 13448 28189 13504 28245
rect 13572 28189 13628 28245
rect 13200 28065 13256 28121
rect 13324 28065 13380 28121
rect 13448 28065 13504 28121
rect 13572 28065 13628 28121
rect 13200 27941 13256 27997
rect 13324 27941 13380 27997
rect 13448 27941 13504 27997
rect 13572 27941 13628 27997
rect 13200 27817 13256 27873
rect 13324 27817 13380 27873
rect 13448 27817 13504 27873
rect 13572 27817 13628 27873
rect 13200 27693 13256 27749
rect 13324 27693 13380 27749
rect 13448 27693 13504 27749
rect 13572 27693 13628 27749
rect 13200 27569 13256 27625
rect 13324 27569 13380 27625
rect 13448 27569 13504 27625
rect 13572 27569 13628 27625
rect 13200 27445 13256 27501
rect 13324 27445 13380 27501
rect 13448 27445 13504 27501
rect 13572 27445 13628 27501
rect 13200 27321 13256 27377
rect 13324 27321 13380 27377
rect 13448 27321 13504 27377
rect 13572 27321 13628 27377
rect 13200 27197 13256 27253
rect 13324 27197 13380 27253
rect 13448 27197 13504 27253
rect 13572 27197 13628 27253
rect 13200 27073 13256 27129
rect 13324 27073 13380 27129
rect 13448 27073 13504 27129
rect 13572 27073 13628 27129
rect 13200 26949 13256 27005
rect 13324 26949 13380 27005
rect 13448 26949 13504 27005
rect 13572 26949 13628 27005
rect 13768 55404 13786 55445
rect 13786 55404 13824 55445
rect 13892 55404 13910 55445
rect 13910 55404 13948 55445
rect 14016 55404 14034 55445
rect 14034 55404 14072 55445
rect 13768 55389 13824 55404
rect 13892 55389 13948 55404
rect 14016 55389 14072 55404
rect 14140 55389 14196 55445
rect 13768 55280 13786 55321
rect 13786 55280 13824 55321
rect 13892 55280 13910 55321
rect 13910 55280 13948 55321
rect 14016 55280 14034 55321
rect 14034 55280 14072 55321
rect 13768 55265 13824 55280
rect 13892 55265 13948 55280
rect 14016 55265 14072 55280
rect 14140 55265 14196 55321
rect 13768 55156 13786 55197
rect 13786 55156 13824 55197
rect 13892 55156 13910 55197
rect 13910 55156 13948 55197
rect 14016 55156 14034 55197
rect 14034 55156 14072 55197
rect 13768 55141 13824 55156
rect 13892 55141 13948 55156
rect 14016 55141 14072 55156
rect 14140 55141 14196 55197
rect 13768 55032 13786 55073
rect 13786 55032 13824 55073
rect 13892 55032 13910 55073
rect 13910 55032 13948 55073
rect 14016 55032 14034 55073
rect 14034 55032 14072 55073
rect 13768 55017 13824 55032
rect 13892 55017 13948 55032
rect 14016 55017 14072 55032
rect 14140 55017 14196 55073
rect 13768 54908 13786 54949
rect 13786 54908 13824 54949
rect 13892 54908 13910 54949
rect 13910 54908 13948 54949
rect 14016 54908 14034 54949
rect 14034 54908 14072 54949
rect 13768 54893 13824 54908
rect 13892 54893 13948 54908
rect 14016 54893 14072 54908
rect 14140 54893 14196 54949
rect 13768 54784 13786 54825
rect 13786 54784 13824 54825
rect 13892 54784 13910 54825
rect 13910 54784 13948 54825
rect 14016 54784 14034 54825
rect 14034 54784 14072 54825
rect 13768 54769 13824 54784
rect 13892 54769 13948 54784
rect 14016 54769 14072 54784
rect 14140 54769 14196 54825
rect 13768 54660 13786 54701
rect 13786 54660 13824 54701
rect 13892 54660 13910 54701
rect 13910 54660 13948 54701
rect 14016 54660 14034 54701
rect 14034 54660 14072 54701
rect 13768 54645 13824 54660
rect 13892 54645 13948 54660
rect 14016 54645 14072 54660
rect 14140 54645 14196 54701
rect 13768 54536 13786 54577
rect 13786 54536 13824 54577
rect 13892 54536 13910 54577
rect 13910 54536 13948 54577
rect 14016 54536 14034 54577
rect 14034 54536 14072 54577
rect 13768 54521 13824 54536
rect 13892 54521 13948 54536
rect 14016 54521 14072 54536
rect 14140 54521 14196 54577
rect 13768 54412 13786 54453
rect 13786 54412 13824 54453
rect 13892 54412 13910 54453
rect 13910 54412 13948 54453
rect 14016 54412 14034 54453
rect 14034 54412 14072 54453
rect 13768 54397 13824 54412
rect 13892 54397 13948 54412
rect 14016 54397 14072 54412
rect 14140 54397 14196 54453
rect 13768 54288 13786 54329
rect 13786 54288 13824 54329
rect 13892 54288 13910 54329
rect 13910 54288 13948 54329
rect 14016 54288 14034 54329
rect 14034 54288 14072 54329
rect 13768 54273 13824 54288
rect 13892 54273 13948 54288
rect 14016 54273 14072 54288
rect 14140 54273 14196 54329
rect 13768 54164 13786 54205
rect 13786 54164 13824 54205
rect 13892 54164 13910 54205
rect 13910 54164 13948 54205
rect 14016 54164 14034 54205
rect 14034 54164 14072 54205
rect 13768 54149 13824 54164
rect 13892 54149 13948 54164
rect 14016 54149 14072 54164
rect 14140 54149 14196 54205
rect 13768 47436 13824 47445
rect 13892 47436 13948 47445
rect 14016 47436 14072 47445
rect 13768 47389 13786 47436
rect 13786 47389 13824 47436
rect 13892 47389 13910 47436
rect 13910 47389 13948 47436
rect 14016 47389 14034 47436
rect 14034 47389 14072 47436
rect 14140 47389 14196 47445
rect 13768 47312 13824 47321
rect 13892 47312 13948 47321
rect 14016 47312 14072 47321
rect 13768 47265 13786 47312
rect 13786 47265 13824 47312
rect 13892 47265 13910 47312
rect 13910 47265 13948 47312
rect 14016 47265 14034 47312
rect 14034 47265 14072 47312
rect 14140 47265 14196 47321
rect 13768 47188 13824 47197
rect 13892 47188 13948 47197
rect 14016 47188 14072 47197
rect 13768 47141 13786 47188
rect 13786 47141 13824 47188
rect 13892 47141 13910 47188
rect 13910 47141 13948 47188
rect 14016 47141 14034 47188
rect 14034 47141 14072 47188
rect 14140 47141 14196 47197
rect 13768 47064 13824 47073
rect 13892 47064 13948 47073
rect 14016 47064 14072 47073
rect 13768 47017 13786 47064
rect 13786 47017 13824 47064
rect 13892 47017 13910 47064
rect 13910 47017 13948 47064
rect 14016 47017 14034 47064
rect 14034 47017 14072 47064
rect 14140 47017 14196 47073
rect 13768 46940 13824 46949
rect 13892 46940 13948 46949
rect 14016 46940 14072 46949
rect 13768 46893 13786 46940
rect 13786 46893 13824 46940
rect 13892 46893 13910 46940
rect 13910 46893 13948 46940
rect 14016 46893 14034 46940
rect 14034 46893 14072 46940
rect 14140 46893 14196 46949
rect 13768 46816 13824 46825
rect 13892 46816 13948 46825
rect 14016 46816 14072 46825
rect 13768 46769 13786 46816
rect 13786 46769 13824 46816
rect 13892 46769 13910 46816
rect 13910 46769 13948 46816
rect 14016 46769 14034 46816
rect 14034 46769 14072 46816
rect 14140 46769 14196 46825
rect 13768 46692 13824 46701
rect 13892 46692 13948 46701
rect 14016 46692 14072 46701
rect 13768 46645 13786 46692
rect 13786 46645 13824 46692
rect 13892 46645 13910 46692
rect 13910 46645 13948 46692
rect 14016 46645 14034 46692
rect 14034 46645 14072 46692
rect 14140 46645 14196 46701
rect 13768 46568 13824 46577
rect 13892 46568 13948 46577
rect 14016 46568 14072 46577
rect 13768 46521 13786 46568
rect 13786 46521 13824 46568
rect 13892 46521 13910 46568
rect 13910 46521 13948 46568
rect 14016 46521 14034 46568
rect 14034 46521 14072 46568
rect 14140 46521 14196 46577
rect 13768 46444 13824 46453
rect 13892 46444 13948 46453
rect 14016 46444 14072 46453
rect 13768 46397 13786 46444
rect 13786 46397 13824 46444
rect 13892 46397 13910 46444
rect 13910 46397 13948 46444
rect 14016 46397 14034 46444
rect 14034 46397 14072 46444
rect 14140 46397 14196 46453
rect 13768 46320 13824 46329
rect 13892 46320 13948 46329
rect 14016 46320 14072 46329
rect 13768 46273 13786 46320
rect 13786 46273 13824 46320
rect 13892 46273 13910 46320
rect 13910 46273 13948 46320
rect 14016 46273 14034 46320
rect 14034 46273 14072 46320
rect 14140 46273 14196 46329
rect 13768 46196 13824 46205
rect 13892 46196 13948 46205
rect 14016 46196 14072 46205
rect 13768 46149 13786 46196
rect 13786 46149 13824 46196
rect 13892 46149 13910 46196
rect 13910 46149 13948 46196
rect 14016 46149 14034 46196
rect 14034 46149 14072 46196
rect 14140 46149 14196 46205
rect 13768 44232 13824 44245
rect 13892 44232 13948 44245
rect 14016 44232 14072 44245
rect 13768 44189 13786 44232
rect 13786 44189 13824 44232
rect 13892 44189 13910 44232
rect 13910 44189 13948 44232
rect 14016 44189 14034 44232
rect 14034 44189 14072 44232
rect 14140 44189 14196 44245
rect 13768 44108 13824 44121
rect 13892 44108 13948 44121
rect 14016 44108 14072 44121
rect 13768 44065 13786 44108
rect 13786 44065 13824 44108
rect 13892 44065 13910 44108
rect 13910 44065 13948 44108
rect 14016 44065 14034 44108
rect 14034 44065 14072 44108
rect 14140 44065 14196 44121
rect 13768 43984 13824 43997
rect 13892 43984 13948 43997
rect 14016 43984 14072 43997
rect 13768 43941 13786 43984
rect 13786 43941 13824 43984
rect 13892 43941 13910 43984
rect 13910 43941 13948 43984
rect 14016 43941 14034 43984
rect 14034 43941 14072 43984
rect 14140 43941 14196 43997
rect 13768 43860 13824 43873
rect 13892 43860 13948 43873
rect 14016 43860 14072 43873
rect 13768 43817 13786 43860
rect 13786 43817 13824 43860
rect 13892 43817 13910 43860
rect 13910 43817 13948 43860
rect 14016 43817 14034 43860
rect 14034 43817 14072 43860
rect 14140 43817 14196 43873
rect 13768 43736 13824 43749
rect 13892 43736 13948 43749
rect 14016 43736 14072 43749
rect 13768 43693 13786 43736
rect 13786 43693 13824 43736
rect 13892 43693 13910 43736
rect 13910 43693 13948 43736
rect 14016 43693 14034 43736
rect 14034 43693 14072 43736
rect 14140 43693 14196 43749
rect 13768 43612 13824 43625
rect 13892 43612 13948 43625
rect 14016 43612 14072 43625
rect 13768 43569 13786 43612
rect 13786 43569 13824 43612
rect 13892 43569 13910 43612
rect 13910 43569 13948 43612
rect 14016 43569 14034 43612
rect 14034 43569 14072 43612
rect 14140 43569 14196 43625
rect 13768 43488 13824 43501
rect 13892 43488 13948 43501
rect 14016 43488 14072 43501
rect 13768 43445 13786 43488
rect 13786 43445 13824 43488
rect 13892 43445 13910 43488
rect 13910 43445 13948 43488
rect 14016 43445 14034 43488
rect 14034 43445 14072 43488
rect 14140 43445 14196 43501
rect 13768 43364 13824 43377
rect 13892 43364 13948 43377
rect 14016 43364 14072 43377
rect 13768 43321 13786 43364
rect 13786 43321 13824 43364
rect 13892 43321 13910 43364
rect 13910 43321 13948 43364
rect 14016 43321 14034 43364
rect 14034 43321 14072 43364
rect 14140 43321 14196 43377
rect 13768 43240 13824 43253
rect 13892 43240 13948 43253
rect 14016 43240 14072 43253
rect 13768 43197 13786 43240
rect 13786 43197 13824 43240
rect 13892 43197 13910 43240
rect 13910 43197 13948 43240
rect 14016 43197 14034 43240
rect 14034 43197 14072 43240
rect 14140 43197 14196 43253
rect 13768 43116 13824 43129
rect 13892 43116 13948 43129
rect 14016 43116 14072 43129
rect 13768 43073 13786 43116
rect 13786 43073 13824 43116
rect 13892 43073 13910 43116
rect 13910 43073 13948 43116
rect 14016 43073 14034 43116
rect 14034 43073 14072 43116
rect 14140 43073 14196 43129
rect 13768 42992 13824 43005
rect 13892 42992 13948 43005
rect 14016 42992 14072 43005
rect 13768 42949 13786 42992
rect 13786 42949 13824 42992
rect 13892 42949 13910 42992
rect 13910 42949 13948 42992
rect 14016 42949 14034 42992
rect 14034 42949 14072 42992
rect 14140 42949 14196 43005
rect 13768 42620 13824 42645
rect 13892 42620 13948 42645
rect 14016 42620 14072 42645
rect 13768 42589 13786 42620
rect 13786 42589 13824 42620
rect 13892 42589 13910 42620
rect 13910 42589 13948 42620
rect 14016 42589 14034 42620
rect 14034 42589 14072 42620
rect 14140 42589 14196 42645
rect 13768 42496 13824 42521
rect 13892 42496 13948 42521
rect 14016 42496 14072 42521
rect 13768 42465 13786 42496
rect 13786 42465 13824 42496
rect 13892 42465 13910 42496
rect 13910 42465 13948 42496
rect 14016 42465 14034 42496
rect 14034 42465 14072 42496
rect 14140 42465 14196 42521
rect 13768 42372 13824 42397
rect 13892 42372 13948 42397
rect 14016 42372 14072 42397
rect 13768 42341 13786 42372
rect 13786 42341 13824 42372
rect 13892 42341 13910 42372
rect 13910 42341 13948 42372
rect 14016 42341 14034 42372
rect 14034 42341 14072 42372
rect 14140 42341 14196 42397
rect 13768 42248 13824 42273
rect 13892 42248 13948 42273
rect 14016 42248 14072 42273
rect 13768 42217 13786 42248
rect 13786 42217 13824 42248
rect 13892 42217 13910 42248
rect 13910 42217 13948 42248
rect 14016 42217 14034 42248
rect 14034 42217 14072 42248
rect 14140 42217 14196 42273
rect 13768 42124 13824 42149
rect 13892 42124 13948 42149
rect 14016 42124 14072 42149
rect 13768 42093 13786 42124
rect 13786 42093 13824 42124
rect 13892 42093 13910 42124
rect 13910 42093 13948 42124
rect 14016 42093 14034 42124
rect 14034 42093 14072 42124
rect 14140 42093 14196 42149
rect 13768 42000 13824 42025
rect 13892 42000 13948 42025
rect 14016 42000 14072 42025
rect 13768 41969 13786 42000
rect 13786 41969 13824 42000
rect 13892 41969 13910 42000
rect 13910 41969 13948 42000
rect 14016 41969 14034 42000
rect 14034 41969 14072 42000
rect 14140 41969 14196 42025
rect 13768 41876 13824 41901
rect 13892 41876 13948 41901
rect 14016 41876 14072 41901
rect 13768 41845 13786 41876
rect 13786 41845 13824 41876
rect 13892 41845 13910 41876
rect 13910 41845 13948 41876
rect 14016 41845 14034 41876
rect 14034 41845 14072 41876
rect 14140 41845 14196 41901
rect 13768 41752 13824 41777
rect 13892 41752 13948 41777
rect 14016 41752 14072 41777
rect 13768 41721 13786 41752
rect 13786 41721 13824 41752
rect 13892 41721 13910 41752
rect 13910 41721 13948 41752
rect 14016 41721 14034 41752
rect 14034 41721 14072 41752
rect 14140 41721 14196 41777
rect 13768 41628 13824 41653
rect 13892 41628 13948 41653
rect 14016 41628 14072 41653
rect 13768 41597 13786 41628
rect 13786 41597 13824 41628
rect 13892 41597 13910 41628
rect 13910 41597 13948 41628
rect 14016 41597 14034 41628
rect 14034 41597 14072 41628
rect 14140 41597 14196 41653
rect 13768 41504 13824 41529
rect 13892 41504 13948 41529
rect 14016 41504 14072 41529
rect 13768 41473 13786 41504
rect 13786 41473 13824 41504
rect 13892 41473 13910 41504
rect 13910 41473 13948 41504
rect 14016 41473 14034 41504
rect 14034 41473 14072 41504
rect 14140 41473 14196 41529
rect 13768 41380 13824 41405
rect 13892 41380 13948 41405
rect 14016 41380 14072 41405
rect 13768 41349 13786 41380
rect 13786 41349 13824 41380
rect 13892 41349 13910 41380
rect 13910 41349 13948 41380
rect 14016 41349 14034 41380
rect 14034 41349 14072 41380
rect 14140 41349 14196 41405
rect 13768 40989 13824 41045
rect 13892 40989 13948 41045
rect 14016 40989 14072 41045
rect 14140 40989 14196 41045
rect 13768 40865 13824 40921
rect 13892 40865 13948 40921
rect 14016 40865 14072 40921
rect 14140 40865 14196 40921
rect 13768 40741 13824 40797
rect 13892 40741 13948 40797
rect 14016 40741 14072 40797
rect 14140 40741 14196 40797
rect 13768 40617 13824 40673
rect 13892 40617 13948 40673
rect 14016 40617 14072 40673
rect 14140 40617 14196 40673
rect 13768 40532 13824 40549
rect 13892 40532 13948 40549
rect 14016 40532 14072 40549
rect 13768 40493 13786 40532
rect 13786 40493 13824 40532
rect 13892 40493 13910 40532
rect 13910 40493 13948 40532
rect 14016 40493 14034 40532
rect 14034 40493 14072 40532
rect 14140 40493 14196 40549
rect 13768 40408 13824 40425
rect 13892 40408 13948 40425
rect 14016 40408 14072 40425
rect 13768 40369 13786 40408
rect 13786 40369 13824 40408
rect 13892 40369 13910 40408
rect 13910 40369 13948 40408
rect 14016 40369 14034 40408
rect 14034 40369 14072 40408
rect 14140 40369 14196 40425
rect 13768 40284 13824 40301
rect 13892 40284 13948 40301
rect 14016 40284 14072 40301
rect 13768 40245 13786 40284
rect 13786 40245 13824 40284
rect 13892 40245 13910 40284
rect 13910 40245 13948 40284
rect 14016 40245 14034 40284
rect 14034 40245 14072 40284
rect 14140 40245 14196 40301
rect 13768 40160 13824 40177
rect 13892 40160 13948 40177
rect 14016 40160 14072 40177
rect 13768 40121 13786 40160
rect 13786 40121 13824 40160
rect 13892 40121 13910 40160
rect 13910 40121 13948 40160
rect 14016 40121 14034 40160
rect 14034 40121 14072 40160
rect 14140 40121 14196 40177
rect 13768 40036 13824 40053
rect 13892 40036 13948 40053
rect 14016 40036 14072 40053
rect 13768 39997 13786 40036
rect 13786 39997 13824 40036
rect 13892 39997 13910 40036
rect 13910 39997 13948 40036
rect 14016 39997 14034 40036
rect 14034 39997 14072 40036
rect 14140 39997 14196 40053
rect 13768 39912 13824 39929
rect 13892 39912 13948 39929
rect 14016 39912 14072 39929
rect 13768 39873 13786 39912
rect 13786 39873 13824 39912
rect 13892 39873 13910 39912
rect 13910 39873 13948 39912
rect 14016 39873 14034 39912
rect 14034 39873 14072 39912
rect 14140 39873 14196 39929
rect 13768 39788 13824 39805
rect 13892 39788 13948 39805
rect 14016 39788 14072 39805
rect 13768 39749 13786 39788
rect 13786 39749 13824 39788
rect 13892 39749 13910 39788
rect 13910 39749 13948 39788
rect 14016 39749 14034 39788
rect 14034 39749 14072 39788
rect 14140 39749 14196 39805
rect 13768 32995 13824 33051
rect 13892 32995 13948 33051
rect 14016 32995 14072 33051
rect 14140 32995 14196 33051
rect 13768 32871 13824 32927
rect 13892 32871 13948 32927
rect 14016 32871 14072 32927
rect 14140 32871 14196 32927
rect 13768 32747 13824 32803
rect 13892 32747 13948 32803
rect 14016 32747 14072 32803
rect 14140 32747 14196 32803
rect 13768 32636 13824 32679
rect 13892 32636 13948 32679
rect 14016 32636 14072 32679
rect 13768 32623 13786 32636
rect 13786 32623 13824 32636
rect 13892 32623 13910 32636
rect 13910 32623 13948 32636
rect 14016 32623 14034 32636
rect 14034 32623 14072 32636
rect 14140 32623 14196 32679
rect 13768 32512 13824 32555
rect 13892 32512 13948 32555
rect 14016 32512 14072 32555
rect 13768 32499 13786 32512
rect 13786 32499 13824 32512
rect 13892 32499 13910 32512
rect 13910 32499 13948 32512
rect 14016 32499 14034 32512
rect 14034 32499 14072 32512
rect 14140 32499 14196 32555
rect 13768 32388 13824 32431
rect 13892 32388 13948 32431
rect 14016 32388 14072 32431
rect 13768 32375 13786 32388
rect 13786 32375 13824 32388
rect 13892 32375 13910 32388
rect 13910 32375 13948 32388
rect 14016 32375 14034 32388
rect 14034 32375 14072 32388
rect 14140 32375 14196 32431
rect 13768 32264 13824 32307
rect 13892 32264 13948 32307
rect 14016 32264 14072 32307
rect 13768 32251 13786 32264
rect 13786 32251 13824 32264
rect 13892 32251 13910 32264
rect 13910 32251 13948 32264
rect 14016 32251 14034 32264
rect 14034 32251 14072 32264
rect 14140 32251 14196 32307
rect 13768 32140 13824 32183
rect 13892 32140 13948 32183
rect 14016 32140 14072 32183
rect 13768 32127 13786 32140
rect 13786 32127 13824 32140
rect 13892 32127 13910 32140
rect 13910 32127 13948 32140
rect 14016 32127 14034 32140
rect 14034 32127 14072 32140
rect 14140 32127 14196 32183
rect 13768 32016 13824 32059
rect 13892 32016 13948 32059
rect 14016 32016 14072 32059
rect 13768 32003 13786 32016
rect 13786 32003 13824 32016
rect 13892 32003 13910 32016
rect 13910 32003 13948 32016
rect 14016 32003 14034 32016
rect 14034 32003 14072 32016
rect 14140 32003 14196 32059
rect 13768 31892 13824 31935
rect 13892 31892 13948 31935
rect 14016 31892 14072 31935
rect 13768 31879 13786 31892
rect 13786 31879 13824 31892
rect 13892 31879 13910 31892
rect 13910 31879 13948 31892
rect 14016 31879 14034 31892
rect 14034 31879 14072 31892
rect 14140 31879 14196 31935
rect 13768 31768 13824 31811
rect 13892 31768 13948 31811
rect 14016 31768 14072 31811
rect 13768 31755 13786 31768
rect 13786 31755 13824 31768
rect 13892 31755 13910 31768
rect 13910 31755 13948 31768
rect 14016 31755 14034 31768
rect 14034 31755 14072 31768
rect 14140 31755 14196 31811
rect 13768 31644 13824 31687
rect 13892 31644 13948 31687
rect 14016 31644 14072 31687
rect 13768 31631 13786 31644
rect 13786 31631 13824 31644
rect 13892 31631 13910 31644
rect 13910 31631 13948 31644
rect 14016 31631 14034 31644
rect 14034 31631 14072 31644
rect 14140 31631 14196 31687
rect 13768 31520 13824 31563
rect 13892 31520 13948 31563
rect 14016 31520 14072 31563
rect 13768 31507 13786 31520
rect 13786 31507 13824 31520
rect 13892 31507 13910 31520
rect 13910 31507 13948 31520
rect 14016 31507 14034 31520
rect 14034 31507 14072 31520
rect 14140 31507 14196 31563
rect 13768 31396 13824 31439
rect 13892 31396 13948 31439
rect 14016 31396 14072 31439
rect 13768 31383 13786 31396
rect 13786 31383 13824 31396
rect 13892 31383 13910 31396
rect 13910 31383 13948 31396
rect 14016 31383 14034 31396
rect 14034 31383 14072 31396
rect 14140 31383 14196 31439
rect 13768 31272 13824 31315
rect 13892 31272 13948 31315
rect 14016 31272 14072 31315
rect 13768 31259 13786 31272
rect 13786 31259 13824 31272
rect 13892 31259 13910 31272
rect 13910 31259 13948 31272
rect 14016 31259 14034 31272
rect 14034 31259 14072 31272
rect 14140 31259 14196 31315
rect 13768 31148 13824 31191
rect 13892 31148 13948 31191
rect 14016 31148 14072 31191
rect 13768 31135 13786 31148
rect 13786 31135 13824 31148
rect 13892 31135 13910 31148
rect 13910 31135 13948 31148
rect 14016 31135 14034 31148
rect 14034 31135 14072 31148
rect 14140 31135 14196 31191
rect 13768 31024 13824 31067
rect 13892 31024 13948 31067
rect 14016 31024 14072 31067
rect 13768 31011 13786 31024
rect 13786 31011 13824 31024
rect 13892 31011 13910 31024
rect 13910 31011 13948 31024
rect 14016 31011 14034 31024
rect 14034 31011 14072 31024
rect 14140 31011 14196 31067
rect 13768 30900 13824 30943
rect 13892 30900 13948 30943
rect 14016 30900 14072 30943
rect 13768 30887 13786 30900
rect 13786 30887 13824 30900
rect 13892 30887 13910 30900
rect 13910 30887 13948 30900
rect 14016 30887 14034 30900
rect 14034 30887 14072 30900
rect 14140 30887 14196 30943
rect 13768 30776 13824 30819
rect 13892 30776 13948 30819
rect 14016 30776 14072 30819
rect 13768 30763 13786 30776
rect 13786 30763 13824 30776
rect 13892 30763 13910 30776
rect 13910 30763 13948 30776
rect 14016 30763 14034 30776
rect 14034 30763 14072 30776
rect 14140 30763 14196 30819
rect 13768 30652 13824 30695
rect 13892 30652 13948 30695
rect 14016 30652 14072 30695
rect 13768 30639 13786 30652
rect 13786 30639 13824 30652
rect 13892 30639 13910 30652
rect 13910 30639 13948 30652
rect 14016 30639 14034 30652
rect 14034 30639 14072 30652
rect 14140 30639 14196 30695
rect 13768 30528 13824 30571
rect 13892 30528 13948 30571
rect 14016 30528 14072 30571
rect 13768 30515 13786 30528
rect 13786 30515 13824 30528
rect 13892 30515 13910 30528
rect 13910 30515 13948 30528
rect 14016 30515 14034 30528
rect 14034 30515 14072 30528
rect 14140 30515 14196 30571
rect 13768 30404 13824 30447
rect 13892 30404 13948 30447
rect 14016 30404 14072 30447
rect 13768 30391 13786 30404
rect 13786 30391 13824 30404
rect 13892 30391 13910 30404
rect 13910 30391 13948 30404
rect 14016 30391 14034 30404
rect 14034 30391 14072 30404
rect 14140 30391 14196 30447
rect 13768 30280 13824 30323
rect 13892 30280 13948 30323
rect 14016 30280 14072 30323
rect 13768 30267 13786 30280
rect 13786 30267 13824 30280
rect 13892 30267 13910 30280
rect 13910 30267 13948 30280
rect 14016 30267 14034 30280
rect 14034 30267 14072 30280
rect 14140 30267 14196 30323
rect 13768 30156 13824 30199
rect 13892 30156 13948 30199
rect 14016 30156 14072 30199
rect 13768 30143 13786 30156
rect 13786 30143 13824 30156
rect 13892 30143 13910 30156
rect 13910 30143 13948 30156
rect 14016 30143 14034 30156
rect 14034 30143 14072 30156
rect 14140 30143 14196 30199
rect 13768 29789 13824 29845
rect 13892 29789 13948 29845
rect 14016 29789 14072 29845
rect 14140 29789 14196 29845
rect 13768 29665 13824 29721
rect 13892 29665 13948 29721
rect 14016 29665 14072 29721
rect 14140 29665 14196 29721
rect 13768 29541 13824 29597
rect 13892 29541 13948 29597
rect 14016 29541 14072 29597
rect 14140 29541 14196 29597
rect 13768 29417 13824 29473
rect 13892 29417 13948 29473
rect 14016 29417 14072 29473
rect 14140 29417 14196 29473
rect 13768 29293 13824 29349
rect 13892 29293 13948 29349
rect 14016 29293 14072 29349
rect 14140 29293 14196 29349
rect 13768 29169 13824 29225
rect 13892 29169 13948 29225
rect 14016 29169 14072 29225
rect 14140 29169 14196 29225
rect 13768 29045 13824 29101
rect 13892 29045 13948 29101
rect 14016 29045 14072 29101
rect 14140 29045 14196 29101
rect 13768 28921 13824 28977
rect 13892 28921 13948 28977
rect 14016 28921 14072 28977
rect 14140 28921 14196 28977
rect 13768 28797 13824 28853
rect 13892 28797 13948 28853
rect 14016 28797 14072 28853
rect 14140 28797 14196 28853
rect 13768 28688 13824 28729
rect 13892 28688 13948 28729
rect 14016 28688 14072 28729
rect 13768 28673 13786 28688
rect 13786 28673 13824 28688
rect 13892 28673 13910 28688
rect 13910 28673 13948 28688
rect 14016 28673 14034 28688
rect 14034 28673 14072 28688
rect 14140 28673 14196 28729
rect 13768 28564 13824 28605
rect 13892 28564 13948 28605
rect 14016 28564 14072 28605
rect 13768 28549 13786 28564
rect 13786 28549 13824 28564
rect 13892 28549 13910 28564
rect 13910 28549 13948 28564
rect 14016 28549 14034 28564
rect 14034 28549 14072 28564
rect 14140 28549 14196 28605
rect 13768 26595 13824 26651
rect 13892 26595 13948 26651
rect 14016 26595 14072 26651
rect 14140 26595 14196 26651
rect 13768 26471 13824 26527
rect 13892 26471 13948 26527
rect 14016 26471 14072 26527
rect 14140 26471 14196 26527
rect 13768 26347 13824 26403
rect 13892 26347 13948 26403
rect 14016 26347 14072 26403
rect 14140 26347 14196 26403
rect 13768 26223 13824 26279
rect 13892 26223 13948 26279
rect 14016 26223 14072 26279
rect 14140 26223 14196 26279
rect 13768 26099 13824 26155
rect 13892 26099 13948 26155
rect 14016 26099 14072 26155
rect 14140 26099 14196 26155
rect 13768 25975 13824 26031
rect 13892 25975 13948 26031
rect 14016 25975 14072 26031
rect 14140 25975 14196 26031
rect 13768 25851 13824 25907
rect 13892 25851 13948 25907
rect 14016 25851 14072 25907
rect 14140 25851 14196 25907
rect 13768 25727 13824 25783
rect 13892 25727 13948 25783
rect 14016 25727 14072 25783
rect 14140 25727 14196 25783
rect 13768 25603 13824 25659
rect 13892 25603 13948 25659
rect 14016 25603 14072 25659
rect 14140 25603 14196 25659
rect 13768 25479 13824 25535
rect 13892 25479 13948 25535
rect 14016 25479 14072 25535
rect 14140 25479 14196 25535
rect 13768 25355 13824 25411
rect 13892 25355 13948 25411
rect 14016 25355 14072 25411
rect 14140 25355 14196 25411
rect 13768 25231 13824 25287
rect 13892 25231 13948 25287
rect 14016 25231 14072 25287
rect 14140 25231 14196 25287
rect 13768 25107 13824 25163
rect 13892 25107 13948 25163
rect 14016 25107 14072 25163
rect 14140 25107 14196 25163
rect 13768 24983 13824 25039
rect 13892 24983 13948 25039
rect 14016 24983 14072 25039
rect 14140 24983 14196 25039
rect 13768 24859 13824 24915
rect 13892 24859 13948 24915
rect 14016 24859 14072 24915
rect 14140 24859 14196 24915
rect 13768 24740 13824 24791
rect 13892 24740 13948 24791
rect 14016 24740 14072 24791
rect 13768 24735 13786 24740
rect 13786 24735 13824 24740
rect 13892 24735 13910 24740
rect 13910 24735 13948 24740
rect 14016 24735 14034 24740
rect 14034 24735 14072 24740
rect 14140 24735 14196 24791
rect 13768 24616 13824 24667
rect 13892 24616 13948 24667
rect 14016 24616 14072 24667
rect 13768 24611 13786 24616
rect 13786 24611 13824 24616
rect 13892 24611 13910 24616
rect 13910 24611 13948 24616
rect 14016 24611 14034 24616
rect 14034 24611 14072 24616
rect 14140 24611 14196 24667
rect 13768 24492 13824 24543
rect 13892 24492 13948 24543
rect 14016 24492 14072 24543
rect 13768 24487 13786 24492
rect 13786 24487 13824 24492
rect 13892 24487 13910 24492
rect 13910 24487 13948 24492
rect 14016 24487 14034 24492
rect 14034 24487 14072 24492
rect 14140 24487 14196 24543
rect 13768 24368 13824 24419
rect 13892 24368 13948 24419
rect 14016 24368 14072 24419
rect 13768 24363 13786 24368
rect 13786 24363 13824 24368
rect 13892 24363 13910 24368
rect 13910 24363 13948 24368
rect 14016 24363 14034 24368
rect 14034 24363 14072 24368
rect 14140 24363 14196 24419
rect 13768 24244 13824 24295
rect 13892 24244 13948 24295
rect 14016 24244 14072 24295
rect 13768 24239 13786 24244
rect 13786 24239 13824 24244
rect 13892 24239 13910 24244
rect 13910 24239 13948 24244
rect 14016 24239 14034 24244
rect 14034 24239 14072 24244
rect 14140 24239 14196 24295
rect 13768 24120 13824 24171
rect 13892 24120 13948 24171
rect 14016 24120 14072 24171
rect 13768 24115 13786 24120
rect 13786 24115 13824 24120
rect 13892 24115 13910 24120
rect 13910 24115 13948 24120
rect 14016 24115 14034 24120
rect 14034 24115 14072 24120
rect 14140 24115 14196 24171
rect 13768 23996 13824 24047
rect 13892 23996 13948 24047
rect 14016 23996 14072 24047
rect 13768 23991 13786 23996
rect 13786 23991 13824 23996
rect 13892 23991 13910 23996
rect 13910 23991 13948 23996
rect 14016 23991 14034 23996
rect 14034 23991 14072 23996
rect 14140 23991 14196 24047
rect 13768 23872 13824 23923
rect 13892 23872 13948 23923
rect 14016 23872 14072 23923
rect 13768 23867 13786 23872
rect 13786 23867 13824 23872
rect 13892 23867 13910 23872
rect 13910 23867 13948 23872
rect 14016 23867 14034 23872
rect 14034 23867 14072 23872
rect 14140 23867 14196 23923
rect 13768 23748 13824 23799
rect 13892 23748 13948 23799
rect 14016 23748 14072 23799
rect 13768 23743 13786 23748
rect 13786 23743 13824 23748
rect 13892 23743 13910 23748
rect 13910 23743 13948 23748
rect 14016 23743 14034 23748
rect 14034 23743 14072 23748
rect 14140 23743 14196 23799
rect 13768 23448 13786 23451
rect 13786 23448 13824 23451
rect 13892 23448 13910 23451
rect 13910 23448 13948 23451
rect 14016 23448 14034 23451
rect 14034 23448 14072 23451
rect 13768 23395 13824 23448
rect 13892 23395 13948 23448
rect 14016 23395 14072 23448
rect 14140 23395 14196 23451
rect 13768 23324 13786 23327
rect 13786 23324 13824 23327
rect 13892 23324 13910 23327
rect 13910 23324 13948 23327
rect 14016 23324 14034 23327
rect 14034 23324 14072 23327
rect 13768 23271 13824 23324
rect 13892 23271 13948 23324
rect 14016 23271 14072 23324
rect 14140 23271 14196 23327
rect 13768 23200 13786 23203
rect 13786 23200 13824 23203
rect 13892 23200 13910 23203
rect 13910 23200 13948 23203
rect 14016 23200 14034 23203
rect 14034 23200 14072 23203
rect 13768 23147 13824 23200
rect 13892 23147 13948 23200
rect 14016 23147 14072 23200
rect 14140 23147 14196 23203
rect 13768 23076 13786 23079
rect 13786 23076 13824 23079
rect 13892 23076 13910 23079
rect 13910 23076 13948 23079
rect 14016 23076 14034 23079
rect 14034 23076 14072 23079
rect 13768 23023 13824 23076
rect 13892 23023 13948 23076
rect 14016 23023 14072 23076
rect 14140 23023 14196 23079
rect 13768 22952 13786 22955
rect 13786 22952 13824 22955
rect 13892 22952 13910 22955
rect 13910 22952 13948 22955
rect 14016 22952 14034 22955
rect 14034 22952 14072 22955
rect 13768 22899 13824 22952
rect 13892 22899 13948 22952
rect 14016 22899 14072 22952
rect 14140 22899 14196 22955
rect 13768 22828 13786 22831
rect 13786 22828 13824 22831
rect 13892 22828 13910 22831
rect 13910 22828 13948 22831
rect 14016 22828 14034 22831
rect 14034 22828 14072 22831
rect 13768 22775 13824 22828
rect 13892 22775 13948 22828
rect 14016 22775 14072 22828
rect 14140 22775 14196 22831
rect 13768 22704 13786 22707
rect 13786 22704 13824 22707
rect 13892 22704 13910 22707
rect 13910 22704 13948 22707
rect 14016 22704 14034 22707
rect 14034 22704 14072 22707
rect 13768 22651 13824 22704
rect 13892 22651 13948 22704
rect 14016 22651 14072 22704
rect 14140 22651 14196 22707
rect 13768 22580 13786 22583
rect 13786 22580 13824 22583
rect 13892 22580 13910 22583
rect 13910 22580 13948 22583
rect 14016 22580 14034 22583
rect 14034 22580 14072 22583
rect 13768 22527 13824 22580
rect 13892 22527 13948 22580
rect 14016 22527 14072 22580
rect 14140 22527 14196 22583
rect 13768 22456 13786 22459
rect 13786 22456 13824 22459
rect 13892 22456 13910 22459
rect 13910 22456 13948 22459
rect 14016 22456 14034 22459
rect 14034 22456 14072 22459
rect 13768 22403 13824 22456
rect 13892 22403 13948 22456
rect 14016 22403 14072 22456
rect 14140 22403 14196 22459
rect 13768 22332 13786 22335
rect 13786 22332 13824 22335
rect 13892 22332 13910 22335
rect 13910 22332 13948 22335
rect 14016 22332 14034 22335
rect 14034 22332 14072 22335
rect 13768 22279 13824 22332
rect 13892 22279 13948 22332
rect 14016 22279 14072 22332
rect 14140 22279 14196 22335
rect 13768 22208 13786 22211
rect 13786 22208 13824 22211
rect 13892 22208 13910 22211
rect 13910 22208 13948 22211
rect 14016 22208 14034 22211
rect 14034 22208 14072 22211
rect 13768 22155 13824 22208
rect 13892 22155 13948 22208
rect 14016 22155 14072 22208
rect 14140 22155 14196 22211
rect 13768 22084 13786 22087
rect 13786 22084 13824 22087
rect 13892 22084 13910 22087
rect 13910 22084 13948 22087
rect 14016 22084 14034 22087
rect 14034 22084 14072 22087
rect 13768 22031 13824 22084
rect 13892 22031 13948 22084
rect 14016 22031 14072 22084
rect 14140 22031 14196 22087
rect 13768 21960 13786 21963
rect 13786 21960 13824 21963
rect 13892 21960 13910 21963
rect 13910 21960 13948 21963
rect 14016 21960 14034 21963
rect 14034 21960 14072 21963
rect 13768 21907 13824 21960
rect 13892 21907 13948 21960
rect 14016 21907 14072 21960
rect 14140 21907 14196 21963
rect 13768 21836 13786 21839
rect 13786 21836 13824 21839
rect 13892 21836 13910 21839
rect 13910 21836 13948 21839
rect 14016 21836 14034 21839
rect 14034 21836 14072 21839
rect 13768 21783 13824 21836
rect 13892 21783 13948 21836
rect 14016 21783 14072 21836
rect 14140 21783 14196 21839
rect 13768 21712 13786 21715
rect 13786 21712 13824 21715
rect 13892 21712 13910 21715
rect 13910 21712 13948 21715
rect 14016 21712 14034 21715
rect 14034 21712 14072 21715
rect 13768 21659 13824 21712
rect 13892 21659 13948 21712
rect 14016 21659 14072 21712
rect 14140 21659 14196 21715
rect 13768 21588 13786 21591
rect 13786 21588 13824 21591
rect 13892 21588 13910 21591
rect 13910 21588 13948 21591
rect 14016 21588 14034 21591
rect 14034 21588 14072 21591
rect 13768 21535 13824 21588
rect 13892 21535 13948 21588
rect 14016 21535 14072 21588
rect 14140 21535 14196 21591
rect 13768 21411 13824 21467
rect 13892 21411 13948 21467
rect 14016 21411 14072 21467
rect 14140 21411 14196 21467
rect 13768 21287 13824 21343
rect 13892 21287 13948 21343
rect 14016 21287 14072 21343
rect 14140 21287 14196 21343
rect 13768 21163 13824 21219
rect 13892 21163 13948 21219
rect 14016 21163 14072 21219
rect 14140 21163 14196 21219
rect 13768 21039 13824 21095
rect 13892 21039 13948 21095
rect 14016 21039 14072 21095
rect 14140 21039 14196 21095
rect 13768 20915 13824 20971
rect 13892 20915 13948 20971
rect 14016 20915 14072 20971
rect 14140 20915 14196 20971
rect 13768 20791 13824 20847
rect 13892 20791 13948 20847
rect 14016 20791 14072 20847
rect 14140 20791 14196 20847
rect 13768 20667 13824 20723
rect 13892 20667 13948 20723
rect 14016 20667 14072 20723
rect 14140 20667 14196 20723
rect 13768 20543 13824 20599
rect 13892 20543 13948 20599
rect 14016 20543 14072 20599
rect 14140 20543 14196 20599
rect 13768 20195 13824 20251
rect 13892 20195 13948 20251
rect 14016 20195 14072 20251
rect 14140 20195 14196 20251
rect 13768 20071 13824 20127
rect 13892 20071 13948 20127
rect 14016 20071 14072 20127
rect 14140 20071 14196 20127
rect 13768 19947 13824 20003
rect 13892 19947 13948 20003
rect 14016 19947 14072 20003
rect 14140 19947 14196 20003
rect 13768 19823 13824 19879
rect 13892 19823 13948 19879
rect 14016 19823 14072 19879
rect 14140 19823 14196 19879
rect 13768 19699 13824 19755
rect 13892 19699 13948 19755
rect 14016 19699 14072 19755
rect 14140 19699 14196 19755
rect 13768 19575 13824 19631
rect 13892 19575 13948 19631
rect 14016 19575 14072 19631
rect 14140 19575 14196 19631
rect 13768 19451 13824 19507
rect 13892 19451 13948 19507
rect 14016 19451 14072 19507
rect 14140 19451 14196 19507
rect 13768 19327 13824 19383
rect 13892 19327 13948 19383
rect 14016 19327 14072 19383
rect 14140 19327 14196 19383
rect 13768 19203 13824 19259
rect 13892 19203 13948 19259
rect 14016 19203 14072 19259
rect 14140 19203 14196 19259
rect 13768 19079 13824 19135
rect 13892 19079 13948 19135
rect 14016 19079 14072 19135
rect 14140 19079 14196 19135
rect 13768 18955 13824 19011
rect 13892 18955 13948 19011
rect 14016 18955 14072 19011
rect 14140 18955 14196 19011
rect 13768 18831 13824 18887
rect 13892 18831 13948 18887
rect 14016 18831 14072 18887
rect 14140 18831 14196 18887
rect 13768 18707 13824 18763
rect 13892 18707 13948 18763
rect 14016 18707 14072 18763
rect 14140 18707 14196 18763
rect 13768 18583 13824 18639
rect 13892 18583 13948 18639
rect 14016 18583 14072 18639
rect 14140 18583 14196 18639
rect 13768 18459 13824 18515
rect 13892 18459 13948 18515
rect 14016 18459 14072 18515
rect 14140 18459 14196 18515
rect 13768 18335 13824 18391
rect 13892 18335 13948 18391
rect 14016 18335 14072 18391
rect 14140 18335 14196 18391
rect 13768 18211 13824 18267
rect 13892 18211 13948 18267
rect 14016 18211 14072 18267
rect 14140 18211 14196 18267
rect 13768 18087 13824 18143
rect 13892 18087 13948 18143
rect 14016 18087 14072 18143
rect 14140 18087 14196 18143
rect 13768 17963 13824 18019
rect 13892 17963 13948 18019
rect 14016 17963 14072 18019
rect 14140 17963 14196 18019
rect 13768 17839 13824 17895
rect 13892 17839 13948 17895
rect 14016 17839 14072 17895
rect 14140 17839 14196 17895
rect 13768 17715 13824 17771
rect 13892 17715 13948 17771
rect 14016 17715 14072 17771
rect 14140 17715 14196 17771
rect 13768 17591 13824 17647
rect 13892 17591 13948 17647
rect 14016 17591 14072 17647
rect 14140 17591 14196 17647
rect 13768 17467 13824 17523
rect 13892 17467 13948 17523
rect 14016 17467 14072 17523
rect 14140 17467 14196 17523
rect 13768 17343 13824 17399
rect 13892 17343 13948 17399
rect 14016 17343 14072 17399
rect 14140 17343 14196 17399
rect 13768 16995 13824 17051
rect 13892 16995 13948 17051
rect 14016 16995 14072 17051
rect 14140 16995 14196 17051
rect 13768 16871 13824 16927
rect 13892 16871 13948 16927
rect 14016 16871 14072 16927
rect 14140 16871 14196 16927
rect 13768 16747 13824 16803
rect 13892 16747 13948 16803
rect 14016 16747 14072 16803
rect 14140 16747 14196 16803
rect 13768 16623 13824 16679
rect 13892 16623 13948 16679
rect 14016 16623 14072 16679
rect 14140 16623 14196 16679
rect 13768 16499 13824 16555
rect 13892 16499 13948 16555
rect 14016 16499 14072 16555
rect 14140 16499 14196 16555
rect 13768 16375 13824 16431
rect 13892 16375 13948 16431
rect 14016 16375 14072 16431
rect 14140 16375 14196 16431
rect 13768 16251 13824 16307
rect 13892 16251 13948 16307
rect 14016 16251 14072 16307
rect 14140 16251 14196 16307
rect 13768 16127 13824 16183
rect 13892 16127 13948 16183
rect 14016 16127 14072 16183
rect 14140 16127 14196 16183
rect 13768 16003 13824 16059
rect 13892 16003 13948 16059
rect 14016 16003 14072 16059
rect 14140 16003 14196 16059
rect 13768 15879 13824 15935
rect 13892 15879 13948 15935
rect 14016 15879 14072 15935
rect 14140 15879 14196 15935
rect 12632 15631 12688 15687
rect 12756 15631 12812 15687
rect 12880 15631 12936 15687
rect 13004 15631 13060 15687
rect 12632 15507 12688 15563
rect 12756 15507 12812 15563
rect 12880 15507 12936 15563
rect 13004 15507 13060 15563
rect 12632 15383 12688 15439
rect 12756 15383 12812 15439
rect 12880 15383 12936 15439
rect 13004 15383 13060 15439
rect 12632 15259 12688 15315
rect 12756 15259 12812 15315
rect 12880 15259 12936 15315
rect 13004 15259 13060 15315
rect 12632 15135 12688 15191
rect 12756 15135 12812 15191
rect 12880 15135 12936 15191
rect 13004 15135 13060 15191
rect 12632 15011 12688 15067
rect 12756 15011 12812 15067
rect 12880 15011 12936 15067
rect 13004 15011 13060 15067
rect 12632 14887 12688 14943
rect 12756 14887 12812 14943
rect 12880 14887 12936 14943
rect 13004 14887 13060 14943
rect 12632 14763 12688 14819
rect 12756 14763 12812 14819
rect 12880 14763 12936 14819
rect 13004 14763 13060 14819
rect 12632 14639 12688 14695
rect 12756 14639 12812 14695
rect 12880 14639 12936 14695
rect 13004 14639 13060 14695
rect 12632 14515 12688 14571
rect 12756 14515 12812 14571
rect 12880 14515 12936 14571
rect 13004 14515 13060 14571
rect 12632 14391 12688 14447
rect 12756 14391 12812 14447
rect 12880 14391 12936 14447
rect 13004 14391 13060 14447
rect 12632 14267 12688 14323
rect 12756 14267 12812 14323
rect 12880 14267 12936 14323
rect 13004 14267 13060 14323
rect 12632 14143 12688 14199
rect 12756 14143 12812 14199
rect 12880 14143 12936 14199
rect 13004 14143 13060 14199
rect 13768 15755 13824 15811
rect 13892 15755 13948 15811
rect 14016 15755 14072 15811
rect 14140 15755 14196 15811
rect 13768 15631 13824 15687
rect 13892 15631 13948 15687
rect 14016 15631 14072 15687
rect 14140 15631 14196 15687
rect 13768 15507 13824 15563
rect 13892 15507 13948 15563
rect 14016 15507 14072 15563
rect 14140 15507 14196 15563
rect 13768 15383 13824 15439
rect 13892 15383 13948 15439
rect 14016 15383 14072 15439
rect 14140 15383 14196 15439
rect 13768 15259 13824 15315
rect 13892 15259 13948 15315
rect 14016 15259 14072 15315
rect 14140 15259 14196 15315
rect 13768 15135 13824 15191
rect 13892 15135 13948 15191
rect 14016 15135 14072 15191
rect 14140 15135 14196 15191
rect 13768 15011 13824 15067
rect 13892 15011 13948 15067
rect 14016 15011 14072 15067
rect 14140 15011 14196 15067
rect 13768 14887 13824 14943
rect 13892 14887 13948 14943
rect 14016 14887 14072 14943
rect 14140 14887 14196 14943
rect 13768 14763 13824 14819
rect 13892 14763 13948 14819
rect 14016 14763 14072 14819
rect 14140 14763 14196 14819
rect 13768 14639 13824 14695
rect 13892 14639 13948 14695
rect 14016 14639 14072 14695
rect 14140 14639 14196 14695
rect 13768 14515 13824 14571
rect 13892 14515 13948 14571
rect 14016 14515 14072 14571
rect 14140 14515 14196 14571
rect 13768 14391 13824 14447
rect 13892 14391 13948 14447
rect 14016 14391 14072 14447
rect 14140 14391 14196 14447
rect 13768 14267 13824 14323
rect 13892 14267 13948 14323
rect 14016 14267 14072 14323
rect 14140 14267 14196 14323
rect 13768 14143 13824 14199
rect 13892 14143 13948 14199
rect 14016 14143 14072 14199
rect 14140 14143 14196 14199
rect 300 13789 356 13845
rect 424 13789 480 13845
rect 548 13789 604 13845
rect 672 13789 728 13845
rect 300 13665 356 13721
rect 424 13665 480 13721
rect 548 13665 604 13721
rect 672 13665 728 13721
rect 300 13541 356 13597
rect 424 13541 480 13597
rect 548 13541 604 13597
rect 672 13541 728 13597
rect 300 13417 356 13473
rect 424 13417 480 13473
rect 548 13417 604 13473
rect 672 13417 728 13473
rect 300 13293 356 13349
rect 424 13293 480 13349
rect 548 13293 604 13349
rect 672 13293 728 13349
rect 300 13169 356 13225
rect 424 13169 480 13225
rect 548 13169 604 13225
rect 672 13169 728 13225
rect 300 13045 356 13101
rect 424 13045 480 13101
rect 548 13045 604 13101
rect 672 13045 728 13101
rect 300 12921 356 12977
rect 424 12921 480 12977
rect 548 12921 604 12977
rect 672 12921 728 12977
rect 300 12797 356 12853
rect 424 12797 480 12853
rect 548 12797 604 12853
rect 672 12797 728 12853
rect 300 12673 356 12729
rect 424 12673 480 12729
rect 548 12673 604 12729
rect 672 12673 728 12729
rect 300 12549 356 12605
rect 424 12549 480 12605
rect 548 12549 604 12605
rect 672 12549 728 12605
rect 1436 13789 1492 13845
rect 1560 13789 1616 13845
rect 1684 13789 1740 13845
rect 1808 13789 1864 13845
rect 1436 13665 1492 13721
rect 1560 13665 1616 13721
rect 1684 13665 1740 13721
rect 1808 13665 1864 13721
rect 1436 13541 1492 13597
rect 1560 13541 1616 13597
rect 1684 13541 1740 13597
rect 1808 13541 1864 13597
rect 1436 13417 1492 13473
rect 1560 13417 1616 13473
rect 1684 13417 1740 13473
rect 1808 13417 1864 13473
rect 1436 13293 1492 13349
rect 1560 13293 1616 13349
rect 1684 13293 1740 13349
rect 1808 13293 1864 13349
rect 1436 13169 1492 13225
rect 1560 13169 1616 13225
rect 1684 13169 1740 13225
rect 1808 13169 1864 13225
rect 1436 13045 1492 13101
rect 1560 13045 1616 13101
rect 1684 13045 1740 13101
rect 1808 13045 1864 13101
rect 1436 12921 1492 12977
rect 1560 12921 1616 12977
rect 1684 12921 1740 12977
rect 1808 12921 1864 12977
rect 1436 12797 1492 12853
rect 1560 12797 1616 12853
rect 1684 12797 1740 12853
rect 1808 12797 1864 12853
rect 1436 12673 1492 12729
rect 1560 12673 1616 12729
rect 1684 12673 1740 12729
rect 1808 12673 1864 12729
rect 1436 12549 1492 12605
rect 1560 12549 1616 12605
rect 1684 12549 1740 12605
rect 1808 12549 1864 12605
rect 2572 13789 2628 13845
rect 2696 13789 2752 13845
rect 2820 13789 2876 13845
rect 2944 13789 3000 13845
rect 2572 13665 2628 13721
rect 2696 13665 2752 13721
rect 2820 13665 2876 13721
rect 2944 13665 3000 13721
rect 2572 13541 2628 13597
rect 2696 13541 2752 13597
rect 2820 13541 2876 13597
rect 2944 13541 3000 13597
rect 2572 13417 2628 13473
rect 2696 13417 2752 13473
rect 2820 13417 2876 13473
rect 2944 13417 3000 13473
rect 2572 13293 2628 13349
rect 2696 13293 2752 13349
rect 2820 13293 2876 13349
rect 2944 13293 3000 13349
rect 2572 13169 2628 13225
rect 2696 13169 2752 13225
rect 2820 13169 2876 13225
rect 2944 13169 3000 13225
rect 2572 13045 2628 13101
rect 2696 13045 2752 13101
rect 2820 13045 2876 13101
rect 2944 13045 3000 13101
rect 2572 12921 2628 12977
rect 2696 12921 2752 12977
rect 2820 12921 2876 12977
rect 2944 12921 3000 12977
rect 2572 12797 2628 12853
rect 2696 12797 2752 12853
rect 2820 12797 2876 12853
rect 2944 12797 3000 12853
rect 2572 12673 2628 12729
rect 2696 12673 2752 12729
rect 2820 12673 2876 12729
rect 2944 12673 3000 12729
rect 2572 12549 2628 12605
rect 2696 12549 2752 12605
rect 2820 12549 2876 12605
rect 2944 12549 3000 12605
rect 4844 13789 4900 13845
rect 4968 13789 5024 13845
rect 5092 13789 5148 13845
rect 5216 13789 5272 13845
rect 4844 13665 4900 13721
rect 4968 13665 5024 13721
rect 5092 13665 5148 13721
rect 5216 13665 5272 13721
rect 4844 13541 4900 13597
rect 4968 13541 5024 13597
rect 5092 13541 5148 13597
rect 5216 13541 5272 13597
rect 4844 13417 4900 13473
rect 4968 13417 5024 13473
rect 5092 13417 5148 13473
rect 5216 13417 5272 13473
rect 4844 13293 4900 13349
rect 4968 13293 5024 13349
rect 5092 13293 5148 13349
rect 5216 13293 5272 13349
rect 4844 13169 4900 13225
rect 4968 13169 5024 13225
rect 5092 13169 5148 13225
rect 5216 13169 5272 13225
rect 4844 13045 4900 13101
rect 4968 13045 5024 13101
rect 5092 13045 5148 13101
rect 5216 13045 5272 13101
rect 4844 12921 4900 12977
rect 4968 12921 5024 12977
rect 5092 12921 5148 12977
rect 5216 12921 5272 12977
rect 4844 12797 4900 12853
rect 4968 12797 5024 12853
rect 5092 12797 5148 12853
rect 5216 12797 5272 12853
rect 4844 12673 4900 12729
rect 4968 12673 5024 12729
rect 5092 12673 5148 12729
rect 5216 12673 5272 12729
rect 4844 12549 4900 12605
rect 4968 12549 5024 12605
rect 5092 12549 5148 12605
rect 5216 12549 5272 12605
rect 7137 13789 7193 13845
rect 7261 13789 7317 13845
rect 7385 13789 7441 13845
rect 7137 13665 7193 13721
rect 7261 13665 7317 13721
rect 7385 13665 7441 13721
rect 7137 13541 7193 13597
rect 7261 13541 7317 13597
rect 7385 13541 7441 13597
rect 7137 13417 7193 13473
rect 7261 13417 7317 13473
rect 7385 13417 7441 13473
rect 7137 13293 7193 13349
rect 7261 13293 7317 13349
rect 7385 13293 7441 13349
rect 7137 13169 7193 13225
rect 7261 13169 7317 13225
rect 7385 13169 7441 13225
rect 7137 13045 7193 13101
rect 7261 13045 7317 13101
rect 7385 13045 7441 13101
rect 7137 12921 7193 12977
rect 7261 12921 7317 12977
rect 7385 12921 7441 12977
rect 7137 12797 7193 12853
rect 7261 12797 7317 12853
rect 7385 12797 7441 12853
rect 7137 12673 7193 12729
rect 7261 12673 7317 12729
rect 7385 12673 7441 12729
rect 7137 12549 7193 12605
rect 7261 12549 7317 12605
rect 7385 12549 7441 12605
rect 7623 13789 7679 13845
rect 7747 13789 7803 13845
rect 7871 13789 7927 13845
rect 7623 13665 7679 13721
rect 7747 13665 7803 13721
rect 7871 13665 7927 13721
rect 7623 13541 7679 13597
rect 7747 13541 7803 13597
rect 7871 13541 7927 13597
rect 7623 13417 7679 13473
rect 7747 13417 7803 13473
rect 7871 13417 7927 13473
rect 7623 13293 7679 13349
rect 7747 13293 7803 13349
rect 7871 13293 7927 13349
rect 7623 13169 7679 13225
rect 7747 13169 7803 13225
rect 7871 13169 7927 13225
rect 7623 13045 7679 13101
rect 7747 13045 7803 13101
rect 7871 13045 7927 13101
rect 7623 12921 7679 12977
rect 7747 12921 7803 12977
rect 7871 12921 7927 12977
rect 7623 12797 7679 12853
rect 7747 12797 7803 12853
rect 7871 12797 7927 12853
rect 7623 12673 7679 12729
rect 7747 12673 7803 12729
rect 7871 12673 7927 12729
rect 7623 12549 7679 12605
rect 7747 12549 7803 12605
rect 7871 12549 7927 12605
rect 9792 13789 9848 13845
rect 9916 13789 9972 13845
rect 10040 13789 10096 13845
rect 10164 13789 10220 13845
rect 9792 13665 9848 13721
rect 9916 13665 9972 13721
rect 10040 13665 10096 13721
rect 10164 13665 10220 13721
rect 9792 13541 9848 13597
rect 9916 13541 9972 13597
rect 10040 13541 10096 13597
rect 10164 13541 10220 13597
rect 9792 13417 9848 13473
rect 9916 13417 9972 13473
rect 10040 13417 10096 13473
rect 10164 13417 10220 13473
rect 9792 13293 9848 13349
rect 9916 13293 9972 13349
rect 10040 13293 10096 13349
rect 10164 13293 10220 13349
rect 9792 13169 9848 13225
rect 9916 13169 9972 13225
rect 10040 13169 10096 13225
rect 10164 13169 10220 13225
rect 9792 13045 9848 13101
rect 9916 13045 9972 13101
rect 10040 13045 10096 13101
rect 10164 13045 10220 13101
rect 9792 12921 9848 12977
rect 9916 12921 9972 12977
rect 10040 12921 10096 12977
rect 10164 12921 10220 12977
rect 9792 12797 9848 12853
rect 9916 12797 9972 12853
rect 10040 12797 10096 12853
rect 10164 12797 10220 12853
rect 9792 12673 9848 12729
rect 9916 12673 9972 12729
rect 10040 12673 10096 12729
rect 10164 12673 10220 12729
rect 9792 12549 9848 12605
rect 9916 12549 9972 12605
rect 10040 12549 10096 12605
rect 10164 12549 10220 12605
rect 12064 13789 12120 13845
rect 12188 13789 12244 13845
rect 12312 13789 12368 13845
rect 12436 13789 12492 13845
rect 12064 13665 12120 13721
rect 12188 13665 12244 13721
rect 12312 13665 12368 13721
rect 12436 13665 12492 13721
rect 12064 13541 12120 13597
rect 12188 13541 12244 13597
rect 12312 13541 12368 13597
rect 12436 13541 12492 13597
rect 12064 13417 12120 13473
rect 12188 13417 12244 13473
rect 12312 13417 12368 13473
rect 12436 13417 12492 13473
rect 12064 13293 12120 13349
rect 12188 13293 12244 13349
rect 12312 13293 12368 13349
rect 12436 13293 12492 13349
rect 12064 13169 12120 13225
rect 12188 13169 12244 13225
rect 12312 13169 12368 13225
rect 12436 13169 12492 13225
rect 12064 13045 12120 13101
rect 12188 13045 12244 13101
rect 12312 13045 12368 13101
rect 12436 13045 12492 13101
rect 12064 12921 12120 12977
rect 12188 12921 12244 12977
rect 12312 12921 12368 12977
rect 12436 12921 12492 12977
rect 12064 12797 12120 12853
rect 12188 12797 12244 12853
rect 12312 12797 12368 12853
rect 12436 12797 12492 12853
rect 12064 12673 12120 12729
rect 12188 12673 12244 12729
rect 12312 12673 12368 12729
rect 12436 12673 12492 12729
rect 12064 12549 12120 12605
rect 12188 12549 12244 12605
rect 12312 12549 12368 12605
rect 12436 12549 12492 12605
rect 13200 13789 13256 13845
rect 13324 13789 13380 13845
rect 13448 13789 13504 13845
rect 13572 13789 13628 13845
rect 13200 13665 13256 13721
rect 13324 13665 13380 13721
rect 13448 13665 13504 13721
rect 13572 13665 13628 13721
rect 13200 13541 13256 13597
rect 13324 13541 13380 13597
rect 13448 13541 13504 13597
rect 13572 13541 13628 13597
rect 13200 13417 13256 13473
rect 13324 13417 13380 13473
rect 13448 13417 13504 13473
rect 13572 13417 13628 13473
rect 13200 13293 13256 13349
rect 13324 13293 13380 13349
rect 13448 13293 13504 13349
rect 13572 13293 13628 13349
rect 13200 13169 13256 13225
rect 13324 13169 13380 13225
rect 13448 13169 13504 13225
rect 13572 13169 13628 13225
rect 13200 13045 13256 13101
rect 13324 13045 13380 13101
rect 13448 13045 13504 13101
rect 13572 13045 13628 13101
rect 13200 12921 13256 12977
rect 13324 12921 13380 12977
rect 13448 12921 13504 12977
rect 13572 12921 13628 12977
rect 13200 12797 13256 12853
rect 13324 12797 13380 12853
rect 13448 12797 13504 12853
rect 13572 12797 13628 12853
rect 13200 12673 13256 12729
rect 13324 12673 13380 12729
rect 13448 12673 13504 12729
rect 13572 12673 13628 12729
rect 13200 12549 13256 12605
rect 13324 12549 13380 12605
rect 13448 12549 13504 12605
rect 13572 12549 13628 12605
rect 868 12189 924 12245
rect 992 12189 1048 12245
rect 1116 12189 1172 12245
rect 1240 12189 1296 12245
rect 868 12065 924 12121
rect 992 12065 1048 12121
rect 1116 12065 1172 12121
rect 1240 12065 1296 12121
rect 868 11941 924 11997
rect 992 11941 1048 11997
rect 1116 11941 1172 11997
rect 1240 11941 1296 11997
rect 868 11817 924 11873
rect 992 11817 1048 11873
rect 1116 11817 1172 11873
rect 1240 11817 1296 11873
rect 868 11693 924 11749
rect 992 11693 1048 11749
rect 1116 11693 1172 11749
rect 1240 11693 1296 11749
rect 868 11569 924 11625
rect 992 11569 1048 11625
rect 1116 11569 1172 11625
rect 1240 11569 1296 11625
rect 868 11445 924 11501
rect 992 11445 1048 11501
rect 1116 11445 1172 11501
rect 1240 11445 1296 11501
rect 868 11321 924 11377
rect 992 11321 1048 11377
rect 1116 11321 1172 11377
rect 1240 11321 1296 11377
rect 868 11197 924 11253
rect 992 11197 1048 11253
rect 1116 11197 1172 11253
rect 1240 11197 1296 11253
rect 868 11073 924 11129
rect 992 11073 1048 11129
rect 1116 11073 1172 11129
rect 1240 11073 1296 11129
rect 868 10949 924 11005
rect 992 10949 1048 11005
rect 1116 10949 1172 11005
rect 1240 10949 1296 11005
rect 2004 12189 2060 12245
rect 2128 12189 2184 12245
rect 2252 12189 2308 12245
rect 2376 12189 2432 12245
rect 2004 12065 2060 12121
rect 2128 12065 2184 12121
rect 2252 12065 2308 12121
rect 2376 12065 2432 12121
rect 2004 11941 2060 11997
rect 2128 11941 2184 11997
rect 2252 11941 2308 11997
rect 2376 11941 2432 11997
rect 2004 11817 2060 11873
rect 2128 11817 2184 11873
rect 2252 11817 2308 11873
rect 2376 11817 2432 11873
rect 2004 11693 2060 11749
rect 2128 11693 2184 11749
rect 2252 11693 2308 11749
rect 2376 11693 2432 11749
rect 2004 11569 2060 11625
rect 2128 11569 2184 11625
rect 2252 11569 2308 11625
rect 2376 11569 2432 11625
rect 2004 11445 2060 11501
rect 2128 11445 2184 11501
rect 2252 11445 2308 11501
rect 2376 11445 2432 11501
rect 2004 11321 2060 11377
rect 2128 11321 2184 11377
rect 2252 11321 2308 11377
rect 2376 11321 2432 11377
rect 2004 11197 2060 11253
rect 2128 11197 2184 11253
rect 2252 11197 2308 11253
rect 2376 11197 2432 11253
rect 2004 11073 2060 11129
rect 2128 11073 2184 11129
rect 2252 11073 2308 11129
rect 2376 11073 2432 11129
rect 2004 10949 2060 11005
rect 2128 10949 2184 11005
rect 2252 10949 2308 11005
rect 2376 10949 2432 11005
rect 3708 12189 3764 12245
rect 3832 12189 3888 12245
rect 3956 12189 4012 12245
rect 4080 12189 4136 12245
rect 3708 12065 3764 12121
rect 3832 12065 3888 12121
rect 3956 12065 4012 12121
rect 4080 12065 4136 12121
rect 3708 11941 3764 11997
rect 3832 11941 3888 11997
rect 3956 11941 4012 11997
rect 4080 11941 4136 11997
rect 3708 11817 3764 11873
rect 3832 11817 3888 11873
rect 3956 11817 4012 11873
rect 4080 11817 4136 11873
rect 3708 11693 3764 11749
rect 3832 11693 3888 11749
rect 3956 11693 4012 11749
rect 4080 11693 4136 11749
rect 3708 11569 3764 11625
rect 3832 11569 3888 11625
rect 3956 11569 4012 11625
rect 4080 11569 4136 11625
rect 3708 11445 3764 11501
rect 3832 11445 3888 11501
rect 3956 11445 4012 11501
rect 4080 11445 4136 11501
rect 3708 11321 3764 11377
rect 3832 11321 3888 11377
rect 3956 11321 4012 11377
rect 4080 11321 4136 11377
rect 3708 11197 3764 11253
rect 3832 11197 3888 11253
rect 3956 11197 4012 11253
rect 4080 11197 4136 11253
rect 3708 11073 3764 11129
rect 3832 11073 3888 11129
rect 3956 11073 4012 11129
rect 4080 11073 4136 11129
rect 3708 10949 3764 11005
rect 3832 10949 3888 11005
rect 3956 10949 4012 11005
rect 4080 10949 4136 11005
rect 5980 12189 6036 12245
rect 6104 12189 6160 12245
rect 6228 12189 6284 12245
rect 6352 12189 6408 12245
rect 5980 12065 6036 12121
rect 6104 12065 6160 12121
rect 6228 12065 6284 12121
rect 6352 12065 6408 12121
rect 5980 11941 6036 11997
rect 6104 11941 6160 11997
rect 6228 11941 6284 11997
rect 6352 11941 6408 11997
rect 5980 11817 6036 11873
rect 6104 11817 6160 11873
rect 6228 11817 6284 11873
rect 6352 11817 6408 11873
rect 5980 11693 6036 11749
rect 6104 11693 6160 11749
rect 6228 11693 6284 11749
rect 6352 11693 6408 11749
rect 5980 11569 6036 11625
rect 6104 11569 6160 11625
rect 6228 11569 6284 11625
rect 6352 11569 6408 11625
rect 5980 11445 6036 11501
rect 6104 11445 6160 11501
rect 6228 11445 6284 11501
rect 6352 11445 6408 11501
rect 5980 11321 6036 11377
rect 6104 11321 6160 11377
rect 6228 11321 6284 11377
rect 6352 11321 6408 11377
rect 5980 11197 6036 11253
rect 6104 11197 6160 11253
rect 6228 11197 6284 11253
rect 6352 11197 6408 11253
rect 5980 11073 6036 11129
rect 6104 11073 6160 11129
rect 6228 11073 6284 11129
rect 6352 11073 6408 11129
rect 5980 10949 6036 11005
rect 6104 10949 6160 11005
rect 6228 10949 6284 11005
rect 6352 10949 6408 11005
rect 8656 12189 8712 12245
rect 8780 12189 8836 12245
rect 8904 12189 8960 12245
rect 9028 12189 9084 12245
rect 8656 12065 8712 12121
rect 8780 12065 8836 12121
rect 8904 12065 8960 12121
rect 9028 12065 9084 12121
rect 8656 11941 8712 11997
rect 8780 11941 8836 11997
rect 8904 11941 8960 11997
rect 9028 11941 9084 11997
rect 8656 11817 8712 11873
rect 8780 11817 8836 11873
rect 8904 11817 8960 11873
rect 9028 11817 9084 11873
rect 8656 11693 8712 11749
rect 8780 11693 8836 11749
rect 8904 11693 8960 11749
rect 9028 11693 9084 11749
rect 8656 11569 8712 11625
rect 8780 11569 8836 11625
rect 8904 11569 8960 11625
rect 9028 11569 9084 11625
rect 8656 11445 8712 11501
rect 8780 11445 8836 11501
rect 8904 11445 8960 11501
rect 9028 11445 9084 11501
rect 8656 11321 8712 11377
rect 8780 11321 8836 11377
rect 8904 11321 8960 11377
rect 9028 11321 9084 11377
rect 8656 11197 8712 11253
rect 8780 11197 8836 11253
rect 8904 11197 8960 11253
rect 9028 11197 9084 11253
rect 8656 11073 8712 11129
rect 8780 11073 8836 11129
rect 8904 11073 8960 11129
rect 9028 11073 9084 11129
rect 8656 10949 8712 11005
rect 8780 10949 8836 11005
rect 8904 10949 8960 11005
rect 9028 10949 9084 11005
rect 10928 12189 10984 12245
rect 11052 12189 11108 12245
rect 11176 12189 11232 12245
rect 11300 12189 11356 12245
rect 10928 12065 10984 12121
rect 11052 12065 11108 12121
rect 11176 12065 11232 12121
rect 11300 12065 11356 12121
rect 10928 11941 10984 11997
rect 11052 11941 11108 11997
rect 11176 11941 11232 11997
rect 11300 11941 11356 11997
rect 10928 11817 10984 11873
rect 11052 11817 11108 11873
rect 11176 11817 11232 11873
rect 11300 11817 11356 11873
rect 10928 11693 10984 11749
rect 11052 11693 11108 11749
rect 11176 11693 11232 11749
rect 11300 11693 11356 11749
rect 10928 11569 10984 11625
rect 11052 11569 11108 11625
rect 11176 11569 11232 11625
rect 11300 11569 11356 11625
rect 10928 11445 10984 11501
rect 11052 11445 11108 11501
rect 11176 11445 11232 11501
rect 11300 11445 11356 11501
rect 10928 11321 10984 11377
rect 11052 11321 11108 11377
rect 11176 11321 11232 11377
rect 11300 11321 11356 11377
rect 10928 11197 10984 11253
rect 11052 11197 11108 11253
rect 11176 11197 11232 11253
rect 11300 11197 11356 11253
rect 10928 11073 10984 11129
rect 11052 11073 11108 11129
rect 11176 11073 11232 11129
rect 11300 11073 11356 11129
rect 10928 10949 10984 11005
rect 11052 10949 11108 11005
rect 11176 10949 11232 11005
rect 11300 10949 11356 11005
rect 12632 12189 12688 12245
rect 12756 12189 12812 12245
rect 12880 12189 12936 12245
rect 13004 12189 13060 12245
rect 12632 12065 12688 12121
rect 12756 12065 12812 12121
rect 12880 12065 12936 12121
rect 13004 12065 13060 12121
rect 12632 11941 12688 11997
rect 12756 11941 12812 11997
rect 12880 11941 12936 11997
rect 13004 11941 13060 11997
rect 12632 11817 12688 11873
rect 12756 11817 12812 11873
rect 12880 11817 12936 11873
rect 13004 11817 13060 11873
rect 12632 11693 12688 11749
rect 12756 11693 12812 11749
rect 12880 11693 12936 11749
rect 13004 11693 13060 11749
rect 12632 11569 12688 11625
rect 12756 11569 12812 11625
rect 12880 11569 12936 11625
rect 13004 11569 13060 11625
rect 12632 11445 12688 11501
rect 12756 11445 12812 11501
rect 12880 11445 12936 11501
rect 13004 11445 13060 11501
rect 12632 11321 12688 11377
rect 12756 11321 12812 11377
rect 12880 11321 12936 11377
rect 13004 11321 13060 11377
rect 12632 11197 12688 11253
rect 12756 11197 12812 11253
rect 12880 11197 12936 11253
rect 13004 11197 13060 11253
rect 12632 11073 12688 11129
rect 12756 11073 12812 11129
rect 12880 11073 12936 11129
rect 13004 11073 13060 11129
rect 12632 10949 12688 11005
rect 12756 10949 12812 11005
rect 12880 10949 12936 11005
rect 13004 10949 13060 11005
rect 13768 12189 13824 12245
rect 13892 12189 13948 12245
rect 14016 12189 14072 12245
rect 14140 12189 14196 12245
rect 13768 12065 13824 12121
rect 13892 12065 13948 12121
rect 14016 12065 14072 12121
rect 14140 12065 14196 12121
rect 13768 11941 13824 11997
rect 13892 11941 13948 11997
rect 14016 11941 14072 11997
rect 14140 11941 14196 11997
rect 13768 11817 13824 11873
rect 13892 11817 13948 11873
rect 14016 11817 14072 11873
rect 14140 11817 14196 11873
rect 13768 11693 13824 11749
rect 13892 11693 13948 11749
rect 14016 11693 14072 11749
rect 14140 11693 14196 11749
rect 13768 11569 13824 11625
rect 13892 11569 13948 11625
rect 14016 11569 14072 11625
rect 14140 11569 14196 11625
rect 13768 11445 13824 11501
rect 13892 11445 13948 11501
rect 14016 11445 14072 11501
rect 14140 11445 14196 11501
rect 13768 11321 13824 11377
rect 13892 11321 13948 11377
rect 14016 11321 14072 11377
rect 14140 11321 14196 11377
rect 13768 11197 13824 11253
rect 13892 11197 13948 11253
rect 14016 11197 14072 11253
rect 14140 11197 14196 11253
rect 13768 11073 13824 11129
rect 13892 11073 13948 11129
rect 14016 11073 14072 11129
rect 14140 11073 14196 11129
rect 13768 10949 13824 11005
rect 13892 10949 13948 11005
rect 14016 10949 14072 11005
rect 14140 10949 14196 11005
rect 300 10595 356 10651
rect 424 10595 480 10651
rect 548 10595 604 10651
rect 672 10595 728 10651
rect 300 10471 356 10527
rect 424 10471 480 10527
rect 548 10471 604 10527
rect 672 10471 728 10527
rect 300 10347 356 10403
rect 424 10347 480 10403
rect 548 10347 604 10403
rect 672 10347 728 10403
rect 300 10223 356 10279
rect 424 10223 480 10279
rect 548 10223 604 10279
rect 672 10223 728 10279
rect 300 10099 356 10155
rect 424 10099 480 10155
rect 548 10099 604 10155
rect 672 10099 728 10155
rect 300 9975 356 10031
rect 424 9975 480 10031
rect 548 9975 604 10031
rect 672 9975 728 10031
rect 300 9851 356 9907
rect 424 9851 480 9907
rect 548 9851 604 9907
rect 672 9851 728 9907
rect 300 9727 356 9783
rect 424 9727 480 9783
rect 548 9727 604 9783
rect 672 9727 728 9783
rect 300 9603 356 9659
rect 424 9603 480 9659
rect 548 9603 604 9659
rect 672 9603 728 9659
rect 300 9479 356 9535
rect 424 9479 480 9535
rect 548 9479 604 9535
rect 672 9479 728 9535
rect 300 9355 356 9411
rect 424 9355 480 9411
rect 548 9355 604 9411
rect 672 9355 728 9411
rect 300 9231 356 9287
rect 424 9231 480 9287
rect 548 9231 604 9287
rect 672 9231 728 9287
rect 300 9107 356 9163
rect 424 9107 480 9163
rect 548 9107 604 9163
rect 672 9107 728 9163
rect 300 8983 356 9039
rect 424 8983 480 9039
rect 548 8983 604 9039
rect 672 8983 728 9039
rect 300 8859 356 8915
rect 424 8859 480 8915
rect 548 8859 604 8915
rect 672 8859 728 8915
rect 300 8735 356 8791
rect 424 8735 480 8791
rect 548 8735 604 8791
rect 672 8735 728 8791
rect 300 8611 356 8667
rect 424 8611 480 8667
rect 548 8611 604 8667
rect 672 8611 728 8667
rect 300 8487 356 8543
rect 424 8487 480 8543
rect 548 8487 604 8543
rect 672 8487 728 8543
rect 300 8363 356 8419
rect 424 8363 480 8419
rect 548 8363 604 8419
rect 672 8363 728 8419
rect 300 8239 356 8295
rect 424 8239 480 8295
rect 548 8239 604 8295
rect 672 8239 728 8295
rect 300 8115 356 8171
rect 424 8115 480 8171
rect 548 8115 604 8171
rect 672 8115 728 8171
rect 300 7991 356 8047
rect 424 7991 480 8047
rect 548 7991 604 8047
rect 672 7991 728 8047
rect 300 7867 356 7923
rect 424 7867 480 7923
rect 548 7867 604 7923
rect 672 7867 728 7923
rect 300 7743 356 7799
rect 424 7743 480 7799
rect 548 7743 604 7799
rect 672 7743 728 7799
rect 300 7395 356 7451
rect 424 7395 480 7451
rect 548 7395 604 7451
rect 672 7395 728 7451
rect 300 7271 356 7327
rect 424 7271 480 7327
rect 548 7271 604 7327
rect 672 7271 728 7327
rect 300 7147 356 7203
rect 424 7147 480 7203
rect 548 7147 604 7203
rect 672 7147 728 7203
rect 300 7023 356 7079
rect 424 7023 480 7079
rect 548 7023 604 7079
rect 672 7023 728 7079
rect 300 6899 356 6955
rect 424 6899 480 6955
rect 548 6899 604 6955
rect 672 6899 728 6955
rect 300 6775 356 6831
rect 424 6775 480 6831
rect 548 6775 604 6831
rect 672 6775 728 6831
rect 300 6651 356 6707
rect 424 6651 480 6707
rect 548 6651 604 6707
rect 672 6651 728 6707
rect 300 6527 356 6583
rect 424 6527 480 6583
rect 548 6527 604 6583
rect 672 6527 728 6583
rect 300 6403 356 6459
rect 424 6403 480 6459
rect 548 6403 604 6459
rect 672 6403 728 6459
rect 300 6279 356 6335
rect 424 6279 480 6335
rect 548 6279 604 6335
rect 672 6279 728 6335
rect 300 6155 356 6211
rect 424 6155 480 6211
rect 548 6155 604 6211
rect 672 6155 728 6211
rect 300 6031 356 6087
rect 424 6031 480 6087
rect 548 6031 604 6087
rect 672 6031 728 6087
rect 300 5907 356 5963
rect 424 5907 480 5963
rect 548 5907 604 5963
rect 672 5907 728 5963
rect 300 5783 356 5839
rect 424 5783 480 5839
rect 548 5783 604 5839
rect 672 5783 728 5839
rect 300 5659 356 5715
rect 424 5659 480 5715
rect 548 5659 604 5715
rect 672 5659 728 5715
rect 300 5535 356 5591
rect 424 5535 480 5591
rect 548 5535 604 5591
rect 672 5535 728 5591
rect 300 5411 356 5467
rect 424 5411 480 5467
rect 548 5411 604 5467
rect 672 5411 728 5467
rect 300 5287 356 5343
rect 424 5287 480 5343
rect 548 5287 604 5343
rect 672 5287 728 5343
rect 300 5163 356 5219
rect 424 5163 480 5219
rect 548 5163 604 5219
rect 672 5163 728 5219
rect 300 5039 356 5095
rect 424 5039 480 5095
rect 548 5039 604 5095
rect 672 5039 728 5095
rect 300 4915 356 4971
rect 424 4915 480 4971
rect 548 4915 604 4971
rect 672 4915 728 4971
rect 300 4791 356 4847
rect 424 4791 480 4847
rect 548 4791 604 4847
rect 672 4791 728 4847
rect 300 4667 356 4723
rect 424 4667 480 4723
rect 548 4667 604 4723
rect 672 4667 728 4723
rect 300 4543 356 4599
rect 424 4543 480 4599
rect 548 4543 604 4599
rect 672 4543 728 4599
rect 300 4195 356 4251
rect 424 4195 480 4251
rect 548 4195 604 4251
rect 672 4195 728 4251
rect 300 4071 356 4127
rect 424 4071 480 4127
rect 548 4071 604 4127
rect 672 4071 728 4127
rect 300 3947 356 4003
rect 424 3947 480 4003
rect 548 3947 604 4003
rect 672 3947 728 4003
rect 300 3823 356 3879
rect 424 3823 480 3879
rect 548 3823 604 3879
rect 672 3823 728 3879
rect 300 3699 356 3755
rect 424 3699 480 3755
rect 548 3699 604 3755
rect 672 3699 728 3755
rect 300 3575 356 3631
rect 424 3575 480 3631
rect 548 3575 604 3631
rect 672 3575 728 3631
rect 300 3451 356 3507
rect 424 3451 480 3507
rect 548 3451 604 3507
rect 672 3451 728 3507
rect 300 3327 356 3383
rect 424 3327 480 3383
rect 548 3327 604 3383
rect 672 3327 728 3383
rect 300 3203 356 3259
rect 424 3203 480 3259
rect 548 3203 604 3259
rect 672 3203 728 3259
rect 300 3079 356 3135
rect 424 3079 480 3135
rect 548 3079 604 3135
rect 672 3079 728 3135
rect 300 2955 356 3011
rect 424 2955 480 3011
rect 548 2955 604 3011
rect 672 2955 728 3011
rect 300 2831 356 2887
rect 424 2831 480 2887
rect 548 2831 604 2887
rect 672 2831 728 2887
rect 300 2707 356 2763
rect 424 2707 480 2763
rect 548 2707 604 2763
rect 672 2707 728 2763
rect 300 2583 356 2639
rect 424 2583 480 2639
rect 548 2583 604 2639
rect 672 2583 728 2639
rect 300 2459 356 2515
rect 424 2459 480 2515
rect 548 2459 604 2515
rect 672 2459 728 2515
rect 300 2335 356 2391
rect 424 2335 480 2391
rect 548 2335 604 2391
rect 672 2335 728 2391
rect 300 2211 356 2267
rect 424 2211 480 2267
rect 548 2211 604 2267
rect 672 2211 728 2267
rect 300 2087 356 2143
rect 424 2087 480 2143
rect 548 2087 604 2143
rect 672 2087 728 2143
rect 300 1963 356 2019
rect 424 1963 480 2019
rect 548 1963 604 2019
rect 672 1963 728 2019
rect 300 1839 356 1895
rect 424 1839 480 1895
rect 548 1839 604 1895
rect 672 1839 728 1895
rect 300 1715 356 1771
rect 424 1715 480 1771
rect 548 1715 604 1771
rect 672 1715 728 1771
rect 300 1591 356 1647
rect 424 1591 480 1647
rect 548 1591 604 1647
rect 672 1591 728 1647
rect 300 1467 356 1523
rect 424 1467 480 1523
rect 548 1467 604 1523
rect 672 1467 728 1523
rect 300 1343 356 1399
rect 424 1343 480 1399
rect 548 1343 604 1399
rect 672 1343 728 1399
rect 1436 10595 1492 10651
rect 1560 10595 1616 10651
rect 1684 10595 1740 10651
rect 1808 10595 1864 10651
rect 1436 10471 1492 10527
rect 1560 10471 1616 10527
rect 1684 10471 1740 10527
rect 1808 10471 1864 10527
rect 1436 10347 1492 10403
rect 1560 10347 1616 10403
rect 1684 10347 1740 10403
rect 1808 10347 1864 10403
rect 1436 10223 1492 10279
rect 1560 10223 1616 10279
rect 1684 10223 1740 10279
rect 1808 10223 1864 10279
rect 1436 10099 1492 10155
rect 1560 10099 1616 10155
rect 1684 10099 1740 10155
rect 1808 10099 1864 10155
rect 1436 9975 1492 10031
rect 1560 9975 1616 10031
rect 1684 9975 1740 10031
rect 1808 9975 1864 10031
rect 1436 9851 1492 9907
rect 1560 9851 1616 9907
rect 1684 9851 1740 9907
rect 1808 9851 1864 9907
rect 1436 9727 1492 9783
rect 1560 9727 1616 9783
rect 1684 9727 1740 9783
rect 1808 9727 1864 9783
rect 1436 9603 1492 9659
rect 1560 9603 1616 9659
rect 1684 9603 1740 9659
rect 1808 9603 1864 9659
rect 1436 9479 1492 9535
rect 1560 9479 1616 9535
rect 1684 9479 1740 9535
rect 1808 9479 1864 9535
rect 1436 9355 1492 9411
rect 1560 9355 1616 9411
rect 1684 9355 1740 9411
rect 1808 9355 1864 9411
rect 1436 9231 1492 9287
rect 1560 9231 1616 9287
rect 1684 9231 1740 9287
rect 1808 9231 1864 9287
rect 1436 9107 1492 9163
rect 1560 9107 1616 9163
rect 1684 9107 1740 9163
rect 1808 9107 1864 9163
rect 1436 8983 1492 9039
rect 1560 8983 1616 9039
rect 1684 8983 1740 9039
rect 1808 8983 1864 9039
rect 1436 8859 1492 8915
rect 1560 8859 1616 8915
rect 1684 8859 1740 8915
rect 1808 8859 1864 8915
rect 1436 8735 1492 8791
rect 1560 8735 1616 8791
rect 1684 8735 1740 8791
rect 1808 8735 1864 8791
rect 1436 8611 1492 8667
rect 1560 8611 1616 8667
rect 1684 8611 1740 8667
rect 1808 8611 1864 8667
rect 1436 8487 1492 8543
rect 1560 8487 1616 8543
rect 1684 8487 1740 8543
rect 1808 8487 1864 8543
rect 1436 8363 1492 8419
rect 1560 8363 1616 8419
rect 1684 8363 1740 8419
rect 1808 8363 1864 8419
rect 1436 8239 1492 8295
rect 1560 8239 1616 8295
rect 1684 8239 1740 8295
rect 1808 8239 1864 8295
rect 1436 8115 1492 8171
rect 1560 8115 1616 8171
rect 1684 8115 1740 8171
rect 1808 8115 1864 8171
rect 1436 7991 1492 8047
rect 1560 7991 1616 8047
rect 1684 7991 1740 8047
rect 1808 7991 1864 8047
rect 1436 7867 1492 7923
rect 1560 7867 1616 7923
rect 1684 7867 1740 7923
rect 1808 7867 1864 7923
rect 1436 7743 1492 7799
rect 1560 7743 1616 7799
rect 1684 7743 1740 7799
rect 1808 7743 1864 7799
rect 2572 10595 2628 10651
rect 2696 10595 2752 10651
rect 2820 10595 2876 10651
rect 2944 10595 3000 10651
rect 2572 10471 2628 10527
rect 2696 10471 2752 10527
rect 2820 10471 2876 10527
rect 2944 10471 3000 10527
rect 2572 10347 2628 10403
rect 2696 10347 2752 10403
rect 2820 10347 2876 10403
rect 2944 10347 3000 10403
rect 2572 10223 2628 10279
rect 2696 10223 2752 10279
rect 2820 10223 2876 10279
rect 2944 10223 3000 10279
rect 2572 10099 2628 10155
rect 2696 10099 2752 10155
rect 2820 10099 2876 10155
rect 2944 10099 3000 10155
rect 2572 9975 2628 10031
rect 2696 9975 2752 10031
rect 2820 9975 2876 10031
rect 2944 9975 3000 10031
rect 2572 9851 2628 9907
rect 2696 9851 2752 9907
rect 2820 9851 2876 9907
rect 2944 9851 3000 9907
rect 2572 9727 2628 9783
rect 2696 9727 2752 9783
rect 2820 9727 2876 9783
rect 2944 9727 3000 9783
rect 2572 9603 2628 9659
rect 2696 9603 2752 9659
rect 2820 9603 2876 9659
rect 2944 9603 3000 9659
rect 2572 9479 2628 9535
rect 2696 9479 2752 9535
rect 2820 9479 2876 9535
rect 2944 9479 3000 9535
rect 2572 9355 2628 9411
rect 2696 9355 2752 9411
rect 2820 9355 2876 9411
rect 2944 9355 3000 9411
rect 2572 9231 2628 9287
rect 2696 9231 2752 9287
rect 2820 9231 2876 9287
rect 2944 9231 3000 9287
rect 2572 9107 2628 9163
rect 2696 9107 2752 9163
rect 2820 9107 2876 9163
rect 2944 9107 3000 9163
rect 2572 8983 2628 9039
rect 2696 8983 2752 9039
rect 2820 8983 2876 9039
rect 2944 8983 3000 9039
rect 2572 8859 2628 8915
rect 2696 8859 2752 8915
rect 2820 8859 2876 8915
rect 2944 8859 3000 8915
rect 2572 8735 2628 8791
rect 2696 8735 2752 8791
rect 2820 8735 2876 8791
rect 2944 8735 3000 8791
rect 2572 8611 2628 8667
rect 2696 8611 2752 8667
rect 2820 8611 2876 8667
rect 2944 8611 3000 8667
rect 2572 8487 2628 8543
rect 2696 8487 2752 8543
rect 2820 8487 2876 8543
rect 2944 8487 3000 8543
rect 2572 8363 2628 8419
rect 2696 8363 2752 8419
rect 2820 8363 2876 8419
rect 2944 8363 3000 8419
rect 2572 8239 2628 8295
rect 2696 8239 2752 8295
rect 2820 8239 2876 8295
rect 2944 8239 3000 8295
rect 2572 8115 2628 8171
rect 2696 8115 2752 8171
rect 2820 8115 2876 8171
rect 2944 8115 3000 8171
rect 2572 7991 2628 8047
rect 2696 7991 2752 8047
rect 2820 7991 2876 8047
rect 2944 7991 3000 8047
rect 2572 7867 2628 7923
rect 2696 7867 2752 7923
rect 2820 7867 2876 7923
rect 2944 7867 3000 7923
rect 2572 7743 2628 7799
rect 2696 7743 2752 7799
rect 2820 7743 2876 7799
rect 2944 7743 3000 7799
rect 4844 10595 4900 10651
rect 4968 10595 5024 10651
rect 5092 10595 5148 10651
rect 5216 10595 5272 10651
rect 4844 10471 4900 10527
rect 4968 10471 5024 10527
rect 5092 10471 5148 10527
rect 5216 10471 5272 10527
rect 4844 10347 4900 10403
rect 4968 10347 5024 10403
rect 5092 10347 5148 10403
rect 5216 10347 5272 10403
rect 4844 10223 4900 10279
rect 4968 10223 5024 10279
rect 5092 10223 5148 10279
rect 5216 10223 5272 10279
rect 4844 10099 4900 10155
rect 4968 10099 5024 10155
rect 5092 10099 5148 10155
rect 5216 10099 5272 10155
rect 4844 9975 4900 10031
rect 4968 9975 5024 10031
rect 5092 9975 5148 10031
rect 5216 9975 5272 10031
rect 4844 9851 4900 9907
rect 4968 9851 5024 9907
rect 5092 9851 5148 9907
rect 5216 9851 5272 9907
rect 4844 9727 4900 9783
rect 4968 9727 5024 9783
rect 5092 9727 5148 9783
rect 5216 9727 5272 9783
rect 4844 9603 4900 9659
rect 4968 9603 5024 9659
rect 5092 9603 5148 9659
rect 5216 9603 5272 9659
rect 4844 9479 4900 9535
rect 4968 9479 5024 9535
rect 5092 9479 5148 9535
rect 5216 9479 5272 9535
rect 4844 9355 4900 9411
rect 4968 9355 5024 9411
rect 5092 9355 5148 9411
rect 5216 9355 5272 9411
rect 4844 9231 4900 9287
rect 4968 9231 5024 9287
rect 5092 9231 5148 9287
rect 5216 9231 5272 9287
rect 4844 9107 4900 9163
rect 4968 9107 5024 9163
rect 5092 9107 5148 9163
rect 5216 9107 5272 9163
rect 4844 8983 4900 9039
rect 4968 8983 5024 9039
rect 5092 8983 5148 9039
rect 5216 8983 5272 9039
rect 4844 8859 4900 8915
rect 4968 8859 5024 8915
rect 5092 8859 5148 8915
rect 5216 8859 5272 8915
rect 4844 8735 4900 8791
rect 4968 8735 5024 8791
rect 5092 8735 5148 8791
rect 5216 8735 5272 8791
rect 4844 8611 4900 8667
rect 4968 8611 5024 8667
rect 5092 8611 5148 8667
rect 5216 8611 5272 8667
rect 4844 8487 4900 8543
rect 4968 8487 5024 8543
rect 5092 8487 5148 8543
rect 5216 8487 5272 8543
rect 4844 8363 4900 8419
rect 4968 8363 5024 8419
rect 5092 8363 5148 8419
rect 5216 8363 5272 8419
rect 4844 8239 4900 8295
rect 4968 8239 5024 8295
rect 5092 8239 5148 8295
rect 5216 8239 5272 8295
rect 4844 8115 4900 8171
rect 4968 8115 5024 8171
rect 5092 8115 5148 8171
rect 5216 8115 5272 8171
rect 4844 7991 4900 8047
rect 4968 7991 5024 8047
rect 5092 7991 5148 8047
rect 5216 7991 5272 8047
rect 4844 7867 4900 7923
rect 4968 7867 5024 7923
rect 5092 7867 5148 7923
rect 5216 7867 5272 7923
rect 4844 7743 4900 7799
rect 4968 7743 5024 7799
rect 5092 7743 5148 7799
rect 5216 7743 5272 7799
rect 7137 10595 7193 10651
rect 7261 10595 7317 10651
rect 7385 10595 7441 10651
rect 7137 10471 7193 10527
rect 7261 10471 7317 10527
rect 7385 10471 7441 10527
rect 7137 10347 7193 10403
rect 7261 10347 7317 10403
rect 7385 10347 7441 10403
rect 7137 10223 7193 10279
rect 7261 10223 7317 10279
rect 7385 10223 7441 10279
rect 7137 10099 7193 10155
rect 7261 10099 7317 10155
rect 7385 10099 7441 10155
rect 7137 9975 7193 10031
rect 7261 9975 7317 10031
rect 7385 9975 7441 10031
rect 7137 9851 7193 9907
rect 7261 9851 7317 9907
rect 7385 9851 7441 9907
rect 7137 9727 7193 9783
rect 7261 9727 7317 9783
rect 7385 9727 7441 9783
rect 7137 9603 7193 9659
rect 7261 9603 7317 9659
rect 7385 9603 7441 9659
rect 7137 9479 7193 9535
rect 7261 9479 7317 9535
rect 7385 9479 7441 9535
rect 7137 9355 7193 9411
rect 7261 9355 7317 9411
rect 7385 9355 7441 9411
rect 7137 9231 7193 9287
rect 7261 9231 7317 9287
rect 7385 9231 7441 9287
rect 7137 9107 7193 9163
rect 7261 9107 7317 9163
rect 7385 9107 7441 9163
rect 7137 8983 7193 9039
rect 7261 8983 7317 9039
rect 7385 8983 7441 9039
rect 7137 8859 7193 8915
rect 7261 8859 7317 8915
rect 7385 8859 7441 8915
rect 7137 8735 7193 8791
rect 7261 8735 7317 8791
rect 7385 8735 7441 8791
rect 7137 8611 7193 8667
rect 7261 8611 7317 8667
rect 7385 8611 7441 8667
rect 7137 8487 7193 8543
rect 7261 8487 7317 8543
rect 7385 8487 7441 8543
rect 7137 8363 7193 8419
rect 7261 8363 7317 8419
rect 7385 8363 7441 8419
rect 7137 8239 7193 8295
rect 7261 8239 7317 8295
rect 7385 8239 7441 8295
rect 7137 8115 7193 8171
rect 7261 8115 7317 8171
rect 7385 8115 7441 8171
rect 7137 7991 7193 8047
rect 7261 7991 7317 8047
rect 7385 7991 7441 8047
rect 7137 7867 7193 7923
rect 7261 7867 7317 7923
rect 7385 7867 7441 7923
rect 7137 7743 7193 7799
rect 7261 7743 7317 7799
rect 7385 7743 7441 7799
rect 7623 10595 7679 10651
rect 7747 10595 7803 10651
rect 7871 10595 7927 10651
rect 7623 10471 7679 10527
rect 7747 10471 7803 10527
rect 7871 10471 7927 10527
rect 7623 10347 7679 10403
rect 7747 10347 7803 10403
rect 7871 10347 7927 10403
rect 7623 10223 7679 10279
rect 7747 10223 7803 10279
rect 7871 10223 7927 10279
rect 7623 10099 7679 10155
rect 7747 10099 7803 10155
rect 7871 10099 7927 10155
rect 7623 9975 7679 10031
rect 7747 9975 7803 10031
rect 7871 9975 7927 10031
rect 7623 9851 7679 9907
rect 7747 9851 7803 9907
rect 7871 9851 7927 9907
rect 7623 9727 7679 9783
rect 7747 9727 7803 9783
rect 7871 9727 7927 9783
rect 7623 9603 7679 9659
rect 7747 9603 7803 9659
rect 7871 9603 7927 9659
rect 7623 9479 7679 9535
rect 7747 9479 7803 9535
rect 7871 9479 7927 9535
rect 7623 9355 7679 9411
rect 7747 9355 7803 9411
rect 7871 9355 7927 9411
rect 7623 9231 7679 9287
rect 7747 9231 7803 9287
rect 7871 9231 7927 9287
rect 7623 9107 7679 9163
rect 7747 9107 7803 9163
rect 7871 9107 7927 9163
rect 7623 8983 7679 9039
rect 7747 8983 7803 9039
rect 7871 8983 7927 9039
rect 7623 8859 7679 8915
rect 7747 8859 7803 8915
rect 7871 8859 7927 8915
rect 7623 8735 7679 8791
rect 7747 8735 7803 8791
rect 7871 8735 7927 8791
rect 7623 8611 7679 8667
rect 7747 8611 7803 8667
rect 7871 8611 7927 8667
rect 7623 8487 7679 8543
rect 7747 8487 7803 8543
rect 7871 8487 7927 8543
rect 7623 8363 7679 8419
rect 7747 8363 7803 8419
rect 7871 8363 7927 8419
rect 7623 8239 7679 8295
rect 7747 8239 7803 8295
rect 7871 8239 7927 8295
rect 7623 8115 7679 8171
rect 7747 8115 7803 8171
rect 7871 8115 7927 8171
rect 7623 7991 7679 8047
rect 7747 7991 7803 8047
rect 7871 7991 7927 8047
rect 7623 7867 7679 7923
rect 7747 7867 7803 7923
rect 7871 7867 7927 7923
rect 7623 7743 7679 7799
rect 7747 7743 7803 7799
rect 7871 7743 7927 7799
rect 9792 10595 9848 10651
rect 9916 10595 9972 10651
rect 10040 10595 10096 10651
rect 10164 10595 10220 10651
rect 9792 10471 9848 10527
rect 9916 10471 9972 10527
rect 10040 10471 10096 10527
rect 10164 10471 10220 10527
rect 9792 10347 9848 10403
rect 9916 10347 9972 10403
rect 10040 10347 10096 10403
rect 10164 10347 10220 10403
rect 9792 10223 9848 10279
rect 9916 10223 9972 10279
rect 10040 10223 10096 10279
rect 10164 10223 10220 10279
rect 9792 10099 9848 10155
rect 9916 10099 9972 10155
rect 10040 10099 10096 10155
rect 10164 10099 10220 10155
rect 9792 9975 9848 10031
rect 9916 9975 9972 10031
rect 10040 9975 10096 10031
rect 10164 9975 10220 10031
rect 9792 9851 9848 9907
rect 9916 9851 9972 9907
rect 10040 9851 10096 9907
rect 10164 9851 10220 9907
rect 9792 9727 9848 9783
rect 9916 9727 9972 9783
rect 10040 9727 10096 9783
rect 10164 9727 10220 9783
rect 9792 9603 9848 9659
rect 9916 9603 9972 9659
rect 10040 9603 10096 9659
rect 10164 9603 10220 9659
rect 9792 9479 9848 9535
rect 9916 9479 9972 9535
rect 10040 9479 10096 9535
rect 10164 9479 10220 9535
rect 9792 9355 9848 9411
rect 9916 9355 9972 9411
rect 10040 9355 10096 9411
rect 10164 9355 10220 9411
rect 9792 9231 9848 9287
rect 9916 9231 9972 9287
rect 10040 9231 10096 9287
rect 10164 9231 10220 9287
rect 9792 9107 9848 9163
rect 9916 9107 9972 9163
rect 10040 9107 10096 9163
rect 10164 9107 10220 9163
rect 9792 8983 9848 9039
rect 9916 8983 9972 9039
rect 10040 8983 10096 9039
rect 10164 8983 10220 9039
rect 9792 8859 9848 8915
rect 9916 8859 9972 8915
rect 10040 8859 10096 8915
rect 10164 8859 10220 8915
rect 9792 8735 9848 8791
rect 9916 8735 9972 8791
rect 10040 8735 10096 8791
rect 10164 8735 10220 8791
rect 9792 8611 9848 8667
rect 9916 8611 9972 8667
rect 10040 8611 10096 8667
rect 10164 8611 10220 8667
rect 9792 8487 9848 8543
rect 9916 8487 9972 8543
rect 10040 8487 10096 8543
rect 10164 8487 10220 8543
rect 9792 8363 9848 8419
rect 9916 8363 9972 8419
rect 10040 8363 10096 8419
rect 10164 8363 10220 8419
rect 9792 8239 9848 8295
rect 9916 8239 9972 8295
rect 10040 8239 10096 8295
rect 10164 8239 10220 8295
rect 9792 8115 9848 8171
rect 9916 8115 9972 8171
rect 10040 8115 10096 8171
rect 10164 8115 10220 8171
rect 9792 7991 9848 8047
rect 9916 7991 9972 8047
rect 10040 7991 10096 8047
rect 10164 7991 10220 8047
rect 9792 7867 9848 7923
rect 9916 7867 9972 7923
rect 10040 7867 10096 7923
rect 10164 7867 10220 7923
rect 9792 7743 9848 7799
rect 9916 7743 9972 7799
rect 10040 7743 10096 7799
rect 10164 7743 10220 7799
rect 12064 10595 12120 10651
rect 12188 10595 12244 10651
rect 12312 10595 12368 10651
rect 12436 10595 12492 10651
rect 12064 10471 12120 10527
rect 12188 10471 12244 10527
rect 12312 10471 12368 10527
rect 12436 10471 12492 10527
rect 12064 10347 12120 10403
rect 12188 10347 12244 10403
rect 12312 10347 12368 10403
rect 12436 10347 12492 10403
rect 12064 10223 12120 10279
rect 12188 10223 12244 10279
rect 12312 10223 12368 10279
rect 12436 10223 12492 10279
rect 12064 10099 12120 10155
rect 12188 10099 12244 10155
rect 12312 10099 12368 10155
rect 12436 10099 12492 10155
rect 12064 9975 12120 10031
rect 12188 9975 12244 10031
rect 12312 9975 12368 10031
rect 12436 9975 12492 10031
rect 12064 9851 12120 9907
rect 12188 9851 12244 9907
rect 12312 9851 12368 9907
rect 12436 9851 12492 9907
rect 12064 9727 12120 9783
rect 12188 9727 12244 9783
rect 12312 9727 12368 9783
rect 12436 9727 12492 9783
rect 12064 9603 12120 9659
rect 12188 9603 12244 9659
rect 12312 9603 12368 9659
rect 12436 9603 12492 9659
rect 12064 9479 12120 9535
rect 12188 9479 12244 9535
rect 12312 9479 12368 9535
rect 12436 9479 12492 9535
rect 12064 9355 12120 9411
rect 12188 9355 12244 9411
rect 12312 9355 12368 9411
rect 12436 9355 12492 9411
rect 12064 9231 12120 9287
rect 12188 9231 12244 9287
rect 12312 9231 12368 9287
rect 12436 9231 12492 9287
rect 12064 9107 12120 9163
rect 12188 9107 12244 9163
rect 12312 9107 12368 9163
rect 12436 9107 12492 9163
rect 12064 8983 12120 9039
rect 12188 8983 12244 9039
rect 12312 8983 12368 9039
rect 12436 8983 12492 9039
rect 12064 8859 12120 8915
rect 12188 8859 12244 8915
rect 12312 8859 12368 8915
rect 12436 8859 12492 8915
rect 12064 8735 12120 8791
rect 12188 8735 12244 8791
rect 12312 8735 12368 8791
rect 12436 8735 12492 8791
rect 12064 8611 12120 8667
rect 12188 8611 12244 8667
rect 12312 8611 12368 8667
rect 12436 8611 12492 8667
rect 12064 8487 12120 8543
rect 12188 8487 12244 8543
rect 12312 8487 12368 8543
rect 12436 8487 12492 8543
rect 12064 8363 12120 8419
rect 12188 8363 12244 8419
rect 12312 8363 12368 8419
rect 12436 8363 12492 8419
rect 12064 8239 12120 8295
rect 12188 8239 12244 8295
rect 12312 8239 12368 8295
rect 12436 8239 12492 8295
rect 12064 8115 12120 8171
rect 12188 8115 12244 8171
rect 12312 8115 12368 8171
rect 12436 8115 12492 8171
rect 12064 7991 12120 8047
rect 12188 7991 12244 8047
rect 12312 7991 12368 8047
rect 12436 7991 12492 8047
rect 12064 7867 12120 7923
rect 12188 7867 12244 7923
rect 12312 7867 12368 7923
rect 12436 7867 12492 7923
rect 12064 7743 12120 7799
rect 12188 7743 12244 7799
rect 12312 7743 12368 7799
rect 12436 7743 12492 7799
rect 13200 10595 13256 10651
rect 13324 10595 13380 10651
rect 13448 10595 13504 10651
rect 13572 10595 13628 10651
rect 13200 10471 13256 10527
rect 13324 10471 13380 10527
rect 13448 10471 13504 10527
rect 13572 10471 13628 10527
rect 13200 10347 13256 10403
rect 13324 10347 13380 10403
rect 13448 10347 13504 10403
rect 13572 10347 13628 10403
rect 13200 10223 13256 10279
rect 13324 10223 13380 10279
rect 13448 10223 13504 10279
rect 13572 10223 13628 10279
rect 13200 10099 13256 10155
rect 13324 10099 13380 10155
rect 13448 10099 13504 10155
rect 13572 10099 13628 10155
rect 13200 9975 13256 10031
rect 13324 9975 13380 10031
rect 13448 9975 13504 10031
rect 13572 9975 13628 10031
rect 13200 9851 13256 9907
rect 13324 9851 13380 9907
rect 13448 9851 13504 9907
rect 13572 9851 13628 9907
rect 13200 9727 13256 9783
rect 13324 9727 13380 9783
rect 13448 9727 13504 9783
rect 13572 9727 13628 9783
rect 13200 9603 13256 9659
rect 13324 9603 13380 9659
rect 13448 9603 13504 9659
rect 13572 9603 13628 9659
rect 13200 9479 13256 9535
rect 13324 9479 13380 9535
rect 13448 9479 13504 9535
rect 13572 9479 13628 9535
rect 13200 9355 13256 9411
rect 13324 9355 13380 9411
rect 13448 9355 13504 9411
rect 13572 9355 13628 9411
rect 13200 9231 13256 9287
rect 13324 9231 13380 9287
rect 13448 9231 13504 9287
rect 13572 9231 13628 9287
rect 13200 9107 13256 9163
rect 13324 9107 13380 9163
rect 13448 9107 13504 9163
rect 13572 9107 13628 9163
rect 13200 8983 13256 9039
rect 13324 8983 13380 9039
rect 13448 8983 13504 9039
rect 13572 8983 13628 9039
rect 13200 8859 13256 8915
rect 13324 8859 13380 8915
rect 13448 8859 13504 8915
rect 13572 8859 13628 8915
rect 13200 8735 13256 8791
rect 13324 8735 13380 8791
rect 13448 8735 13504 8791
rect 13572 8735 13628 8791
rect 13200 8611 13256 8667
rect 13324 8611 13380 8667
rect 13448 8611 13504 8667
rect 13572 8611 13628 8667
rect 13200 8487 13256 8543
rect 13324 8487 13380 8543
rect 13448 8487 13504 8543
rect 13572 8487 13628 8543
rect 13200 8363 13256 8419
rect 13324 8363 13380 8419
rect 13448 8363 13504 8419
rect 13572 8363 13628 8419
rect 13200 8239 13256 8295
rect 13324 8239 13380 8295
rect 13448 8239 13504 8295
rect 13572 8239 13628 8295
rect 13200 8115 13256 8171
rect 13324 8115 13380 8171
rect 13448 8115 13504 8171
rect 13572 8115 13628 8171
rect 13200 7991 13256 8047
rect 13324 7991 13380 8047
rect 13448 7991 13504 8047
rect 13572 7991 13628 8047
rect 13200 7867 13256 7923
rect 13324 7867 13380 7923
rect 13448 7867 13504 7923
rect 13572 7867 13628 7923
rect 13200 7743 13256 7799
rect 13324 7743 13380 7799
rect 13448 7743 13504 7799
rect 13572 7743 13628 7799
rect 1436 7395 1492 7451
rect 1560 7395 1616 7451
rect 1684 7395 1740 7451
rect 1808 7395 1864 7451
rect 1436 7271 1492 7327
rect 1560 7271 1616 7327
rect 1684 7271 1740 7327
rect 1808 7271 1864 7327
rect 1436 7147 1492 7203
rect 1560 7147 1616 7203
rect 1684 7147 1740 7203
rect 1808 7147 1864 7203
rect 1436 7023 1492 7079
rect 1560 7023 1616 7079
rect 1684 7023 1740 7079
rect 1808 7023 1864 7079
rect 1436 6899 1492 6955
rect 1560 6899 1616 6955
rect 1684 6899 1740 6955
rect 1808 6899 1864 6955
rect 1436 6775 1492 6831
rect 1560 6775 1616 6831
rect 1684 6775 1740 6831
rect 1808 6775 1864 6831
rect 1436 6651 1492 6707
rect 1560 6651 1616 6707
rect 1684 6651 1740 6707
rect 1808 6651 1864 6707
rect 1436 6527 1492 6583
rect 1560 6527 1616 6583
rect 1684 6527 1740 6583
rect 1808 6527 1864 6583
rect 1436 6403 1492 6459
rect 1560 6403 1616 6459
rect 1684 6403 1740 6459
rect 1808 6403 1864 6459
rect 1436 6279 1492 6335
rect 1560 6279 1616 6335
rect 1684 6279 1740 6335
rect 1808 6279 1864 6335
rect 1436 6155 1492 6211
rect 1560 6155 1616 6211
rect 1684 6155 1740 6211
rect 1808 6155 1864 6211
rect 1436 6031 1492 6087
rect 1560 6031 1616 6087
rect 1684 6031 1740 6087
rect 1808 6031 1864 6087
rect 1436 5907 1492 5963
rect 1560 5907 1616 5963
rect 1684 5907 1740 5963
rect 1808 5907 1864 5963
rect 1436 5783 1492 5839
rect 1560 5783 1616 5839
rect 1684 5783 1740 5839
rect 1808 5783 1864 5839
rect 1436 5659 1492 5715
rect 1560 5659 1616 5715
rect 1684 5659 1740 5715
rect 1808 5659 1864 5715
rect 1436 5535 1492 5591
rect 1560 5535 1616 5591
rect 1684 5535 1740 5591
rect 1808 5535 1864 5591
rect 1436 5411 1492 5467
rect 1560 5411 1616 5467
rect 1684 5411 1740 5467
rect 1808 5411 1864 5467
rect 1436 5287 1492 5343
rect 1560 5287 1616 5343
rect 1684 5287 1740 5343
rect 1808 5287 1864 5343
rect 1436 5163 1492 5219
rect 1560 5163 1616 5219
rect 1684 5163 1740 5219
rect 1808 5163 1864 5219
rect 1436 5039 1492 5095
rect 1560 5039 1616 5095
rect 1684 5039 1740 5095
rect 1808 5039 1864 5095
rect 1436 4915 1492 4971
rect 1560 4915 1616 4971
rect 1684 4915 1740 4971
rect 1808 4915 1864 4971
rect 1436 4791 1492 4847
rect 1560 4791 1616 4847
rect 1684 4791 1740 4847
rect 1808 4791 1864 4847
rect 1436 4667 1492 4723
rect 1560 4667 1616 4723
rect 1684 4667 1740 4723
rect 1808 4667 1864 4723
rect 1436 4543 1492 4599
rect 1560 4543 1616 4599
rect 1684 4543 1740 4599
rect 1808 4543 1864 4599
rect 2572 7395 2628 7451
rect 2696 7395 2752 7451
rect 2820 7395 2876 7451
rect 2944 7395 3000 7451
rect 2572 7271 2628 7327
rect 2696 7271 2752 7327
rect 2820 7271 2876 7327
rect 2944 7271 3000 7327
rect 2572 7147 2628 7203
rect 2696 7147 2752 7203
rect 2820 7147 2876 7203
rect 2944 7147 3000 7203
rect 2572 7023 2628 7079
rect 2696 7023 2752 7079
rect 2820 7023 2876 7079
rect 2944 7023 3000 7079
rect 2572 6899 2628 6955
rect 2696 6899 2752 6955
rect 2820 6899 2876 6955
rect 2944 6899 3000 6955
rect 2572 6775 2628 6831
rect 2696 6775 2752 6831
rect 2820 6775 2876 6831
rect 2944 6775 3000 6831
rect 2572 6651 2628 6707
rect 2696 6651 2752 6707
rect 2820 6651 2876 6707
rect 2944 6651 3000 6707
rect 2572 6527 2628 6583
rect 2696 6527 2752 6583
rect 2820 6527 2876 6583
rect 2944 6527 3000 6583
rect 2572 6403 2628 6459
rect 2696 6403 2752 6459
rect 2820 6403 2876 6459
rect 2944 6403 3000 6459
rect 2572 6279 2628 6335
rect 2696 6279 2752 6335
rect 2820 6279 2876 6335
rect 2944 6279 3000 6335
rect 2572 6155 2628 6211
rect 2696 6155 2752 6211
rect 2820 6155 2876 6211
rect 2944 6155 3000 6211
rect 2572 6031 2628 6087
rect 2696 6031 2752 6087
rect 2820 6031 2876 6087
rect 2944 6031 3000 6087
rect 2572 5907 2628 5963
rect 2696 5907 2752 5963
rect 2820 5907 2876 5963
rect 2944 5907 3000 5963
rect 2572 5783 2628 5839
rect 2696 5783 2752 5839
rect 2820 5783 2876 5839
rect 2944 5783 3000 5839
rect 2572 5659 2628 5715
rect 2696 5659 2752 5715
rect 2820 5659 2876 5715
rect 2944 5659 3000 5715
rect 2572 5535 2628 5591
rect 2696 5535 2752 5591
rect 2820 5535 2876 5591
rect 2944 5535 3000 5591
rect 2572 5411 2628 5467
rect 2696 5411 2752 5467
rect 2820 5411 2876 5467
rect 2944 5411 3000 5467
rect 2572 5287 2628 5343
rect 2696 5287 2752 5343
rect 2820 5287 2876 5343
rect 2944 5287 3000 5343
rect 2572 5163 2628 5219
rect 2696 5163 2752 5219
rect 2820 5163 2876 5219
rect 2944 5163 3000 5219
rect 2572 5039 2628 5095
rect 2696 5039 2752 5095
rect 2820 5039 2876 5095
rect 2944 5039 3000 5095
rect 2572 4915 2628 4971
rect 2696 4915 2752 4971
rect 2820 4915 2876 4971
rect 2944 4915 3000 4971
rect 2572 4791 2628 4847
rect 2696 4791 2752 4847
rect 2820 4791 2876 4847
rect 2944 4791 3000 4847
rect 2572 4667 2628 4723
rect 2696 4667 2752 4723
rect 2820 4667 2876 4723
rect 2944 4667 3000 4723
rect 2572 4543 2628 4599
rect 2696 4543 2752 4599
rect 2820 4543 2876 4599
rect 2944 4543 3000 4599
rect 4844 7395 4900 7451
rect 4968 7395 5024 7451
rect 5092 7395 5148 7451
rect 5216 7395 5272 7451
rect 4844 7271 4900 7327
rect 4968 7271 5024 7327
rect 5092 7271 5148 7327
rect 5216 7271 5272 7327
rect 4844 7147 4900 7203
rect 4968 7147 5024 7203
rect 5092 7147 5148 7203
rect 5216 7147 5272 7203
rect 4844 7023 4900 7079
rect 4968 7023 5024 7079
rect 5092 7023 5148 7079
rect 5216 7023 5272 7079
rect 4844 6899 4900 6955
rect 4968 6899 5024 6955
rect 5092 6899 5148 6955
rect 5216 6899 5272 6955
rect 4844 6775 4900 6831
rect 4968 6775 5024 6831
rect 5092 6775 5148 6831
rect 5216 6775 5272 6831
rect 4844 6651 4900 6707
rect 4968 6651 5024 6707
rect 5092 6651 5148 6707
rect 5216 6651 5272 6707
rect 4844 6527 4900 6583
rect 4968 6527 5024 6583
rect 5092 6527 5148 6583
rect 5216 6527 5272 6583
rect 4844 6403 4900 6459
rect 4968 6403 5024 6459
rect 5092 6403 5148 6459
rect 5216 6403 5272 6459
rect 4844 6279 4900 6335
rect 4968 6279 5024 6335
rect 5092 6279 5148 6335
rect 5216 6279 5272 6335
rect 4844 6155 4900 6211
rect 4968 6155 5024 6211
rect 5092 6155 5148 6211
rect 5216 6155 5272 6211
rect 4844 6031 4900 6087
rect 4968 6031 5024 6087
rect 5092 6031 5148 6087
rect 5216 6031 5272 6087
rect 4844 5907 4900 5963
rect 4968 5907 5024 5963
rect 5092 5907 5148 5963
rect 5216 5907 5272 5963
rect 4844 5783 4900 5839
rect 4968 5783 5024 5839
rect 5092 5783 5148 5839
rect 5216 5783 5272 5839
rect 4844 5659 4900 5715
rect 4968 5659 5024 5715
rect 5092 5659 5148 5715
rect 5216 5659 5272 5715
rect 4844 5535 4900 5591
rect 4968 5535 5024 5591
rect 5092 5535 5148 5591
rect 5216 5535 5272 5591
rect 4844 5411 4900 5467
rect 4968 5411 5024 5467
rect 5092 5411 5148 5467
rect 5216 5411 5272 5467
rect 4844 5287 4900 5343
rect 4968 5287 5024 5343
rect 5092 5287 5148 5343
rect 5216 5287 5272 5343
rect 4844 5163 4900 5219
rect 4968 5163 5024 5219
rect 5092 5163 5148 5219
rect 5216 5163 5272 5219
rect 4844 5039 4900 5095
rect 4968 5039 5024 5095
rect 5092 5039 5148 5095
rect 5216 5039 5272 5095
rect 4844 4915 4900 4971
rect 4968 4915 5024 4971
rect 5092 4915 5148 4971
rect 5216 4915 5272 4971
rect 4844 4791 4900 4847
rect 4968 4791 5024 4847
rect 5092 4791 5148 4847
rect 5216 4791 5272 4847
rect 4844 4667 4900 4723
rect 4968 4667 5024 4723
rect 5092 4667 5148 4723
rect 5216 4667 5272 4723
rect 4844 4543 4900 4599
rect 4968 4543 5024 4599
rect 5092 4543 5148 4599
rect 5216 4543 5272 4599
rect 7137 7395 7193 7451
rect 7261 7395 7317 7451
rect 7385 7395 7441 7451
rect 7137 7271 7193 7327
rect 7261 7271 7317 7327
rect 7385 7271 7441 7327
rect 7137 7147 7193 7203
rect 7261 7147 7317 7203
rect 7385 7147 7441 7203
rect 7137 7023 7193 7079
rect 7261 7023 7317 7079
rect 7385 7023 7441 7079
rect 7137 6899 7193 6955
rect 7261 6899 7317 6955
rect 7385 6899 7441 6955
rect 7137 6775 7193 6831
rect 7261 6775 7317 6831
rect 7385 6775 7441 6831
rect 7137 6651 7193 6707
rect 7261 6651 7317 6707
rect 7385 6651 7441 6707
rect 7137 6527 7193 6583
rect 7261 6527 7317 6583
rect 7385 6527 7441 6583
rect 7137 6403 7193 6459
rect 7261 6403 7317 6459
rect 7385 6403 7441 6459
rect 7137 6279 7193 6335
rect 7261 6279 7317 6335
rect 7385 6279 7441 6335
rect 7137 6155 7193 6211
rect 7261 6155 7317 6211
rect 7385 6155 7441 6211
rect 7137 6031 7193 6087
rect 7261 6031 7317 6087
rect 7385 6031 7441 6087
rect 7137 5907 7193 5963
rect 7261 5907 7317 5963
rect 7385 5907 7441 5963
rect 7137 5783 7193 5839
rect 7261 5783 7317 5839
rect 7385 5783 7441 5839
rect 7137 5659 7193 5715
rect 7261 5659 7317 5715
rect 7385 5659 7441 5715
rect 7137 5535 7193 5591
rect 7261 5535 7317 5591
rect 7385 5535 7441 5591
rect 7137 5411 7193 5467
rect 7261 5411 7317 5467
rect 7385 5411 7441 5467
rect 7137 5287 7193 5343
rect 7261 5287 7317 5343
rect 7385 5287 7441 5343
rect 7137 5163 7193 5219
rect 7261 5163 7317 5219
rect 7385 5163 7441 5219
rect 7137 5039 7193 5095
rect 7261 5039 7317 5095
rect 7385 5039 7441 5095
rect 7137 4915 7193 4971
rect 7261 4915 7317 4971
rect 7385 4915 7441 4971
rect 7137 4791 7193 4847
rect 7261 4791 7317 4847
rect 7385 4791 7441 4847
rect 7137 4667 7193 4723
rect 7261 4667 7317 4723
rect 7385 4667 7441 4723
rect 7137 4543 7193 4599
rect 7261 4543 7317 4599
rect 7385 4543 7441 4599
rect 7623 7395 7679 7451
rect 7747 7395 7803 7451
rect 7871 7395 7927 7451
rect 7623 7271 7679 7327
rect 7747 7271 7803 7327
rect 7871 7271 7927 7327
rect 7623 7147 7679 7203
rect 7747 7147 7803 7203
rect 7871 7147 7927 7203
rect 7623 7023 7679 7079
rect 7747 7023 7803 7079
rect 7871 7023 7927 7079
rect 7623 6899 7679 6955
rect 7747 6899 7803 6955
rect 7871 6899 7927 6955
rect 7623 6775 7679 6831
rect 7747 6775 7803 6831
rect 7871 6775 7927 6831
rect 7623 6651 7679 6707
rect 7747 6651 7803 6707
rect 7871 6651 7927 6707
rect 7623 6527 7679 6583
rect 7747 6527 7803 6583
rect 7871 6527 7927 6583
rect 7623 6403 7679 6459
rect 7747 6403 7803 6459
rect 7871 6403 7927 6459
rect 7623 6279 7679 6335
rect 7747 6279 7803 6335
rect 7871 6279 7927 6335
rect 7623 6155 7679 6211
rect 7747 6155 7803 6211
rect 7871 6155 7927 6211
rect 7623 6031 7679 6087
rect 7747 6031 7803 6087
rect 7871 6031 7927 6087
rect 7623 5907 7679 5963
rect 7747 5907 7803 5963
rect 7871 5907 7927 5963
rect 7623 5783 7679 5839
rect 7747 5783 7803 5839
rect 7871 5783 7927 5839
rect 7623 5659 7679 5715
rect 7747 5659 7803 5715
rect 7871 5659 7927 5715
rect 7623 5535 7679 5591
rect 7747 5535 7803 5591
rect 7871 5535 7927 5591
rect 7623 5411 7679 5467
rect 7747 5411 7803 5467
rect 7871 5411 7927 5467
rect 7623 5287 7679 5343
rect 7747 5287 7803 5343
rect 7871 5287 7927 5343
rect 7623 5163 7679 5219
rect 7747 5163 7803 5219
rect 7871 5163 7927 5219
rect 7623 5039 7679 5095
rect 7747 5039 7803 5095
rect 7871 5039 7927 5095
rect 7623 4915 7679 4971
rect 7747 4915 7803 4971
rect 7871 4915 7927 4971
rect 7623 4791 7679 4847
rect 7747 4791 7803 4847
rect 7871 4791 7927 4847
rect 7623 4667 7679 4723
rect 7747 4667 7803 4723
rect 7871 4667 7927 4723
rect 7623 4543 7679 4599
rect 7747 4543 7803 4599
rect 7871 4543 7927 4599
rect 9792 7395 9848 7451
rect 9916 7395 9972 7451
rect 10040 7395 10096 7451
rect 10164 7395 10220 7451
rect 9792 7271 9848 7327
rect 9916 7271 9972 7327
rect 10040 7271 10096 7327
rect 10164 7271 10220 7327
rect 9792 7147 9848 7203
rect 9916 7147 9972 7203
rect 10040 7147 10096 7203
rect 10164 7147 10220 7203
rect 9792 7023 9848 7079
rect 9916 7023 9972 7079
rect 10040 7023 10096 7079
rect 10164 7023 10220 7079
rect 9792 6899 9848 6955
rect 9916 6899 9972 6955
rect 10040 6899 10096 6955
rect 10164 6899 10220 6955
rect 9792 6775 9848 6831
rect 9916 6775 9972 6831
rect 10040 6775 10096 6831
rect 10164 6775 10220 6831
rect 9792 6651 9848 6707
rect 9916 6651 9972 6707
rect 10040 6651 10096 6707
rect 10164 6651 10220 6707
rect 9792 6527 9848 6583
rect 9916 6527 9972 6583
rect 10040 6527 10096 6583
rect 10164 6527 10220 6583
rect 9792 6403 9848 6459
rect 9916 6403 9972 6459
rect 10040 6403 10096 6459
rect 10164 6403 10220 6459
rect 9792 6279 9848 6335
rect 9916 6279 9972 6335
rect 10040 6279 10096 6335
rect 10164 6279 10220 6335
rect 9792 6155 9848 6211
rect 9916 6155 9972 6211
rect 10040 6155 10096 6211
rect 10164 6155 10220 6211
rect 9792 6031 9848 6087
rect 9916 6031 9972 6087
rect 10040 6031 10096 6087
rect 10164 6031 10220 6087
rect 9792 5907 9848 5963
rect 9916 5907 9972 5963
rect 10040 5907 10096 5963
rect 10164 5907 10220 5963
rect 9792 5783 9848 5839
rect 9916 5783 9972 5839
rect 10040 5783 10096 5839
rect 10164 5783 10220 5839
rect 9792 5659 9848 5715
rect 9916 5659 9972 5715
rect 10040 5659 10096 5715
rect 10164 5659 10220 5715
rect 9792 5535 9848 5591
rect 9916 5535 9972 5591
rect 10040 5535 10096 5591
rect 10164 5535 10220 5591
rect 9792 5411 9848 5467
rect 9916 5411 9972 5467
rect 10040 5411 10096 5467
rect 10164 5411 10220 5467
rect 9792 5287 9848 5343
rect 9916 5287 9972 5343
rect 10040 5287 10096 5343
rect 10164 5287 10220 5343
rect 9792 5163 9848 5219
rect 9916 5163 9972 5219
rect 10040 5163 10096 5219
rect 10164 5163 10220 5219
rect 9792 5039 9848 5095
rect 9916 5039 9972 5095
rect 10040 5039 10096 5095
rect 10164 5039 10220 5095
rect 9792 4915 9848 4971
rect 9916 4915 9972 4971
rect 10040 4915 10096 4971
rect 10164 4915 10220 4971
rect 9792 4791 9848 4847
rect 9916 4791 9972 4847
rect 10040 4791 10096 4847
rect 10164 4791 10220 4847
rect 9792 4667 9848 4723
rect 9916 4667 9972 4723
rect 10040 4667 10096 4723
rect 10164 4667 10220 4723
rect 9792 4543 9848 4599
rect 9916 4543 9972 4599
rect 10040 4543 10096 4599
rect 10164 4543 10220 4599
rect 12064 7395 12120 7451
rect 12188 7395 12244 7451
rect 12312 7395 12368 7451
rect 12436 7395 12492 7451
rect 12064 7271 12120 7327
rect 12188 7271 12244 7327
rect 12312 7271 12368 7327
rect 12436 7271 12492 7327
rect 12064 7147 12120 7203
rect 12188 7147 12244 7203
rect 12312 7147 12368 7203
rect 12436 7147 12492 7203
rect 12064 7023 12120 7079
rect 12188 7023 12244 7079
rect 12312 7023 12368 7079
rect 12436 7023 12492 7079
rect 12064 6899 12120 6955
rect 12188 6899 12244 6955
rect 12312 6899 12368 6955
rect 12436 6899 12492 6955
rect 12064 6775 12120 6831
rect 12188 6775 12244 6831
rect 12312 6775 12368 6831
rect 12436 6775 12492 6831
rect 12064 6651 12120 6707
rect 12188 6651 12244 6707
rect 12312 6651 12368 6707
rect 12436 6651 12492 6707
rect 12064 6527 12120 6583
rect 12188 6527 12244 6583
rect 12312 6527 12368 6583
rect 12436 6527 12492 6583
rect 12064 6403 12120 6459
rect 12188 6403 12244 6459
rect 12312 6403 12368 6459
rect 12436 6403 12492 6459
rect 12064 6279 12120 6335
rect 12188 6279 12244 6335
rect 12312 6279 12368 6335
rect 12436 6279 12492 6335
rect 12064 6155 12120 6211
rect 12188 6155 12244 6211
rect 12312 6155 12368 6211
rect 12436 6155 12492 6211
rect 12064 6031 12120 6087
rect 12188 6031 12244 6087
rect 12312 6031 12368 6087
rect 12436 6031 12492 6087
rect 12064 5907 12120 5963
rect 12188 5907 12244 5963
rect 12312 5907 12368 5963
rect 12436 5907 12492 5963
rect 12064 5783 12120 5839
rect 12188 5783 12244 5839
rect 12312 5783 12368 5839
rect 12436 5783 12492 5839
rect 12064 5659 12120 5715
rect 12188 5659 12244 5715
rect 12312 5659 12368 5715
rect 12436 5659 12492 5715
rect 12064 5535 12120 5591
rect 12188 5535 12244 5591
rect 12312 5535 12368 5591
rect 12436 5535 12492 5591
rect 12064 5411 12120 5467
rect 12188 5411 12244 5467
rect 12312 5411 12368 5467
rect 12436 5411 12492 5467
rect 12064 5287 12120 5343
rect 12188 5287 12244 5343
rect 12312 5287 12368 5343
rect 12436 5287 12492 5343
rect 12064 5163 12120 5219
rect 12188 5163 12244 5219
rect 12312 5163 12368 5219
rect 12436 5163 12492 5219
rect 12064 5039 12120 5095
rect 12188 5039 12244 5095
rect 12312 5039 12368 5095
rect 12436 5039 12492 5095
rect 12064 4915 12120 4971
rect 12188 4915 12244 4971
rect 12312 4915 12368 4971
rect 12436 4915 12492 4971
rect 12064 4791 12120 4847
rect 12188 4791 12244 4847
rect 12312 4791 12368 4847
rect 12436 4791 12492 4847
rect 12064 4667 12120 4723
rect 12188 4667 12244 4723
rect 12312 4667 12368 4723
rect 12436 4667 12492 4723
rect 12064 4543 12120 4599
rect 12188 4543 12244 4599
rect 12312 4543 12368 4599
rect 12436 4543 12492 4599
rect 13200 7395 13256 7451
rect 13324 7395 13380 7451
rect 13448 7395 13504 7451
rect 13572 7395 13628 7451
rect 13200 7271 13256 7327
rect 13324 7271 13380 7327
rect 13448 7271 13504 7327
rect 13572 7271 13628 7327
rect 13200 7147 13256 7203
rect 13324 7147 13380 7203
rect 13448 7147 13504 7203
rect 13572 7147 13628 7203
rect 13200 7023 13256 7079
rect 13324 7023 13380 7079
rect 13448 7023 13504 7079
rect 13572 7023 13628 7079
rect 13200 6899 13256 6955
rect 13324 6899 13380 6955
rect 13448 6899 13504 6955
rect 13572 6899 13628 6955
rect 13200 6775 13256 6831
rect 13324 6775 13380 6831
rect 13448 6775 13504 6831
rect 13572 6775 13628 6831
rect 13200 6651 13256 6707
rect 13324 6651 13380 6707
rect 13448 6651 13504 6707
rect 13572 6651 13628 6707
rect 13200 6527 13256 6583
rect 13324 6527 13380 6583
rect 13448 6527 13504 6583
rect 13572 6527 13628 6583
rect 13200 6403 13256 6459
rect 13324 6403 13380 6459
rect 13448 6403 13504 6459
rect 13572 6403 13628 6459
rect 13200 6279 13256 6335
rect 13324 6279 13380 6335
rect 13448 6279 13504 6335
rect 13572 6279 13628 6335
rect 13200 6155 13256 6211
rect 13324 6155 13380 6211
rect 13448 6155 13504 6211
rect 13572 6155 13628 6211
rect 13200 6031 13256 6087
rect 13324 6031 13380 6087
rect 13448 6031 13504 6087
rect 13572 6031 13628 6087
rect 13200 5907 13256 5963
rect 13324 5907 13380 5963
rect 13448 5907 13504 5963
rect 13572 5907 13628 5963
rect 13200 5783 13256 5839
rect 13324 5783 13380 5839
rect 13448 5783 13504 5839
rect 13572 5783 13628 5839
rect 13200 5659 13256 5715
rect 13324 5659 13380 5715
rect 13448 5659 13504 5715
rect 13572 5659 13628 5715
rect 13200 5535 13256 5591
rect 13324 5535 13380 5591
rect 13448 5535 13504 5591
rect 13572 5535 13628 5591
rect 13200 5411 13256 5467
rect 13324 5411 13380 5467
rect 13448 5411 13504 5467
rect 13572 5411 13628 5467
rect 13200 5287 13256 5343
rect 13324 5287 13380 5343
rect 13448 5287 13504 5343
rect 13572 5287 13628 5343
rect 13200 5163 13256 5219
rect 13324 5163 13380 5219
rect 13448 5163 13504 5219
rect 13572 5163 13628 5219
rect 13200 5039 13256 5095
rect 13324 5039 13380 5095
rect 13448 5039 13504 5095
rect 13572 5039 13628 5095
rect 13200 4915 13256 4971
rect 13324 4915 13380 4971
rect 13448 4915 13504 4971
rect 13572 4915 13628 4971
rect 13200 4791 13256 4847
rect 13324 4791 13380 4847
rect 13448 4791 13504 4847
rect 13572 4791 13628 4847
rect 13200 4667 13256 4723
rect 13324 4667 13380 4723
rect 13448 4667 13504 4723
rect 13572 4667 13628 4723
rect 13200 4543 13256 4599
rect 13324 4543 13380 4599
rect 13448 4543 13504 4599
rect 13572 4543 13628 4599
rect 1436 4195 1492 4251
rect 1560 4195 1616 4251
rect 1684 4195 1740 4251
rect 1808 4195 1864 4251
rect 1436 4071 1492 4127
rect 1560 4071 1616 4127
rect 1684 4071 1740 4127
rect 1808 4071 1864 4127
rect 1436 3947 1492 4003
rect 1560 3947 1616 4003
rect 1684 3947 1740 4003
rect 1808 3947 1864 4003
rect 1436 3823 1492 3879
rect 1560 3823 1616 3879
rect 1684 3823 1740 3879
rect 1808 3823 1864 3879
rect 1436 3699 1492 3755
rect 1560 3699 1616 3755
rect 1684 3699 1740 3755
rect 1808 3699 1864 3755
rect 1436 3575 1492 3631
rect 1560 3575 1616 3631
rect 1684 3575 1740 3631
rect 1808 3575 1864 3631
rect 1436 3451 1492 3507
rect 1560 3451 1616 3507
rect 1684 3451 1740 3507
rect 1808 3451 1864 3507
rect 1436 3327 1492 3383
rect 1560 3327 1616 3383
rect 1684 3327 1740 3383
rect 1808 3327 1864 3383
rect 1436 3203 1492 3259
rect 1560 3203 1616 3259
rect 1684 3203 1740 3259
rect 1808 3203 1864 3259
rect 1436 3079 1492 3135
rect 1560 3079 1616 3135
rect 1684 3079 1740 3135
rect 1808 3079 1864 3135
rect 1436 2955 1492 3011
rect 1560 2955 1616 3011
rect 1684 2955 1740 3011
rect 1808 2955 1864 3011
rect 1436 2831 1492 2887
rect 1560 2831 1616 2887
rect 1684 2831 1740 2887
rect 1808 2831 1864 2887
rect 1436 2707 1492 2763
rect 1560 2707 1616 2763
rect 1684 2707 1740 2763
rect 1808 2707 1864 2763
rect 1436 2583 1492 2639
rect 1560 2583 1616 2639
rect 1684 2583 1740 2639
rect 1808 2583 1864 2639
rect 1436 2459 1492 2515
rect 1560 2459 1616 2515
rect 1684 2459 1740 2515
rect 1808 2459 1864 2515
rect 1436 2335 1492 2391
rect 1560 2335 1616 2391
rect 1684 2335 1740 2391
rect 1808 2335 1864 2391
rect 1436 2211 1492 2267
rect 1560 2211 1616 2267
rect 1684 2211 1740 2267
rect 1808 2211 1864 2267
rect 1436 2087 1492 2143
rect 1560 2087 1616 2143
rect 1684 2087 1740 2143
rect 1808 2087 1864 2143
rect 1436 1963 1492 2019
rect 1560 1963 1616 2019
rect 1684 1963 1740 2019
rect 1808 1963 1864 2019
rect 1436 1839 1492 1895
rect 1560 1839 1616 1895
rect 1684 1839 1740 1895
rect 1808 1839 1864 1895
rect 1436 1715 1492 1771
rect 1560 1715 1616 1771
rect 1684 1715 1740 1771
rect 1808 1715 1864 1771
rect 1436 1591 1492 1647
rect 1560 1591 1616 1647
rect 1684 1591 1740 1647
rect 1808 1591 1864 1647
rect 1436 1467 1492 1523
rect 1560 1467 1616 1523
rect 1684 1467 1740 1523
rect 1808 1467 1864 1523
rect 1436 1343 1492 1399
rect 1560 1343 1616 1399
rect 1684 1343 1740 1399
rect 1808 1343 1864 1399
rect 2572 4195 2628 4251
rect 2696 4195 2752 4251
rect 2820 4195 2876 4251
rect 2944 4195 3000 4251
rect 2572 4071 2628 4127
rect 2696 4071 2752 4127
rect 2820 4071 2876 4127
rect 2944 4071 3000 4127
rect 2572 3947 2628 4003
rect 2696 3947 2752 4003
rect 2820 3947 2876 4003
rect 2944 3947 3000 4003
rect 2572 3823 2628 3879
rect 2696 3823 2752 3879
rect 2820 3823 2876 3879
rect 2944 3823 3000 3879
rect 2572 3699 2628 3755
rect 2696 3699 2752 3755
rect 2820 3699 2876 3755
rect 2944 3699 3000 3755
rect 2572 3575 2628 3631
rect 2696 3575 2752 3631
rect 2820 3575 2876 3631
rect 2944 3575 3000 3631
rect 2572 3451 2628 3507
rect 2696 3451 2752 3507
rect 2820 3451 2876 3507
rect 2944 3451 3000 3507
rect 2572 3327 2628 3383
rect 2696 3327 2752 3383
rect 2820 3327 2876 3383
rect 2944 3327 3000 3383
rect 2572 3203 2628 3259
rect 2696 3203 2752 3259
rect 2820 3203 2876 3259
rect 2944 3203 3000 3259
rect 2572 3079 2628 3135
rect 2696 3079 2752 3135
rect 2820 3079 2876 3135
rect 2944 3079 3000 3135
rect 2572 2955 2628 3011
rect 2696 2955 2752 3011
rect 2820 2955 2876 3011
rect 2944 2955 3000 3011
rect 2572 2831 2628 2887
rect 2696 2831 2752 2887
rect 2820 2831 2876 2887
rect 2944 2831 3000 2887
rect 2572 2707 2628 2763
rect 2696 2707 2752 2763
rect 2820 2707 2876 2763
rect 2944 2707 3000 2763
rect 2572 2583 2628 2639
rect 2696 2583 2752 2639
rect 2820 2583 2876 2639
rect 2944 2583 3000 2639
rect 2572 2459 2628 2515
rect 2696 2459 2752 2515
rect 2820 2459 2876 2515
rect 2944 2459 3000 2515
rect 2572 2335 2628 2391
rect 2696 2335 2752 2391
rect 2820 2335 2876 2391
rect 2944 2335 3000 2391
rect 2572 2211 2628 2267
rect 2696 2211 2752 2267
rect 2820 2211 2876 2267
rect 2944 2211 3000 2267
rect 2572 2087 2628 2143
rect 2696 2087 2752 2143
rect 2820 2087 2876 2143
rect 2944 2087 3000 2143
rect 2572 1963 2628 2019
rect 2696 1963 2752 2019
rect 2820 1963 2876 2019
rect 2944 1963 3000 2019
rect 2572 1839 2628 1895
rect 2696 1839 2752 1895
rect 2820 1839 2876 1895
rect 2944 1839 3000 1895
rect 2572 1715 2628 1771
rect 2696 1715 2752 1771
rect 2820 1715 2876 1771
rect 2944 1715 3000 1771
rect 2572 1591 2628 1647
rect 2696 1591 2752 1647
rect 2820 1591 2876 1647
rect 2944 1591 3000 1647
rect 2572 1467 2628 1523
rect 2696 1467 2752 1523
rect 2820 1467 2876 1523
rect 2944 1467 3000 1523
rect 2572 1343 2628 1399
rect 2696 1343 2752 1399
rect 2820 1343 2876 1399
rect 2944 1343 3000 1399
rect 4844 4195 4900 4251
rect 4968 4195 5024 4251
rect 5092 4195 5148 4251
rect 5216 4195 5272 4251
rect 4844 4071 4900 4127
rect 4968 4071 5024 4127
rect 5092 4071 5148 4127
rect 5216 4071 5272 4127
rect 4844 3947 4900 4003
rect 4968 3947 5024 4003
rect 5092 3947 5148 4003
rect 5216 3947 5272 4003
rect 4844 3823 4900 3879
rect 4968 3823 5024 3879
rect 5092 3823 5148 3879
rect 5216 3823 5272 3879
rect 4844 3699 4900 3755
rect 4968 3699 5024 3755
rect 5092 3699 5148 3755
rect 5216 3699 5272 3755
rect 4844 3575 4900 3631
rect 4968 3575 5024 3631
rect 5092 3575 5148 3631
rect 5216 3575 5272 3631
rect 4844 3451 4900 3507
rect 4968 3451 5024 3507
rect 5092 3451 5148 3507
rect 5216 3451 5272 3507
rect 4844 3327 4900 3383
rect 4968 3327 5024 3383
rect 5092 3327 5148 3383
rect 5216 3327 5272 3383
rect 4844 3203 4900 3259
rect 4968 3203 5024 3259
rect 5092 3203 5148 3259
rect 5216 3203 5272 3259
rect 4844 3079 4900 3135
rect 4968 3079 5024 3135
rect 5092 3079 5148 3135
rect 5216 3079 5272 3135
rect 4844 2955 4900 3011
rect 4968 2955 5024 3011
rect 5092 2955 5148 3011
rect 5216 2955 5272 3011
rect 4844 2831 4900 2887
rect 4968 2831 5024 2887
rect 5092 2831 5148 2887
rect 5216 2831 5272 2887
rect 4844 2707 4900 2763
rect 4968 2707 5024 2763
rect 5092 2707 5148 2763
rect 5216 2707 5272 2763
rect 4844 2583 4900 2639
rect 4968 2583 5024 2639
rect 5092 2583 5148 2639
rect 5216 2583 5272 2639
rect 4844 2459 4900 2515
rect 4968 2459 5024 2515
rect 5092 2459 5148 2515
rect 5216 2459 5272 2515
rect 4844 2335 4900 2391
rect 4968 2335 5024 2391
rect 5092 2335 5148 2391
rect 5216 2335 5272 2391
rect 4844 2211 4900 2267
rect 4968 2211 5024 2267
rect 5092 2211 5148 2267
rect 5216 2211 5272 2267
rect 4844 2087 4900 2143
rect 4968 2087 5024 2143
rect 5092 2087 5148 2143
rect 5216 2087 5272 2143
rect 4844 1963 4900 2019
rect 4968 1963 5024 2019
rect 5092 1963 5148 2019
rect 5216 1963 5272 2019
rect 4844 1839 4900 1895
rect 4968 1839 5024 1895
rect 5092 1839 5148 1895
rect 5216 1839 5272 1895
rect 4844 1715 4900 1771
rect 4968 1715 5024 1771
rect 5092 1715 5148 1771
rect 5216 1715 5272 1771
rect 4844 1591 4900 1647
rect 4968 1591 5024 1647
rect 5092 1591 5148 1647
rect 5216 1591 5272 1647
rect 4844 1467 4900 1523
rect 4968 1467 5024 1523
rect 5092 1467 5148 1523
rect 5216 1467 5272 1523
rect 4844 1343 4900 1399
rect 4968 1343 5024 1399
rect 5092 1343 5148 1399
rect 5216 1343 5272 1399
rect 7137 4195 7193 4251
rect 7261 4195 7317 4251
rect 7385 4195 7441 4251
rect 7137 4071 7193 4127
rect 7261 4071 7317 4127
rect 7385 4071 7441 4127
rect 7137 3947 7193 4003
rect 7261 3947 7317 4003
rect 7385 3947 7441 4003
rect 7137 3823 7193 3879
rect 7261 3823 7317 3879
rect 7385 3823 7441 3879
rect 7137 3699 7193 3755
rect 7261 3699 7317 3755
rect 7385 3699 7441 3755
rect 7137 3575 7193 3631
rect 7261 3575 7317 3631
rect 7385 3575 7441 3631
rect 7137 3451 7193 3507
rect 7261 3451 7317 3507
rect 7385 3451 7441 3507
rect 7137 3327 7193 3383
rect 7261 3327 7317 3383
rect 7385 3327 7441 3383
rect 7137 3203 7193 3259
rect 7261 3203 7317 3259
rect 7385 3203 7441 3259
rect 7137 3079 7193 3135
rect 7261 3079 7317 3135
rect 7385 3079 7441 3135
rect 7137 2955 7193 3011
rect 7261 2955 7317 3011
rect 7385 2955 7441 3011
rect 7137 2831 7193 2887
rect 7261 2831 7317 2887
rect 7385 2831 7441 2887
rect 7137 2707 7193 2763
rect 7261 2707 7317 2763
rect 7385 2707 7441 2763
rect 7137 2583 7193 2639
rect 7261 2583 7317 2639
rect 7385 2583 7441 2639
rect 7137 2459 7193 2515
rect 7261 2459 7317 2515
rect 7385 2459 7441 2515
rect 7137 2335 7193 2391
rect 7261 2335 7317 2391
rect 7385 2335 7441 2391
rect 7137 2211 7193 2267
rect 7261 2211 7317 2267
rect 7385 2211 7441 2267
rect 7137 2087 7193 2143
rect 7261 2087 7317 2143
rect 7385 2087 7441 2143
rect 7137 1963 7193 2019
rect 7261 1963 7317 2019
rect 7385 1963 7441 2019
rect 7137 1839 7193 1895
rect 7261 1839 7317 1895
rect 7385 1839 7441 1895
rect 7137 1715 7193 1771
rect 7261 1715 7317 1771
rect 7385 1715 7441 1771
rect 7137 1591 7193 1647
rect 7261 1591 7317 1647
rect 7385 1591 7441 1647
rect 7137 1467 7193 1523
rect 7261 1467 7317 1523
rect 7385 1467 7441 1523
rect 7137 1343 7193 1399
rect 7261 1343 7317 1399
rect 7385 1343 7441 1399
rect 7623 4195 7679 4251
rect 7747 4195 7803 4251
rect 7871 4195 7927 4251
rect 7623 4071 7679 4127
rect 7747 4071 7803 4127
rect 7871 4071 7927 4127
rect 7623 3947 7679 4003
rect 7747 3947 7803 4003
rect 7871 3947 7927 4003
rect 7623 3823 7679 3879
rect 7747 3823 7803 3879
rect 7871 3823 7927 3879
rect 7623 3699 7679 3755
rect 7747 3699 7803 3755
rect 7871 3699 7927 3755
rect 7623 3575 7679 3631
rect 7747 3575 7803 3631
rect 7871 3575 7927 3631
rect 7623 3451 7679 3507
rect 7747 3451 7803 3507
rect 7871 3451 7927 3507
rect 7623 3327 7679 3383
rect 7747 3327 7803 3383
rect 7871 3327 7927 3383
rect 7623 3203 7679 3259
rect 7747 3203 7803 3259
rect 7871 3203 7927 3259
rect 7623 3079 7679 3135
rect 7747 3079 7803 3135
rect 7871 3079 7927 3135
rect 7623 2955 7679 3011
rect 7747 2955 7803 3011
rect 7871 2955 7927 3011
rect 7623 2831 7679 2887
rect 7747 2831 7803 2887
rect 7871 2831 7927 2887
rect 7623 2707 7679 2763
rect 7747 2707 7803 2763
rect 7871 2707 7927 2763
rect 7623 2583 7679 2639
rect 7747 2583 7803 2639
rect 7871 2583 7927 2639
rect 7623 2459 7679 2515
rect 7747 2459 7803 2515
rect 7871 2459 7927 2515
rect 7623 2335 7679 2391
rect 7747 2335 7803 2391
rect 7871 2335 7927 2391
rect 7623 2211 7679 2267
rect 7747 2211 7803 2267
rect 7871 2211 7927 2267
rect 7623 2087 7679 2143
rect 7747 2087 7803 2143
rect 7871 2087 7927 2143
rect 7623 1963 7679 2019
rect 7747 1963 7803 2019
rect 7871 1963 7927 2019
rect 7623 1839 7679 1895
rect 7747 1839 7803 1895
rect 7871 1839 7927 1895
rect 7623 1715 7679 1771
rect 7747 1715 7803 1771
rect 7871 1715 7927 1771
rect 7623 1591 7679 1647
rect 7747 1591 7803 1647
rect 7871 1591 7927 1647
rect 7623 1467 7679 1523
rect 7747 1467 7803 1523
rect 7871 1467 7927 1523
rect 7623 1343 7679 1399
rect 7747 1343 7803 1399
rect 7871 1343 7927 1399
rect 9792 4195 9848 4251
rect 9916 4195 9972 4251
rect 10040 4195 10096 4251
rect 10164 4195 10220 4251
rect 9792 4071 9848 4127
rect 9916 4071 9972 4127
rect 10040 4071 10096 4127
rect 10164 4071 10220 4127
rect 9792 3947 9848 4003
rect 9916 3947 9972 4003
rect 10040 3947 10096 4003
rect 10164 3947 10220 4003
rect 9792 3823 9848 3879
rect 9916 3823 9972 3879
rect 10040 3823 10096 3879
rect 10164 3823 10220 3879
rect 9792 3699 9848 3755
rect 9916 3699 9972 3755
rect 10040 3699 10096 3755
rect 10164 3699 10220 3755
rect 9792 3575 9848 3631
rect 9916 3575 9972 3631
rect 10040 3575 10096 3631
rect 10164 3575 10220 3631
rect 9792 3451 9848 3507
rect 9916 3451 9972 3507
rect 10040 3451 10096 3507
rect 10164 3451 10220 3507
rect 9792 3327 9848 3383
rect 9916 3327 9972 3383
rect 10040 3327 10096 3383
rect 10164 3327 10220 3383
rect 9792 3203 9848 3259
rect 9916 3203 9972 3259
rect 10040 3203 10096 3259
rect 10164 3203 10220 3259
rect 9792 3079 9848 3135
rect 9916 3079 9972 3135
rect 10040 3079 10096 3135
rect 10164 3079 10220 3135
rect 9792 2955 9848 3011
rect 9916 2955 9972 3011
rect 10040 2955 10096 3011
rect 10164 2955 10220 3011
rect 9792 2831 9848 2887
rect 9916 2831 9972 2887
rect 10040 2831 10096 2887
rect 10164 2831 10220 2887
rect 9792 2707 9848 2763
rect 9916 2707 9972 2763
rect 10040 2707 10096 2763
rect 10164 2707 10220 2763
rect 9792 2583 9848 2639
rect 9916 2583 9972 2639
rect 10040 2583 10096 2639
rect 10164 2583 10220 2639
rect 9792 2459 9848 2515
rect 9916 2459 9972 2515
rect 10040 2459 10096 2515
rect 10164 2459 10220 2515
rect 9792 2335 9848 2391
rect 9916 2335 9972 2391
rect 10040 2335 10096 2391
rect 10164 2335 10220 2391
rect 9792 2211 9848 2267
rect 9916 2211 9972 2267
rect 10040 2211 10096 2267
rect 10164 2211 10220 2267
rect 9792 2087 9848 2143
rect 9916 2087 9972 2143
rect 10040 2087 10096 2143
rect 10164 2087 10220 2143
rect 9792 1963 9848 2019
rect 9916 1963 9972 2019
rect 10040 1963 10096 2019
rect 10164 1963 10220 2019
rect 9792 1839 9848 1895
rect 9916 1839 9972 1895
rect 10040 1839 10096 1895
rect 10164 1839 10220 1895
rect 9792 1715 9848 1771
rect 9916 1715 9972 1771
rect 10040 1715 10096 1771
rect 10164 1715 10220 1771
rect 9792 1591 9848 1647
rect 9916 1591 9972 1647
rect 10040 1591 10096 1647
rect 10164 1591 10220 1647
rect 9792 1467 9848 1523
rect 9916 1467 9972 1523
rect 10040 1467 10096 1523
rect 10164 1467 10220 1523
rect 9792 1343 9848 1399
rect 9916 1343 9972 1399
rect 10040 1343 10096 1399
rect 10164 1343 10220 1399
rect 12064 4195 12120 4251
rect 12188 4195 12244 4251
rect 12312 4195 12368 4251
rect 12436 4195 12492 4251
rect 12064 4071 12120 4127
rect 12188 4071 12244 4127
rect 12312 4071 12368 4127
rect 12436 4071 12492 4127
rect 12064 3947 12120 4003
rect 12188 3947 12244 4003
rect 12312 3947 12368 4003
rect 12436 3947 12492 4003
rect 12064 3823 12120 3879
rect 12188 3823 12244 3879
rect 12312 3823 12368 3879
rect 12436 3823 12492 3879
rect 12064 3699 12120 3755
rect 12188 3699 12244 3755
rect 12312 3699 12368 3755
rect 12436 3699 12492 3755
rect 12064 3575 12120 3631
rect 12188 3575 12244 3631
rect 12312 3575 12368 3631
rect 12436 3575 12492 3631
rect 12064 3451 12120 3507
rect 12188 3451 12244 3507
rect 12312 3451 12368 3507
rect 12436 3451 12492 3507
rect 12064 3327 12120 3383
rect 12188 3327 12244 3383
rect 12312 3327 12368 3383
rect 12436 3327 12492 3383
rect 12064 3203 12120 3259
rect 12188 3203 12244 3259
rect 12312 3203 12368 3259
rect 12436 3203 12492 3259
rect 12064 3079 12120 3135
rect 12188 3079 12244 3135
rect 12312 3079 12368 3135
rect 12436 3079 12492 3135
rect 12064 2955 12120 3011
rect 12188 2955 12244 3011
rect 12312 2955 12368 3011
rect 12436 2955 12492 3011
rect 12064 2831 12120 2887
rect 12188 2831 12244 2887
rect 12312 2831 12368 2887
rect 12436 2831 12492 2887
rect 12064 2707 12120 2763
rect 12188 2707 12244 2763
rect 12312 2707 12368 2763
rect 12436 2707 12492 2763
rect 12064 2583 12120 2639
rect 12188 2583 12244 2639
rect 12312 2583 12368 2639
rect 12436 2583 12492 2639
rect 12064 2459 12120 2515
rect 12188 2459 12244 2515
rect 12312 2459 12368 2515
rect 12436 2459 12492 2515
rect 12064 2335 12120 2391
rect 12188 2335 12244 2391
rect 12312 2335 12368 2391
rect 12436 2335 12492 2391
rect 12064 2211 12120 2267
rect 12188 2211 12244 2267
rect 12312 2211 12368 2267
rect 12436 2211 12492 2267
rect 12064 2087 12120 2143
rect 12188 2087 12244 2143
rect 12312 2087 12368 2143
rect 12436 2087 12492 2143
rect 12064 1963 12120 2019
rect 12188 1963 12244 2019
rect 12312 1963 12368 2019
rect 12436 1963 12492 2019
rect 12064 1839 12120 1895
rect 12188 1839 12244 1895
rect 12312 1839 12368 1895
rect 12436 1839 12492 1895
rect 12064 1715 12120 1771
rect 12188 1715 12244 1771
rect 12312 1715 12368 1771
rect 12436 1715 12492 1771
rect 12064 1591 12120 1647
rect 12188 1591 12244 1647
rect 12312 1591 12368 1647
rect 12436 1591 12492 1647
rect 12064 1467 12120 1523
rect 12188 1467 12244 1523
rect 12312 1467 12368 1523
rect 12436 1467 12492 1523
rect 12064 1343 12120 1399
rect 12188 1343 12244 1399
rect 12312 1343 12368 1399
rect 12436 1343 12492 1399
rect 13200 4195 13256 4251
rect 13324 4195 13380 4251
rect 13448 4195 13504 4251
rect 13572 4195 13628 4251
rect 13200 4071 13256 4127
rect 13324 4071 13380 4127
rect 13448 4071 13504 4127
rect 13572 4071 13628 4127
rect 13200 3947 13256 4003
rect 13324 3947 13380 4003
rect 13448 3947 13504 4003
rect 13572 3947 13628 4003
rect 13200 3823 13256 3879
rect 13324 3823 13380 3879
rect 13448 3823 13504 3879
rect 13572 3823 13628 3879
rect 13200 3699 13256 3755
rect 13324 3699 13380 3755
rect 13448 3699 13504 3755
rect 13572 3699 13628 3755
rect 13200 3575 13256 3631
rect 13324 3575 13380 3631
rect 13448 3575 13504 3631
rect 13572 3575 13628 3631
rect 13200 3451 13256 3507
rect 13324 3451 13380 3507
rect 13448 3451 13504 3507
rect 13572 3451 13628 3507
rect 13200 3327 13256 3383
rect 13324 3327 13380 3383
rect 13448 3327 13504 3383
rect 13572 3327 13628 3383
rect 13200 3203 13256 3259
rect 13324 3203 13380 3259
rect 13448 3203 13504 3259
rect 13572 3203 13628 3259
rect 13200 3079 13256 3135
rect 13324 3079 13380 3135
rect 13448 3079 13504 3135
rect 13572 3079 13628 3135
rect 13200 2955 13256 3011
rect 13324 2955 13380 3011
rect 13448 2955 13504 3011
rect 13572 2955 13628 3011
rect 13200 2831 13256 2887
rect 13324 2831 13380 2887
rect 13448 2831 13504 2887
rect 13572 2831 13628 2887
rect 13200 2707 13256 2763
rect 13324 2707 13380 2763
rect 13448 2707 13504 2763
rect 13572 2707 13628 2763
rect 13200 2583 13256 2639
rect 13324 2583 13380 2639
rect 13448 2583 13504 2639
rect 13572 2583 13628 2639
rect 13200 2459 13256 2515
rect 13324 2459 13380 2515
rect 13448 2459 13504 2515
rect 13572 2459 13628 2515
rect 13200 2335 13256 2391
rect 13324 2335 13380 2391
rect 13448 2335 13504 2391
rect 13572 2335 13628 2391
rect 13200 2211 13256 2267
rect 13324 2211 13380 2267
rect 13448 2211 13504 2267
rect 13572 2211 13628 2267
rect 13200 2087 13256 2143
rect 13324 2087 13380 2143
rect 13448 2087 13504 2143
rect 13572 2087 13628 2143
rect 13200 1963 13256 2019
rect 13324 1963 13380 2019
rect 13448 1963 13504 2019
rect 13572 1963 13628 2019
rect 13200 1839 13256 1895
rect 13324 1839 13380 1895
rect 13448 1839 13504 1895
rect 13572 1839 13628 1895
rect 13200 1715 13256 1771
rect 13324 1715 13380 1771
rect 13448 1715 13504 1771
rect 13572 1715 13628 1771
rect 13200 1591 13256 1647
rect 13324 1591 13380 1647
rect 13448 1591 13504 1647
rect 13572 1591 13628 1647
rect 13200 1467 13256 1523
rect 13324 1467 13380 1523
rect 13448 1467 13504 1523
rect 13572 1467 13628 1523
rect 13200 1343 13256 1399
rect 13324 1343 13380 1399
rect 13448 1343 13504 1399
rect 13572 1343 13628 1399
rect 14336 56866 14392 56922
rect 14460 56866 14516 56922
rect 14584 56866 14640 56922
rect 14708 56866 14764 56922
rect 14336 56742 14392 56798
rect 14460 56742 14516 56798
rect 14584 56742 14640 56798
rect 14708 56742 14764 56798
rect 14336 56659 14352 56674
rect 14352 56659 14392 56674
rect 14460 56659 14512 56674
rect 14512 56659 14516 56674
rect 14584 56659 14620 56674
rect 14620 56659 14640 56674
rect 14336 56618 14392 56659
rect 14460 56618 14516 56659
rect 14584 56618 14640 56659
rect 14708 56618 14764 56674
rect 14336 56495 14392 56550
rect 14460 56495 14516 56550
rect 14584 56495 14640 56550
rect 14336 56494 14352 56495
rect 14352 56494 14392 56495
rect 14460 56494 14512 56495
rect 14512 56494 14516 56495
rect 14584 56494 14620 56495
rect 14620 56494 14640 56495
rect 14708 56494 14764 56550
rect 14336 56370 14392 56426
rect 14460 56370 14516 56426
rect 14584 56370 14640 56426
rect 14708 56370 14764 56426
rect 14336 56246 14392 56302
rect 14460 56246 14516 56302
rect 14584 56246 14640 56302
rect 14708 56246 14764 56302
rect 14336 56122 14392 56178
rect 14460 56122 14516 56178
rect 14584 56122 14640 56178
rect 14708 56122 14764 56178
rect 14336 55998 14392 56054
rect 14460 55998 14516 56054
rect 14584 55998 14640 56054
rect 14708 55998 14764 56054
rect 14336 55874 14392 55930
rect 14460 55874 14516 55930
rect 14584 55874 14640 55930
rect 14708 55874 14764 55930
rect 14336 55750 14392 55806
rect 14460 55750 14516 55806
rect 14584 55750 14640 55806
rect 14708 55750 14764 55806
rect 14336 53789 14392 53845
rect 14460 53789 14516 53845
rect 14584 53789 14640 53845
rect 14708 53789 14764 53845
rect 14336 53665 14392 53721
rect 14460 53665 14516 53721
rect 14584 53665 14640 53721
rect 14708 53665 14764 53721
rect 14336 53541 14392 53597
rect 14460 53541 14516 53597
rect 14584 53541 14640 53597
rect 14708 53541 14764 53597
rect 14336 53417 14392 53473
rect 14460 53417 14516 53473
rect 14584 53417 14640 53473
rect 14708 53417 14764 53473
rect 14336 53293 14392 53349
rect 14460 53293 14516 53349
rect 14584 53293 14640 53349
rect 14708 53293 14764 53349
rect 14336 53169 14392 53225
rect 14460 53169 14516 53225
rect 14584 53169 14640 53225
rect 14708 53169 14764 53225
rect 14336 53045 14392 53101
rect 14460 53045 14516 53101
rect 14584 53045 14640 53101
rect 14708 53045 14764 53101
rect 14336 52964 14352 52977
rect 14352 52964 14392 52977
rect 14460 52964 14512 52977
rect 14512 52964 14516 52977
rect 14584 52964 14620 52977
rect 14620 52964 14640 52977
rect 14336 52921 14392 52964
rect 14460 52921 14516 52964
rect 14584 52921 14640 52964
rect 14708 52921 14764 52977
rect 14336 52800 14392 52853
rect 14460 52800 14516 52853
rect 14584 52800 14640 52853
rect 14336 52797 14352 52800
rect 14352 52797 14392 52800
rect 14460 52797 14512 52800
rect 14512 52797 14516 52800
rect 14584 52797 14620 52800
rect 14620 52797 14640 52800
rect 14708 52797 14764 52853
rect 14336 52692 14392 52729
rect 14460 52692 14516 52729
rect 14584 52692 14640 52729
rect 14336 52673 14352 52692
rect 14352 52673 14392 52692
rect 14460 52673 14512 52692
rect 14512 52673 14516 52692
rect 14584 52673 14620 52692
rect 14620 52673 14640 52692
rect 14708 52673 14764 52729
rect 14336 52584 14392 52605
rect 14460 52584 14516 52605
rect 14584 52584 14640 52605
rect 14336 52549 14352 52584
rect 14352 52549 14392 52584
rect 14460 52549 14512 52584
rect 14512 52549 14516 52584
rect 14584 52549 14620 52584
rect 14620 52549 14640 52584
rect 14708 52549 14764 52605
rect 14952 52271 15008 52273
rect 14952 52219 14954 52271
rect 14954 52219 15006 52271
rect 15006 52219 15008 52271
rect 14952 52163 15008 52219
rect 14952 52111 14954 52163
rect 14954 52111 15006 52163
rect 15006 52111 15008 52163
rect 14952 52055 15008 52111
rect 14952 52003 14954 52055
rect 14954 52003 15006 52055
rect 15006 52003 15008 52055
rect 14952 51947 15008 52003
rect 14952 51895 14954 51947
rect 14954 51895 15006 51947
rect 15006 51895 15008 51947
rect 14952 51839 15008 51895
rect 14952 51787 14954 51839
rect 14954 51787 15006 51839
rect 15006 51787 15008 51839
rect 14952 51731 15008 51787
rect 14952 51679 14954 51731
rect 14954 51679 15006 51731
rect 15006 51679 15008 51731
rect 14952 51623 15008 51679
rect 14952 51571 14954 51623
rect 14954 51571 15006 51623
rect 15006 51571 15008 51623
rect 14952 51515 15008 51571
rect 14952 51463 14954 51515
rect 14954 51463 15006 51515
rect 15006 51463 15008 51515
rect 14952 51407 15008 51463
rect 14952 51355 14954 51407
rect 14954 51355 15006 51407
rect 15006 51355 15008 51407
rect 14952 51299 15008 51355
rect 14952 51247 14954 51299
rect 14954 51247 15006 51299
rect 15006 51247 15008 51299
rect 14952 51191 15008 51247
rect 14952 51139 14954 51191
rect 14954 51139 15006 51191
rect 15006 51139 15008 51191
rect 14952 51083 15008 51139
rect 14952 51031 14954 51083
rect 14954 51031 15006 51083
rect 15006 51031 15008 51083
rect 14952 50975 15008 51031
rect 14952 50923 14954 50975
rect 14954 50923 15006 50975
rect 15006 50923 15008 50975
rect 14952 50921 15008 50923
rect 14336 49016 14352 49045
rect 14352 49016 14392 49045
rect 14460 49016 14512 49045
rect 14512 49016 14516 49045
rect 14584 49016 14620 49045
rect 14620 49016 14640 49045
rect 14336 48989 14392 49016
rect 14460 48989 14516 49016
rect 14584 48989 14640 49016
rect 14708 48989 14764 49045
rect 14336 48908 14352 48921
rect 14352 48908 14392 48921
rect 14460 48908 14512 48921
rect 14512 48908 14516 48921
rect 14584 48908 14620 48921
rect 14620 48908 14640 48921
rect 14336 48865 14392 48908
rect 14460 48865 14516 48908
rect 14584 48865 14640 48908
rect 14708 48865 14764 48921
rect 14336 48744 14392 48797
rect 14460 48744 14516 48797
rect 14584 48744 14640 48797
rect 14336 48741 14352 48744
rect 14352 48741 14392 48744
rect 14460 48741 14512 48744
rect 14512 48741 14516 48744
rect 14584 48741 14620 48744
rect 14620 48741 14640 48744
rect 14708 48741 14764 48797
rect 14336 48636 14392 48673
rect 14460 48636 14516 48673
rect 14584 48636 14640 48673
rect 14336 48617 14352 48636
rect 14352 48617 14392 48636
rect 14460 48617 14512 48636
rect 14512 48617 14516 48636
rect 14584 48617 14620 48636
rect 14620 48617 14640 48636
rect 14708 48617 14764 48673
rect 14336 48493 14392 48549
rect 14460 48493 14516 48549
rect 14584 48493 14640 48549
rect 14708 48493 14764 48549
rect 14336 48369 14392 48425
rect 14460 48369 14516 48425
rect 14584 48369 14640 48425
rect 14708 48369 14764 48425
rect 14336 48245 14392 48301
rect 14460 48245 14516 48301
rect 14584 48245 14640 48301
rect 14708 48245 14764 48301
rect 14336 48121 14392 48177
rect 14460 48121 14516 48177
rect 14584 48121 14640 48177
rect 14708 48121 14764 48177
rect 14336 47997 14392 48053
rect 14460 47997 14516 48053
rect 14584 47997 14640 48053
rect 14708 47997 14764 48053
rect 14336 47873 14392 47929
rect 14460 47873 14516 47929
rect 14584 47873 14640 47929
rect 14708 47873 14764 47929
rect 14336 47749 14392 47805
rect 14460 47749 14516 47805
rect 14584 47749 14640 47805
rect 14708 47749 14764 47805
rect 14336 45789 14392 45845
rect 14460 45789 14516 45845
rect 14584 45789 14640 45845
rect 14708 45789 14764 45845
rect 14336 45665 14392 45721
rect 14460 45665 14516 45721
rect 14584 45665 14640 45721
rect 14708 45665 14764 45721
rect 14336 45541 14392 45597
rect 14460 45541 14516 45597
rect 14584 45541 14640 45597
rect 14708 45541 14764 45597
rect 14336 45417 14392 45473
rect 14460 45417 14516 45473
rect 14584 45417 14640 45473
rect 14708 45417 14764 45473
rect 14336 45293 14392 45349
rect 14460 45293 14516 45349
rect 14584 45293 14640 45349
rect 14708 45293 14764 45349
rect 14336 45169 14392 45225
rect 14460 45169 14516 45225
rect 14584 45169 14640 45225
rect 14708 45169 14764 45225
rect 14336 45068 14352 45101
rect 14352 45068 14392 45101
rect 14460 45068 14512 45101
rect 14512 45068 14516 45101
rect 14584 45068 14620 45101
rect 14620 45068 14640 45101
rect 14336 45045 14392 45068
rect 14460 45045 14516 45068
rect 14584 45045 14640 45068
rect 14708 45045 14764 45101
rect 14336 44960 14352 44977
rect 14352 44960 14392 44977
rect 14460 44960 14512 44977
rect 14512 44960 14516 44977
rect 14584 44960 14620 44977
rect 14620 44960 14640 44977
rect 14336 44921 14392 44960
rect 14460 44921 14516 44960
rect 14584 44921 14640 44960
rect 14708 44921 14764 44977
rect 14336 44852 14352 44853
rect 14352 44852 14392 44853
rect 14460 44852 14512 44853
rect 14512 44852 14516 44853
rect 14584 44852 14620 44853
rect 14620 44852 14640 44853
rect 14336 44797 14392 44852
rect 14460 44797 14516 44852
rect 14584 44797 14640 44852
rect 14708 44797 14764 44853
rect 14336 44688 14392 44729
rect 14460 44688 14516 44729
rect 14584 44688 14640 44729
rect 14336 44673 14352 44688
rect 14352 44673 14392 44688
rect 14460 44673 14512 44688
rect 14512 44673 14516 44688
rect 14584 44673 14620 44688
rect 14620 44673 14640 44688
rect 14708 44673 14764 44729
rect 14336 44549 14392 44605
rect 14460 44549 14516 44605
rect 14584 44549 14640 44605
rect 14708 44549 14764 44605
rect 14952 37871 15008 37873
rect 14952 37819 14954 37871
rect 14954 37819 15006 37871
rect 15006 37819 15008 37871
rect 14952 37763 15008 37819
rect 14952 37711 14954 37763
rect 14954 37711 15006 37763
rect 15006 37711 15008 37763
rect 14952 37655 15008 37711
rect 14952 37603 14954 37655
rect 14954 37603 15006 37655
rect 15006 37603 15008 37655
rect 14952 37547 15008 37603
rect 14952 37495 14954 37547
rect 14954 37495 15006 37547
rect 15006 37495 15008 37547
rect 14952 37439 15008 37495
rect 14952 37387 14954 37439
rect 14954 37387 15006 37439
rect 15006 37387 15008 37439
rect 14952 37331 15008 37387
rect 14952 37279 14954 37331
rect 14954 37279 15006 37331
rect 15006 37279 15008 37331
rect 14952 37223 15008 37279
rect 14952 37171 14954 37223
rect 14954 37171 15006 37223
rect 15006 37171 15008 37223
rect 14952 37115 15008 37171
rect 14952 37063 14954 37115
rect 14954 37063 15006 37115
rect 15006 37063 15008 37115
rect 14952 37007 15008 37063
rect 14952 36955 14954 37007
rect 14954 36955 15006 37007
rect 15006 36955 15008 37007
rect 14952 36899 15008 36955
rect 14952 36847 14954 36899
rect 14954 36847 15006 36899
rect 15006 36847 15008 36899
rect 14952 36791 15008 36847
rect 14952 36739 14954 36791
rect 14954 36739 15006 36791
rect 15006 36739 15008 36791
rect 14952 36683 15008 36739
rect 14952 36631 14954 36683
rect 14954 36631 15006 36683
rect 15006 36631 15008 36683
rect 14952 36575 15008 36631
rect 14952 36523 14954 36575
rect 14954 36523 15006 36575
rect 15006 36523 15008 36575
rect 14952 36521 15008 36523
rect 14336 36195 14392 36251
rect 14460 36195 14516 36251
rect 14584 36195 14640 36251
rect 14708 36195 14764 36251
rect 14336 36071 14392 36127
rect 14460 36071 14516 36127
rect 14584 36071 14640 36127
rect 14708 36071 14764 36127
rect 14336 35947 14392 36003
rect 14460 35947 14516 36003
rect 14584 35947 14640 36003
rect 14708 35947 14764 36003
rect 14336 35823 14392 35879
rect 14460 35823 14516 35879
rect 14584 35823 14640 35879
rect 14708 35823 14764 35879
rect 14336 35699 14392 35755
rect 14460 35699 14516 35755
rect 14584 35699 14640 35755
rect 14708 35699 14764 35755
rect 14336 35575 14392 35631
rect 14460 35575 14516 35631
rect 14584 35575 14640 35631
rect 14708 35575 14764 35631
rect 14336 35451 14392 35507
rect 14460 35451 14516 35507
rect 14584 35451 14640 35507
rect 14708 35451 14764 35507
rect 14336 35327 14392 35383
rect 14460 35327 14516 35383
rect 14584 35327 14640 35383
rect 14708 35327 14764 35383
rect 14336 35203 14392 35259
rect 14460 35203 14516 35259
rect 14584 35203 14640 35259
rect 14708 35203 14764 35259
rect 14336 35079 14392 35135
rect 14460 35079 14516 35135
rect 14584 35079 14640 35135
rect 14708 35079 14764 35135
rect 14336 34955 14392 35011
rect 14460 34955 14516 35011
rect 14584 34955 14640 35011
rect 14708 34955 14764 35011
rect 14336 34831 14392 34887
rect 14460 34831 14516 34887
rect 14584 34831 14640 34887
rect 14708 34831 14764 34887
rect 14336 34707 14392 34763
rect 14460 34707 14516 34763
rect 14584 34707 14640 34763
rect 14708 34707 14764 34763
rect 14336 34583 14392 34639
rect 14460 34583 14516 34639
rect 14584 34583 14640 34639
rect 14708 34583 14764 34639
rect 14336 34459 14392 34515
rect 14460 34459 14516 34515
rect 14584 34459 14640 34515
rect 14708 34459 14764 34515
rect 14336 34335 14392 34391
rect 14460 34335 14516 34391
rect 14584 34335 14640 34391
rect 14708 34335 14764 34391
rect 14336 34211 14392 34267
rect 14460 34211 14516 34267
rect 14584 34211 14640 34267
rect 14708 34211 14764 34267
rect 14336 34087 14392 34143
rect 14460 34087 14516 34143
rect 14584 34087 14640 34143
rect 14708 34087 14764 34143
rect 14336 33963 14392 34019
rect 14460 33963 14516 34019
rect 14584 33963 14640 34019
rect 14708 33963 14764 34019
rect 14336 33839 14392 33895
rect 14460 33839 14516 33895
rect 14584 33839 14640 33895
rect 14708 33839 14764 33895
rect 14336 33715 14392 33771
rect 14460 33715 14516 33771
rect 14584 33715 14640 33771
rect 14708 33715 14764 33771
rect 14336 33591 14392 33647
rect 14460 33591 14516 33647
rect 14584 33591 14640 33647
rect 14708 33591 14764 33647
rect 14336 33467 14392 33523
rect 14460 33467 14516 33523
rect 14584 33467 14640 33523
rect 14708 33467 14764 33523
rect 14336 33343 14392 33399
rect 14460 33343 14516 33399
rect 14584 33343 14640 33399
rect 14708 33343 14764 33399
rect 14336 28189 14392 28245
rect 14460 28189 14516 28245
rect 14584 28189 14640 28245
rect 14708 28189 14764 28245
rect 14336 28065 14392 28121
rect 14460 28065 14516 28121
rect 14584 28065 14640 28121
rect 14708 28065 14764 28121
rect 14336 27941 14392 27997
rect 14460 27941 14516 27997
rect 14584 27941 14640 27997
rect 14708 27941 14764 27997
rect 14336 27817 14392 27873
rect 14460 27817 14516 27873
rect 14584 27817 14640 27873
rect 14708 27817 14764 27873
rect 14336 27693 14392 27749
rect 14460 27693 14516 27749
rect 14584 27693 14640 27749
rect 14708 27693 14764 27749
rect 14336 27569 14392 27625
rect 14460 27569 14516 27625
rect 14584 27569 14640 27625
rect 14708 27569 14764 27625
rect 14336 27445 14392 27501
rect 14460 27445 14516 27501
rect 14584 27445 14640 27501
rect 14708 27445 14764 27501
rect 14336 27321 14392 27377
rect 14460 27321 14516 27377
rect 14584 27321 14640 27377
rect 14708 27321 14764 27377
rect 14336 27197 14392 27253
rect 14460 27197 14516 27253
rect 14584 27197 14640 27253
rect 14708 27197 14764 27253
rect 14336 27073 14392 27129
rect 14460 27073 14516 27129
rect 14584 27073 14640 27129
rect 14708 27073 14764 27129
rect 14336 26949 14392 27005
rect 14460 26949 14516 27005
rect 14584 26949 14640 27005
rect 14708 26949 14764 27005
rect 14336 13789 14392 13845
rect 14460 13789 14516 13845
rect 14584 13789 14640 13845
rect 14708 13789 14764 13845
rect 14336 13665 14392 13721
rect 14460 13665 14516 13721
rect 14584 13665 14640 13721
rect 14708 13665 14764 13721
rect 14336 13541 14392 13597
rect 14460 13541 14516 13597
rect 14584 13541 14640 13597
rect 14708 13541 14764 13597
rect 14336 13417 14392 13473
rect 14460 13417 14516 13473
rect 14584 13417 14640 13473
rect 14708 13417 14764 13473
rect 14336 13293 14392 13349
rect 14460 13293 14516 13349
rect 14584 13293 14640 13349
rect 14708 13293 14764 13349
rect 14336 13169 14392 13225
rect 14460 13169 14516 13225
rect 14584 13169 14640 13225
rect 14708 13169 14764 13225
rect 14336 13045 14392 13101
rect 14460 13045 14516 13101
rect 14584 13045 14640 13101
rect 14708 13045 14764 13101
rect 14336 12921 14392 12977
rect 14460 12921 14516 12977
rect 14584 12921 14640 12977
rect 14708 12921 14764 12977
rect 14336 12797 14392 12853
rect 14460 12797 14516 12853
rect 14584 12797 14640 12853
rect 14708 12797 14764 12853
rect 14336 12673 14392 12729
rect 14460 12673 14516 12729
rect 14584 12673 14640 12729
rect 14708 12673 14764 12729
rect 14336 12549 14392 12605
rect 14460 12549 14516 12605
rect 14584 12549 14640 12605
rect 14708 12549 14764 12605
rect 14336 10595 14392 10651
rect 14460 10595 14516 10651
rect 14584 10595 14640 10651
rect 14708 10595 14764 10651
rect 14336 10471 14392 10527
rect 14460 10471 14516 10527
rect 14584 10471 14640 10527
rect 14708 10471 14764 10527
rect 14336 10347 14392 10403
rect 14460 10347 14516 10403
rect 14584 10347 14640 10403
rect 14708 10347 14764 10403
rect 14336 10223 14392 10279
rect 14460 10223 14516 10279
rect 14584 10223 14640 10279
rect 14708 10223 14764 10279
rect 14336 10099 14392 10155
rect 14460 10099 14516 10155
rect 14584 10099 14640 10155
rect 14708 10099 14764 10155
rect 14336 9975 14392 10031
rect 14460 9975 14516 10031
rect 14584 9975 14640 10031
rect 14708 9975 14764 10031
rect 14336 9851 14392 9907
rect 14460 9851 14516 9907
rect 14584 9851 14640 9907
rect 14708 9851 14764 9907
rect 14336 9727 14392 9783
rect 14460 9727 14516 9783
rect 14584 9727 14640 9783
rect 14708 9727 14764 9783
rect 14336 9603 14392 9659
rect 14460 9603 14516 9659
rect 14584 9603 14640 9659
rect 14708 9603 14764 9659
rect 14336 9479 14392 9535
rect 14460 9479 14516 9535
rect 14584 9479 14640 9535
rect 14708 9479 14764 9535
rect 14336 9355 14392 9411
rect 14460 9355 14516 9411
rect 14584 9355 14640 9411
rect 14708 9355 14764 9411
rect 14336 9231 14392 9287
rect 14460 9231 14516 9287
rect 14584 9231 14640 9287
rect 14708 9231 14764 9287
rect 14336 9107 14392 9163
rect 14460 9107 14516 9163
rect 14584 9107 14640 9163
rect 14708 9107 14764 9163
rect 14336 8983 14392 9039
rect 14460 8983 14516 9039
rect 14584 8983 14640 9039
rect 14708 8983 14764 9039
rect 14336 8859 14392 8915
rect 14460 8859 14516 8915
rect 14584 8859 14640 8915
rect 14708 8859 14764 8915
rect 14336 8735 14392 8791
rect 14460 8735 14516 8791
rect 14584 8735 14640 8791
rect 14708 8735 14764 8791
rect 14336 8611 14392 8667
rect 14460 8611 14516 8667
rect 14584 8611 14640 8667
rect 14708 8611 14764 8667
rect 14336 8487 14392 8543
rect 14460 8487 14516 8543
rect 14584 8487 14640 8543
rect 14708 8487 14764 8543
rect 14336 8363 14392 8419
rect 14460 8363 14516 8419
rect 14584 8363 14640 8419
rect 14708 8363 14764 8419
rect 14336 8239 14392 8295
rect 14460 8239 14516 8295
rect 14584 8239 14640 8295
rect 14708 8239 14764 8295
rect 14336 8115 14392 8171
rect 14460 8115 14516 8171
rect 14584 8115 14640 8171
rect 14708 8115 14764 8171
rect 14336 7991 14392 8047
rect 14460 7991 14516 8047
rect 14584 7991 14640 8047
rect 14708 7991 14764 8047
rect 14336 7867 14392 7923
rect 14460 7867 14516 7923
rect 14584 7867 14640 7923
rect 14708 7867 14764 7923
rect 14336 7743 14392 7799
rect 14460 7743 14516 7799
rect 14584 7743 14640 7799
rect 14708 7743 14764 7799
rect 14336 7395 14392 7451
rect 14460 7395 14516 7451
rect 14584 7395 14640 7451
rect 14708 7395 14764 7451
rect 14336 7271 14392 7327
rect 14460 7271 14516 7327
rect 14584 7271 14640 7327
rect 14708 7271 14764 7327
rect 14336 7147 14392 7203
rect 14460 7147 14516 7203
rect 14584 7147 14640 7203
rect 14708 7147 14764 7203
rect 14336 7023 14392 7079
rect 14460 7023 14516 7079
rect 14584 7023 14640 7079
rect 14708 7023 14764 7079
rect 14336 6899 14392 6955
rect 14460 6899 14516 6955
rect 14584 6899 14640 6955
rect 14708 6899 14764 6955
rect 14336 6775 14392 6831
rect 14460 6775 14516 6831
rect 14584 6775 14640 6831
rect 14708 6775 14764 6831
rect 14336 6651 14392 6707
rect 14460 6651 14516 6707
rect 14584 6651 14640 6707
rect 14708 6651 14764 6707
rect 14336 6527 14392 6583
rect 14460 6527 14516 6583
rect 14584 6527 14640 6583
rect 14708 6527 14764 6583
rect 14336 6403 14392 6459
rect 14460 6403 14516 6459
rect 14584 6403 14640 6459
rect 14708 6403 14764 6459
rect 14336 6279 14392 6335
rect 14460 6279 14516 6335
rect 14584 6279 14640 6335
rect 14708 6279 14764 6335
rect 14336 6155 14392 6211
rect 14460 6155 14516 6211
rect 14584 6155 14640 6211
rect 14708 6155 14764 6211
rect 14336 6031 14392 6087
rect 14460 6031 14516 6087
rect 14584 6031 14640 6087
rect 14708 6031 14764 6087
rect 14336 5907 14392 5963
rect 14460 5907 14516 5963
rect 14584 5907 14640 5963
rect 14708 5907 14764 5963
rect 14336 5783 14392 5839
rect 14460 5783 14516 5839
rect 14584 5783 14640 5839
rect 14708 5783 14764 5839
rect 14336 5659 14392 5715
rect 14460 5659 14516 5715
rect 14584 5659 14640 5715
rect 14708 5659 14764 5715
rect 14336 5535 14392 5591
rect 14460 5535 14516 5591
rect 14584 5535 14640 5591
rect 14708 5535 14764 5591
rect 14336 5411 14392 5467
rect 14460 5411 14516 5467
rect 14584 5411 14640 5467
rect 14708 5411 14764 5467
rect 14336 5287 14392 5343
rect 14460 5287 14516 5343
rect 14584 5287 14640 5343
rect 14708 5287 14764 5343
rect 14336 5163 14392 5219
rect 14460 5163 14516 5219
rect 14584 5163 14640 5219
rect 14708 5163 14764 5219
rect 14336 5039 14392 5095
rect 14460 5039 14516 5095
rect 14584 5039 14640 5095
rect 14708 5039 14764 5095
rect 14336 4915 14392 4971
rect 14460 4915 14516 4971
rect 14584 4915 14640 4971
rect 14708 4915 14764 4971
rect 14336 4791 14392 4847
rect 14460 4791 14516 4847
rect 14584 4791 14640 4847
rect 14708 4791 14764 4847
rect 14336 4667 14392 4723
rect 14460 4667 14516 4723
rect 14584 4667 14640 4723
rect 14708 4667 14764 4723
rect 14336 4543 14392 4599
rect 14460 4543 14516 4599
rect 14584 4543 14640 4599
rect 14708 4543 14764 4599
rect 14336 4195 14392 4251
rect 14460 4195 14516 4251
rect 14584 4195 14640 4251
rect 14708 4195 14764 4251
rect 14336 4071 14392 4127
rect 14460 4071 14516 4127
rect 14584 4071 14640 4127
rect 14708 4071 14764 4127
rect 14336 3947 14392 4003
rect 14460 3947 14516 4003
rect 14584 3947 14640 4003
rect 14708 3947 14764 4003
rect 14336 3823 14392 3879
rect 14460 3823 14516 3879
rect 14584 3823 14640 3879
rect 14708 3823 14764 3879
rect 14336 3699 14392 3755
rect 14460 3699 14516 3755
rect 14584 3699 14640 3755
rect 14708 3699 14764 3755
rect 14336 3575 14392 3631
rect 14460 3575 14516 3631
rect 14584 3575 14640 3631
rect 14708 3575 14764 3631
rect 14336 3451 14392 3507
rect 14460 3451 14516 3507
rect 14584 3451 14640 3507
rect 14708 3451 14764 3507
rect 14336 3327 14392 3383
rect 14460 3327 14516 3383
rect 14584 3327 14640 3383
rect 14708 3327 14764 3383
rect 14336 3203 14392 3259
rect 14460 3203 14516 3259
rect 14584 3203 14640 3259
rect 14708 3203 14764 3259
rect 14336 3079 14392 3135
rect 14460 3079 14516 3135
rect 14584 3079 14640 3135
rect 14708 3079 14764 3135
rect 14336 2955 14392 3011
rect 14460 2955 14516 3011
rect 14584 2955 14640 3011
rect 14708 2955 14764 3011
rect 14336 2831 14392 2887
rect 14460 2831 14516 2887
rect 14584 2831 14640 2887
rect 14708 2831 14764 2887
rect 14336 2707 14392 2763
rect 14460 2707 14516 2763
rect 14584 2707 14640 2763
rect 14708 2707 14764 2763
rect 14336 2583 14392 2639
rect 14460 2583 14516 2639
rect 14584 2583 14640 2639
rect 14708 2583 14764 2639
rect 14336 2459 14392 2515
rect 14460 2459 14516 2515
rect 14584 2459 14640 2515
rect 14708 2459 14764 2515
rect 14336 2335 14392 2391
rect 14460 2335 14516 2391
rect 14584 2335 14640 2391
rect 14708 2335 14764 2391
rect 14336 2211 14392 2267
rect 14460 2211 14516 2267
rect 14584 2211 14640 2267
rect 14708 2211 14764 2267
rect 14336 2087 14392 2143
rect 14460 2087 14516 2143
rect 14584 2087 14640 2143
rect 14708 2087 14764 2143
rect 14336 1963 14392 2019
rect 14460 1963 14516 2019
rect 14584 1963 14640 2019
rect 14708 1963 14764 2019
rect 14336 1839 14392 1895
rect 14460 1839 14516 1895
rect 14584 1839 14640 1895
rect 14708 1839 14764 1895
rect 14336 1715 14392 1771
rect 14460 1715 14516 1771
rect 14584 1715 14640 1771
rect 14708 1715 14764 1771
rect 14336 1591 14392 1647
rect 14460 1591 14516 1647
rect 14584 1591 14640 1647
rect 14708 1591 14764 1647
rect 14336 1467 14392 1523
rect 14460 1467 14516 1523
rect 14584 1467 14640 1523
rect 14708 1467 14764 1523
rect 14336 1343 14392 1399
rect 14460 1343 14516 1399
rect 14584 1343 14640 1399
rect 14708 1343 14764 1399
<< metal3 >>
rect 290 56922 738 56932
rect 290 56866 300 56922
rect 356 56866 424 56922
rect 480 56866 548 56922
rect 604 56866 672 56922
rect 728 56866 738 56922
rect 290 56798 738 56866
rect 290 56742 300 56798
rect 356 56742 424 56798
rect 480 56742 548 56798
rect 604 56742 672 56798
rect 728 56742 738 56798
rect 290 56674 738 56742
rect 290 56618 300 56674
rect 356 56618 424 56674
rect 480 56618 548 56674
rect 604 56618 672 56674
rect 728 56618 738 56674
rect 290 56550 738 56618
rect 290 56494 300 56550
rect 356 56494 424 56550
rect 480 56494 548 56550
rect 604 56494 672 56550
rect 728 56494 738 56550
rect 290 56426 738 56494
rect 290 56370 300 56426
rect 356 56370 424 56426
rect 480 56370 548 56426
rect 604 56370 672 56426
rect 728 56370 738 56426
rect 290 56302 738 56370
rect 290 56246 300 56302
rect 356 56246 424 56302
rect 480 56246 548 56302
rect 604 56246 672 56302
rect 728 56246 738 56302
rect 290 56178 738 56246
rect 290 56122 300 56178
rect 356 56122 424 56178
rect 480 56122 548 56178
rect 604 56122 672 56178
rect 728 56122 738 56178
rect 290 56054 738 56122
rect 290 55998 300 56054
rect 356 55998 424 56054
rect 480 55998 548 56054
rect 604 55998 672 56054
rect 728 55998 738 56054
rect 290 55930 738 55998
rect 290 55874 300 55930
rect 356 55874 424 55930
rect 480 55874 548 55930
rect 604 55874 672 55930
rect 728 55874 738 55930
rect 290 55806 738 55874
rect 290 55750 300 55806
rect 356 55750 424 55806
rect 480 55750 548 55806
rect 604 55750 672 55806
rect 728 55750 738 55806
rect 290 55740 738 55750
rect 1426 56922 1874 56932
rect 1426 56866 1436 56922
rect 1492 56866 1560 56922
rect 1616 56866 1684 56922
rect 1740 56866 1808 56922
rect 1864 56866 1874 56922
rect 1426 56798 1874 56866
rect 1426 56742 1436 56798
rect 1492 56742 1560 56798
rect 1616 56742 1684 56798
rect 1740 56742 1808 56798
rect 1864 56742 1874 56798
rect 1426 56674 1874 56742
rect 1426 56618 1436 56674
rect 1492 56618 1560 56674
rect 1616 56618 1684 56674
rect 1740 56618 1808 56674
rect 1864 56618 1874 56674
rect 1426 56550 1874 56618
rect 1426 56494 1436 56550
rect 1492 56494 1560 56550
rect 1616 56494 1684 56550
rect 1740 56494 1808 56550
rect 1864 56494 1874 56550
rect 1426 56426 1874 56494
rect 1426 56370 1436 56426
rect 1492 56370 1560 56426
rect 1616 56370 1684 56426
rect 1740 56370 1808 56426
rect 1864 56370 1874 56426
rect 1426 56302 1874 56370
rect 1426 56246 1436 56302
rect 1492 56246 1560 56302
rect 1616 56246 1684 56302
rect 1740 56246 1808 56302
rect 1864 56246 1874 56302
rect 1426 56178 1874 56246
rect 1426 56122 1436 56178
rect 1492 56122 1560 56178
rect 1616 56122 1684 56178
rect 1740 56122 1808 56178
rect 1864 56122 1874 56178
rect 1426 56054 1874 56122
rect 1426 55998 1436 56054
rect 1492 55998 1560 56054
rect 1616 55998 1684 56054
rect 1740 55998 1808 56054
rect 1864 55998 1874 56054
rect 1426 55930 1874 55998
rect 1426 55874 1436 55930
rect 1492 55874 1560 55930
rect 1616 55874 1684 55930
rect 1740 55874 1808 55930
rect 1864 55874 1874 55930
rect 1426 55806 1874 55874
rect 1426 55750 1436 55806
rect 1492 55750 1560 55806
rect 1616 55750 1684 55806
rect 1740 55750 1808 55806
rect 1864 55750 1874 55806
rect 1426 55740 1874 55750
rect 2562 56922 3010 56932
rect 2562 56866 2572 56922
rect 2628 56866 2696 56922
rect 2752 56866 2820 56922
rect 2876 56866 2944 56922
rect 3000 56866 3010 56922
rect 2562 56798 3010 56866
rect 2562 56742 2572 56798
rect 2628 56742 2696 56798
rect 2752 56742 2820 56798
rect 2876 56742 2944 56798
rect 3000 56742 3010 56798
rect 2562 56674 3010 56742
rect 2562 56618 2572 56674
rect 2628 56618 2696 56674
rect 2752 56618 2820 56674
rect 2876 56618 2944 56674
rect 3000 56618 3010 56674
rect 2562 56550 3010 56618
rect 2562 56494 2572 56550
rect 2628 56494 2696 56550
rect 2752 56494 2820 56550
rect 2876 56494 2944 56550
rect 3000 56494 3010 56550
rect 2562 56426 3010 56494
rect 2562 56370 2572 56426
rect 2628 56370 2696 56426
rect 2752 56370 2820 56426
rect 2876 56370 2944 56426
rect 3000 56370 3010 56426
rect 2562 56302 3010 56370
rect 2562 56246 2572 56302
rect 2628 56246 2696 56302
rect 2752 56246 2820 56302
rect 2876 56246 2944 56302
rect 3000 56246 3010 56302
rect 2562 56178 3010 56246
rect 2562 56122 2572 56178
rect 2628 56122 2696 56178
rect 2752 56122 2820 56178
rect 2876 56122 2944 56178
rect 3000 56122 3010 56178
rect 2562 56054 3010 56122
rect 2562 55998 2572 56054
rect 2628 55998 2696 56054
rect 2752 55998 2820 56054
rect 2876 55998 2944 56054
rect 3000 55998 3010 56054
rect 2562 55930 3010 55998
rect 2562 55874 2572 55930
rect 2628 55874 2696 55930
rect 2752 55874 2820 55930
rect 2876 55874 2944 55930
rect 3000 55874 3010 55930
rect 2562 55806 3010 55874
rect 2562 55750 2572 55806
rect 2628 55750 2696 55806
rect 2752 55750 2820 55806
rect 2876 55750 2944 55806
rect 3000 55750 3010 55806
rect 2562 55740 3010 55750
rect 4834 56922 5282 56932
rect 4834 56866 4844 56922
rect 4900 56866 4968 56922
rect 5024 56866 5092 56922
rect 5148 56866 5216 56922
rect 5272 56866 5282 56922
rect 4834 56798 5282 56866
rect 4834 56742 4844 56798
rect 4900 56742 4968 56798
rect 5024 56742 5092 56798
rect 5148 56742 5216 56798
rect 5272 56742 5282 56798
rect 4834 56674 5282 56742
rect 4834 56618 4844 56674
rect 4900 56618 4968 56674
rect 5024 56618 5092 56674
rect 5148 56618 5216 56674
rect 5272 56618 5282 56674
rect 4834 56550 5282 56618
rect 4834 56494 4844 56550
rect 4900 56494 4968 56550
rect 5024 56494 5092 56550
rect 5148 56494 5216 56550
rect 5272 56494 5282 56550
rect 4834 56426 5282 56494
rect 4834 56370 4844 56426
rect 4900 56370 4968 56426
rect 5024 56370 5092 56426
rect 5148 56370 5216 56426
rect 5272 56370 5282 56426
rect 4834 56302 5282 56370
rect 4834 56246 4844 56302
rect 4900 56246 4968 56302
rect 5024 56246 5092 56302
rect 5148 56246 5216 56302
rect 5272 56246 5282 56302
rect 4834 56178 5282 56246
rect 4834 56122 4844 56178
rect 4900 56122 4968 56178
rect 5024 56122 5092 56178
rect 5148 56122 5216 56178
rect 5272 56122 5282 56178
rect 4834 56054 5282 56122
rect 4834 55998 4844 56054
rect 4900 55998 4968 56054
rect 5024 55998 5092 56054
rect 5148 55998 5216 56054
rect 5272 55998 5282 56054
rect 4834 55930 5282 55998
rect 4834 55874 4844 55930
rect 4900 55874 4968 55930
rect 5024 55874 5092 55930
rect 5148 55874 5216 55930
rect 5272 55874 5282 55930
rect 4834 55806 5282 55874
rect 4834 55750 4844 55806
rect 4900 55750 4968 55806
rect 5024 55750 5092 55806
rect 5148 55750 5216 55806
rect 5272 55750 5282 55806
rect 4834 55740 5282 55750
rect 7127 56922 7451 56932
rect 7127 56866 7137 56922
rect 7193 56866 7261 56922
rect 7317 56866 7385 56922
rect 7441 56866 7451 56922
rect 7127 56798 7451 56866
rect 7127 56742 7137 56798
rect 7193 56742 7261 56798
rect 7317 56742 7385 56798
rect 7441 56742 7451 56798
rect 7127 56674 7451 56742
rect 7127 56618 7137 56674
rect 7193 56618 7261 56674
rect 7317 56618 7385 56674
rect 7441 56618 7451 56674
rect 7127 56550 7451 56618
rect 7127 56494 7137 56550
rect 7193 56494 7261 56550
rect 7317 56494 7385 56550
rect 7441 56494 7451 56550
rect 7127 56426 7451 56494
rect 7127 56370 7137 56426
rect 7193 56370 7261 56426
rect 7317 56370 7385 56426
rect 7441 56370 7451 56426
rect 7127 56302 7451 56370
rect 7127 56246 7137 56302
rect 7193 56246 7261 56302
rect 7317 56246 7385 56302
rect 7441 56246 7451 56302
rect 7127 56178 7451 56246
rect 7127 56122 7137 56178
rect 7193 56122 7261 56178
rect 7317 56122 7385 56178
rect 7441 56122 7451 56178
rect 7127 56054 7451 56122
rect 7127 55998 7137 56054
rect 7193 55998 7261 56054
rect 7317 55998 7385 56054
rect 7441 55998 7451 56054
rect 7127 55930 7451 55998
rect 7127 55874 7137 55930
rect 7193 55874 7261 55930
rect 7317 55874 7385 55930
rect 7441 55874 7451 55930
rect 7127 55806 7451 55874
rect 7127 55750 7137 55806
rect 7193 55750 7261 55806
rect 7317 55750 7385 55806
rect 7441 55750 7451 55806
rect 7127 55740 7451 55750
rect 7613 56922 7937 56932
rect 7613 56866 7623 56922
rect 7679 56866 7747 56922
rect 7803 56866 7871 56922
rect 7927 56866 7937 56922
rect 7613 56798 7937 56866
rect 7613 56742 7623 56798
rect 7679 56742 7747 56798
rect 7803 56742 7871 56798
rect 7927 56742 7937 56798
rect 7613 56674 7937 56742
rect 7613 56618 7623 56674
rect 7679 56618 7747 56674
rect 7803 56618 7871 56674
rect 7927 56618 7937 56674
rect 7613 56550 7937 56618
rect 7613 56494 7623 56550
rect 7679 56494 7747 56550
rect 7803 56494 7871 56550
rect 7927 56494 7937 56550
rect 7613 56426 7937 56494
rect 7613 56370 7623 56426
rect 7679 56370 7747 56426
rect 7803 56370 7871 56426
rect 7927 56370 7937 56426
rect 7613 56302 7937 56370
rect 7613 56246 7623 56302
rect 7679 56246 7747 56302
rect 7803 56246 7871 56302
rect 7927 56246 7937 56302
rect 7613 56178 7937 56246
rect 7613 56122 7623 56178
rect 7679 56122 7747 56178
rect 7803 56122 7871 56178
rect 7927 56122 7937 56178
rect 7613 56054 7937 56122
rect 7613 55998 7623 56054
rect 7679 55998 7747 56054
rect 7803 55998 7871 56054
rect 7927 55998 7937 56054
rect 7613 55930 7937 55998
rect 7613 55874 7623 55930
rect 7679 55874 7747 55930
rect 7803 55874 7871 55930
rect 7927 55874 7937 55930
rect 7613 55806 7937 55874
rect 7613 55750 7623 55806
rect 7679 55750 7747 55806
rect 7803 55750 7871 55806
rect 7927 55750 7937 55806
rect 7613 55740 7937 55750
rect 9782 56922 10230 56932
rect 9782 56866 9792 56922
rect 9848 56866 9916 56922
rect 9972 56866 10040 56922
rect 10096 56866 10164 56922
rect 10220 56866 10230 56922
rect 9782 56798 10230 56866
rect 9782 56742 9792 56798
rect 9848 56742 9916 56798
rect 9972 56742 10040 56798
rect 10096 56742 10164 56798
rect 10220 56742 10230 56798
rect 9782 56674 10230 56742
rect 9782 56618 9792 56674
rect 9848 56618 9916 56674
rect 9972 56618 10040 56674
rect 10096 56618 10164 56674
rect 10220 56618 10230 56674
rect 9782 56550 10230 56618
rect 9782 56494 9792 56550
rect 9848 56494 9916 56550
rect 9972 56494 10040 56550
rect 10096 56494 10164 56550
rect 10220 56494 10230 56550
rect 9782 56426 10230 56494
rect 9782 56370 9792 56426
rect 9848 56370 9916 56426
rect 9972 56370 10040 56426
rect 10096 56370 10164 56426
rect 10220 56370 10230 56426
rect 9782 56302 10230 56370
rect 9782 56246 9792 56302
rect 9848 56246 9916 56302
rect 9972 56246 10040 56302
rect 10096 56246 10164 56302
rect 10220 56246 10230 56302
rect 9782 56178 10230 56246
rect 9782 56122 9792 56178
rect 9848 56122 9916 56178
rect 9972 56122 10040 56178
rect 10096 56122 10164 56178
rect 10220 56122 10230 56178
rect 9782 56054 10230 56122
rect 9782 55998 9792 56054
rect 9848 55998 9916 56054
rect 9972 55998 10040 56054
rect 10096 55998 10164 56054
rect 10220 55998 10230 56054
rect 9782 55930 10230 55998
rect 9782 55874 9792 55930
rect 9848 55874 9916 55930
rect 9972 55874 10040 55930
rect 10096 55874 10164 55930
rect 10220 55874 10230 55930
rect 9782 55806 10230 55874
rect 9782 55750 9792 55806
rect 9848 55750 9916 55806
rect 9972 55750 10040 55806
rect 10096 55750 10164 55806
rect 10220 55750 10230 55806
rect 9782 55740 10230 55750
rect 12054 56922 12502 56932
rect 12054 56866 12064 56922
rect 12120 56866 12188 56922
rect 12244 56866 12312 56922
rect 12368 56866 12436 56922
rect 12492 56866 12502 56922
rect 12054 56798 12502 56866
rect 12054 56742 12064 56798
rect 12120 56742 12188 56798
rect 12244 56742 12312 56798
rect 12368 56742 12436 56798
rect 12492 56742 12502 56798
rect 12054 56674 12502 56742
rect 12054 56618 12064 56674
rect 12120 56618 12188 56674
rect 12244 56618 12312 56674
rect 12368 56618 12436 56674
rect 12492 56618 12502 56674
rect 12054 56550 12502 56618
rect 12054 56494 12064 56550
rect 12120 56494 12188 56550
rect 12244 56494 12312 56550
rect 12368 56494 12436 56550
rect 12492 56494 12502 56550
rect 12054 56426 12502 56494
rect 12054 56370 12064 56426
rect 12120 56370 12188 56426
rect 12244 56370 12312 56426
rect 12368 56370 12436 56426
rect 12492 56370 12502 56426
rect 12054 56302 12502 56370
rect 12054 56246 12064 56302
rect 12120 56246 12188 56302
rect 12244 56246 12312 56302
rect 12368 56246 12436 56302
rect 12492 56246 12502 56302
rect 12054 56178 12502 56246
rect 12054 56122 12064 56178
rect 12120 56122 12188 56178
rect 12244 56122 12312 56178
rect 12368 56122 12436 56178
rect 12492 56122 12502 56178
rect 12054 56054 12502 56122
rect 12054 55998 12064 56054
rect 12120 55998 12188 56054
rect 12244 55998 12312 56054
rect 12368 55998 12436 56054
rect 12492 55998 12502 56054
rect 12054 55930 12502 55998
rect 12054 55874 12064 55930
rect 12120 55874 12188 55930
rect 12244 55874 12312 55930
rect 12368 55874 12436 55930
rect 12492 55874 12502 55930
rect 12054 55806 12502 55874
rect 12054 55750 12064 55806
rect 12120 55750 12188 55806
rect 12244 55750 12312 55806
rect 12368 55750 12436 55806
rect 12492 55750 12502 55806
rect 12054 55740 12502 55750
rect 13190 56922 13638 56932
rect 13190 56866 13200 56922
rect 13256 56866 13324 56922
rect 13380 56866 13448 56922
rect 13504 56866 13572 56922
rect 13628 56866 13638 56922
rect 13190 56798 13638 56866
rect 13190 56742 13200 56798
rect 13256 56742 13324 56798
rect 13380 56742 13448 56798
rect 13504 56742 13572 56798
rect 13628 56742 13638 56798
rect 13190 56674 13638 56742
rect 13190 56618 13200 56674
rect 13256 56618 13324 56674
rect 13380 56618 13448 56674
rect 13504 56618 13572 56674
rect 13628 56618 13638 56674
rect 13190 56550 13638 56618
rect 13190 56494 13200 56550
rect 13256 56494 13324 56550
rect 13380 56494 13448 56550
rect 13504 56494 13572 56550
rect 13628 56494 13638 56550
rect 13190 56426 13638 56494
rect 13190 56370 13200 56426
rect 13256 56370 13324 56426
rect 13380 56370 13448 56426
rect 13504 56370 13572 56426
rect 13628 56370 13638 56426
rect 13190 56302 13638 56370
rect 13190 56246 13200 56302
rect 13256 56246 13324 56302
rect 13380 56246 13448 56302
rect 13504 56246 13572 56302
rect 13628 56246 13638 56302
rect 13190 56178 13638 56246
rect 13190 56122 13200 56178
rect 13256 56122 13324 56178
rect 13380 56122 13448 56178
rect 13504 56122 13572 56178
rect 13628 56122 13638 56178
rect 13190 56054 13638 56122
rect 13190 55998 13200 56054
rect 13256 55998 13324 56054
rect 13380 55998 13448 56054
rect 13504 55998 13572 56054
rect 13628 55998 13638 56054
rect 13190 55930 13638 55998
rect 13190 55874 13200 55930
rect 13256 55874 13324 55930
rect 13380 55874 13448 55930
rect 13504 55874 13572 55930
rect 13628 55874 13638 55930
rect 13190 55806 13638 55874
rect 13190 55750 13200 55806
rect 13256 55750 13324 55806
rect 13380 55750 13448 55806
rect 13504 55750 13572 55806
rect 13628 55750 13638 55806
rect 13190 55740 13638 55750
rect 14326 56922 14774 56932
rect 14326 56866 14336 56922
rect 14392 56866 14460 56922
rect 14516 56866 14584 56922
rect 14640 56866 14708 56922
rect 14764 56866 14774 56922
rect 14326 56798 14774 56866
rect 14326 56742 14336 56798
rect 14392 56742 14460 56798
rect 14516 56742 14584 56798
rect 14640 56742 14708 56798
rect 14764 56742 14774 56798
rect 14326 56674 14774 56742
rect 14326 56618 14336 56674
rect 14392 56618 14460 56674
rect 14516 56618 14584 56674
rect 14640 56618 14708 56674
rect 14764 56618 14774 56674
rect 14326 56550 14774 56618
rect 14326 56494 14336 56550
rect 14392 56494 14460 56550
rect 14516 56494 14584 56550
rect 14640 56494 14708 56550
rect 14764 56494 14774 56550
rect 14326 56426 14774 56494
rect 14326 56370 14336 56426
rect 14392 56370 14460 56426
rect 14516 56370 14584 56426
rect 14640 56370 14708 56426
rect 14764 56370 14774 56426
rect 14326 56302 14774 56370
rect 14326 56246 14336 56302
rect 14392 56246 14460 56302
rect 14516 56246 14584 56302
rect 14640 56246 14708 56302
rect 14764 56246 14774 56302
rect 14326 56178 14774 56246
rect 14326 56122 14336 56178
rect 14392 56122 14460 56178
rect 14516 56122 14584 56178
rect 14640 56122 14708 56178
rect 14764 56122 14774 56178
rect 14326 56054 14774 56122
rect 14326 55998 14336 56054
rect 14392 55998 14460 56054
rect 14516 55998 14584 56054
rect 14640 55998 14708 56054
rect 14764 55998 14774 56054
rect 14326 55930 14774 55998
rect 14326 55874 14336 55930
rect 14392 55874 14460 55930
rect 14516 55874 14584 55930
rect 14640 55874 14708 55930
rect 14764 55874 14774 55930
rect 14326 55806 14774 55874
rect 14326 55750 14336 55806
rect 14392 55750 14460 55806
rect 14516 55750 14584 55806
rect 14640 55750 14708 55806
rect 14764 55750 14774 55806
rect 14326 55740 14774 55750
rect 858 55445 1306 55455
rect 858 55389 868 55445
rect 924 55389 992 55445
rect 1048 55389 1116 55445
rect 1172 55389 1240 55445
rect 1296 55389 1306 55445
rect 858 55321 1306 55389
rect 858 55265 868 55321
rect 924 55265 992 55321
rect 1048 55265 1116 55321
rect 1172 55265 1240 55321
rect 1296 55265 1306 55321
rect 858 55197 1306 55265
rect 858 55141 868 55197
rect 924 55141 992 55197
rect 1048 55141 1116 55197
rect 1172 55141 1240 55197
rect 1296 55141 1306 55197
rect 858 55073 1306 55141
rect 858 55017 868 55073
rect 924 55017 992 55073
rect 1048 55017 1116 55073
rect 1172 55017 1240 55073
rect 1296 55017 1306 55073
rect 858 54949 1306 55017
rect 858 54893 868 54949
rect 924 54893 992 54949
rect 1048 54893 1116 54949
rect 1172 54893 1240 54949
rect 1296 54893 1306 54949
rect 858 54825 1306 54893
rect 858 54769 868 54825
rect 924 54769 992 54825
rect 1048 54769 1116 54825
rect 1172 54769 1240 54825
rect 1296 54769 1306 54825
rect 858 54701 1306 54769
rect 858 54645 868 54701
rect 924 54645 992 54701
rect 1048 54645 1116 54701
rect 1172 54645 1240 54701
rect 1296 54645 1306 54701
rect 858 54577 1306 54645
rect 858 54521 868 54577
rect 924 54521 992 54577
rect 1048 54521 1116 54577
rect 1172 54521 1240 54577
rect 1296 54521 1306 54577
rect 858 54453 1306 54521
rect 858 54397 868 54453
rect 924 54397 992 54453
rect 1048 54397 1116 54453
rect 1172 54397 1240 54453
rect 1296 54397 1306 54453
rect 858 54329 1306 54397
rect 858 54273 868 54329
rect 924 54273 992 54329
rect 1048 54273 1116 54329
rect 1172 54273 1240 54329
rect 1296 54273 1306 54329
rect 858 54205 1306 54273
rect 858 54149 868 54205
rect 924 54149 992 54205
rect 1048 54149 1116 54205
rect 1172 54149 1240 54205
rect 1296 54149 1306 54205
rect 858 54139 1306 54149
rect 1994 55445 2442 55455
rect 1994 55389 2004 55445
rect 2060 55389 2128 55445
rect 2184 55389 2252 55445
rect 2308 55389 2376 55445
rect 2432 55389 2442 55445
rect 1994 55321 2442 55389
rect 1994 55265 2004 55321
rect 2060 55265 2128 55321
rect 2184 55265 2252 55321
rect 2308 55265 2376 55321
rect 2432 55265 2442 55321
rect 1994 55197 2442 55265
rect 1994 55141 2004 55197
rect 2060 55141 2128 55197
rect 2184 55141 2252 55197
rect 2308 55141 2376 55197
rect 2432 55141 2442 55197
rect 1994 55073 2442 55141
rect 1994 55017 2004 55073
rect 2060 55017 2128 55073
rect 2184 55017 2252 55073
rect 2308 55017 2376 55073
rect 2432 55017 2442 55073
rect 1994 54949 2442 55017
rect 1994 54893 2004 54949
rect 2060 54893 2128 54949
rect 2184 54893 2252 54949
rect 2308 54893 2376 54949
rect 2432 54893 2442 54949
rect 1994 54825 2442 54893
rect 1994 54769 2004 54825
rect 2060 54769 2128 54825
rect 2184 54769 2252 54825
rect 2308 54769 2376 54825
rect 2432 54769 2442 54825
rect 1994 54701 2442 54769
rect 1994 54645 2004 54701
rect 2060 54645 2128 54701
rect 2184 54645 2252 54701
rect 2308 54645 2376 54701
rect 2432 54645 2442 54701
rect 1994 54577 2442 54645
rect 1994 54521 2004 54577
rect 2060 54521 2128 54577
rect 2184 54521 2252 54577
rect 2308 54521 2376 54577
rect 2432 54521 2442 54577
rect 1994 54453 2442 54521
rect 1994 54397 2004 54453
rect 2060 54397 2128 54453
rect 2184 54397 2252 54453
rect 2308 54397 2376 54453
rect 2432 54397 2442 54453
rect 1994 54329 2442 54397
rect 1994 54273 2004 54329
rect 2060 54273 2128 54329
rect 2184 54273 2252 54329
rect 2308 54273 2376 54329
rect 2432 54273 2442 54329
rect 1994 54205 2442 54273
rect 1994 54149 2004 54205
rect 2060 54149 2128 54205
rect 2184 54149 2252 54205
rect 2308 54149 2376 54205
rect 2432 54149 2442 54205
rect 1994 54139 2442 54149
rect 3698 55445 4146 55455
rect 3698 55389 3708 55445
rect 3764 55389 3832 55445
rect 3888 55389 3956 55445
rect 4012 55389 4080 55445
rect 4136 55389 4146 55445
rect 3698 55321 4146 55389
rect 3698 55265 3708 55321
rect 3764 55265 3832 55321
rect 3888 55265 3956 55321
rect 4012 55265 4080 55321
rect 4136 55265 4146 55321
rect 3698 55197 4146 55265
rect 3698 55141 3708 55197
rect 3764 55141 3832 55197
rect 3888 55141 3956 55197
rect 4012 55141 4080 55197
rect 4136 55141 4146 55197
rect 3698 55073 4146 55141
rect 3698 55017 3708 55073
rect 3764 55017 3832 55073
rect 3888 55017 3956 55073
rect 4012 55017 4080 55073
rect 4136 55017 4146 55073
rect 3698 54949 4146 55017
rect 3698 54893 3708 54949
rect 3764 54893 3832 54949
rect 3888 54893 3956 54949
rect 4012 54893 4080 54949
rect 4136 54893 4146 54949
rect 3698 54825 4146 54893
rect 3698 54769 3708 54825
rect 3764 54769 3832 54825
rect 3888 54769 3956 54825
rect 4012 54769 4080 54825
rect 4136 54769 4146 54825
rect 3698 54701 4146 54769
rect 3698 54645 3708 54701
rect 3764 54645 3832 54701
rect 3888 54645 3956 54701
rect 4012 54645 4080 54701
rect 4136 54645 4146 54701
rect 3698 54577 4146 54645
rect 3698 54521 3708 54577
rect 3764 54521 3832 54577
rect 3888 54521 3956 54577
rect 4012 54521 4080 54577
rect 4136 54521 4146 54577
rect 3698 54453 4146 54521
rect 3698 54397 3708 54453
rect 3764 54397 3832 54453
rect 3888 54397 3956 54453
rect 4012 54397 4080 54453
rect 4136 54397 4146 54453
rect 3698 54329 4146 54397
rect 3698 54273 3708 54329
rect 3764 54273 3832 54329
rect 3888 54273 3956 54329
rect 4012 54273 4080 54329
rect 4136 54273 4146 54329
rect 3698 54205 4146 54273
rect 3698 54149 3708 54205
rect 3764 54149 3832 54205
rect 3888 54149 3956 54205
rect 4012 54149 4080 54205
rect 4136 54149 4146 54205
rect 3698 54139 4146 54149
rect 5970 55445 6418 55455
rect 5970 55389 5980 55445
rect 6036 55389 6104 55445
rect 6160 55389 6228 55445
rect 6284 55389 6352 55445
rect 6408 55389 6418 55445
rect 5970 55321 6418 55389
rect 5970 55265 5980 55321
rect 6036 55265 6104 55321
rect 6160 55265 6228 55321
rect 6284 55265 6352 55321
rect 6408 55265 6418 55321
rect 5970 55197 6418 55265
rect 5970 55141 5980 55197
rect 6036 55141 6104 55197
rect 6160 55141 6228 55197
rect 6284 55141 6352 55197
rect 6408 55141 6418 55197
rect 5970 55073 6418 55141
rect 5970 55017 5980 55073
rect 6036 55017 6104 55073
rect 6160 55017 6228 55073
rect 6284 55017 6352 55073
rect 6408 55017 6418 55073
rect 5970 54949 6418 55017
rect 5970 54893 5980 54949
rect 6036 54893 6104 54949
rect 6160 54893 6228 54949
rect 6284 54893 6352 54949
rect 6408 54893 6418 54949
rect 5970 54825 6418 54893
rect 5970 54769 5980 54825
rect 6036 54769 6104 54825
rect 6160 54769 6228 54825
rect 6284 54769 6352 54825
rect 6408 54769 6418 54825
rect 5970 54701 6418 54769
rect 5970 54645 5980 54701
rect 6036 54645 6104 54701
rect 6160 54645 6228 54701
rect 6284 54645 6352 54701
rect 6408 54645 6418 54701
rect 5970 54577 6418 54645
rect 5970 54521 5980 54577
rect 6036 54521 6104 54577
rect 6160 54521 6228 54577
rect 6284 54521 6352 54577
rect 6408 54521 6418 54577
rect 5970 54453 6418 54521
rect 5970 54397 5980 54453
rect 6036 54397 6104 54453
rect 6160 54397 6228 54453
rect 6284 54397 6352 54453
rect 6408 54397 6418 54453
rect 5970 54329 6418 54397
rect 5970 54273 5980 54329
rect 6036 54273 6104 54329
rect 6160 54273 6228 54329
rect 6284 54273 6352 54329
rect 6408 54273 6418 54329
rect 5970 54205 6418 54273
rect 5970 54149 5980 54205
rect 6036 54149 6104 54205
rect 6160 54149 6228 54205
rect 6284 54149 6352 54205
rect 6408 54149 6418 54205
rect 5970 54139 6418 54149
rect 8646 55445 9094 55455
rect 8646 55389 8656 55445
rect 8712 55389 8780 55445
rect 8836 55389 8904 55445
rect 8960 55389 9028 55445
rect 9084 55389 9094 55445
rect 8646 55321 9094 55389
rect 8646 55265 8656 55321
rect 8712 55265 8780 55321
rect 8836 55265 8904 55321
rect 8960 55265 9028 55321
rect 9084 55265 9094 55321
rect 8646 55197 9094 55265
rect 8646 55141 8656 55197
rect 8712 55141 8780 55197
rect 8836 55141 8904 55197
rect 8960 55141 9028 55197
rect 9084 55141 9094 55197
rect 8646 55073 9094 55141
rect 8646 55017 8656 55073
rect 8712 55017 8780 55073
rect 8836 55017 8904 55073
rect 8960 55017 9028 55073
rect 9084 55017 9094 55073
rect 8646 54949 9094 55017
rect 8646 54893 8656 54949
rect 8712 54893 8780 54949
rect 8836 54893 8904 54949
rect 8960 54893 9028 54949
rect 9084 54893 9094 54949
rect 8646 54825 9094 54893
rect 8646 54769 8656 54825
rect 8712 54769 8780 54825
rect 8836 54769 8904 54825
rect 8960 54769 9028 54825
rect 9084 54769 9094 54825
rect 8646 54701 9094 54769
rect 8646 54645 8656 54701
rect 8712 54645 8780 54701
rect 8836 54645 8904 54701
rect 8960 54645 9028 54701
rect 9084 54645 9094 54701
rect 8646 54577 9094 54645
rect 8646 54521 8656 54577
rect 8712 54521 8780 54577
rect 8836 54521 8904 54577
rect 8960 54521 9028 54577
rect 9084 54521 9094 54577
rect 8646 54453 9094 54521
rect 8646 54397 8656 54453
rect 8712 54397 8780 54453
rect 8836 54397 8904 54453
rect 8960 54397 9028 54453
rect 9084 54397 9094 54453
rect 8646 54329 9094 54397
rect 8646 54273 8656 54329
rect 8712 54273 8780 54329
rect 8836 54273 8904 54329
rect 8960 54273 9028 54329
rect 9084 54273 9094 54329
rect 8646 54205 9094 54273
rect 8646 54149 8656 54205
rect 8712 54149 8780 54205
rect 8836 54149 8904 54205
rect 8960 54149 9028 54205
rect 9084 54149 9094 54205
rect 8646 54139 9094 54149
rect 10918 55445 11366 55455
rect 10918 55389 10928 55445
rect 10984 55389 11052 55445
rect 11108 55389 11176 55445
rect 11232 55389 11300 55445
rect 11356 55389 11366 55445
rect 10918 55321 11366 55389
rect 10918 55265 10928 55321
rect 10984 55265 11052 55321
rect 11108 55265 11176 55321
rect 11232 55265 11300 55321
rect 11356 55265 11366 55321
rect 10918 55197 11366 55265
rect 10918 55141 10928 55197
rect 10984 55141 11052 55197
rect 11108 55141 11176 55197
rect 11232 55141 11300 55197
rect 11356 55141 11366 55197
rect 10918 55073 11366 55141
rect 10918 55017 10928 55073
rect 10984 55017 11052 55073
rect 11108 55017 11176 55073
rect 11232 55017 11300 55073
rect 11356 55017 11366 55073
rect 10918 54949 11366 55017
rect 10918 54893 10928 54949
rect 10984 54893 11052 54949
rect 11108 54893 11176 54949
rect 11232 54893 11300 54949
rect 11356 54893 11366 54949
rect 10918 54825 11366 54893
rect 10918 54769 10928 54825
rect 10984 54769 11052 54825
rect 11108 54769 11176 54825
rect 11232 54769 11300 54825
rect 11356 54769 11366 54825
rect 10918 54701 11366 54769
rect 10918 54645 10928 54701
rect 10984 54645 11052 54701
rect 11108 54645 11176 54701
rect 11232 54645 11300 54701
rect 11356 54645 11366 54701
rect 10918 54577 11366 54645
rect 10918 54521 10928 54577
rect 10984 54521 11052 54577
rect 11108 54521 11176 54577
rect 11232 54521 11300 54577
rect 11356 54521 11366 54577
rect 10918 54453 11366 54521
rect 10918 54397 10928 54453
rect 10984 54397 11052 54453
rect 11108 54397 11176 54453
rect 11232 54397 11300 54453
rect 11356 54397 11366 54453
rect 10918 54329 11366 54397
rect 10918 54273 10928 54329
rect 10984 54273 11052 54329
rect 11108 54273 11176 54329
rect 11232 54273 11300 54329
rect 11356 54273 11366 54329
rect 10918 54205 11366 54273
rect 10918 54149 10928 54205
rect 10984 54149 11052 54205
rect 11108 54149 11176 54205
rect 11232 54149 11300 54205
rect 11356 54149 11366 54205
rect 10918 54139 11366 54149
rect 12622 55445 13070 55455
rect 12622 55389 12632 55445
rect 12688 55389 12756 55445
rect 12812 55389 12880 55445
rect 12936 55389 13004 55445
rect 13060 55389 13070 55445
rect 12622 55321 13070 55389
rect 12622 55265 12632 55321
rect 12688 55265 12756 55321
rect 12812 55265 12880 55321
rect 12936 55265 13004 55321
rect 13060 55265 13070 55321
rect 12622 55197 13070 55265
rect 12622 55141 12632 55197
rect 12688 55141 12756 55197
rect 12812 55141 12880 55197
rect 12936 55141 13004 55197
rect 13060 55141 13070 55197
rect 12622 55073 13070 55141
rect 12622 55017 12632 55073
rect 12688 55017 12756 55073
rect 12812 55017 12880 55073
rect 12936 55017 13004 55073
rect 13060 55017 13070 55073
rect 12622 54949 13070 55017
rect 12622 54893 12632 54949
rect 12688 54893 12756 54949
rect 12812 54893 12880 54949
rect 12936 54893 13004 54949
rect 13060 54893 13070 54949
rect 12622 54825 13070 54893
rect 12622 54769 12632 54825
rect 12688 54769 12756 54825
rect 12812 54769 12880 54825
rect 12936 54769 13004 54825
rect 13060 54769 13070 54825
rect 12622 54701 13070 54769
rect 12622 54645 12632 54701
rect 12688 54645 12756 54701
rect 12812 54645 12880 54701
rect 12936 54645 13004 54701
rect 13060 54645 13070 54701
rect 12622 54577 13070 54645
rect 12622 54521 12632 54577
rect 12688 54521 12756 54577
rect 12812 54521 12880 54577
rect 12936 54521 13004 54577
rect 13060 54521 13070 54577
rect 12622 54453 13070 54521
rect 12622 54397 12632 54453
rect 12688 54397 12756 54453
rect 12812 54397 12880 54453
rect 12936 54397 13004 54453
rect 13060 54397 13070 54453
rect 12622 54329 13070 54397
rect 12622 54273 12632 54329
rect 12688 54273 12756 54329
rect 12812 54273 12880 54329
rect 12936 54273 13004 54329
rect 13060 54273 13070 54329
rect 12622 54205 13070 54273
rect 12622 54149 12632 54205
rect 12688 54149 12756 54205
rect 12812 54149 12880 54205
rect 12936 54149 13004 54205
rect 13060 54149 13070 54205
rect 12622 54139 13070 54149
rect 13758 55445 14206 55455
rect 13758 55389 13768 55445
rect 13824 55389 13892 55445
rect 13948 55389 14016 55445
rect 14072 55389 14140 55445
rect 14196 55389 14206 55445
rect 13758 55321 14206 55389
rect 13758 55265 13768 55321
rect 13824 55265 13892 55321
rect 13948 55265 14016 55321
rect 14072 55265 14140 55321
rect 14196 55265 14206 55321
rect 13758 55197 14206 55265
rect 13758 55141 13768 55197
rect 13824 55141 13892 55197
rect 13948 55141 14016 55197
rect 14072 55141 14140 55197
rect 14196 55141 14206 55197
rect 13758 55073 14206 55141
rect 13758 55017 13768 55073
rect 13824 55017 13892 55073
rect 13948 55017 14016 55073
rect 14072 55017 14140 55073
rect 14196 55017 14206 55073
rect 13758 54949 14206 55017
rect 13758 54893 13768 54949
rect 13824 54893 13892 54949
rect 13948 54893 14016 54949
rect 14072 54893 14140 54949
rect 14196 54893 14206 54949
rect 13758 54825 14206 54893
rect 13758 54769 13768 54825
rect 13824 54769 13892 54825
rect 13948 54769 14016 54825
rect 14072 54769 14140 54825
rect 14196 54769 14206 54825
rect 13758 54701 14206 54769
rect 13758 54645 13768 54701
rect 13824 54645 13892 54701
rect 13948 54645 14016 54701
rect 14072 54645 14140 54701
rect 14196 54645 14206 54701
rect 13758 54577 14206 54645
rect 13758 54521 13768 54577
rect 13824 54521 13892 54577
rect 13948 54521 14016 54577
rect 14072 54521 14140 54577
rect 14196 54521 14206 54577
rect 13758 54453 14206 54521
rect 13758 54397 13768 54453
rect 13824 54397 13892 54453
rect 13948 54397 14016 54453
rect 14072 54397 14140 54453
rect 14196 54397 14206 54453
rect 13758 54329 14206 54397
rect 13758 54273 13768 54329
rect 13824 54273 13892 54329
rect 13948 54273 14016 54329
rect 14072 54273 14140 54329
rect 14196 54273 14206 54329
rect 13758 54205 14206 54273
rect 13758 54149 13768 54205
rect 13824 54149 13892 54205
rect 13948 54149 14016 54205
rect 14072 54149 14140 54205
rect 14196 54149 14206 54205
rect 13758 54139 14206 54149
rect 290 53845 738 53855
rect 290 53789 300 53845
rect 356 53789 424 53845
rect 480 53789 548 53845
rect 604 53789 672 53845
rect 728 53789 738 53845
rect 290 53721 738 53789
rect 290 53665 300 53721
rect 356 53665 424 53721
rect 480 53665 548 53721
rect 604 53665 672 53721
rect 728 53665 738 53721
rect 290 53597 738 53665
rect 290 53541 300 53597
rect 356 53541 424 53597
rect 480 53541 548 53597
rect 604 53541 672 53597
rect 728 53541 738 53597
rect 290 53473 738 53541
rect 290 53417 300 53473
rect 356 53417 424 53473
rect 480 53417 548 53473
rect 604 53417 672 53473
rect 728 53417 738 53473
rect 290 53349 738 53417
rect 290 53293 300 53349
rect 356 53293 424 53349
rect 480 53293 548 53349
rect 604 53293 672 53349
rect 728 53293 738 53349
rect 290 53225 738 53293
rect 290 53169 300 53225
rect 356 53169 424 53225
rect 480 53169 548 53225
rect 604 53169 672 53225
rect 728 53169 738 53225
rect 290 53101 738 53169
rect 290 53045 300 53101
rect 356 53045 424 53101
rect 480 53045 548 53101
rect 604 53045 672 53101
rect 728 53045 738 53101
rect 290 52977 738 53045
rect 290 52921 300 52977
rect 356 52921 424 52977
rect 480 52921 548 52977
rect 604 52921 672 52977
rect 728 52921 738 52977
rect 290 52853 738 52921
rect 290 52797 300 52853
rect 356 52797 424 52853
rect 480 52797 548 52853
rect 604 52797 672 52853
rect 728 52797 738 52853
rect 290 52729 738 52797
rect 290 52673 300 52729
rect 356 52673 424 52729
rect 480 52673 548 52729
rect 604 52673 672 52729
rect 728 52673 738 52729
rect 290 52605 738 52673
rect 290 52549 300 52605
rect 356 52549 424 52605
rect 480 52549 548 52605
rect 604 52549 672 52605
rect 728 52549 738 52605
rect 290 52539 738 52549
rect 1426 53845 1874 53855
rect 1426 53789 1436 53845
rect 1492 53789 1560 53845
rect 1616 53789 1684 53845
rect 1740 53789 1808 53845
rect 1864 53789 1874 53845
rect 1426 53721 1874 53789
rect 1426 53665 1436 53721
rect 1492 53665 1560 53721
rect 1616 53665 1684 53721
rect 1740 53665 1808 53721
rect 1864 53665 1874 53721
rect 1426 53597 1874 53665
rect 1426 53541 1436 53597
rect 1492 53541 1560 53597
rect 1616 53541 1684 53597
rect 1740 53541 1808 53597
rect 1864 53541 1874 53597
rect 1426 53473 1874 53541
rect 1426 53417 1436 53473
rect 1492 53417 1560 53473
rect 1616 53417 1684 53473
rect 1740 53417 1808 53473
rect 1864 53417 1874 53473
rect 1426 53349 1874 53417
rect 1426 53293 1436 53349
rect 1492 53293 1560 53349
rect 1616 53293 1684 53349
rect 1740 53293 1808 53349
rect 1864 53293 1874 53349
rect 1426 53225 1874 53293
rect 1426 53169 1436 53225
rect 1492 53169 1560 53225
rect 1616 53169 1684 53225
rect 1740 53169 1808 53225
rect 1864 53169 1874 53225
rect 1426 53101 1874 53169
rect 1426 53045 1436 53101
rect 1492 53045 1560 53101
rect 1616 53045 1684 53101
rect 1740 53045 1808 53101
rect 1864 53045 1874 53101
rect 1426 52977 1874 53045
rect 1426 52921 1436 52977
rect 1492 52921 1560 52977
rect 1616 52921 1684 52977
rect 1740 52921 1808 52977
rect 1864 52921 1874 52977
rect 1426 52853 1874 52921
rect 1426 52797 1436 52853
rect 1492 52797 1560 52853
rect 1616 52797 1684 52853
rect 1740 52797 1808 52853
rect 1864 52797 1874 52853
rect 1426 52729 1874 52797
rect 1426 52673 1436 52729
rect 1492 52673 1560 52729
rect 1616 52673 1684 52729
rect 1740 52673 1808 52729
rect 1864 52673 1874 52729
rect 1426 52605 1874 52673
rect 1426 52549 1436 52605
rect 1492 52549 1560 52605
rect 1616 52549 1684 52605
rect 1740 52549 1808 52605
rect 1864 52549 1874 52605
rect 1426 52539 1874 52549
rect 2562 53845 3010 53855
rect 2562 53789 2572 53845
rect 2628 53789 2696 53845
rect 2752 53789 2820 53845
rect 2876 53789 2944 53845
rect 3000 53789 3010 53845
rect 2562 53721 3010 53789
rect 2562 53665 2572 53721
rect 2628 53665 2696 53721
rect 2752 53665 2820 53721
rect 2876 53665 2944 53721
rect 3000 53665 3010 53721
rect 2562 53597 3010 53665
rect 2562 53541 2572 53597
rect 2628 53541 2696 53597
rect 2752 53541 2820 53597
rect 2876 53541 2944 53597
rect 3000 53541 3010 53597
rect 2562 53473 3010 53541
rect 2562 53417 2572 53473
rect 2628 53417 2696 53473
rect 2752 53417 2820 53473
rect 2876 53417 2944 53473
rect 3000 53417 3010 53473
rect 2562 53349 3010 53417
rect 2562 53293 2572 53349
rect 2628 53293 2696 53349
rect 2752 53293 2820 53349
rect 2876 53293 2944 53349
rect 3000 53293 3010 53349
rect 2562 53225 3010 53293
rect 2562 53169 2572 53225
rect 2628 53169 2696 53225
rect 2752 53169 2820 53225
rect 2876 53169 2944 53225
rect 3000 53169 3010 53225
rect 2562 53101 3010 53169
rect 2562 53045 2572 53101
rect 2628 53045 2696 53101
rect 2752 53045 2820 53101
rect 2876 53045 2944 53101
rect 3000 53045 3010 53101
rect 2562 52977 3010 53045
rect 2562 52921 2572 52977
rect 2628 52921 2696 52977
rect 2752 52921 2820 52977
rect 2876 52921 2944 52977
rect 3000 52921 3010 52977
rect 2562 52853 3010 52921
rect 2562 52797 2572 52853
rect 2628 52797 2696 52853
rect 2752 52797 2820 52853
rect 2876 52797 2944 52853
rect 3000 52797 3010 52853
rect 2562 52729 3010 52797
rect 2562 52673 2572 52729
rect 2628 52673 2696 52729
rect 2752 52673 2820 52729
rect 2876 52673 2944 52729
rect 3000 52673 3010 52729
rect 2562 52605 3010 52673
rect 2562 52549 2572 52605
rect 2628 52549 2696 52605
rect 2752 52549 2820 52605
rect 2876 52549 2944 52605
rect 3000 52549 3010 52605
rect 2562 52539 3010 52549
rect 4834 53845 5282 53855
rect 4834 53789 4844 53845
rect 4900 53789 4968 53845
rect 5024 53789 5092 53845
rect 5148 53789 5216 53845
rect 5272 53789 5282 53845
rect 4834 53721 5282 53789
rect 4834 53665 4844 53721
rect 4900 53665 4968 53721
rect 5024 53665 5092 53721
rect 5148 53665 5216 53721
rect 5272 53665 5282 53721
rect 4834 53597 5282 53665
rect 4834 53541 4844 53597
rect 4900 53541 4968 53597
rect 5024 53541 5092 53597
rect 5148 53541 5216 53597
rect 5272 53541 5282 53597
rect 4834 53473 5282 53541
rect 4834 53417 4844 53473
rect 4900 53417 4968 53473
rect 5024 53417 5092 53473
rect 5148 53417 5216 53473
rect 5272 53417 5282 53473
rect 4834 53349 5282 53417
rect 4834 53293 4844 53349
rect 4900 53293 4968 53349
rect 5024 53293 5092 53349
rect 5148 53293 5216 53349
rect 5272 53293 5282 53349
rect 4834 53225 5282 53293
rect 4834 53169 4844 53225
rect 4900 53169 4968 53225
rect 5024 53169 5092 53225
rect 5148 53169 5216 53225
rect 5272 53169 5282 53225
rect 4834 53101 5282 53169
rect 4834 53045 4844 53101
rect 4900 53045 4968 53101
rect 5024 53045 5092 53101
rect 5148 53045 5216 53101
rect 5272 53045 5282 53101
rect 4834 52977 5282 53045
rect 4834 52921 4844 52977
rect 4900 52921 4968 52977
rect 5024 52921 5092 52977
rect 5148 52921 5216 52977
rect 5272 52921 5282 52977
rect 4834 52853 5282 52921
rect 4834 52797 4844 52853
rect 4900 52797 4968 52853
rect 5024 52797 5092 52853
rect 5148 52797 5216 52853
rect 5272 52797 5282 52853
rect 4834 52729 5282 52797
rect 4834 52673 4844 52729
rect 4900 52673 4968 52729
rect 5024 52673 5092 52729
rect 5148 52673 5216 52729
rect 5272 52673 5282 52729
rect 4834 52605 5282 52673
rect 4834 52549 4844 52605
rect 4900 52549 4968 52605
rect 5024 52549 5092 52605
rect 5148 52549 5216 52605
rect 5272 52549 5282 52605
rect 4834 52539 5282 52549
rect 7127 53845 7451 53855
rect 7127 53789 7137 53845
rect 7193 53789 7261 53845
rect 7317 53789 7385 53845
rect 7441 53789 7451 53845
rect 7127 53721 7451 53789
rect 7127 53665 7137 53721
rect 7193 53665 7261 53721
rect 7317 53665 7385 53721
rect 7441 53665 7451 53721
rect 7127 53597 7451 53665
rect 7127 53541 7137 53597
rect 7193 53541 7261 53597
rect 7317 53541 7385 53597
rect 7441 53541 7451 53597
rect 7127 53473 7451 53541
rect 7127 53417 7137 53473
rect 7193 53417 7261 53473
rect 7317 53417 7385 53473
rect 7441 53417 7451 53473
rect 7127 53349 7451 53417
rect 7127 53293 7137 53349
rect 7193 53293 7261 53349
rect 7317 53293 7385 53349
rect 7441 53293 7451 53349
rect 7127 53225 7451 53293
rect 7127 53169 7137 53225
rect 7193 53169 7261 53225
rect 7317 53169 7385 53225
rect 7441 53169 7451 53225
rect 7127 53101 7451 53169
rect 7127 53045 7137 53101
rect 7193 53045 7261 53101
rect 7317 53045 7385 53101
rect 7441 53045 7451 53101
rect 7127 52977 7451 53045
rect 7127 52921 7137 52977
rect 7193 52921 7261 52977
rect 7317 52921 7385 52977
rect 7441 52921 7451 52977
rect 7127 52853 7451 52921
rect 7127 52797 7137 52853
rect 7193 52797 7261 52853
rect 7317 52797 7385 52853
rect 7441 52797 7451 52853
rect 7127 52729 7451 52797
rect 7127 52673 7137 52729
rect 7193 52673 7261 52729
rect 7317 52673 7385 52729
rect 7441 52673 7451 52729
rect 7127 52605 7451 52673
rect 7127 52549 7137 52605
rect 7193 52549 7261 52605
rect 7317 52549 7385 52605
rect 7441 52549 7451 52605
rect 7127 52539 7451 52549
rect 7613 53845 7937 53855
rect 7613 53789 7623 53845
rect 7679 53789 7747 53845
rect 7803 53789 7871 53845
rect 7927 53789 7937 53845
rect 7613 53721 7937 53789
rect 7613 53665 7623 53721
rect 7679 53665 7747 53721
rect 7803 53665 7871 53721
rect 7927 53665 7937 53721
rect 7613 53597 7937 53665
rect 7613 53541 7623 53597
rect 7679 53541 7747 53597
rect 7803 53541 7871 53597
rect 7927 53541 7937 53597
rect 7613 53473 7937 53541
rect 7613 53417 7623 53473
rect 7679 53417 7747 53473
rect 7803 53417 7871 53473
rect 7927 53417 7937 53473
rect 7613 53349 7937 53417
rect 7613 53293 7623 53349
rect 7679 53293 7747 53349
rect 7803 53293 7871 53349
rect 7927 53293 7937 53349
rect 7613 53225 7937 53293
rect 7613 53169 7623 53225
rect 7679 53169 7747 53225
rect 7803 53169 7871 53225
rect 7927 53169 7937 53225
rect 7613 53101 7937 53169
rect 7613 53045 7623 53101
rect 7679 53045 7747 53101
rect 7803 53045 7871 53101
rect 7927 53045 7937 53101
rect 7613 52977 7937 53045
rect 7613 52921 7623 52977
rect 7679 52921 7747 52977
rect 7803 52921 7871 52977
rect 7927 52921 7937 52977
rect 7613 52853 7937 52921
rect 7613 52797 7623 52853
rect 7679 52797 7747 52853
rect 7803 52797 7871 52853
rect 7927 52797 7937 52853
rect 7613 52729 7937 52797
rect 7613 52673 7623 52729
rect 7679 52673 7747 52729
rect 7803 52673 7871 52729
rect 7927 52673 7937 52729
rect 7613 52605 7937 52673
rect 7613 52549 7623 52605
rect 7679 52549 7747 52605
rect 7803 52549 7871 52605
rect 7927 52549 7937 52605
rect 7613 52539 7937 52549
rect 9782 53845 10230 53855
rect 9782 53789 9792 53845
rect 9848 53789 9916 53845
rect 9972 53789 10040 53845
rect 10096 53789 10164 53845
rect 10220 53789 10230 53845
rect 9782 53721 10230 53789
rect 9782 53665 9792 53721
rect 9848 53665 9916 53721
rect 9972 53665 10040 53721
rect 10096 53665 10164 53721
rect 10220 53665 10230 53721
rect 9782 53597 10230 53665
rect 9782 53541 9792 53597
rect 9848 53541 9916 53597
rect 9972 53541 10040 53597
rect 10096 53541 10164 53597
rect 10220 53541 10230 53597
rect 9782 53473 10230 53541
rect 9782 53417 9792 53473
rect 9848 53417 9916 53473
rect 9972 53417 10040 53473
rect 10096 53417 10164 53473
rect 10220 53417 10230 53473
rect 9782 53349 10230 53417
rect 9782 53293 9792 53349
rect 9848 53293 9916 53349
rect 9972 53293 10040 53349
rect 10096 53293 10164 53349
rect 10220 53293 10230 53349
rect 9782 53225 10230 53293
rect 9782 53169 9792 53225
rect 9848 53169 9916 53225
rect 9972 53169 10040 53225
rect 10096 53169 10164 53225
rect 10220 53169 10230 53225
rect 9782 53101 10230 53169
rect 9782 53045 9792 53101
rect 9848 53045 9916 53101
rect 9972 53045 10040 53101
rect 10096 53045 10164 53101
rect 10220 53045 10230 53101
rect 9782 52977 10230 53045
rect 9782 52921 9792 52977
rect 9848 52921 9916 52977
rect 9972 52921 10040 52977
rect 10096 52921 10164 52977
rect 10220 52921 10230 52977
rect 9782 52853 10230 52921
rect 9782 52797 9792 52853
rect 9848 52797 9916 52853
rect 9972 52797 10040 52853
rect 10096 52797 10164 52853
rect 10220 52797 10230 52853
rect 9782 52729 10230 52797
rect 9782 52673 9792 52729
rect 9848 52673 9916 52729
rect 9972 52673 10040 52729
rect 10096 52673 10164 52729
rect 10220 52673 10230 52729
rect 9782 52605 10230 52673
rect 9782 52549 9792 52605
rect 9848 52549 9916 52605
rect 9972 52549 10040 52605
rect 10096 52549 10164 52605
rect 10220 52549 10230 52605
rect 9782 52539 10230 52549
rect 12054 53845 12502 53855
rect 12054 53789 12064 53845
rect 12120 53789 12188 53845
rect 12244 53789 12312 53845
rect 12368 53789 12436 53845
rect 12492 53789 12502 53845
rect 12054 53721 12502 53789
rect 12054 53665 12064 53721
rect 12120 53665 12188 53721
rect 12244 53665 12312 53721
rect 12368 53665 12436 53721
rect 12492 53665 12502 53721
rect 12054 53597 12502 53665
rect 12054 53541 12064 53597
rect 12120 53541 12188 53597
rect 12244 53541 12312 53597
rect 12368 53541 12436 53597
rect 12492 53541 12502 53597
rect 12054 53473 12502 53541
rect 12054 53417 12064 53473
rect 12120 53417 12188 53473
rect 12244 53417 12312 53473
rect 12368 53417 12436 53473
rect 12492 53417 12502 53473
rect 12054 53349 12502 53417
rect 12054 53293 12064 53349
rect 12120 53293 12188 53349
rect 12244 53293 12312 53349
rect 12368 53293 12436 53349
rect 12492 53293 12502 53349
rect 12054 53225 12502 53293
rect 12054 53169 12064 53225
rect 12120 53169 12188 53225
rect 12244 53169 12312 53225
rect 12368 53169 12436 53225
rect 12492 53169 12502 53225
rect 12054 53101 12502 53169
rect 12054 53045 12064 53101
rect 12120 53045 12188 53101
rect 12244 53045 12312 53101
rect 12368 53045 12436 53101
rect 12492 53045 12502 53101
rect 12054 52977 12502 53045
rect 12054 52921 12064 52977
rect 12120 52921 12188 52977
rect 12244 52921 12312 52977
rect 12368 52921 12436 52977
rect 12492 52921 12502 52977
rect 12054 52853 12502 52921
rect 12054 52797 12064 52853
rect 12120 52797 12188 52853
rect 12244 52797 12312 52853
rect 12368 52797 12436 52853
rect 12492 52797 12502 52853
rect 12054 52729 12502 52797
rect 12054 52673 12064 52729
rect 12120 52673 12188 52729
rect 12244 52673 12312 52729
rect 12368 52673 12436 52729
rect 12492 52673 12502 52729
rect 12054 52605 12502 52673
rect 12054 52549 12064 52605
rect 12120 52549 12188 52605
rect 12244 52549 12312 52605
rect 12368 52549 12436 52605
rect 12492 52549 12502 52605
rect 12054 52539 12502 52549
rect 13190 53845 13638 53855
rect 13190 53789 13200 53845
rect 13256 53789 13324 53845
rect 13380 53789 13448 53845
rect 13504 53789 13572 53845
rect 13628 53789 13638 53845
rect 13190 53721 13638 53789
rect 13190 53665 13200 53721
rect 13256 53665 13324 53721
rect 13380 53665 13448 53721
rect 13504 53665 13572 53721
rect 13628 53665 13638 53721
rect 13190 53597 13638 53665
rect 13190 53541 13200 53597
rect 13256 53541 13324 53597
rect 13380 53541 13448 53597
rect 13504 53541 13572 53597
rect 13628 53541 13638 53597
rect 13190 53473 13638 53541
rect 13190 53417 13200 53473
rect 13256 53417 13324 53473
rect 13380 53417 13448 53473
rect 13504 53417 13572 53473
rect 13628 53417 13638 53473
rect 13190 53349 13638 53417
rect 13190 53293 13200 53349
rect 13256 53293 13324 53349
rect 13380 53293 13448 53349
rect 13504 53293 13572 53349
rect 13628 53293 13638 53349
rect 13190 53225 13638 53293
rect 13190 53169 13200 53225
rect 13256 53169 13324 53225
rect 13380 53169 13448 53225
rect 13504 53169 13572 53225
rect 13628 53169 13638 53225
rect 13190 53101 13638 53169
rect 13190 53045 13200 53101
rect 13256 53045 13324 53101
rect 13380 53045 13448 53101
rect 13504 53045 13572 53101
rect 13628 53045 13638 53101
rect 13190 52977 13638 53045
rect 13190 52921 13200 52977
rect 13256 52921 13324 52977
rect 13380 52921 13448 52977
rect 13504 52921 13572 52977
rect 13628 52921 13638 52977
rect 13190 52853 13638 52921
rect 13190 52797 13200 52853
rect 13256 52797 13324 52853
rect 13380 52797 13448 52853
rect 13504 52797 13572 52853
rect 13628 52797 13638 52853
rect 13190 52729 13638 52797
rect 13190 52673 13200 52729
rect 13256 52673 13324 52729
rect 13380 52673 13448 52729
rect 13504 52673 13572 52729
rect 13628 52673 13638 52729
rect 13190 52605 13638 52673
rect 13190 52549 13200 52605
rect 13256 52549 13324 52605
rect 13380 52549 13448 52605
rect 13504 52549 13572 52605
rect 13628 52549 13638 52605
rect 13190 52539 13638 52549
rect 14326 53845 14774 53855
rect 14326 53789 14336 53845
rect 14392 53789 14460 53845
rect 14516 53789 14584 53845
rect 14640 53789 14708 53845
rect 14764 53789 14774 53845
rect 14326 53721 14774 53789
rect 14326 53665 14336 53721
rect 14392 53665 14460 53721
rect 14516 53665 14584 53721
rect 14640 53665 14708 53721
rect 14764 53665 14774 53721
rect 14326 53597 14774 53665
rect 14326 53541 14336 53597
rect 14392 53541 14460 53597
rect 14516 53541 14584 53597
rect 14640 53541 14708 53597
rect 14764 53541 14774 53597
rect 14326 53473 14774 53541
rect 14326 53417 14336 53473
rect 14392 53417 14460 53473
rect 14516 53417 14584 53473
rect 14640 53417 14708 53473
rect 14764 53417 14774 53473
rect 14326 53349 14774 53417
rect 14326 53293 14336 53349
rect 14392 53293 14460 53349
rect 14516 53293 14584 53349
rect 14640 53293 14708 53349
rect 14764 53293 14774 53349
rect 14326 53225 14774 53293
rect 14326 53169 14336 53225
rect 14392 53169 14460 53225
rect 14516 53169 14584 53225
rect 14640 53169 14708 53225
rect 14764 53169 14774 53225
rect 14326 53101 14774 53169
rect 14326 53045 14336 53101
rect 14392 53045 14460 53101
rect 14516 53045 14584 53101
rect 14640 53045 14708 53101
rect 14764 53045 14774 53101
rect 14326 52977 14774 53045
rect 14326 52921 14336 52977
rect 14392 52921 14460 52977
rect 14516 52921 14584 52977
rect 14640 52921 14708 52977
rect 14764 52921 14774 52977
rect 14326 52853 14774 52921
rect 14326 52797 14336 52853
rect 14392 52797 14460 52853
rect 14516 52797 14584 52853
rect 14640 52797 14708 52853
rect 14764 52797 14774 52853
rect 14326 52729 14774 52797
rect 14326 52673 14336 52729
rect 14392 52673 14460 52729
rect 14516 52673 14584 52729
rect 14640 52673 14708 52729
rect 14764 52673 14774 52729
rect 14326 52605 14774 52673
rect 14326 52549 14336 52605
rect 14392 52549 14460 52605
rect 14516 52549 14584 52605
rect 14640 52549 14708 52605
rect 14764 52549 14774 52605
rect 14326 52539 14774 52549
rect 46 52273 122 52283
rect 46 50921 56 52273
rect 112 50921 122 52273
rect 14942 52273 15018 52283
rect 13160 52245 13360 52255
rect 13160 52189 13170 52245
rect 13226 52189 13294 52245
rect 13350 52189 13360 52245
rect 13160 52121 13360 52189
rect 13160 52065 13170 52121
rect 13226 52065 13294 52121
rect 13350 52065 13360 52121
rect 13160 51997 13360 52065
rect 13160 51941 13170 51997
rect 13226 51941 13294 51997
rect 13350 51941 13360 51997
rect 13160 51873 13360 51941
rect 13160 51817 13170 51873
rect 13226 51817 13294 51873
rect 13350 51817 13360 51873
rect 13160 51749 13360 51817
rect 13160 51693 13170 51749
rect 13226 51693 13294 51749
rect 13350 51693 13360 51749
rect 13160 51625 13360 51693
rect 13160 51569 13170 51625
rect 13226 51569 13294 51625
rect 13350 51569 13360 51625
rect 13160 51501 13360 51569
rect 13160 51445 13170 51501
rect 13226 51445 13294 51501
rect 13350 51445 13360 51501
rect 13160 51377 13360 51445
rect 13160 51321 13170 51377
rect 13226 51321 13294 51377
rect 13350 51321 13360 51377
rect 13160 51253 13360 51321
rect 13160 51197 13170 51253
rect 13226 51197 13294 51253
rect 13350 51197 13360 51253
rect 13160 51129 13360 51197
rect 13160 51073 13170 51129
rect 13226 51073 13294 51129
rect 13350 51073 13360 51129
rect 13160 51005 13360 51073
rect 13160 50949 13170 51005
rect 13226 50949 13294 51005
rect 13350 50949 13360 51005
rect 13160 50939 13360 50949
rect 46 50911 122 50921
rect 14942 50921 14952 52273
rect 15008 50921 15018 52273
rect 14942 50911 15018 50921
rect 828 50645 1028 50655
rect 828 50589 838 50645
rect 894 50589 962 50645
rect 1018 50589 1028 50645
rect 828 50521 1028 50589
rect 828 50465 838 50521
rect 894 50465 962 50521
rect 1018 50465 1028 50521
rect 828 50397 1028 50465
rect 828 50341 838 50397
rect 894 50341 962 50397
rect 1018 50341 1028 50397
rect 828 50273 1028 50341
rect 828 50217 838 50273
rect 894 50217 962 50273
rect 1018 50217 1028 50273
rect 828 50149 1028 50217
rect 828 50093 838 50149
rect 894 50093 962 50149
rect 1018 50093 1028 50149
rect 828 50025 1028 50093
rect 828 49969 838 50025
rect 894 49969 962 50025
rect 1018 49969 1028 50025
rect 828 49901 1028 49969
rect 828 49845 838 49901
rect 894 49845 962 49901
rect 1018 49845 1028 49901
rect 828 49777 1028 49845
rect 828 49721 838 49777
rect 894 49721 962 49777
rect 1018 49721 1028 49777
rect 828 49653 1028 49721
rect 828 49597 838 49653
rect 894 49597 962 49653
rect 1018 49597 1028 49653
rect 828 49529 1028 49597
rect 828 49473 838 49529
rect 894 49473 962 49529
rect 1018 49473 1028 49529
rect 828 49405 1028 49473
rect 828 49349 838 49405
rect 894 49349 962 49405
rect 1018 49349 1028 49405
rect 828 49339 1028 49349
rect 290 49045 738 49055
rect 290 48989 300 49045
rect 356 48989 424 49045
rect 480 48989 548 49045
rect 604 48989 672 49045
rect 728 48989 738 49045
rect 290 48921 738 48989
rect 290 48865 300 48921
rect 356 48865 424 48921
rect 480 48865 548 48921
rect 604 48865 672 48921
rect 728 48865 738 48921
rect 290 48797 738 48865
rect 290 48741 300 48797
rect 356 48741 424 48797
rect 480 48741 548 48797
rect 604 48741 672 48797
rect 728 48741 738 48797
rect 290 48673 738 48741
rect 290 48617 300 48673
rect 356 48617 424 48673
rect 480 48617 548 48673
rect 604 48617 672 48673
rect 728 48617 738 48673
rect 290 48549 738 48617
rect 290 48493 300 48549
rect 356 48493 424 48549
rect 480 48493 548 48549
rect 604 48493 672 48549
rect 728 48493 738 48549
rect 290 48425 738 48493
rect 290 48369 300 48425
rect 356 48369 424 48425
rect 480 48369 548 48425
rect 604 48369 672 48425
rect 728 48369 738 48425
rect 290 48301 738 48369
rect 290 48245 300 48301
rect 356 48245 424 48301
rect 480 48245 548 48301
rect 604 48245 672 48301
rect 728 48245 738 48301
rect 290 48177 738 48245
rect 290 48121 300 48177
rect 356 48121 424 48177
rect 480 48121 548 48177
rect 604 48121 672 48177
rect 728 48121 738 48177
rect 290 48053 738 48121
rect 290 47997 300 48053
rect 356 47997 424 48053
rect 480 47997 548 48053
rect 604 47997 672 48053
rect 728 47997 738 48053
rect 290 47929 738 47997
rect 290 47873 300 47929
rect 356 47873 424 47929
rect 480 47873 548 47929
rect 604 47873 672 47929
rect 728 47873 738 47929
rect 290 47805 738 47873
rect 290 47749 300 47805
rect 356 47749 424 47805
rect 480 47749 548 47805
rect 604 47749 672 47805
rect 728 47749 738 47805
rect 290 47739 738 47749
rect 1426 49045 1874 49055
rect 1426 48989 1436 49045
rect 1492 48989 1560 49045
rect 1616 48989 1684 49045
rect 1740 48989 1808 49045
rect 1864 48989 1874 49045
rect 1426 48921 1874 48989
rect 1426 48865 1436 48921
rect 1492 48865 1560 48921
rect 1616 48865 1684 48921
rect 1740 48865 1808 48921
rect 1864 48865 1874 48921
rect 1426 48797 1874 48865
rect 1426 48741 1436 48797
rect 1492 48741 1560 48797
rect 1616 48741 1684 48797
rect 1740 48741 1808 48797
rect 1864 48741 1874 48797
rect 1426 48673 1874 48741
rect 1426 48617 1436 48673
rect 1492 48617 1560 48673
rect 1616 48617 1684 48673
rect 1740 48617 1808 48673
rect 1864 48617 1874 48673
rect 1426 48549 1874 48617
rect 1426 48493 1436 48549
rect 1492 48493 1560 48549
rect 1616 48493 1684 48549
rect 1740 48493 1808 48549
rect 1864 48493 1874 48549
rect 1426 48425 1874 48493
rect 1426 48369 1436 48425
rect 1492 48369 1560 48425
rect 1616 48369 1684 48425
rect 1740 48369 1808 48425
rect 1864 48369 1874 48425
rect 1426 48301 1874 48369
rect 1426 48245 1436 48301
rect 1492 48245 1560 48301
rect 1616 48245 1684 48301
rect 1740 48245 1808 48301
rect 1864 48245 1874 48301
rect 1426 48177 1874 48245
rect 1426 48121 1436 48177
rect 1492 48121 1560 48177
rect 1616 48121 1684 48177
rect 1740 48121 1808 48177
rect 1864 48121 1874 48177
rect 1426 48053 1874 48121
rect 1426 47997 1436 48053
rect 1492 47997 1560 48053
rect 1616 47997 1684 48053
rect 1740 47997 1808 48053
rect 1864 47997 1874 48053
rect 1426 47929 1874 47997
rect 1426 47873 1436 47929
rect 1492 47873 1560 47929
rect 1616 47873 1684 47929
rect 1740 47873 1808 47929
rect 1864 47873 1874 47929
rect 1426 47805 1874 47873
rect 1426 47749 1436 47805
rect 1492 47749 1560 47805
rect 1616 47749 1684 47805
rect 1740 47749 1808 47805
rect 1864 47749 1874 47805
rect 1426 47739 1874 47749
rect 2562 49045 3010 49055
rect 2562 48989 2572 49045
rect 2628 48989 2696 49045
rect 2752 48989 2820 49045
rect 2876 48989 2944 49045
rect 3000 48989 3010 49045
rect 2562 48921 3010 48989
rect 2562 48865 2572 48921
rect 2628 48865 2696 48921
rect 2752 48865 2820 48921
rect 2876 48865 2944 48921
rect 3000 48865 3010 48921
rect 2562 48797 3010 48865
rect 2562 48741 2572 48797
rect 2628 48741 2696 48797
rect 2752 48741 2820 48797
rect 2876 48741 2944 48797
rect 3000 48741 3010 48797
rect 2562 48673 3010 48741
rect 2562 48617 2572 48673
rect 2628 48617 2696 48673
rect 2752 48617 2820 48673
rect 2876 48617 2944 48673
rect 3000 48617 3010 48673
rect 2562 48549 3010 48617
rect 2562 48493 2572 48549
rect 2628 48493 2696 48549
rect 2752 48493 2820 48549
rect 2876 48493 2944 48549
rect 3000 48493 3010 48549
rect 2562 48425 3010 48493
rect 2562 48369 2572 48425
rect 2628 48369 2696 48425
rect 2752 48369 2820 48425
rect 2876 48369 2944 48425
rect 3000 48369 3010 48425
rect 2562 48301 3010 48369
rect 2562 48245 2572 48301
rect 2628 48245 2696 48301
rect 2752 48245 2820 48301
rect 2876 48245 2944 48301
rect 3000 48245 3010 48301
rect 2562 48177 3010 48245
rect 2562 48121 2572 48177
rect 2628 48121 2696 48177
rect 2752 48121 2820 48177
rect 2876 48121 2944 48177
rect 3000 48121 3010 48177
rect 2562 48053 3010 48121
rect 2562 47997 2572 48053
rect 2628 47997 2696 48053
rect 2752 47997 2820 48053
rect 2876 47997 2944 48053
rect 3000 47997 3010 48053
rect 2562 47929 3010 47997
rect 2562 47873 2572 47929
rect 2628 47873 2696 47929
rect 2752 47873 2820 47929
rect 2876 47873 2944 47929
rect 3000 47873 3010 47929
rect 2562 47805 3010 47873
rect 2562 47749 2572 47805
rect 2628 47749 2696 47805
rect 2752 47749 2820 47805
rect 2876 47749 2944 47805
rect 3000 47749 3010 47805
rect 2562 47739 3010 47749
rect 4834 49045 5282 49055
rect 4834 48989 4844 49045
rect 4900 48989 4968 49045
rect 5024 48989 5092 49045
rect 5148 48989 5216 49045
rect 5272 48989 5282 49045
rect 4834 48921 5282 48989
rect 4834 48865 4844 48921
rect 4900 48865 4968 48921
rect 5024 48865 5092 48921
rect 5148 48865 5216 48921
rect 5272 48865 5282 48921
rect 4834 48797 5282 48865
rect 4834 48741 4844 48797
rect 4900 48741 4968 48797
rect 5024 48741 5092 48797
rect 5148 48741 5216 48797
rect 5272 48741 5282 48797
rect 4834 48673 5282 48741
rect 4834 48617 4844 48673
rect 4900 48617 4968 48673
rect 5024 48617 5092 48673
rect 5148 48617 5216 48673
rect 5272 48617 5282 48673
rect 4834 48549 5282 48617
rect 4834 48493 4844 48549
rect 4900 48493 4968 48549
rect 5024 48493 5092 48549
rect 5148 48493 5216 48549
rect 5272 48493 5282 48549
rect 4834 48425 5282 48493
rect 4834 48369 4844 48425
rect 4900 48369 4968 48425
rect 5024 48369 5092 48425
rect 5148 48369 5216 48425
rect 5272 48369 5282 48425
rect 4834 48301 5282 48369
rect 4834 48245 4844 48301
rect 4900 48245 4968 48301
rect 5024 48245 5092 48301
rect 5148 48245 5216 48301
rect 5272 48245 5282 48301
rect 4834 48177 5282 48245
rect 4834 48121 4844 48177
rect 4900 48121 4968 48177
rect 5024 48121 5092 48177
rect 5148 48121 5216 48177
rect 5272 48121 5282 48177
rect 4834 48053 5282 48121
rect 4834 47997 4844 48053
rect 4900 47997 4968 48053
rect 5024 47997 5092 48053
rect 5148 47997 5216 48053
rect 5272 47997 5282 48053
rect 4834 47929 5282 47997
rect 4834 47873 4844 47929
rect 4900 47873 4968 47929
rect 5024 47873 5092 47929
rect 5148 47873 5216 47929
rect 5272 47873 5282 47929
rect 4834 47805 5282 47873
rect 4834 47749 4844 47805
rect 4900 47749 4968 47805
rect 5024 47749 5092 47805
rect 5148 47749 5216 47805
rect 5272 47749 5282 47805
rect 4834 47739 5282 47749
rect 7127 49045 7451 49055
rect 7127 48989 7137 49045
rect 7193 48989 7261 49045
rect 7317 48989 7385 49045
rect 7441 48989 7451 49045
rect 7127 48921 7451 48989
rect 7127 48865 7137 48921
rect 7193 48865 7261 48921
rect 7317 48865 7385 48921
rect 7441 48865 7451 48921
rect 7127 48797 7451 48865
rect 7127 48741 7137 48797
rect 7193 48741 7261 48797
rect 7317 48741 7385 48797
rect 7441 48741 7451 48797
rect 7127 48673 7451 48741
rect 7127 48617 7137 48673
rect 7193 48617 7261 48673
rect 7317 48617 7385 48673
rect 7441 48617 7451 48673
rect 7127 48549 7451 48617
rect 7127 48493 7137 48549
rect 7193 48493 7261 48549
rect 7317 48493 7385 48549
rect 7441 48493 7451 48549
rect 7127 48425 7451 48493
rect 7127 48369 7137 48425
rect 7193 48369 7261 48425
rect 7317 48369 7385 48425
rect 7441 48369 7451 48425
rect 7127 48301 7451 48369
rect 7127 48245 7137 48301
rect 7193 48245 7261 48301
rect 7317 48245 7385 48301
rect 7441 48245 7451 48301
rect 7127 48177 7451 48245
rect 7127 48121 7137 48177
rect 7193 48121 7261 48177
rect 7317 48121 7385 48177
rect 7441 48121 7451 48177
rect 7127 48053 7451 48121
rect 7127 47997 7137 48053
rect 7193 47997 7261 48053
rect 7317 47997 7385 48053
rect 7441 47997 7451 48053
rect 7127 47929 7451 47997
rect 7127 47873 7137 47929
rect 7193 47873 7261 47929
rect 7317 47873 7385 47929
rect 7441 47873 7451 47929
rect 7127 47805 7451 47873
rect 7127 47749 7137 47805
rect 7193 47749 7261 47805
rect 7317 47749 7385 47805
rect 7441 47749 7451 47805
rect 7127 47739 7451 47749
rect 7613 49045 7937 49055
rect 7613 48989 7623 49045
rect 7679 48989 7747 49045
rect 7803 48989 7871 49045
rect 7927 48989 7937 49045
rect 7613 48921 7937 48989
rect 7613 48865 7623 48921
rect 7679 48865 7747 48921
rect 7803 48865 7871 48921
rect 7927 48865 7937 48921
rect 7613 48797 7937 48865
rect 7613 48741 7623 48797
rect 7679 48741 7747 48797
rect 7803 48741 7871 48797
rect 7927 48741 7937 48797
rect 7613 48673 7937 48741
rect 7613 48617 7623 48673
rect 7679 48617 7747 48673
rect 7803 48617 7871 48673
rect 7927 48617 7937 48673
rect 7613 48549 7937 48617
rect 7613 48493 7623 48549
rect 7679 48493 7747 48549
rect 7803 48493 7871 48549
rect 7927 48493 7937 48549
rect 7613 48425 7937 48493
rect 7613 48369 7623 48425
rect 7679 48369 7747 48425
rect 7803 48369 7871 48425
rect 7927 48369 7937 48425
rect 7613 48301 7937 48369
rect 7613 48245 7623 48301
rect 7679 48245 7747 48301
rect 7803 48245 7871 48301
rect 7927 48245 7937 48301
rect 7613 48177 7937 48245
rect 7613 48121 7623 48177
rect 7679 48121 7747 48177
rect 7803 48121 7871 48177
rect 7927 48121 7937 48177
rect 7613 48053 7937 48121
rect 7613 47997 7623 48053
rect 7679 47997 7747 48053
rect 7803 47997 7871 48053
rect 7927 47997 7937 48053
rect 7613 47929 7937 47997
rect 7613 47873 7623 47929
rect 7679 47873 7747 47929
rect 7803 47873 7871 47929
rect 7927 47873 7937 47929
rect 7613 47805 7937 47873
rect 7613 47749 7623 47805
rect 7679 47749 7747 47805
rect 7803 47749 7871 47805
rect 7927 47749 7937 47805
rect 7613 47739 7937 47749
rect 9782 49045 10230 49055
rect 9782 48989 9792 49045
rect 9848 48989 9916 49045
rect 9972 48989 10040 49045
rect 10096 48989 10164 49045
rect 10220 48989 10230 49045
rect 9782 48921 10230 48989
rect 9782 48865 9792 48921
rect 9848 48865 9916 48921
rect 9972 48865 10040 48921
rect 10096 48865 10164 48921
rect 10220 48865 10230 48921
rect 9782 48797 10230 48865
rect 9782 48741 9792 48797
rect 9848 48741 9916 48797
rect 9972 48741 10040 48797
rect 10096 48741 10164 48797
rect 10220 48741 10230 48797
rect 9782 48673 10230 48741
rect 9782 48617 9792 48673
rect 9848 48617 9916 48673
rect 9972 48617 10040 48673
rect 10096 48617 10164 48673
rect 10220 48617 10230 48673
rect 9782 48549 10230 48617
rect 9782 48493 9792 48549
rect 9848 48493 9916 48549
rect 9972 48493 10040 48549
rect 10096 48493 10164 48549
rect 10220 48493 10230 48549
rect 9782 48425 10230 48493
rect 9782 48369 9792 48425
rect 9848 48369 9916 48425
rect 9972 48369 10040 48425
rect 10096 48369 10164 48425
rect 10220 48369 10230 48425
rect 9782 48301 10230 48369
rect 9782 48245 9792 48301
rect 9848 48245 9916 48301
rect 9972 48245 10040 48301
rect 10096 48245 10164 48301
rect 10220 48245 10230 48301
rect 9782 48177 10230 48245
rect 9782 48121 9792 48177
rect 9848 48121 9916 48177
rect 9972 48121 10040 48177
rect 10096 48121 10164 48177
rect 10220 48121 10230 48177
rect 9782 48053 10230 48121
rect 9782 47997 9792 48053
rect 9848 47997 9916 48053
rect 9972 47997 10040 48053
rect 10096 47997 10164 48053
rect 10220 47997 10230 48053
rect 9782 47929 10230 47997
rect 9782 47873 9792 47929
rect 9848 47873 9916 47929
rect 9972 47873 10040 47929
rect 10096 47873 10164 47929
rect 10220 47873 10230 47929
rect 9782 47805 10230 47873
rect 9782 47749 9792 47805
rect 9848 47749 9916 47805
rect 9972 47749 10040 47805
rect 10096 47749 10164 47805
rect 10220 47749 10230 47805
rect 9782 47739 10230 47749
rect 12054 49045 12502 49055
rect 12054 48989 12064 49045
rect 12120 48989 12188 49045
rect 12244 48989 12312 49045
rect 12368 48989 12436 49045
rect 12492 48989 12502 49045
rect 12054 48921 12502 48989
rect 12054 48865 12064 48921
rect 12120 48865 12188 48921
rect 12244 48865 12312 48921
rect 12368 48865 12436 48921
rect 12492 48865 12502 48921
rect 12054 48797 12502 48865
rect 12054 48741 12064 48797
rect 12120 48741 12188 48797
rect 12244 48741 12312 48797
rect 12368 48741 12436 48797
rect 12492 48741 12502 48797
rect 12054 48673 12502 48741
rect 12054 48617 12064 48673
rect 12120 48617 12188 48673
rect 12244 48617 12312 48673
rect 12368 48617 12436 48673
rect 12492 48617 12502 48673
rect 12054 48549 12502 48617
rect 12054 48493 12064 48549
rect 12120 48493 12188 48549
rect 12244 48493 12312 48549
rect 12368 48493 12436 48549
rect 12492 48493 12502 48549
rect 12054 48425 12502 48493
rect 12054 48369 12064 48425
rect 12120 48369 12188 48425
rect 12244 48369 12312 48425
rect 12368 48369 12436 48425
rect 12492 48369 12502 48425
rect 12054 48301 12502 48369
rect 12054 48245 12064 48301
rect 12120 48245 12188 48301
rect 12244 48245 12312 48301
rect 12368 48245 12436 48301
rect 12492 48245 12502 48301
rect 12054 48177 12502 48245
rect 12054 48121 12064 48177
rect 12120 48121 12188 48177
rect 12244 48121 12312 48177
rect 12368 48121 12436 48177
rect 12492 48121 12502 48177
rect 12054 48053 12502 48121
rect 12054 47997 12064 48053
rect 12120 47997 12188 48053
rect 12244 47997 12312 48053
rect 12368 47997 12436 48053
rect 12492 47997 12502 48053
rect 12054 47929 12502 47997
rect 12054 47873 12064 47929
rect 12120 47873 12188 47929
rect 12244 47873 12312 47929
rect 12368 47873 12436 47929
rect 12492 47873 12502 47929
rect 12054 47805 12502 47873
rect 12054 47749 12064 47805
rect 12120 47749 12188 47805
rect 12244 47749 12312 47805
rect 12368 47749 12436 47805
rect 12492 47749 12502 47805
rect 12054 47739 12502 47749
rect 13468 49045 13668 49055
rect 13468 48989 13478 49045
rect 13534 48989 13602 49045
rect 13658 48989 13668 49045
rect 13468 48921 13668 48989
rect 13468 48865 13478 48921
rect 13534 48865 13602 48921
rect 13658 48865 13668 48921
rect 13468 48797 13668 48865
rect 13468 48741 13478 48797
rect 13534 48741 13602 48797
rect 13658 48741 13668 48797
rect 13468 48673 13668 48741
rect 13468 48617 13478 48673
rect 13534 48617 13602 48673
rect 13658 48617 13668 48673
rect 13468 48549 13668 48617
rect 13468 48493 13478 48549
rect 13534 48493 13602 48549
rect 13658 48493 13668 48549
rect 13468 48425 13668 48493
rect 13468 48369 13478 48425
rect 13534 48369 13602 48425
rect 13658 48369 13668 48425
rect 13468 48301 13668 48369
rect 13468 48245 13478 48301
rect 13534 48245 13602 48301
rect 13658 48245 13668 48301
rect 13468 48177 13668 48245
rect 13468 48121 13478 48177
rect 13534 48121 13602 48177
rect 13658 48121 13668 48177
rect 13468 48053 13668 48121
rect 13468 47997 13478 48053
rect 13534 47997 13602 48053
rect 13658 47997 13668 48053
rect 13468 47929 13668 47997
rect 13468 47873 13478 47929
rect 13534 47873 13602 47929
rect 13658 47873 13668 47929
rect 13468 47805 13668 47873
rect 13468 47749 13478 47805
rect 13534 47749 13602 47805
rect 13658 47749 13668 47805
rect 13468 47739 13668 47749
rect 14326 49045 14774 49055
rect 14326 48989 14336 49045
rect 14392 48989 14460 49045
rect 14516 48989 14584 49045
rect 14640 48989 14708 49045
rect 14764 48989 14774 49045
rect 14326 48921 14774 48989
rect 14326 48865 14336 48921
rect 14392 48865 14460 48921
rect 14516 48865 14584 48921
rect 14640 48865 14708 48921
rect 14764 48865 14774 48921
rect 14326 48797 14774 48865
rect 14326 48741 14336 48797
rect 14392 48741 14460 48797
rect 14516 48741 14584 48797
rect 14640 48741 14708 48797
rect 14764 48741 14774 48797
rect 14326 48673 14774 48741
rect 14326 48617 14336 48673
rect 14392 48617 14460 48673
rect 14516 48617 14584 48673
rect 14640 48617 14708 48673
rect 14764 48617 14774 48673
rect 14326 48549 14774 48617
rect 14326 48493 14336 48549
rect 14392 48493 14460 48549
rect 14516 48493 14584 48549
rect 14640 48493 14708 48549
rect 14764 48493 14774 48549
rect 14326 48425 14774 48493
rect 14326 48369 14336 48425
rect 14392 48369 14460 48425
rect 14516 48369 14584 48425
rect 14640 48369 14708 48425
rect 14764 48369 14774 48425
rect 14326 48301 14774 48369
rect 14326 48245 14336 48301
rect 14392 48245 14460 48301
rect 14516 48245 14584 48301
rect 14640 48245 14708 48301
rect 14764 48245 14774 48301
rect 14326 48177 14774 48245
rect 14326 48121 14336 48177
rect 14392 48121 14460 48177
rect 14516 48121 14584 48177
rect 14640 48121 14708 48177
rect 14764 48121 14774 48177
rect 14326 48053 14774 48121
rect 14326 47997 14336 48053
rect 14392 47997 14460 48053
rect 14516 47997 14584 48053
rect 14640 47997 14708 48053
rect 14764 47997 14774 48053
rect 14326 47929 14774 47997
rect 14326 47873 14336 47929
rect 14392 47873 14460 47929
rect 14516 47873 14584 47929
rect 14640 47873 14708 47929
rect 14764 47873 14774 47929
rect 14326 47805 14774 47873
rect 14326 47749 14336 47805
rect 14392 47749 14460 47805
rect 14516 47749 14584 47805
rect 14640 47749 14708 47805
rect 14764 47749 14774 47805
rect 14326 47739 14774 47749
rect 1136 47445 1336 47455
rect 1136 47389 1146 47445
rect 1202 47389 1270 47445
rect 1326 47389 1336 47445
rect 1136 47321 1336 47389
rect 1136 47265 1146 47321
rect 1202 47265 1270 47321
rect 1326 47265 1336 47321
rect 1136 47197 1336 47265
rect 1136 47141 1146 47197
rect 1202 47141 1270 47197
rect 1326 47141 1336 47197
rect 1136 47073 1336 47141
rect 1136 47017 1146 47073
rect 1202 47017 1270 47073
rect 1326 47017 1336 47073
rect 1136 46949 1336 47017
rect 1136 46893 1146 46949
rect 1202 46893 1270 46949
rect 1326 46893 1336 46949
rect 1136 46825 1336 46893
rect 1136 46769 1146 46825
rect 1202 46769 1270 46825
rect 1326 46769 1336 46825
rect 1136 46701 1336 46769
rect 1136 46645 1146 46701
rect 1202 46645 1270 46701
rect 1326 46645 1336 46701
rect 1136 46577 1336 46645
rect 1136 46521 1146 46577
rect 1202 46521 1270 46577
rect 1326 46521 1336 46577
rect 1136 46453 1336 46521
rect 1136 46397 1146 46453
rect 1202 46397 1270 46453
rect 1326 46397 1336 46453
rect 1136 46329 1336 46397
rect 1136 46273 1146 46329
rect 1202 46273 1270 46329
rect 1326 46273 1336 46329
rect 1136 46205 1336 46273
rect 1136 46149 1146 46205
rect 1202 46149 1270 46205
rect 1326 46149 1336 46205
rect 1136 46139 1336 46149
rect 1994 47445 2442 47455
rect 1994 47389 2004 47445
rect 2060 47389 2128 47445
rect 2184 47389 2252 47445
rect 2308 47389 2376 47445
rect 2432 47389 2442 47445
rect 1994 47321 2442 47389
rect 1994 47265 2004 47321
rect 2060 47265 2128 47321
rect 2184 47265 2252 47321
rect 2308 47265 2376 47321
rect 2432 47265 2442 47321
rect 1994 47197 2442 47265
rect 1994 47141 2004 47197
rect 2060 47141 2128 47197
rect 2184 47141 2252 47197
rect 2308 47141 2376 47197
rect 2432 47141 2442 47197
rect 1994 47073 2442 47141
rect 1994 47017 2004 47073
rect 2060 47017 2128 47073
rect 2184 47017 2252 47073
rect 2308 47017 2376 47073
rect 2432 47017 2442 47073
rect 1994 46949 2442 47017
rect 1994 46893 2004 46949
rect 2060 46893 2128 46949
rect 2184 46893 2252 46949
rect 2308 46893 2376 46949
rect 2432 46893 2442 46949
rect 1994 46825 2442 46893
rect 1994 46769 2004 46825
rect 2060 46769 2128 46825
rect 2184 46769 2252 46825
rect 2308 46769 2376 46825
rect 2432 46769 2442 46825
rect 1994 46701 2442 46769
rect 1994 46645 2004 46701
rect 2060 46645 2128 46701
rect 2184 46645 2252 46701
rect 2308 46645 2376 46701
rect 2432 46645 2442 46701
rect 1994 46577 2442 46645
rect 1994 46521 2004 46577
rect 2060 46521 2128 46577
rect 2184 46521 2252 46577
rect 2308 46521 2376 46577
rect 2432 46521 2442 46577
rect 1994 46453 2442 46521
rect 1994 46397 2004 46453
rect 2060 46397 2128 46453
rect 2184 46397 2252 46453
rect 2308 46397 2376 46453
rect 2432 46397 2442 46453
rect 1994 46329 2442 46397
rect 1994 46273 2004 46329
rect 2060 46273 2128 46329
rect 2184 46273 2252 46329
rect 2308 46273 2376 46329
rect 2432 46273 2442 46329
rect 1994 46205 2442 46273
rect 1994 46149 2004 46205
rect 2060 46149 2128 46205
rect 2184 46149 2252 46205
rect 2308 46149 2376 46205
rect 2432 46149 2442 46205
rect 1994 46139 2442 46149
rect 3698 47445 4146 47455
rect 3698 47389 3708 47445
rect 3764 47389 3832 47445
rect 3888 47389 3956 47445
rect 4012 47389 4080 47445
rect 4136 47389 4146 47445
rect 3698 47321 4146 47389
rect 3698 47265 3708 47321
rect 3764 47265 3832 47321
rect 3888 47265 3956 47321
rect 4012 47265 4080 47321
rect 4136 47265 4146 47321
rect 3698 47197 4146 47265
rect 3698 47141 3708 47197
rect 3764 47141 3832 47197
rect 3888 47141 3956 47197
rect 4012 47141 4080 47197
rect 4136 47141 4146 47197
rect 3698 47073 4146 47141
rect 3698 47017 3708 47073
rect 3764 47017 3832 47073
rect 3888 47017 3956 47073
rect 4012 47017 4080 47073
rect 4136 47017 4146 47073
rect 3698 46949 4146 47017
rect 3698 46893 3708 46949
rect 3764 46893 3832 46949
rect 3888 46893 3956 46949
rect 4012 46893 4080 46949
rect 4136 46893 4146 46949
rect 3698 46825 4146 46893
rect 3698 46769 3708 46825
rect 3764 46769 3832 46825
rect 3888 46769 3956 46825
rect 4012 46769 4080 46825
rect 4136 46769 4146 46825
rect 3698 46701 4146 46769
rect 3698 46645 3708 46701
rect 3764 46645 3832 46701
rect 3888 46645 3956 46701
rect 4012 46645 4080 46701
rect 4136 46645 4146 46701
rect 3698 46577 4146 46645
rect 3698 46521 3708 46577
rect 3764 46521 3832 46577
rect 3888 46521 3956 46577
rect 4012 46521 4080 46577
rect 4136 46521 4146 46577
rect 3698 46453 4146 46521
rect 3698 46397 3708 46453
rect 3764 46397 3832 46453
rect 3888 46397 3956 46453
rect 4012 46397 4080 46453
rect 4136 46397 4146 46453
rect 3698 46329 4146 46397
rect 3698 46273 3708 46329
rect 3764 46273 3832 46329
rect 3888 46273 3956 46329
rect 4012 46273 4080 46329
rect 4136 46273 4146 46329
rect 3698 46205 4146 46273
rect 3698 46149 3708 46205
rect 3764 46149 3832 46205
rect 3888 46149 3956 46205
rect 4012 46149 4080 46205
rect 4136 46149 4146 46205
rect 3698 46139 4146 46149
rect 5970 47445 6418 47455
rect 5970 47389 5980 47445
rect 6036 47389 6104 47445
rect 6160 47389 6228 47445
rect 6284 47389 6352 47445
rect 6408 47389 6418 47445
rect 5970 47321 6418 47389
rect 5970 47265 5980 47321
rect 6036 47265 6104 47321
rect 6160 47265 6228 47321
rect 6284 47265 6352 47321
rect 6408 47265 6418 47321
rect 5970 47197 6418 47265
rect 5970 47141 5980 47197
rect 6036 47141 6104 47197
rect 6160 47141 6228 47197
rect 6284 47141 6352 47197
rect 6408 47141 6418 47197
rect 5970 47073 6418 47141
rect 5970 47017 5980 47073
rect 6036 47017 6104 47073
rect 6160 47017 6228 47073
rect 6284 47017 6352 47073
rect 6408 47017 6418 47073
rect 5970 46949 6418 47017
rect 5970 46893 5980 46949
rect 6036 46893 6104 46949
rect 6160 46893 6228 46949
rect 6284 46893 6352 46949
rect 6408 46893 6418 46949
rect 5970 46825 6418 46893
rect 5970 46769 5980 46825
rect 6036 46769 6104 46825
rect 6160 46769 6228 46825
rect 6284 46769 6352 46825
rect 6408 46769 6418 46825
rect 5970 46701 6418 46769
rect 5970 46645 5980 46701
rect 6036 46645 6104 46701
rect 6160 46645 6228 46701
rect 6284 46645 6352 46701
rect 6408 46645 6418 46701
rect 5970 46577 6418 46645
rect 5970 46521 5980 46577
rect 6036 46521 6104 46577
rect 6160 46521 6228 46577
rect 6284 46521 6352 46577
rect 6408 46521 6418 46577
rect 5970 46453 6418 46521
rect 5970 46397 5980 46453
rect 6036 46397 6104 46453
rect 6160 46397 6228 46453
rect 6284 46397 6352 46453
rect 6408 46397 6418 46453
rect 5970 46329 6418 46397
rect 5970 46273 5980 46329
rect 6036 46273 6104 46329
rect 6160 46273 6228 46329
rect 6284 46273 6352 46329
rect 6408 46273 6418 46329
rect 5970 46205 6418 46273
rect 5970 46149 5980 46205
rect 6036 46149 6104 46205
rect 6160 46149 6228 46205
rect 6284 46149 6352 46205
rect 6408 46149 6418 46205
rect 5970 46139 6418 46149
rect 8646 47445 9094 47455
rect 8646 47389 8656 47445
rect 8712 47389 8780 47445
rect 8836 47389 8904 47445
rect 8960 47389 9028 47445
rect 9084 47389 9094 47445
rect 8646 47321 9094 47389
rect 8646 47265 8656 47321
rect 8712 47265 8780 47321
rect 8836 47265 8904 47321
rect 8960 47265 9028 47321
rect 9084 47265 9094 47321
rect 8646 47197 9094 47265
rect 8646 47141 8656 47197
rect 8712 47141 8780 47197
rect 8836 47141 8904 47197
rect 8960 47141 9028 47197
rect 9084 47141 9094 47197
rect 8646 47073 9094 47141
rect 8646 47017 8656 47073
rect 8712 47017 8780 47073
rect 8836 47017 8904 47073
rect 8960 47017 9028 47073
rect 9084 47017 9094 47073
rect 8646 46949 9094 47017
rect 8646 46893 8656 46949
rect 8712 46893 8780 46949
rect 8836 46893 8904 46949
rect 8960 46893 9028 46949
rect 9084 46893 9094 46949
rect 8646 46825 9094 46893
rect 8646 46769 8656 46825
rect 8712 46769 8780 46825
rect 8836 46769 8904 46825
rect 8960 46769 9028 46825
rect 9084 46769 9094 46825
rect 8646 46701 9094 46769
rect 8646 46645 8656 46701
rect 8712 46645 8780 46701
rect 8836 46645 8904 46701
rect 8960 46645 9028 46701
rect 9084 46645 9094 46701
rect 8646 46577 9094 46645
rect 8646 46521 8656 46577
rect 8712 46521 8780 46577
rect 8836 46521 8904 46577
rect 8960 46521 9028 46577
rect 9084 46521 9094 46577
rect 8646 46453 9094 46521
rect 8646 46397 8656 46453
rect 8712 46397 8780 46453
rect 8836 46397 8904 46453
rect 8960 46397 9028 46453
rect 9084 46397 9094 46453
rect 8646 46329 9094 46397
rect 8646 46273 8656 46329
rect 8712 46273 8780 46329
rect 8836 46273 8904 46329
rect 8960 46273 9028 46329
rect 9084 46273 9094 46329
rect 8646 46205 9094 46273
rect 8646 46149 8656 46205
rect 8712 46149 8780 46205
rect 8836 46149 8904 46205
rect 8960 46149 9028 46205
rect 9084 46149 9094 46205
rect 8646 46139 9094 46149
rect 10918 47445 11366 47455
rect 10918 47389 10928 47445
rect 10984 47389 11052 47445
rect 11108 47389 11176 47445
rect 11232 47389 11300 47445
rect 11356 47389 11366 47445
rect 10918 47321 11366 47389
rect 10918 47265 10928 47321
rect 10984 47265 11052 47321
rect 11108 47265 11176 47321
rect 11232 47265 11300 47321
rect 11356 47265 11366 47321
rect 10918 47197 11366 47265
rect 10918 47141 10928 47197
rect 10984 47141 11052 47197
rect 11108 47141 11176 47197
rect 11232 47141 11300 47197
rect 11356 47141 11366 47197
rect 10918 47073 11366 47141
rect 10918 47017 10928 47073
rect 10984 47017 11052 47073
rect 11108 47017 11176 47073
rect 11232 47017 11300 47073
rect 11356 47017 11366 47073
rect 10918 46949 11366 47017
rect 10918 46893 10928 46949
rect 10984 46893 11052 46949
rect 11108 46893 11176 46949
rect 11232 46893 11300 46949
rect 11356 46893 11366 46949
rect 10918 46825 11366 46893
rect 10918 46769 10928 46825
rect 10984 46769 11052 46825
rect 11108 46769 11176 46825
rect 11232 46769 11300 46825
rect 11356 46769 11366 46825
rect 10918 46701 11366 46769
rect 10918 46645 10928 46701
rect 10984 46645 11052 46701
rect 11108 46645 11176 46701
rect 11232 46645 11300 46701
rect 11356 46645 11366 46701
rect 10918 46577 11366 46645
rect 10918 46521 10928 46577
rect 10984 46521 11052 46577
rect 11108 46521 11176 46577
rect 11232 46521 11300 46577
rect 11356 46521 11366 46577
rect 10918 46453 11366 46521
rect 10918 46397 10928 46453
rect 10984 46397 11052 46453
rect 11108 46397 11176 46453
rect 11232 46397 11300 46453
rect 11356 46397 11366 46453
rect 10918 46329 11366 46397
rect 10918 46273 10928 46329
rect 10984 46273 11052 46329
rect 11108 46273 11176 46329
rect 11232 46273 11300 46329
rect 11356 46273 11366 46329
rect 10918 46205 11366 46273
rect 10918 46149 10928 46205
rect 10984 46149 11052 46205
rect 11108 46149 11176 46205
rect 11232 46149 11300 46205
rect 11356 46149 11366 46205
rect 10918 46139 11366 46149
rect 12622 47445 13070 47455
rect 12622 47389 12632 47445
rect 12688 47389 12756 47445
rect 12812 47389 12880 47445
rect 12936 47389 13004 47445
rect 13060 47389 13070 47445
rect 12622 47321 13070 47389
rect 12622 47265 12632 47321
rect 12688 47265 12756 47321
rect 12812 47265 12880 47321
rect 12936 47265 13004 47321
rect 13060 47265 13070 47321
rect 12622 47197 13070 47265
rect 12622 47141 12632 47197
rect 12688 47141 12756 47197
rect 12812 47141 12880 47197
rect 12936 47141 13004 47197
rect 13060 47141 13070 47197
rect 12622 47073 13070 47141
rect 12622 47017 12632 47073
rect 12688 47017 12756 47073
rect 12812 47017 12880 47073
rect 12936 47017 13004 47073
rect 13060 47017 13070 47073
rect 12622 46949 13070 47017
rect 12622 46893 12632 46949
rect 12688 46893 12756 46949
rect 12812 46893 12880 46949
rect 12936 46893 13004 46949
rect 13060 46893 13070 46949
rect 12622 46825 13070 46893
rect 12622 46769 12632 46825
rect 12688 46769 12756 46825
rect 12812 46769 12880 46825
rect 12936 46769 13004 46825
rect 13060 46769 13070 46825
rect 12622 46701 13070 46769
rect 12622 46645 12632 46701
rect 12688 46645 12756 46701
rect 12812 46645 12880 46701
rect 12936 46645 13004 46701
rect 13060 46645 13070 46701
rect 12622 46577 13070 46645
rect 12622 46521 12632 46577
rect 12688 46521 12756 46577
rect 12812 46521 12880 46577
rect 12936 46521 13004 46577
rect 13060 46521 13070 46577
rect 12622 46453 13070 46521
rect 12622 46397 12632 46453
rect 12688 46397 12756 46453
rect 12812 46397 12880 46453
rect 12936 46397 13004 46453
rect 13060 46397 13070 46453
rect 12622 46329 13070 46397
rect 12622 46273 12632 46329
rect 12688 46273 12756 46329
rect 12812 46273 12880 46329
rect 12936 46273 13004 46329
rect 13060 46273 13070 46329
rect 12622 46205 13070 46273
rect 12622 46149 12632 46205
rect 12688 46149 12756 46205
rect 12812 46149 12880 46205
rect 12936 46149 13004 46205
rect 13060 46149 13070 46205
rect 12622 46139 13070 46149
rect 13758 47445 14206 47455
rect 13758 47389 13768 47445
rect 13824 47389 13892 47445
rect 13948 47389 14016 47445
rect 14072 47389 14140 47445
rect 14196 47389 14206 47445
rect 13758 47321 14206 47389
rect 13758 47265 13768 47321
rect 13824 47265 13892 47321
rect 13948 47265 14016 47321
rect 14072 47265 14140 47321
rect 14196 47265 14206 47321
rect 13758 47197 14206 47265
rect 13758 47141 13768 47197
rect 13824 47141 13892 47197
rect 13948 47141 14016 47197
rect 14072 47141 14140 47197
rect 14196 47141 14206 47197
rect 13758 47073 14206 47141
rect 13758 47017 13768 47073
rect 13824 47017 13892 47073
rect 13948 47017 14016 47073
rect 14072 47017 14140 47073
rect 14196 47017 14206 47073
rect 13758 46949 14206 47017
rect 13758 46893 13768 46949
rect 13824 46893 13892 46949
rect 13948 46893 14016 46949
rect 14072 46893 14140 46949
rect 14196 46893 14206 46949
rect 13758 46825 14206 46893
rect 13758 46769 13768 46825
rect 13824 46769 13892 46825
rect 13948 46769 14016 46825
rect 14072 46769 14140 46825
rect 14196 46769 14206 46825
rect 13758 46701 14206 46769
rect 13758 46645 13768 46701
rect 13824 46645 13892 46701
rect 13948 46645 14016 46701
rect 14072 46645 14140 46701
rect 14196 46645 14206 46701
rect 13758 46577 14206 46645
rect 13758 46521 13768 46577
rect 13824 46521 13892 46577
rect 13948 46521 14016 46577
rect 14072 46521 14140 46577
rect 14196 46521 14206 46577
rect 13758 46453 14206 46521
rect 13758 46397 13768 46453
rect 13824 46397 13892 46453
rect 13948 46397 14016 46453
rect 14072 46397 14140 46453
rect 14196 46397 14206 46453
rect 13758 46329 14206 46397
rect 13758 46273 13768 46329
rect 13824 46273 13892 46329
rect 13948 46273 14016 46329
rect 14072 46273 14140 46329
rect 14196 46273 14206 46329
rect 13758 46205 14206 46273
rect 13758 46149 13768 46205
rect 13824 46149 13892 46205
rect 13948 46149 14016 46205
rect 14072 46149 14140 46205
rect 14196 46149 14206 46205
rect 13758 46139 14206 46149
rect 290 45845 738 45855
rect 290 45789 300 45845
rect 356 45789 424 45845
rect 480 45789 548 45845
rect 604 45789 672 45845
rect 728 45789 738 45845
rect 290 45721 738 45789
rect 290 45665 300 45721
rect 356 45665 424 45721
rect 480 45665 548 45721
rect 604 45665 672 45721
rect 728 45665 738 45721
rect 290 45597 738 45665
rect 290 45541 300 45597
rect 356 45541 424 45597
rect 480 45541 548 45597
rect 604 45541 672 45597
rect 728 45541 738 45597
rect 290 45473 738 45541
rect 290 45417 300 45473
rect 356 45417 424 45473
rect 480 45417 548 45473
rect 604 45417 672 45473
rect 728 45417 738 45473
rect 290 45349 738 45417
rect 290 45293 300 45349
rect 356 45293 424 45349
rect 480 45293 548 45349
rect 604 45293 672 45349
rect 728 45293 738 45349
rect 290 45225 738 45293
rect 290 45169 300 45225
rect 356 45169 424 45225
rect 480 45169 548 45225
rect 604 45169 672 45225
rect 728 45169 738 45225
rect 290 45101 738 45169
rect 290 45045 300 45101
rect 356 45045 424 45101
rect 480 45045 548 45101
rect 604 45045 672 45101
rect 728 45045 738 45101
rect 290 44977 738 45045
rect 290 44921 300 44977
rect 356 44921 424 44977
rect 480 44921 548 44977
rect 604 44921 672 44977
rect 728 44921 738 44977
rect 290 44853 738 44921
rect 290 44797 300 44853
rect 356 44797 424 44853
rect 480 44797 548 44853
rect 604 44797 672 44853
rect 728 44797 738 44853
rect 290 44729 738 44797
rect 290 44673 300 44729
rect 356 44673 424 44729
rect 480 44673 548 44729
rect 604 44673 672 44729
rect 728 44673 738 44729
rect 290 44605 738 44673
rect 290 44549 300 44605
rect 356 44549 424 44605
rect 480 44549 548 44605
rect 604 44549 672 44605
rect 728 44549 738 44605
rect 290 44539 738 44549
rect 1426 45845 1874 45855
rect 1426 45789 1436 45845
rect 1492 45789 1560 45845
rect 1616 45789 1684 45845
rect 1740 45789 1808 45845
rect 1864 45789 1874 45845
rect 1426 45721 1874 45789
rect 1426 45665 1436 45721
rect 1492 45665 1560 45721
rect 1616 45665 1684 45721
rect 1740 45665 1808 45721
rect 1864 45665 1874 45721
rect 1426 45597 1874 45665
rect 1426 45541 1436 45597
rect 1492 45541 1560 45597
rect 1616 45541 1684 45597
rect 1740 45541 1808 45597
rect 1864 45541 1874 45597
rect 1426 45473 1874 45541
rect 1426 45417 1436 45473
rect 1492 45417 1560 45473
rect 1616 45417 1684 45473
rect 1740 45417 1808 45473
rect 1864 45417 1874 45473
rect 1426 45349 1874 45417
rect 1426 45293 1436 45349
rect 1492 45293 1560 45349
rect 1616 45293 1684 45349
rect 1740 45293 1808 45349
rect 1864 45293 1874 45349
rect 1426 45225 1874 45293
rect 1426 45169 1436 45225
rect 1492 45169 1560 45225
rect 1616 45169 1684 45225
rect 1740 45169 1808 45225
rect 1864 45169 1874 45225
rect 1426 45101 1874 45169
rect 1426 45045 1436 45101
rect 1492 45045 1560 45101
rect 1616 45045 1684 45101
rect 1740 45045 1808 45101
rect 1864 45045 1874 45101
rect 1426 44977 1874 45045
rect 1426 44921 1436 44977
rect 1492 44921 1560 44977
rect 1616 44921 1684 44977
rect 1740 44921 1808 44977
rect 1864 44921 1874 44977
rect 1426 44853 1874 44921
rect 1426 44797 1436 44853
rect 1492 44797 1560 44853
rect 1616 44797 1684 44853
rect 1740 44797 1808 44853
rect 1864 44797 1874 44853
rect 1426 44729 1874 44797
rect 1426 44673 1436 44729
rect 1492 44673 1560 44729
rect 1616 44673 1684 44729
rect 1740 44673 1808 44729
rect 1864 44673 1874 44729
rect 1426 44605 1874 44673
rect 1426 44549 1436 44605
rect 1492 44549 1560 44605
rect 1616 44549 1684 44605
rect 1740 44549 1808 44605
rect 1864 44549 1874 44605
rect 1426 44539 1874 44549
rect 2562 45845 3010 45855
rect 2562 45789 2572 45845
rect 2628 45789 2696 45845
rect 2752 45789 2820 45845
rect 2876 45789 2944 45845
rect 3000 45789 3010 45845
rect 2562 45721 3010 45789
rect 2562 45665 2572 45721
rect 2628 45665 2696 45721
rect 2752 45665 2820 45721
rect 2876 45665 2944 45721
rect 3000 45665 3010 45721
rect 2562 45597 3010 45665
rect 2562 45541 2572 45597
rect 2628 45541 2696 45597
rect 2752 45541 2820 45597
rect 2876 45541 2944 45597
rect 3000 45541 3010 45597
rect 2562 45473 3010 45541
rect 2562 45417 2572 45473
rect 2628 45417 2696 45473
rect 2752 45417 2820 45473
rect 2876 45417 2944 45473
rect 3000 45417 3010 45473
rect 2562 45349 3010 45417
rect 2562 45293 2572 45349
rect 2628 45293 2696 45349
rect 2752 45293 2820 45349
rect 2876 45293 2944 45349
rect 3000 45293 3010 45349
rect 2562 45225 3010 45293
rect 2562 45169 2572 45225
rect 2628 45169 2696 45225
rect 2752 45169 2820 45225
rect 2876 45169 2944 45225
rect 3000 45169 3010 45225
rect 2562 45101 3010 45169
rect 2562 45045 2572 45101
rect 2628 45045 2696 45101
rect 2752 45045 2820 45101
rect 2876 45045 2944 45101
rect 3000 45045 3010 45101
rect 2562 44977 3010 45045
rect 2562 44921 2572 44977
rect 2628 44921 2696 44977
rect 2752 44921 2820 44977
rect 2876 44921 2944 44977
rect 3000 44921 3010 44977
rect 2562 44853 3010 44921
rect 2562 44797 2572 44853
rect 2628 44797 2696 44853
rect 2752 44797 2820 44853
rect 2876 44797 2944 44853
rect 3000 44797 3010 44853
rect 2562 44729 3010 44797
rect 2562 44673 2572 44729
rect 2628 44673 2696 44729
rect 2752 44673 2820 44729
rect 2876 44673 2944 44729
rect 3000 44673 3010 44729
rect 2562 44605 3010 44673
rect 2562 44549 2572 44605
rect 2628 44549 2696 44605
rect 2752 44549 2820 44605
rect 2876 44549 2944 44605
rect 3000 44549 3010 44605
rect 2562 44539 3010 44549
rect 4834 45845 5282 45855
rect 4834 45789 4844 45845
rect 4900 45789 4968 45845
rect 5024 45789 5092 45845
rect 5148 45789 5216 45845
rect 5272 45789 5282 45845
rect 4834 45721 5282 45789
rect 4834 45665 4844 45721
rect 4900 45665 4968 45721
rect 5024 45665 5092 45721
rect 5148 45665 5216 45721
rect 5272 45665 5282 45721
rect 4834 45597 5282 45665
rect 4834 45541 4844 45597
rect 4900 45541 4968 45597
rect 5024 45541 5092 45597
rect 5148 45541 5216 45597
rect 5272 45541 5282 45597
rect 4834 45473 5282 45541
rect 4834 45417 4844 45473
rect 4900 45417 4968 45473
rect 5024 45417 5092 45473
rect 5148 45417 5216 45473
rect 5272 45417 5282 45473
rect 4834 45349 5282 45417
rect 4834 45293 4844 45349
rect 4900 45293 4968 45349
rect 5024 45293 5092 45349
rect 5148 45293 5216 45349
rect 5272 45293 5282 45349
rect 4834 45225 5282 45293
rect 4834 45169 4844 45225
rect 4900 45169 4968 45225
rect 5024 45169 5092 45225
rect 5148 45169 5216 45225
rect 5272 45169 5282 45225
rect 4834 45101 5282 45169
rect 4834 45045 4844 45101
rect 4900 45045 4968 45101
rect 5024 45045 5092 45101
rect 5148 45045 5216 45101
rect 5272 45045 5282 45101
rect 4834 44977 5282 45045
rect 4834 44921 4844 44977
rect 4900 44921 4968 44977
rect 5024 44921 5092 44977
rect 5148 44921 5216 44977
rect 5272 44921 5282 44977
rect 4834 44853 5282 44921
rect 4834 44797 4844 44853
rect 4900 44797 4968 44853
rect 5024 44797 5092 44853
rect 5148 44797 5216 44853
rect 5272 44797 5282 44853
rect 4834 44729 5282 44797
rect 4834 44673 4844 44729
rect 4900 44673 4968 44729
rect 5024 44673 5092 44729
rect 5148 44673 5216 44729
rect 5272 44673 5282 44729
rect 4834 44605 5282 44673
rect 4834 44549 4844 44605
rect 4900 44549 4968 44605
rect 5024 44549 5092 44605
rect 5148 44549 5216 44605
rect 5272 44549 5282 44605
rect 4834 44539 5282 44549
rect 7127 45845 7451 45855
rect 7127 45789 7137 45845
rect 7193 45789 7261 45845
rect 7317 45789 7385 45845
rect 7441 45789 7451 45845
rect 7127 45721 7451 45789
rect 7127 45665 7137 45721
rect 7193 45665 7261 45721
rect 7317 45665 7385 45721
rect 7441 45665 7451 45721
rect 7127 45597 7451 45665
rect 7127 45541 7137 45597
rect 7193 45541 7261 45597
rect 7317 45541 7385 45597
rect 7441 45541 7451 45597
rect 7127 45473 7451 45541
rect 7127 45417 7137 45473
rect 7193 45417 7261 45473
rect 7317 45417 7385 45473
rect 7441 45417 7451 45473
rect 7127 45349 7451 45417
rect 7127 45293 7137 45349
rect 7193 45293 7261 45349
rect 7317 45293 7385 45349
rect 7441 45293 7451 45349
rect 7127 45225 7451 45293
rect 7127 45169 7137 45225
rect 7193 45169 7261 45225
rect 7317 45169 7385 45225
rect 7441 45169 7451 45225
rect 7127 45101 7451 45169
rect 7127 45045 7137 45101
rect 7193 45045 7261 45101
rect 7317 45045 7385 45101
rect 7441 45045 7451 45101
rect 7127 44977 7451 45045
rect 7127 44921 7137 44977
rect 7193 44921 7261 44977
rect 7317 44921 7385 44977
rect 7441 44921 7451 44977
rect 7127 44853 7451 44921
rect 7127 44797 7137 44853
rect 7193 44797 7261 44853
rect 7317 44797 7385 44853
rect 7441 44797 7451 44853
rect 7127 44729 7451 44797
rect 7127 44673 7137 44729
rect 7193 44673 7261 44729
rect 7317 44673 7385 44729
rect 7441 44673 7451 44729
rect 7127 44605 7451 44673
rect 7127 44549 7137 44605
rect 7193 44549 7261 44605
rect 7317 44549 7385 44605
rect 7441 44549 7451 44605
rect 7127 44539 7451 44549
rect 7613 45845 7937 45855
rect 7613 45789 7623 45845
rect 7679 45789 7747 45845
rect 7803 45789 7871 45845
rect 7927 45789 7937 45845
rect 7613 45721 7937 45789
rect 7613 45665 7623 45721
rect 7679 45665 7747 45721
rect 7803 45665 7871 45721
rect 7927 45665 7937 45721
rect 7613 45597 7937 45665
rect 7613 45541 7623 45597
rect 7679 45541 7747 45597
rect 7803 45541 7871 45597
rect 7927 45541 7937 45597
rect 7613 45473 7937 45541
rect 7613 45417 7623 45473
rect 7679 45417 7747 45473
rect 7803 45417 7871 45473
rect 7927 45417 7937 45473
rect 7613 45349 7937 45417
rect 7613 45293 7623 45349
rect 7679 45293 7747 45349
rect 7803 45293 7871 45349
rect 7927 45293 7937 45349
rect 7613 45225 7937 45293
rect 7613 45169 7623 45225
rect 7679 45169 7747 45225
rect 7803 45169 7871 45225
rect 7927 45169 7937 45225
rect 7613 45101 7937 45169
rect 7613 45045 7623 45101
rect 7679 45045 7747 45101
rect 7803 45045 7871 45101
rect 7927 45045 7937 45101
rect 7613 44977 7937 45045
rect 7613 44921 7623 44977
rect 7679 44921 7747 44977
rect 7803 44921 7871 44977
rect 7927 44921 7937 44977
rect 7613 44853 7937 44921
rect 7613 44797 7623 44853
rect 7679 44797 7747 44853
rect 7803 44797 7871 44853
rect 7927 44797 7937 44853
rect 7613 44729 7937 44797
rect 7613 44673 7623 44729
rect 7679 44673 7747 44729
rect 7803 44673 7871 44729
rect 7927 44673 7937 44729
rect 7613 44605 7937 44673
rect 7613 44549 7623 44605
rect 7679 44549 7747 44605
rect 7803 44549 7871 44605
rect 7927 44549 7937 44605
rect 7613 44539 7937 44549
rect 9782 45845 10230 45855
rect 9782 45789 9792 45845
rect 9848 45789 9916 45845
rect 9972 45789 10040 45845
rect 10096 45789 10164 45845
rect 10220 45789 10230 45845
rect 9782 45721 10230 45789
rect 9782 45665 9792 45721
rect 9848 45665 9916 45721
rect 9972 45665 10040 45721
rect 10096 45665 10164 45721
rect 10220 45665 10230 45721
rect 9782 45597 10230 45665
rect 9782 45541 9792 45597
rect 9848 45541 9916 45597
rect 9972 45541 10040 45597
rect 10096 45541 10164 45597
rect 10220 45541 10230 45597
rect 9782 45473 10230 45541
rect 9782 45417 9792 45473
rect 9848 45417 9916 45473
rect 9972 45417 10040 45473
rect 10096 45417 10164 45473
rect 10220 45417 10230 45473
rect 9782 45349 10230 45417
rect 9782 45293 9792 45349
rect 9848 45293 9916 45349
rect 9972 45293 10040 45349
rect 10096 45293 10164 45349
rect 10220 45293 10230 45349
rect 9782 45225 10230 45293
rect 9782 45169 9792 45225
rect 9848 45169 9916 45225
rect 9972 45169 10040 45225
rect 10096 45169 10164 45225
rect 10220 45169 10230 45225
rect 9782 45101 10230 45169
rect 9782 45045 9792 45101
rect 9848 45045 9916 45101
rect 9972 45045 10040 45101
rect 10096 45045 10164 45101
rect 10220 45045 10230 45101
rect 9782 44977 10230 45045
rect 9782 44921 9792 44977
rect 9848 44921 9916 44977
rect 9972 44921 10040 44977
rect 10096 44921 10164 44977
rect 10220 44921 10230 44977
rect 9782 44853 10230 44921
rect 9782 44797 9792 44853
rect 9848 44797 9916 44853
rect 9972 44797 10040 44853
rect 10096 44797 10164 44853
rect 10220 44797 10230 44853
rect 9782 44729 10230 44797
rect 9782 44673 9792 44729
rect 9848 44673 9916 44729
rect 9972 44673 10040 44729
rect 10096 44673 10164 44729
rect 10220 44673 10230 44729
rect 9782 44605 10230 44673
rect 9782 44549 9792 44605
rect 9848 44549 9916 44605
rect 9972 44549 10040 44605
rect 10096 44549 10164 44605
rect 10220 44549 10230 44605
rect 9782 44539 10230 44549
rect 12054 45845 12502 45855
rect 12054 45789 12064 45845
rect 12120 45789 12188 45845
rect 12244 45789 12312 45845
rect 12368 45789 12436 45845
rect 12492 45789 12502 45845
rect 12054 45721 12502 45789
rect 12054 45665 12064 45721
rect 12120 45665 12188 45721
rect 12244 45665 12312 45721
rect 12368 45665 12436 45721
rect 12492 45665 12502 45721
rect 12054 45597 12502 45665
rect 12054 45541 12064 45597
rect 12120 45541 12188 45597
rect 12244 45541 12312 45597
rect 12368 45541 12436 45597
rect 12492 45541 12502 45597
rect 12054 45473 12502 45541
rect 12054 45417 12064 45473
rect 12120 45417 12188 45473
rect 12244 45417 12312 45473
rect 12368 45417 12436 45473
rect 12492 45417 12502 45473
rect 12054 45349 12502 45417
rect 12054 45293 12064 45349
rect 12120 45293 12188 45349
rect 12244 45293 12312 45349
rect 12368 45293 12436 45349
rect 12492 45293 12502 45349
rect 12054 45225 12502 45293
rect 12054 45169 12064 45225
rect 12120 45169 12188 45225
rect 12244 45169 12312 45225
rect 12368 45169 12436 45225
rect 12492 45169 12502 45225
rect 12054 45101 12502 45169
rect 12054 45045 12064 45101
rect 12120 45045 12188 45101
rect 12244 45045 12312 45101
rect 12368 45045 12436 45101
rect 12492 45045 12502 45101
rect 12054 44977 12502 45045
rect 12054 44921 12064 44977
rect 12120 44921 12188 44977
rect 12244 44921 12312 44977
rect 12368 44921 12436 44977
rect 12492 44921 12502 44977
rect 12054 44853 12502 44921
rect 12054 44797 12064 44853
rect 12120 44797 12188 44853
rect 12244 44797 12312 44853
rect 12368 44797 12436 44853
rect 12492 44797 12502 44853
rect 12054 44729 12502 44797
rect 12054 44673 12064 44729
rect 12120 44673 12188 44729
rect 12244 44673 12312 44729
rect 12368 44673 12436 44729
rect 12492 44673 12502 44729
rect 12054 44605 12502 44673
rect 12054 44549 12064 44605
rect 12120 44549 12188 44605
rect 12244 44549 12312 44605
rect 12368 44549 12436 44605
rect 12492 44549 12502 44605
rect 12054 44539 12502 44549
rect 13468 45845 13668 45855
rect 13468 45789 13478 45845
rect 13534 45789 13602 45845
rect 13658 45789 13668 45845
rect 13468 45721 13668 45789
rect 13468 45665 13478 45721
rect 13534 45665 13602 45721
rect 13658 45665 13668 45721
rect 13468 45597 13668 45665
rect 13468 45541 13478 45597
rect 13534 45541 13602 45597
rect 13658 45541 13668 45597
rect 13468 45473 13668 45541
rect 13468 45417 13478 45473
rect 13534 45417 13602 45473
rect 13658 45417 13668 45473
rect 13468 45349 13668 45417
rect 13468 45293 13478 45349
rect 13534 45293 13602 45349
rect 13658 45293 13668 45349
rect 13468 45225 13668 45293
rect 13468 45169 13478 45225
rect 13534 45169 13602 45225
rect 13658 45169 13668 45225
rect 13468 45101 13668 45169
rect 13468 45045 13478 45101
rect 13534 45045 13602 45101
rect 13658 45045 13668 45101
rect 13468 44977 13668 45045
rect 13468 44921 13478 44977
rect 13534 44921 13602 44977
rect 13658 44921 13668 44977
rect 13468 44853 13668 44921
rect 13468 44797 13478 44853
rect 13534 44797 13602 44853
rect 13658 44797 13668 44853
rect 13468 44729 13668 44797
rect 13468 44673 13478 44729
rect 13534 44673 13602 44729
rect 13658 44673 13668 44729
rect 13468 44605 13668 44673
rect 13468 44549 13478 44605
rect 13534 44549 13602 44605
rect 13658 44549 13668 44605
rect 13468 44539 13668 44549
rect 14326 45845 14774 45855
rect 14326 45789 14336 45845
rect 14392 45789 14460 45845
rect 14516 45789 14584 45845
rect 14640 45789 14708 45845
rect 14764 45789 14774 45845
rect 14326 45721 14774 45789
rect 14326 45665 14336 45721
rect 14392 45665 14460 45721
rect 14516 45665 14584 45721
rect 14640 45665 14708 45721
rect 14764 45665 14774 45721
rect 14326 45597 14774 45665
rect 14326 45541 14336 45597
rect 14392 45541 14460 45597
rect 14516 45541 14584 45597
rect 14640 45541 14708 45597
rect 14764 45541 14774 45597
rect 14326 45473 14774 45541
rect 14326 45417 14336 45473
rect 14392 45417 14460 45473
rect 14516 45417 14584 45473
rect 14640 45417 14708 45473
rect 14764 45417 14774 45473
rect 14326 45349 14774 45417
rect 14326 45293 14336 45349
rect 14392 45293 14460 45349
rect 14516 45293 14584 45349
rect 14640 45293 14708 45349
rect 14764 45293 14774 45349
rect 14326 45225 14774 45293
rect 14326 45169 14336 45225
rect 14392 45169 14460 45225
rect 14516 45169 14584 45225
rect 14640 45169 14708 45225
rect 14764 45169 14774 45225
rect 14326 45101 14774 45169
rect 14326 45045 14336 45101
rect 14392 45045 14460 45101
rect 14516 45045 14584 45101
rect 14640 45045 14708 45101
rect 14764 45045 14774 45101
rect 14326 44977 14774 45045
rect 14326 44921 14336 44977
rect 14392 44921 14460 44977
rect 14516 44921 14584 44977
rect 14640 44921 14708 44977
rect 14764 44921 14774 44977
rect 14326 44853 14774 44921
rect 14326 44797 14336 44853
rect 14392 44797 14460 44853
rect 14516 44797 14584 44853
rect 14640 44797 14708 44853
rect 14764 44797 14774 44853
rect 14326 44729 14774 44797
rect 14326 44673 14336 44729
rect 14392 44673 14460 44729
rect 14516 44673 14584 44729
rect 14640 44673 14708 44729
rect 14764 44673 14774 44729
rect 14326 44605 14774 44673
rect 14326 44549 14336 44605
rect 14392 44549 14460 44605
rect 14516 44549 14584 44605
rect 14640 44549 14708 44605
rect 14764 44549 14774 44605
rect 14326 44539 14774 44549
rect 1136 44245 1336 44255
rect 1136 44189 1146 44245
rect 1202 44189 1270 44245
rect 1326 44189 1336 44245
rect 1136 44121 1336 44189
rect 1136 44065 1146 44121
rect 1202 44065 1270 44121
rect 1326 44065 1336 44121
rect 1136 43997 1336 44065
rect 1136 43941 1146 43997
rect 1202 43941 1270 43997
rect 1326 43941 1336 43997
rect 1136 43873 1336 43941
rect 1136 43817 1146 43873
rect 1202 43817 1270 43873
rect 1326 43817 1336 43873
rect 1136 43749 1336 43817
rect 1136 43693 1146 43749
rect 1202 43693 1270 43749
rect 1326 43693 1336 43749
rect 1136 43625 1336 43693
rect 1136 43569 1146 43625
rect 1202 43569 1270 43625
rect 1326 43569 1336 43625
rect 1136 43501 1336 43569
rect 1136 43445 1146 43501
rect 1202 43445 1270 43501
rect 1326 43445 1336 43501
rect 1136 43377 1336 43445
rect 1136 43321 1146 43377
rect 1202 43321 1270 43377
rect 1326 43321 1336 43377
rect 1136 43253 1336 43321
rect 1136 43197 1146 43253
rect 1202 43197 1270 43253
rect 1326 43197 1336 43253
rect 1136 43129 1336 43197
rect 1136 43073 1146 43129
rect 1202 43073 1270 43129
rect 1326 43073 1336 43129
rect 1136 43005 1336 43073
rect 1136 42949 1146 43005
rect 1202 42949 1270 43005
rect 1326 42949 1336 43005
rect 1136 42939 1336 42949
rect 1994 44245 2442 44255
rect 1994 44189 2004 44245
rect 2060 44189 2128 44245
rect 2184 44189 2252 44245
rect 2308 44189 2376 44245
rect 2432 44189 2442 44245
rect 1994 44121 2442 44189
rect 1994 44065 2004 44121
rect 2060 44065 2128 44121
rect 2184 44065 2252 44121
rect 2308 44065 2376 44121
rect 2432 44065 2442 44121
rect 1994 43997 2442 44065
rect 1994 43941 2004 43997
rect 2060 43941 2128 43997
rect 2184 43941 2252 43997
rect 2308 43941 2376 43997
rect 2432 43941 2442 43997
rect 1994 43873 2442 43941
rect 1994 43817 2004 43873
rect 2060 43817 2128 43873
rect 2184 43817 2252 43873
rect 2308 43817 2376 43873
rect 2432 43817 2442 43873
rect 1994 43749 2442 43817
rect 1994 43693 2004 43749
rect 2060 43693 2128 43749
rect 2184 43693 2252 43749
rect 2308 43693 2376 43749
rect 2432 43693 2442 43749
rect 1994 43625 2442 43693
rect 1994 43569 2004 43625
rect 2060 43569 2128 43625
rect 2184 43569 2252 43625
rect 2308 43569 2376 43625
rect 2432 43569 2442 43625
rect 1994 43501 2442 43569
rect 1994 43445 2004 43501
rect 2060 43445 2128 43501
rect 2184 43445 2252 43501
rect 2308 43445 2376 43501
rect 2432 43445 2442 43501
rect 1994 43377 2442 43445
rect 1994 43321 2004 43377
rect 2060 43321 2128 43377
rect 2184 43321 2252 43377
rect 2308 43321 2376 43377
rect 2432 43321 2442 43377
rect 1994 43253 2442 43321
rect 1994 43197 2004 43253
rect 2060 43197 2128 43253
rect 2184 43197 2252 43253
rect 2308 43197 2376 43253
rect 2432 43197 2442 43253
rect 1994 43129 2442 43197
rect 1994 43073 2004 43129
rect 2060 43073 2128 43129
rect 2184 43073 2252 43129
rect 2308 43073 2376 43129
rect 2432 43073 2442 43129
rect 1994 43005 2442 43073
rect 1994 42949 2004 43005
rect 2060 42949 2128 43005
rect 2184 42949 2252 43005
rect 2308 42949 2376 43005
rect 2432 42949 2442 43005
rect 1994 42939 2442 42949
rect 3698 44245 4146 44255
rect 3698 44189 3708 44245
rect 3764 44189 3832 44245
rect 3888 44189 3956 44245
rect 4012 44189 4080 44245
rect 4136 44189 4146 44245
rect 3698 44121 4146 44189
rect 3698 44065 3708 44121
rect 3764 44065 3832 44121
rect 3888 44065 3956 44121
rect 4012 44065 4080 44121
rect 4136 44065 4146 44121
rect 3698 43997 4146 44065
rect 3698 43941 3708 43997
rect 3764 43941 3832 43997
rect 3888 43941 3956 43997
rect 4012 43941 4080 43997
rect 4136 43941 4146 43997
rect 3698 43873 4146 43941
rect 3698 43817 3708 43873
rect 3764 43817 3832 43873
rect 3888 43817 3956 43873
rect 4012 43817 4080 43873
rect 4136 43817 4146 43873
rect 3698 43749 4146 43817
rect 3698 43693 3708 43749
rect 3764 43693 3832 43749
rect 3888 43693 3956 43749
rect 4012 43693 4080 43749
rect 4136 43693 4146 43749
rect 3698 43625 4146 43693
rect 3698 43569 3708 43625
rect 3764 43569 3832 43625
rect 3888 43569 3956 43625
rect 4012 43569 4080 43625
rect 4136 43569 4146 43625
rect 3698 43501 4146 43569
rect 3698 43445 3708 43501
rect 3764 43445 3832 43501
rect 3888 43445 3956 43501
rect 4012 43445 4080 43501
rect 4136 43445 4146 43501
rect 3698 43377 4146 43445
rect 3698 43321 3708 43377
rect 3764 43321 3832 43377
rect 3888 43321 3956 43377
rect 4012 43321 4080 43377
rect 4136 43321 4146 43377
rect 3698 43253 4146 43321
rect 3698 43197 3708 43253
rect 3764 43197 3832 43253
rect 3888 43197 3956 43253
rect 4012 43197 4080 43253
rect 4136 43197 4146 43253
rect 3698 43129 4146 43197
rect 3698 43073 3708 43129
rect 3764 43073 3832 43129
rect 3888 43073 3956 43129
rect 4012 43073 4080 43129
rect 4136 43073 4146 43129
rect 3698 43005 4146 43073
rect 3698 42949 3708 43005
rect 3764 42949 3832 43005
rect 3888 42949 3956 43005
rect 4012 42949 4080 43005
rect 4136 42949 4146 43005
rect 3698 42939 4146 42949
rect 5970 44245 6418 44255
rect 5970 44189 5980 44245
rect 6036 44189 6104 44245
rect 6160 44189 6228 44245
rect 6284 44189 6352 44245
rect 6408 44189 6418 44245
rect 5970 44121 6418 44189
rect 5970 44065 5980 44121
rect 6036 44065 6104 44121
rect 6160 44065 6228 44121
rect 6284 44065 6352 44121
rect 6408 44065 6418 44121
rect 5970 43997 6418 44065
rect 5970 43941 5980 43997
rect 6036 43941 6104 43997
rect 6160 43941 6228 43997
rect 6284 43941 6352 43997
rect 6408 43941 6418 43997
rect 5970 43873 6418 43941
rect 5970 43817 5980 43873
rect 6036 43817 6104 43873
rect 6160 43817 6228 43873
rect 6284 43817 6352 43873
rect 6408 43817 6418 43873
rect 5970 43749 6418 43817
rect 5970 43693 5980 43749
rect 6036 43693 6104 43749
rect 6160 43693 6228 43749
rect 6284 43693 6352 43749
rect 6408 43693 6418 43749
rect 5970 43625 6418 43693
rect 5970 43569 5980 43625
rect 6036 43569 6104 43625
rect 6160 43569 6228 43625
rect 6284 43569 6352 43625
rect 6408 43569 6418 43625
rect 5970 43501 6418 43569
rect 5970 43445 5980 43501
rect 6036 43445 6104 43501
rect 6160 43445 6228 43501
rect 6284 43445 6352 43501
rect 6408 43445 6418 43501
rect 5970 43377 6418 43445
rect 5970 43321 5980 43377
rect 6036 43321 6104 43377
rect 6160 43321 6228 43377
rect 6284 43321 6352 43377
rect 6408 43321 6418 43377
rect 5970 43253 6418 43321
rect 5970 43197 5980 43253
rect 6036 43197 6104 43253
rect 6160 43197 6228 43253
rect 6284 43197 6352 43253
rect 6408 43197 6418 43253
rect 5970 43129 6418 43197
rect 5970 43073 5980 43129
rect 6036 43073 6104 43129
rect 6160 43073 6228 43129
rect 6284 43073 6352 43129
rect 6408 43073 6418 43129
rect 5970 43005 6418 43073
rect 5970 42949 5980 43005
rect 6036 42949 6104 43005
rect 6160 42949 6228 43005
rect 6284 42949 6352 43005
rect 6408 42949 6418 43005
rect 5970 42939 6418 42949
rect 8646 44245 9094 44255
rect 8646 44189 8656 44245
rect 8712 44189 8780 44245
rect 8836 44189 8904 44245
rect 8960 44189 9028 44245
rect 9084 44189 9094 44245
rect 8646 44121 9094 44189
rect 8646 44065 8656 44121
rect 8712 44065 8780 44121
rect 8836 44065 8904 44121
rect 8960 44065 9028 44121
rect 9084 44065 9094 44121
rect 8646 43997 9094 44065
rect 8646 43941 8656 43997
rect 8712 43941 8780 43997
rect 8836 43941 8904 43997
rect 8960 43941 9028 43997
rect 9084 43941 9094 43997
rect 8646 43873 9094 43941
rect 8646 43817 8656 43873
rect 8712 43817 8780 43873
rect 8836 43817 8904 43873
rect 8960 43817 9028 43873
rect 9084 43817 9094 43873
rect 8646 43749 9094 43817
rect 8646 43693 8656 43749
rect 8712 43693 8780 43749
rect 8836 43693 8904 43749
rect 8960 43693 9028 43749
rect 9084 43693 9094 43749
rect 8646 43625 9094 43693
rect 8646 43569 8656 43625
rect 8712 43569 8780 43625
rect 8836 43569 8904 43625
rect 8960 43569 9028 43625
rect 9084 43569 9094 43625
rect 8646 43501 9094 43569
rect 8646 43445 8656 43501
rect 8712 43445 8780 43501
rect 8836 43445 8904 43501
rect 8960 43445 9028 43501
rect 9084 43445 9094 43501
rect 8646 43377 9094 43445
rect 8646 43321 8656 43377
rect 8712 43321 8780 43377
rect 8836 43321 8904 43377
rect 8960 43321 9028 43377
rect 9084 43321 9094 43377
rect 8646 43253 9094 43321
rect 8646 43197 8656 43253
rect 8712 43197 8780 43253
rect 8836 43197 8904 43253
rect 8960 43197 9028 43253
rect 9084 43197 9094 43253
rect 8646 43129 9094 43197
rect 8646 43073 8656 43129
rect 8712 43073 8780 43129
rect 8836 43073 8904 43129
rect 8960 43073 9028 43129
rect 9084 43073 9094 43129
rect 8646 43005 9094 43073
rect 8646 42949 8656 43005
rect 8712 42949 8780 43005
rect 8836 42949 8904 43005
rect 8960 42949 9028 43005
rect 9084 42949 9094 43005
rect 8646 42939 9094 42949
rect 10918 44245 11366 44255
rect 10918 44189 10928 44245
rect 10984 44189 11052 44245
rect 11108 44189 11176 44245
rect 11232 44189 11300 44245
rect 11356 44189 11366 44245
rect 10918 44121 11366 44189
rect 10918 44065 10928 44121
rect 10984 44065 11052 44121
rect 11108 44065 11176 44121
rect 11232 44065 11300 44121
rect 11356 44065 11366 44121
rect 10918 43997 11366 44065
rect 10918 43941 10928 43997
rect 10984 43941 11052 43997
rect 11108 43941 11176 43997
rect 11232 43941 11300 43997
rect 11356 43941 11366 43997
rect 10918 43873 11366 43941
rect 10918 43817 10928 43873
rect 10984 43817 11052 43873
rect 11108 43817 11176 43873
rect 11232 43817 11300 43873
rect 11356 43817 11366 43873
rect 10918 43749 11366 43817
rect 10918 43693 10928 43749
rect 10984 43693 11052 43749
rect 11108 43693 11176 43749
rect 11232 43693 11300 43749
rect 11356 43693 11366 43749
rect 10918 43625 11366 43693
rect 10918 43569 10928 43625
rect 10984 43569 11052 43625
rect 11108 43569 11176 43625
rect 11232 43569 11300 43625
rect 11356 43569 11366 43625
rect 10918 43501 11366 43569
rect 10918 43445 10928 43501
rect 10984 43445 11052 43501
rect 11108 43445 11176 43501
rect 11232 43445 11300 43501
rect 11356 43445 11366 43501
rect 10918 43377 11366 43445
rect 10918 43321 10928 43377
rect 10984 43321 11052 43377
rect 11108 43321 11176 43377
rect 11232 43321 11300 43377
rect 11356 43321 11366 43377
rect 10918 43253 11366 43321
rect 10918 43197 10928 43253
rect 10984 43197 11052 43253
rect 11108 43197 11176 43253
rect 11232 43197 11300 43253
rect 11356 43197 11366 43253
rect 10918 43129 11366 43197
rect 10918 43073 10928 43129
rect 10984 43073 11052 43129
rect 11108 43073 11176 43129
rect 11232 43073 11300 43129
rect 11356 43073 11366 43129
rect 10918 43005 11366 43073
rect 10918 42949 10928 43005
rect 10984 42949 11052 43005
rect 11108 42949 11176 43005
rect 11232 42949 11300 43005
rect 11356 42949 11366 43005
rect 10918 42939 11366 42949
rect 12622 44245 13070 44255
rect 12622 44189 12632 44245
rect 12688 44189 12756 44245
rect 12812 44189 12880 44245
rect 12936 44189 13004 44245
rect 13060 44189 13070 44245
rect 12622 44121 13070 44189
rect 12622 44065 12632 44121
rect 12688 44065 12756 44121
rect 12812 44065 12880 44121
rect 12936 44065 13004 44121
rect 13060 44065 13070 44121
rect 12622 43997 13070 44065
rect 12622 43941 12632 43997
rect 12688 43941 12756 43997
rect 12812 43941 12880 43997
rect 12936 43941 13004 43997
rect 13060 43941 13070 43997
rect 12622 43873 13070 43941
rect 12622 43817 12632 43873
rect 12688 43817 12756 43873
rect 12812 43817 12880 43873
rect 12936 43817 13004 43873
rect 13060 43817 13070 43873
rect 12622 43749 13070 43817
rect 12622 43693 12632 43749
rect 12688 43693 12756 43749
rect 12812 43693 12880 43749
rect 12936 43693 13004 43749
rect 13060 43693 13070 43749
rect 12622 43625 13070 43693
rect 12622 43569 12632 43625
rect 12688 43569 12756 43625
rect 12812 43569 12880 43625
rect 12936 43569 13004 43625
rect 13060 43569 13070 43625
rect 12622 43501 13070 43569
rect 12622 43445 12632 43501
rect 12688 43445 12756 43501
rect 12812 43445 12880 43501
rect 12936 43445 13004 43501
rect 13060 43445 13070 43501
rect 12622 43377 13070 43445
rect 12622 43321 12632 43377
rect 12688 43321 12756 43377
rect 12812 43321 12880 43377
rect 12936 43321 13004 43377
rect 13060 43321 13070 43377
rect 12622 43253 13070 43321
rect 12622 43197 12632 43253
rect 12688 43197 12756 43253
rect 12812 43197 12880 43253
rect 12936 43197 13004 43253
rect 13060 43197 13070 43253
rect 12622 43129 13070 43197
rect 12622 43073 12632 43129
rect 12688 43073 12756 43129
rect 12812 43073 12880 43129
rect 12936 43073 13004 43129
rect 13060 43073 13070 43129
rect 12622 43005 13070 43073
rect 12622 42949 12632 43005
rect 12688 42949 12756 43005
rect 12812 42949 12880 43005
rect 12936 42949 13004 43005
rect 13060 42949 13070 43005
rect 12622 42939 13070 42949
rect 13758 44245 14206 44255
rect 13758 44189 13768 44245
rect 13824 44189 13892 44245
rect 13948 44189 14016 44245
rect 14072 44189 14140 44245
rect 14196 44189 14206 44245
rect 13758 44121 14206 44189
rect 13758 44065 13768 44121
rect 13824 44065 13892 44121
rect 13948 44065 14016 44121
rect 14072 44065 14140 44121
rect 14196 44065 14206 44121
rect 13758 43997 14206 44065
rect 13758 43941 13768 43997
rect 13824 43941 13892 43997
rect 13948 43941 14016 43997
rect 14072 43941 14140 43997
rect 14196 43941 14206 43997
rect 13758 43873 14206 43941
rect 13758 43817 13768 43873
rect 13824 43817 13892 43873
rect 13948 43817 14016 43873
rect 14072 43817 14140 43873
rect 14196 43817 14206 43873
rect 13758 43749 14206 43817
rect 13758 43693 13768 43749
rect 13824 43693 13892 43749
rect 13948 43693 14016 43749
rect 14072 43693 14140 43749
rect 14196 43693 14206 43749
rect 13758 43625 14206 43693
rect 13758 43569 13768 43625
rect 13824 43569 13892 43625
rect 13948 43569 14016 43625
rect 14072 43569 14140 43625
rect 14196 43569 14206 43625
rect 13758 43501 14206 43569
rect 13758 43445 13768 43501
rect 13824 43445 13892 43501
rect 13948 43445 14016 43501
rect 14072 43445 14140 43501
rect 14196 43445 14206 43501
rect 13758 43377 14206 43445
rect 13758 43321 13768 43377
rect 13824 43321 13892 43377
rect 13948 43321 14016 43377
rect 14072 43321 14140 43377
rect 14196 43321 14206 43377
rect 13758 43253 14206 43321
rect 13758 43197 13768 43253
rect 13824 43197 13892 43253
rect 13948 43197 14016 43253
rect 14072 43197 14140 43253
rect 14196 43197 14206 43253
rect 13758 43129 14206 43197
rect 13758 43073 13768 43129
rect 13824 43073 13892 43129
rect 13948 43073 14016 43129
rect 14072 43073 14140 43129
rect 14196 43073 14206 43129
rect 13758 43005 14206 43073
rect 13758 42949 13768 43005
rect 13824 42949 13892 43005
rect 13948 42949 14016 43005
rect 14072 42949 14140 43005
rect 14196 42949 14206 43005
rect 13758 42939 14206 42949
rect 1136 42645 1336 42655
rect 1136 42589 1146 42645
rect 1202 42589 1270 42645
rect 1326 42589 1336 42645
rect 1136 42521 1336 42589
rect 1136 42465 1146 42521
rect 1202 42465 1270 42521
rect 1326 42465 1336 42521
rect 1136 42397 1336 42465
rect 1136 42341 1146 42397
rect 1202 42341 1270 42397
rect 1326 42341 1336 42397
rect 1136 42273 1336 42341
rect 1136 42217 1146 42273
rect 1202 42217 1270 42273
rect 1326 42217 1336 42273
rect 1136 42149 1336 42217
rect 1136 42093 1146 42149
rect 1202 42093 1270 42149
rect 1326 42093 1336 42149
rect 1136 42025 1336 42093
rect 1136 41969 1146 42025
rect 1202 41969 1270 42025
rect 1326 41969 1336 42025
rect 1136 41901 1336 41969
rect 1136 41845 1146 41901
rect 1202 41845 1270 41901
rect 1326 41845 1336 41901
rect 1136 41777 1336 41845
rect 1136 41721 1146 41777
rect 1202 41721 1270 41777
rect 1326 41721 1336 41777
rect 1136 41653 1336 41721
rect 1136 41597 1146 41653
rect 1202 41597 1270 41653
rect 1326 41597 1336 41653
rect 1136 41529 1336 41597
rect 1136 41473 1146 41529
rect 1202 41473 1270 41529
rect 1326 41473 1336 41529
rect 1136 41405 1336 41473
rect 1136 41349 1146 41405
rect 1202 41349 1270 41405
rect 1326 41349 1336 41405
rect 1136 41339 1336 41349
rect 1994 42645 2442 42655
rect 1994 42589 2004 42645
rect 2060 42589 2128 42645
rect 2184 42589 2252 42645
rect 2308 42589 2376 42645
rect 2432 42589 2442 42645
rect 1994 42521 2442 42589
rect 1994 42465 2004 42521
rect 2060 42465 2128 42521
rect 2184 42465 2252 42521
rect 2308 42465 2376 42521
rect 2432 42465 2442 42521
rect 1994 42397 2442 42465
rect 1994 42341 2004 42397
rect 2060 42341 2128 42397
rect 2184 42341 2252 42397
rect 2308 42341 2376 42397
rect 2432 42341 2442 42397
rect 1994 42273 2442 42341
rect 1994 42217 2004 42273
rect 2060 42217 2128 42273
rect 2184 42217 2252 42273
rect 2308 42217 2376 42273
rect 2432 42217 2442 42273
rect 1994 42149 2442 42217
rect 1994 42093 2004 42149
rect 2060 42093 2128 42149
rect 2184 42093 2252 42149
rect 2308 42093 2376 42149
rect 2432 42093 2442 42149
rect 1994 42025 2442 42093
rect 1994 41969 2004 42025
rect 2060 41969 2128 42025
rect 2184 41969 2252 42025
rect 2308 41969 2376 42025
rect 2432 41969 2442 42025
rect 1994 41901 2442 41969
rect 1994 41845 2004 41901
rect 2060 41845 2128 41901
rect 2184 41845 2252 41901
rect 2308 41845 2376 41901
rect 2432 41845 2442 41901
rect 1994 41777 2442 41845
rect 1994 41721 2004 41777
rect 2060 41721 2128 41777
rect 2184 41721 2252 41777
rect 2308 41721 2376 41777
rect 2432 41721 2442 41777
rect 1994 41653 2442 41721
rect 1994 41597 2004 41653
rect 2060 41597 2128 41653
rect 2184 41597 2252 41653
rect 2308 41597 2376 41653
rect 2432 41597 2442 41653
rect 1994 41529 2442 41597
rect 1994 41473 2004 41529
rect 2060 41473 2128 41529
rect 2184 41473 2252 41529
rect 2308 41473 2376 41529
rect 2432 41473 2442 41529
rect 1994 41405 2442 41473
rect 1994 41349 2004 41405
rect 2060 41349 2128 41405
rect 2184 41349 2252 41405
rect 2308 41349 2376 41405
rect 2432 41349 2442 41405
rect 1994 41339 2442 41349
rect 3698 42645 4146 42655
rect 3698 42589 3708 42645
rect 3764 42589 3832 42645
rect 3888 42589 3956 42645
rect 4012 42589 4080 42645
rect 4136 42589 4146 42645
rect 3698 42521 4146 42589
rect 3698 42465 3708 42521
rect 3764 42465 3832 42521
rect 3888 42465 3956 42521
rect 4012 42465 4080 42521
rect 4136 42465 4146 42521
rect 3698 42397 4146 42465
rect 3698 42341 3708 42397
rect 3764 42341 3832 42397
rect 3888 42341 3956 42397
rect 4012 42341 4080 42397
rect 4136 42341 4146 42397
rect 3698 42273 4146 42341
rect 3698 42217 3708 42273
rect 3764 42217 3832 42273
rect 3888 42217 3956 42273
rect 4012 42217 4080 42273
rect 4136 42217 4146 42273
rect 3698 42149 4146 42217
rect 3698 42093 3708 42149
rect 3764 42093 3832 42149
rect 3888 42093 3956 42149
rect 4012 42093 4080 42149
rect 4136 42093 4146 42149
rect 3698 42025 4146 42093
rect 3698 41969 3708 42025
rect 3764 41969 3832 42025
rect 3888 41969 3956 42025
rect 4012 41969 4080 42025
rect 4136 41969 4146 42025
rect 3698 41901 4146 41969
rect 3698 41845 3708 41901
rect 3764 41845 3832 41901
rect 3888 41845 3956 41901
rect 4012 41845 4080 41901
rect 4136 41845 4146 41901
rect 3698 41777 4146 41845
rect 3698 41721 3708 41777
rect 3764 41721 3832 41777
rect 3888 41721 3956 41777
rect 4012 41721 4080 41777
rect 4136 41721 4146 41777
rect 3698 41653 4146 41721
rect 3698 41597 3708 41653
rect 3764 41597 3832 41653
rect 3888 41597 3956 41653
rect 4012 41597 4080 41653
rect 4136 41597 4146 41653
rect 3698 41529 4146 41597
rect 3698 41473 3708 41529
rect 3764 41473 3832 41529
rect 3888 41473 3956 41529
rect 4012 41473 4080 41529
rect 4136 41473 4146 41529
rect 3698 41405 4146 41473
rect 3698 41349 3708 41405
rect 3764 41349 3832 41405
rect 3888 41349 3956 41405
rect 4012 41349 4080 41405
rect 4136 41349 4146 41405
rect 3698 41339 4146 41349
rect 5970 42645 6418 42655
rect 5970 42589 5980 42645
rect 6036 42589 6104 42645
rect 6160 42589 6228 42645
rect 6284 42589 6352 42645
rect 6408 42589 6418 42645
rect 5970 42521 6418 42589
rect 5970 42465 5980 42521
rect 6036 42465 6104 42521
rect 6160 42465 6228 42521
rect 6284 42465 6352 42521
rect 6408 42465 6418 42521
rect 5970 42397 6418 42465
rect 5970 42341 5980 42397
rect 6036 42341 6104 42397
rect 6160 42341 6228 42397
rect 6284 42341 6352 42397
rect 6408 42341 6418 42397
rect 5970 42273 6418 42341
rect 5970 42217 5980 42273
rect 6036 42217 6104 42273
rect 6160 42217 6228 42273
rect 6284 42217 6352 42273
rect 6408 42217 6418 42273
rect 5970 42149 6418 42217
rect 5970 42093 5980 42149
rect 6036 42093 6104 42149
rect 6160 42093 6228 42149
rect 6284 42093 6352 42149
rect 6408 42093 6418 42149
rect 5970 42025 6418 42093
rect 5970 41969 5980 42025
rect 6036 41969 6104 42025
rect 6160 41969 6228 42025
rect 6284 41969 6352 42025
rect 6408 41969 6418 42025
rect 5970 41901 6418 41969
rect 5970 41845 5980 41901
rect 6036 41845 6104 41901
rect 6160 41845 6228 41901
rect 6284 41845 6352 41901
rect 6408 41845 6418 41901
rect 5970 41777 6418 41845
rect 5970 41721 5980 41777
rect 6036 41721 6104 41777
rect 6160 41721 6228 41777
rect 6284 41721 6352 41777
rect 6408 41721 6418 41777
rect 5970 41653 6418 41721
rect 5970 41597 5980 41653
rect 6036 41597 6104 41653
rect 6160 41597 6228 41653
rect 6284 41597 6352 41653
rect 6408 41597 6418 41653
rect 5970 41529 6418 41597
rect 5970 41473 5980 41529
rect 6036 41473 6104 41529
rect 6160 41473 6228 41529
rect 6284 41473 6352 41529
rect 6408 41473 6418 41529
rect 5970 41405 6418 41473
rect 5970 41349 5980 41405
rect 6036 41349 6104 41405
rect 6160 41349 6228 41405
rect 6284 41349 6352 41405
rect 6408 41349 6418 41405
rect 5970 41339 6418 41349
rect 8646 42645 9094 42655
rect 8646 42589 8656 42645
rect 8712 42589 8780 42645
rect 8836 42589 8904 42645
rect 8960 42589 9028 42645
rect 9084 42589 9094 42645
rect 8646 42521 9094 42589
rect 8646 42465 8656 42521
rect 8712 42465 8780 42521
rect 8836 42465 8904 42521
rect 8960 42465 9028 42521
rect 9084 42465 9094 42521
rect 8646 42397 9094 42465
rect 8646 42341 8656 42397
rect 8712 42341 8780 42397
rect 8836 42341 8904 42397
rect 8960 42341 9028 42397
rect 9084 42341 9094 42397
rect 8646 42273 9094 42341
rect 8646 42217 8656 42273
rect 8712 42217 8780 42273
rect 8836 42217 8904 42273
rect 8960 42217 9028 42273
rect 9084 42217 9094 42273
rect 8646 42149 9094 42217
rect 8646 42093 8656 42149
rect 8712 42093 8780 42149
rect 8836 42093 8904 42149
rect 8960 42093 9028 42149
rect 9084 42093 9094 42149
rect 8646 42025 9094 42093
rect 8646 41969 8656 42025
rect 8712 41969 8780 42025
rect 8836 41969 8904 42025
rect 8960 41969 9028 42025
rect 9084 41969 9094 42025
rect 8646 41901 9094 41969
rect 8646 41845 8656 41901
rect 8712 41845 8780 41901
rect 8836 41845 8904 41901
rect 8960 41845 9028 41901
rect 9084 41845 9094 41901
rect 8646 41777 9094 41845
rect 8646 41721 8656 41777
rect 8712 41721 8780 41777
rect 8836 41721 8904 41777
rect 8960 41721 9028 41777
rect 9084 41721 9094 41777
rect 8646 41653 9094 41721
rect 8646 41597 8656 41653
rect 8712 41597 8780 41653
rect 8836 41597 8904 41653
rect 8960 41597 9028 41653
rect 9084 41597 9094 41653
rect 8646 41529 9094 41597
rect 8646 41473 8656 41529
rect 8712 41473 8780 41529
rect 8836 41473 8904 41529
rect 8960 41473 9028 41529
rect 9084 41473 9094 41529
rect 8646 41405 9094 41473
rect 8646 41349 8656 41405
rect 8712 41349 8780 41405
rect 8836 41349 8904 41405
rect 8960 41349 9028 41405
rect 9084 41349 9094 41405
rect 8646 41339 9094 41349
rect 10918 42645 11366 42655
rect 10918 42589 10928 42645
rect 10984 42589 11052 42645
rect 11108 42589 11176 42645
rect 11232 42589 11300 42645
rect 11356 42589 11366 42645
rect 10918 42521 11366 42589
rect 10918 42465 10928 42521
rect 10984 42465 11052 42521
rect 11108 42465 11176 42521
rect 11232 42465 11300 42521
rect 11356 42465 11366 42521
rect 10918 42397 11366 42465
rect 10918 42341 10928 42397
rect 10984 42341 11052 42397
rect 11108 42341 11176 42397
rect 11232 42341 11300 42397
rect 11356 42341 11366 42397
rect 10918 42273 11366 42341
rect 10918 42217 10928 42273
rect 10984 42217 11052 42273
rect 11108 42217 11176 42273
rect 11232 42217 11300 42273
rect 11356 42217 11366 42273
rect 10918 42149 11366 42217
rect 10918 42093 10928 42149
rect 10984 42093 11052 42149
rect 11108 42093 11176 42149
rect 11232 42093 11300 42149
rect 11356 42093 11366 42149
rect 10918 42025 11366 42093
rect 10918 41969 10928 42025
rect 10984 41969 11052 42025
rect 11108 41969 11176 42025
rect 11232 41969 11300 42025
rect 11356 41969 11366 42025
rect 10918 41901 11366 41969
rect 10918 41845 10928 41901
rect 10984 41845 11052 41901
rect 11108 41845 11176 41901
rect 11232 41845 11300 41901
rect 11356 41845 11366 41901
rect 10918 41777 11366 41845
rect 10918 41721 10928 41777
rect 10984 41721 11052 41777
rect 11108 41721 11176 41777
rect 11232 41721 11300 41777
rect 11356 41721 11366 41777
rect 10918 41653 11366 41721
rect 10918 41597 10928 41653
rect 10984 41597 11052 41653
rect 11108 41597 11176 41653
rect 11232 41597 11300 41653
rect 11356 41597 11366 41653
rect 10918 41529 11366 41597
rect 10918 41473 10928 41529
rect 10984 41473 11052 41529
rect 11108 41473 11176 41529
rect 11232 41473 11300 41529
rect 11356 41473 11366 41529
rect 10918 41405 11366 41473
rect 10918 41349 10928 41405
rect 10984 41349 11052 41405
rect 11108 41349 11176 41405
rect 11232 41349 11300 41405
rect 11356 41349 11366 41405
rect 10918 41339 11366 41349
rect 12622 42645 13070 42655
rect 12622 42589 12632 42645
rect 12688 42589 12756 42645
rect 12812 42589 12880 42645
rect 12936 42589 13004 42645
rect 13060 42589 13070 42645
rect 12622 42521 13070 42589
rect 12622 42465 12632 42521
rect 12688 42465 12756 42521
rect 12812 42465 12880 42521
rect 12936 42465 13004 42521
rect 13060 42465 13070 42521
rect 12622 42397 13070 42465
rect 12622 42341 12632 42397
rect 12688 42341 12756 42397
rect 12812 42341 12880 42397
rect 12936 42341 13004 42397
rect 13060 42341 13070 42397
rect 12622 42273 13070 42341
rect 12622 42217 12632 42273
rect 12688 42217 12756 42273
rect 12812 42217 12880 42273
rect 12936 42217 13004 42273
rect 13060 42217 13070 42273
rect 12622 42149 13070 42217
rect 12622 42093 12632 42149
rect 12688 42093 12756 42149
rect 12812 42093 12880 42149
rect 12936 42093 13004 42149
rect 13060 42093 13070 42149
rect 12622 42025 13070 42093
rect 12622 41969 12632 42025
rect 12688 41969 12756 42025
rect 12812 41969 12880 42025
rect 12936 41969 13004 42025
rect 13060 41969 13070 42025
rect 12622 41901 13070 41969
rect 12622 41845 12632 41901
rect 12688 41845 12756 41901
rect 12812 41845 12880 41901
rect 12936 41845 13004 41901
rect 13060 41845 13070 41901
rect 12622 41777 13070 41845
rect 12622 41721 12632 41777
rect 12688 41721 12756 41777
rect 12812 41721 12880 41777
rect 12936 41721 13004 41777
rect 13060 41721 13070 41777
rect 12622 41653 13070 41721
rect 12622 41597 12632 41653
rect 12688 41597 12756 41653
rect 12812 41597 12880 41653
rect 12936 41597 13004 41653
rect 13060 41597 13070 41653
rect 12622 41529 13070 41597
rect 12622 41473 12632 41529
rect 12688 41473 12756 41529
rect 12812 41473 12880 41529
rect 12936 41473 13004 41529
rect 13060 41473 13070 41529
rect 12622 41405 13070 41473
rect 12622 41349 12632 41405
rect 12688 41349 12756 41405
rect 12812 41349 12880 41405
rect 12936 41349 13004 41405
rect 13060 41349 13070 41405
rect 12622 41339 13070 41349
rect 13758 42645 14206 42655
rect 13758 42589 13768 42645
rect 13824 42589 13892 42645
rect 13948 42589 14016 42645
rect 14072 42589 14140 42645
rect 14196 42589 14206 42645
rect 13758 42521 14206 42589
rect 13758 42465 13768 42521
rect 13824 42465 13892 42521
rect 13948 42465 14016 42521
rect 14072 42465 14140 42521
rect 14196 42465 14206 42521
rect 13758 42397 14206 42465
rect 13758 42341 13768 42397
rect 13824 42341 13892 42397
rect 13948 42341 14016 42397
rect 14072 42341 14140 42397
rect 14196 42341 14206 42397
rect 13758 42273 14206 42341
rect 13758 42217 13768 42273
rect 13824 42217 13892 42273
rect 13948 42217 14016 42273
rect 14072 42217 14140 42273
rect 14196 42217 14206 42273
rect 13758 42149 14206 42217
rect 13758 42093 13768 42149
rect 13824 42093 13892 42149
rect 13948 42093 14016 42149
rect 14072 42093 14140 42149
rect 14196 42093 14206 42149
rect 13758 42025 14206 42093
rect 13758 41969 13768 42025
rect 13824 41969 13892 42025
rect 13948 41969 14016 42025
rect 14072 41969 14140 42025
rect 14196 41969 14206 42025
rect 13758 41901 14206 41969
rect 13758 41845 13768 41901
rect 13824 41845 13892 41901
rect 13948 41845 14016 41901
rect 14072 41845 14140 41901
rect 14196 41845 14206 41901
rect 13758 41777 14206 41845
rect 13758 41721 13768 41777
rect 13824 41721 13892 41777
rect 13948 41721 14016 41777
rect 14072 41721 14140 41777
rect 14196 41721 14206 41777
rect 13758 41653 14206 41721
rect 13758 41597 13768 41653
rect 13824 41597 13892 41653
rect 13948 41597 14016 41653
rect 14072 41597 14140 41653
rect 14196 41597 14206 41653
rect 13758 41529 14206 41597
rect 13758 41473 13768 41529
rect 13824 41473 13892 41529
rect 13948 41473 14016 41529
rect 14072 41473 14140 41529
rect 14196 41473 14206 41529
rect 13758 41405 14206 41473
rect 13758 41349 13768 41405
rect 13824 41349 13892 41405
rect 13948 41349 14016 41405
rect 14072 41349 14140 41405
rect 14196 41349 14206 41405
rect 13758 41339 14206 41349
rect 1136 41045 1336 41055
rect 1136 40989 1146 41045
rect 1202 40989 1270 41045
rect 1326 40989 1336 41045
rect 1136 40921 1336 40989
rect 1136 40865 1146 40921
rect 1202 40865 1270 40921
rect 1326 40865 1336 40921
rect 1136 40797 1336 40865
rect 1136 40741 1146 40797
rect 1202 40741 1270 40797
rect 1326 40741 1336 40797
rect 1136 40673 1336 40741
rect 1136 40617 1146 40673
rect 1202 40617 1270 40673
rect 1326 40617 1336 40673
rect 1136 40549 1336 40617
rect 1136 40493 1146 40549
rect 1202 40493 1270 40549
rect 1326 40493 1336 40549
rect 1136 40425 1336 40493
rect 1136 40369 1146 40425
rect 1202 40369 1270 40425
rect 1326 40369 1336 40425
rect 1136 40301 1336 40369
rect 1136 40245 1146 40301
rect 1202 40245 1270 40301
rect 1326 40245 1336 40301
rect 1136 40177 1336 40245
rect 1136 40121 1146 40177
rect 1202 40121 1270 40177
rect 1326 40121 1336 40177
rect 1136 40053 1336 40121
rect 1136 39997 1146 40053
rect 1202 39997 1270 40053
rect 1326 39997 1336 40053
rect 1136 39929 1336 39997
rect 1136 39873 1146 39929
rect 1202 39873 1270 39929
rect 1326 39873 1336 39929
rect 1136 39805 1336 39873
rect 1136 39749 1146 39805
rect 1202 39749 1270 39805
rect 1326 39749 1336 39805
rect 1136 39739 1336 39749
rect 1994 41045 2442 41055
rect 1994 40989 2004 41045
rect 2060 40989 2128 41045
rect 2184 40989 2252 41045
rect 2308 40989 2376 41045
rect 2432 40989 2442 41045
rect 1994 40921 2442 40989
rect 1994 40865 2004 40921
rect 2060 40865 2128 40921
rect 2184 40865 2252 40921
rect 2308 40865 2376 40921
rect 2432 40865 2442 40921
rect 1994 40797 2442 40865
rect 1994 40741 2004 40797
rect 2060 40741 2128 40797
rect 2184 40741 2252 40797
rect 2308 40741 2376 40797
rect 2432 40741 2442 40797
rect 1994 40673 2442 40741
rect 1994 40617 2004 40673
rect 2060 40617 2128 40673
rect 2184 40617 2252 40673
rect 2308 40617 2376 40673
rect 2432 40617 2442 40673
rect 1994 40549 2442 40617
rect 1994 40493 2004 40549
rect 2060 40493 2128 40549
rect 2184 40493 2252 40549
rect 2308 40493 2376 40549
rect 2432 40493 2442 40549
rect 1994 40425 2442 40493
rect 1994 40369 2004 40425
rect 2060 40369 2128 40425
rect 2184 40369 2252 40425
rect 2308 40369 2376 40425
rect 2432 40369 2442 40425
rect 1994 40301 2442 40369
rect 1994 40245 2004 40301
rect 2060 40245 2128 40301
rect 2184 40245 2252 40301
rect 2308 40245 2376 40301
rect 2432 40245 2442 40301
rect 1994 40177 2442 40245
rect 1994 40121 2004 40177
rect 2060 40121 2128 40177
rect 2184 40121 2252 40177
rect 2308 40121 2376 40177
rect 2432 40121 2442 40177
rect 1994 40053 2442 40121
rect 1994 39997 2004 40053
rect 2060 39997 2128 40053
rect 2184 39997 2252 40053
rect 2308 39997 2376 40053
rect 2432 39997 2442 40053
rect 1994 39929 2442 39997
rect 1994 39873 2004 39929
rect 2060 39873 2128 39929
rect 2184 39873 2252 39929
rect 2308 39873 2376 39929
rect 2432 39873 2442 39929
rect 1994 39805 2442 39873
rect 1994 39749 2004 39805
rect 2060 39749 2128 39805
rect 2184 39749 2252 39805
rect 2308 39749 2376 39805
rect 2432 39749 2442 39805
rect 1994 39739 2442 39749
rect 3698 41045 4146 41055
rect 3698 40989 3708 41045
rect 3764 40989 3832 41045
rect 3888 40989 3956 41045
rect 4012 40989 4080 41045
rect 4136 40989 4146 41045
rect 3698 40921 4146 40989
rect 3698 40865 3708 40921
rect 3764 40865 3832 40921
rect 3888 40865 3956 40921
rect 4012 40865 4080 40921
rect 4136 40865 4146 40921
rect 3698 40797 4146 40865
rect 3698 40741 3708 40797
rect 3764 40741 3832 40797
rect 3888 40741 3956 40797
rect 4012 40741 4080 40797
rect 4136 40741 4146 40797
rect 3698 40673 4146 40741
rect 3698 40617 3708 40673
rect 3764 40617 3832 40673
rect 3888 40617 3956 40673
rect 4012 40617 4080 40673
rect 4136 40617 4146 40673
rect 3698 40549 4146 40617
rect 3698 40493 3708 40549
rect 3764 40493 3832 40549
rect 3888 40493 3956 40549
rect 4012 40493 4080 40549
rect 4136 40493 4146 40549
rect 3698 40425 4146 40493
rect 3698 40369 3708 40425
rect 3764 40369 3832 40425
rect 3888 40369 3956 40425
rect 4012 40369 4080 40425
rect 4136 40369 4146 40425
rect 3698 40301 4146 40369
rect 3698 40245 3708 40301
rect 3764 40245 3832 40301
rect 3888 40245 3956 40301
rect 4012 40245 4080 40301
rect 4136 40245 4146 40301
rect 3698 40177 4146 40245
rect 3698 40121 3708 40177
rect 3764 40121 3832 40177
rect 3888 40121 3956 40177
rect 4012 40121 4080 40177
rect 4136 40121 4146 40177
rect 3698 40053 4146 40121
rect 3698 39997 3708 40053
rect 3764 39997 3832 40053
rect 3888 39997 3956 40053
rect 4012 39997 4080 40053
rect 4136 39997 4146 40053
rect 3698 39929 4146 39997
rect 3698 39873 3708 39929
rect 3764 39873 3832 39929
rect 3888 39873 3956 39929
rect 4012 39873 4080 39929
rect 4136 39873 4146 39929
rect 3698 39805 4146 39873
rect 3698 39749 3708 39805
rect 3764 39749 3832 39805
rect 3888 39749 3956 39805
rect 4012 39749 4080 39805
rect 4136 39749 4146 39805
rect 3698 39739 4146 39749
rect 5970 41045 6418 41055
rect 5970 40989 5980 41045
rect 6036 40989 6104 41045
rect 6160 40989 6228 41045
rect 6284 40989 6352 41045
rect 6408 40989 6418 41045
rect 5970 40921 6418 40989
rect 5970 40865 5980 40921
rect 6036 40865 6104 40921
rect 6160 40865 6228 40921
rect 6284 40865 6352 40921
rect 6408 40865 6418 40921
rect 5970 40797 6418 40865
rect 5970 40741 5980 40797
rect 6036 40741 6104 40797
rect 6160 40741 6228 40797
rect 6284 40741 6352 40797
rect 6408 40741 6418 40797
rect 5970 40673 6418 40741
rect 5970 40617 5980 40673
rect 6036 40617 6104 40673
rect 6160 40617 6228 40673
rect 6284 40617 6352 40673
rect 6408 40617 6418 40673
rect 5970 40549 6418 40617
rect 5970 40493 5980 40549
rect 6036 40493 6104 40549
rect 6160 40493 6228 40549
rect 6284 40493 6352 40549
rect 6408 40493 6418 40549
rect 5970 40425 6418 40493
rect 5970 40369 5980 40425
rect 6036 40369 6104 40425
rect 6160 40369 6228 40425
rect 6284 40369 6352 40425
rect 6408 40369 6418 40425
rect 5970 40301 6418 40369
rect 5970 40245 5980 40301
rect 6036 40245 6104 40301
rect 6160 40245 6228 40301
rect 6284 40245 6352 40301
rect 6408 40245 6418 40301
rect 5970 40177 6418 40245
rect 5970 40121 5980 40177
rect 6036 40121 6104 40177
rect 6160 40121 6228 40177
rect 6284 40121 6352 40177
rect 6408 40121 6418 40177
rect 5970 40053 6418 40121
rect 5970 39997 5980 40053
rect 6036 39997 6104 40053
rect 6160 39997 6228 40053
rect 6284 39997 6352 40053
rect 6408 39997 6418 40053
rect 5970 39929 6418 39997
rect 5970 39873 5980 39929
rect 6036 39873 6104 39929
rect 6160 39873 6228 39929
rect 6284 39873 6352 39929
rect 6408 39873 6418 39929
rect 5970 39805 6418 39873
rect 5970 39749 5980 39805
rect 6036 39749 6104 39805
rect 6160 39749 6228 39805
rect 6284 39749 6352 39805
rect 6408 39749 6418 39805
rect 5970 39739 6418 39749
rect 8646 41045 9094 41055
rect 8646 40989 8656 41045
rect 8712 40989 8780 41045
rect 8836 40989 8904 41045
rect 8960 40989 9028 41045
rect 9084 40989 9094 41045
rect 8646 40921 9094 40989
rect 8646 40865 8656 40921
rect 8712 40865 8780 40921
rect 8836 40865 8904 40921
rect 8960 40865 9028 40921
rect 9084 40865 9094 40921
rect 8646 40797 9094 40865
rect 8646 40741 8656 40797
rect 8712 40741 8780 40797
rect 8836 40741 8904 40797
rect 8960 40741 9028 40797
rect 9084 40741 9094 40797
rect 8646 40673 9094 40741
rect 8646 40617 8656 40673
rect 8712 40617 8780 40673
rect 8836 40617 8904 40673
rect 8960 40617 9028 40673
rect 9084 40617 9094 40673
rect 8646 40549 9094 40617
rect 8646 40493 8656 40549
rect 8712 40493 8780 40549
rect 8836 40493 8904 40549
rect 8960 40493 9028 40549
rect 9084 40493 9094 40549
rect 8646 40425 9094 40493
rect 8646 40369 8656 40425
rect 8712 40369 8780 40425
rect 8836 40369 8904 40425
rect 8960 40369 9028 40425
rect 9084 40369 9094 40425
rect 8646 40301 9094 40369
rect 8646 40245 8656 40301
rect 8712 40245 8780 40301
rect 8836 40245 8904 40301
rect 8960 40245 9028 40301
rect 9084 40245 9094 40301
rect 8646 40177 9094 40245
rect 8646 40121 8656 40177
rect 8712 40121 8780 40177
rect 8836 40121 8904 40177
rect 8960 40121 9028 40177
rect 9084 40121 9094 40177
rect 8646 40053 9094 40121
rect 8646 39997 8656 40053
rect 8712 39997 8780 40053
rect 8836 39997 8904 40053
rect 8960 39997 9028 40053
rect 9084 39997 9094 40053
rect 8646 39929 9094 39997
rect 8646 39873 8656 39929
rect 8712 39873 8780 39929
rect 8836 39873 8904 39929
rect 8960 39873 9028 39929
rect 9084 39873 9094 39929
rect 8646 39805 9094 39873
rect 8646 39749 8656 39805
rect 8712 39749 8780 39805
rect 8836 39749 8904 39805
rect 8960 39749 9028 39805
rect 9084 39749 9094 39805
rect 8646 39739 9094 39749
rect 10918 41045 11366 41055
rect 10918 40989 10928 41045
rect 10984 40989 11052 41045
rect 11108 40989 11176 41045
rect 11232 40989 11300 41045
rect 11356 40989 11366 41045
rect 10918 40921 11366 40989
rect 10918 40865 10928 40921
rect 10984 40865 11052 40921
rect 11108 40865 11176 40921
rect 11232 40865 11300 40921
rect 11356 40865 11366 40921
rect 10918 40797 11366 40865
rect 10918 40741 10928 40797
rect 10984 40741 11052 40797
rect 11108 40741 11176 40797
rect 11232 40741 11300 40797
rect 11356 40741 11366 40797
rect 10918 40673 11366 40741
rect 10918 40617 10928 40673
rect 10984 40617 11052 40673
rect 11108 40617 11176 40673
rect 11232 40617 11300 40673
rect 11356 40617 11366 40673
rect 10918 40549 11366 40617
rect 10918 40493 10928 40549
rect 10984 40493 11052 40549
rect 11108 40493 11176 40549
rect 11232 40493 11300 40549
rect 11356 40493 11366 40549
rect 10918 40425 11366 40493
rect 10918 40369 10928 40425
rect 10984 40369 11052 40425
rect 11108 40369 11176 40425
rect 11232 40369 11300 40425
rect 11356 40369 11366 40425
rect 10918 40301 11366 40369
rect 10918 40245 10928 40301
rect 10984 40245 11052 40301
rect 11108 40245 11176 40301
rect 11232 40245 11300 40301
rect 11356 40245 11366 40301
rect 10918 40177 11366 40245
rect 10918 40121 10928 40177
rect 10984 40121 11052 40177
rect 11108 40121 11176 40177
rect 11232 40121 11300 40177
rect 11356 40121 11366 40177
rect 10918 40053 11366 40121
rect 10918 39997 10928 40053
rect 10984 39997 11052 40053
rect 11108 39997 11176 40053
rect 11232 39997 11300 40053
rect 11356 39997 11366 40053
rect 10918 39929 11366 39997
rect 10918 39873 10928 39929
rect 10984 39873 11052 39929
rect 11108 39873 11176 39929
rect 11232 39873 11300 39929
rect 11356 39873 11366 39929
rect 10918 39805 11366 39873
rect 10918 39749 10928 39805
rect 10984 39749 11052 39805
rect 11108 39749 11176 39805
rect 11232 39749 11300 39805
rect 11356 39749 11366 39805
rect 10918 39739 11366 39749
rect 12622 41045 13070 41055
rect 12622 40989 12632 41045
rect 12688 40989 12756 41045
rect 12812 40989 12880 41045
rect 12936 40989 13004 41045
rect 13060 40989 13070 41045
rect 12622 40921 13070 40989
rect 12622 40865 12632 40921
rect 12688 40865 12756 40921
rect 12812 40865 12880 40921
rect 12936 40865 13004 40921
rect 13060 40865 13070 40921
rect 12622 40797 13070 40865
rect 12622 40741 12632 40797
rect 12688 40741 12756 40797
rect 12812 40741 12880 40797
rect 12936 40741 13004 40797
rect 13060 40741 13070 40797
rect 12622 40673 13070 40741
rect 12622 40617 12632 40673
rect 12688 40617 12756 40673
rect 12812 40617 12880 40673
rect 12936 40617 13004 40673
rect 13060 40617 13070 40673
rect 12622 40549 13070 40617
rect 12622 40493 12632 40549
rect 12688 40493 12756 40549
rect 12812 40493 12880 40549
rect 12936 40493 13004 40549
rect 13060 40493 13070 40549
rect 12622 40425 13070 40493
rect 12622 40369 12632 40425
rect 12688 40369 12756 40425
rect 12812 40369 12880 40425
rect 12936 40369 13004 40425
rect 13060 40369 13070 40425
rect 12622 40301 13070 40369
rect 12622 40245 12632 40301
rect 12688 40245 12756 40301
rect 12812 40245 12880 40301
rect 12936 40245 13004 40301
rect 13060 40245 13070 40301
rect 12622 40177 13070 40245
rect 12622 40121 12632 40177
rect 12688 40121 12756 40177
rect 12812 40121 12880 40177
rect 12936 40121 13004 40177
rect 13060 40121 13070 40177
rect 12622 40053 13070 40121
rect 12622 39997 12632 40053
rect 12688 39997 12756 40053
rect 12812 39997 12880 40053
rect 12936 39997 13004 40053
rect 13060 39997 13070 40053
rect 12622 39929 13070 39997
rect 12622 39873 12632 39929
rect 12688 39873 12756 39929
rect 12812 39873 12880 39929
rect 12936 39873 13004 39929
rect 13060 39873 13070 39929
rect 12622 39805 13070 39873
rect 12622 39749 12632 39805
rect 12688 39749 12756 39805
rect 12812 39749 12880 39805
rect 12936 39749 13004 39805
rect 13060 39749 13070 39805
rect 12622 39739 13070 39749
rect 13758 41045 14206 41055
rect 13758 40989 13768 41045
rect 13824 40989 13892 41045
rect 13948 40989 14016 41045
rect 14072 40989 14140 41045
rect 14196 40989 14206 41045
rect 13758 40921 14206 40989
rect 13758 40865 13768 40921
rect 13824 40865 13892 40921
rect 13948 40865 14016 40921
rect 14072 40865 14140 40921
rect 14196 40865 14206 40921
rect 13758 40797 14206 40865
rect 13758 40741 13768 40797
rect 13824 40741 13892 40797
rect 13948 40741 14016 40797
rect 14072 40741 14140 40797
rect 14196 40741 14206 40797
rect 13758 40673 14206 40741
rect 13758 40617 13768 40673
rect 13824 40617 13892 40673
rect 13948 40617 14016 40673
rect 14072 40617 14140 40673
rect 14196 40617 14206 40673
rect 13758 40549 14206 40617
rect 13758 40493 13768 40549
rect 13824 40493 13892 40549
rect 13948 40493 14016 40549
rect 14072 40493 14140 40549
rect 14196 40493 14206 40549
rect 13758 40425 14206 40493
rect 13758 40369 13768 40425
rect 13824 40369 13892 40425
rect 13948 40369 14016 40425
rect 14072 40369 14140 40425
rect 14196 40369 14206 40425
rect 13758 40301 14206 40369
rect 13758 40245 13768 40301
rect 13824 40245 13892 40301
rect 13948 40245 14016 40301
rect 14072 40245 14140 40301
rect 14196 40245 14206 40301
rect 13758 40177 14206 40245
rect 13758 40121 13768 40177
rect 13824 40121 13892 40177
rect 13948 40121 14016 40177
rect 14072 40121 14140 40177
rect 14196 40121 14206 40177
rect 13758 40053 14206 40121
rect 13758 39997 13768 40053
rect 13824 39997 13892 40053
rect 13948 39997 14016 40053
rect 14072 39997 14140 40053
rect 14196 39997 14206 40053
rect 13758 39929 14206 39997
rect 13758 39873 13768 39929
rect 13824 39873 13892 39929
rect 13948 39873 14016 39929
rect 14072 39873 14140 39929
rect 14196 39873 14206 39929
rect 13758 39805 14206 39873
rect 13758 39749 13768 39805
rect 13824 39749 13892 39805
rect 13948 39749 14016 39805
rect 14072 39749 14140 39805
rect 14196 39749 14206 39805
rect 13758 39739 14206 39749
rect 828 39445 1028 39455
rect 828 39389 838 39445
rect 894 39389 962 39445
rect 1018 39389 1028 39445
rect 828 39321 1028 39389
rect 828 39265 838 39321
rect 894 39265 962 39321
rect 1018 39265 1028 39321
rect 828 39197 1028 39265
rect 828 39141 838 39197
rect 894 39141 962 39197
rect 1018 39141 1028 39197
rect 828 39073 1028 39141
rect 828 39017 838 39073
rect 894 39017 962 39073
rect 1018 39017 1028 39073
rect 828 38949 1028 39017
rect 828 38893 838 38949
rect 894 38893 962 38949
rect 1018 38893 1028 38949
rect 828 38825 1028 38893
rect 828 38769 838 38825
rect 894 38769 962 38825
rect 1018 38769 1028 38825
rect 828 38701 1028 38769
rect 828 38645 838 38701
rect 894 38645 962 38701
rect 1018 38645 1028 38701
rect 828 38577 1028 38645
rect 828 38521 838 38577
rect 894 38521 962 38577
rect 1018 38521 1028 38577
rect 828 38453 1028 38521
rect 828 38397 838 38453
rect 894 38397 962 38453
rect 1018 38397 1028 38453
rect 828 38329 1028 38397
rect 828 38273 838 38329
rect 894 38273 962 38329
rect 1018 38273 1028 38329
rect 828 38205 1028 38273
rect 828 38149 838 38205
rect 894 38149 962 38205
rect 1018 38149 1028 38205
rect 828 38139 1028 38149
rect 46 37873 122 37883
rect 46 36521 56 37873
rect 112 36521 122 37873
rect 14942 37873 15018 37883
rect 13160 37845 13360 37855
rect 13160 37789 13170 37845
rect 13226 37789 13294 37845
rect 13350 37789 13360 37845
rect 13160 37721 13360 37789
rect 13160 37665 13170 37721
rect 13226 37665 13294 37721
rect 13350 37665 13360 37721
rect 13160 37597 13360 37665
rect 13160 37541 13170 37597
rect 13226 37541 13294 37597
rect 13350 37541 13360 37597
rect 13160 37473 13360 37541
rect 13160 37417 13170 37473
rect 13226 37417 13294 37473
rect 13350 37417 13360 37473
rect 13160 37349 13360 37417
rect 13160 37293 13170 37349
rect 13226 37293 13294 37349
rect 13350 37293 13360 37349
rect 13160 37225 13360 37293
rect 13160 37169 13170 37225
rect 13226 37169 13294 37225
rect 13350 37169 13360 37225
rect 13160 37101 13360 37169
rect 13160 37045 13170 37101
rect 13226 37045 13294 37101
rect 13350 37045 13360 37101
rect 13160 36977 13360 37045
rect 13160 36921 13170 36977
rect 13226 36921 13294 36977
rect 13350 36921 13360 36977
rect 13160 36853 13360 36921
rect 13160 36797 13170 36853
rect 13226 36797 13294 36853
rect 13350 36797 13360 36853
rect 13160 36729 13360 36797
rect 13160 36673 13170 36729
rect 13226 36673 13294 36729
rect 13350 36673 13360 36729
rect 13160 36605 13360 36673
rect 13160 36549 13170 36605
rect 13226 36549 13294 36605
rect 13350 36549 13360 36605
rect 13160 36539 13360 36549
rect 46 36511 122 36521
rect 14942 36521 14952 37873
rect 15008 36521 15018 37873
rect 14942 36511 15018 36521
rect 290 36251 738 36261
rect 290 36195 300 36251
rect 356 36195 424 36251
rect 480 36195 548 36251
rect 604 36195 672 36251
rect 728 36195 738 36251
rect 290 36127 738 36195
rect 290 36071 300 36127
rect 356 36071 424 36127
rect 480 36071 548 36127
rect 604 36071 672 36127
rect 728 36071 738 36127
rect 290 36003 738 36071
rect 290 35947 300 36003
rect 356 35947 424 36003
rect 480 35947 548 36003
rect 604 35947 672 36003
rect 728 35947 738 36003
rect 290 35879 738 35947
rect 290 35823 300 35879
rect 356 35823 424 35879
rect 480 35823 548 35879
rect 604 35823 672 35879
rect 728 35823 738 35879
rect 290 35755 738 35823
rect 290 35699 300 35755
rect 356 35699 424 35755
rect 480 35699 548 35755
rect 604 35699 672 35755
rect 728 35699 738 35755
rect 290 35631 738 35699
rect 290 35575 300 35631
rect 356 35575 424 35631
rect 480 35575 548 35631
rect 604 35575 672 35631
rect 728 35575 738 35631
rect 290 35507 738 35575
rect 290 35451 300 35507
rect 356 35451 424 35507
rect 480 35451 548 35507
rect 604 35451 672 35507
rect 728 35451 738 35507
rect 290 35383 738 35451
rect 290 35327 300 35383
rect 356 35327 424 35383
rect 480 35327 548 35383
rect 604 35327 672 35383
rect 728 35327 738 35383
rect 290 35259 738 35327
rect 290 35203 300 35259
rect 356 35203 424 35259
rect 480 35203 548 35259
rect 604 35203 672 35259
rect 728 35203 738 35259
rect 290 35135 738 35203
rect 290 35079 300 35135
rect 356 35079 424 35135
rect 480 35079 548 35135
rect 604 35079 672 35135
rect 728 35079 738 35135
rect 290 35011 738 35079
rect 290 34955 300 35011
rect 356 34955 424 35011
rect 480 34955 548 35011
rect 604 34955 672 35011
rect 728 34955 738 35011
rect 290 34887 738 34955
rect 290 34831 300 34887
rect 356 34831 424 34887
rect 480 34831 548 34887
rect 604 34831 672 34887
rect 728 34831 738 34887
rect 290 34763 738 34831
rect 290 34707 300 34763
rect 356 34707 424 34763
rect 480 34707 548 34763
rect 604 34707 672 34763
rect 728 34707 738 34763
rect 290 34639 738 34707
rect 290 34583 300 34639
rect 356 34583 424 34639
rect 480 34583 548 34639
rect 604 34583 672 34639
rect 728 34583 738 34639
rect 290 34515 738 34583
rect 290 34459 300 34515
rect 356 34459 424 34515
rect 480 34459 548 34515
rect 604 34459 672 34515
rect 728 34459 738 34515
rect 290 34391 738 34459
rect 290 34335 300 34391
rect 356 34335 424 34391
rect 480 34335 548 34391
rect 604 34335 672 34391
rect 728 34335 738 34391
rect 290 34267 738 34335
rect 290 34211 300 34267
rect 356 34211 424 34267
rect 480 34211 548 34267
rect 604 34211 672 34267
rect 728 34211 738 34267
rect 290 34143 738 34211
rect 290 34087 300 34143
rect 356 34087 424 34143
rect 480 34087 548 34143
rect 604 34087 672 34143
rect 728 34087 738 34143
rect 290 34019 738 34087
rect 290 33963 300 34019
rect 356 33963 424 34019
rect 480 33963 548 34019
rect 604 33963 672 34019
rect 728 33963 738 34019
rect 290 33895 738 33963
rect 290 33839 300 33895
rect 356 33839 424 33895
rect 480 33839 548 33895
rect 604 33839 672 33895
rect 728 33839 738 33895
rect 290 33771 738 33839
rect 290 33715 300 33771
rect 356 33715 424 33771
rect 480 33715 548 33771
rect 604 33715 672 33771
rect 728 33715 738 33771
rect 290 33647 738 33715
rect 290 33591 300 33647
rect 356 33591 424 33647
rect 480 33591 548 33647
rect 604 33591 672 33647
rect 728 33591 738 33647
rect 290 33523 738 33591
rect 290 33467 300 33523
rect 356 33467 424 33523
rect 480 33467 548 33523
rect 604 33467 672 33523
rect 728 33467 738 33523
rect 290 33399 738 33467
rect 290 33343 300 33399
rect 356 33343 424 33399
rect 480 33343 548 33399
rect 604 33343 672 33399
rect 728 33343 738 33399
rect 290 33333 738 33343
rect 1426 36251 1874 36261
rect 1426 36195 1436 36251
rect 1492 36195 1560 36251
rect 1616 36195 1684 36251
rect 1740 36195 1808 36251
rect 1864 36195 1874 36251
rect 1426 36127 1874 36195
rect 1426 36071 1436 36127
rect 1492 36071 1560 36127
rect 1616 36071 1684 36127
rect 1740 36071 1808 36127
rect 1864 36071 1874 36127
rect 1426 36003 1874 36071
rect 1426 35947 1436 36003
rect 1492 35947 1560 36003
rect 1616 35947 1684 36003
rect 1740 35947 1808 36003
rect 1864 35947 1874 36003
rect 1426 35879 1874 35947
rect 1426 35823 1436 35879
rect 1492 35823 1560 35879
rect 1616 35823 1684 35879
rect 1740 35823 1808 35879
rect 1864 35823 1874 35879
rect 1426 35755 1874 35823
rect 1426 35699 1436 35755
rect 1492 35699 1560 35755
rect 1616 35699 1684 35755
rect 1740 35699 1808 35755
rect 1864 35699 1874 35755
rect 1426 35631 1874 35699
rect 1426 35575 1436 35631
rect 1492 35575 1560 35631
rect 1616 35575 1684 35631
rect 1740 35575 1808 35631
rect 1864 35575 1874 35631
rect 1426 35507 1874 35575
rect 1426 35451 1436 35507
rect 1492 35451 1560 35507
rect 1616 35451 1684 35507
rect 1740 35451 1808 35507
rect 1864 35451 1874 35507
rect 1426 35383 1874 35451
rect 1426 35327 1436 35383
rect 1492 35327 1560 35383
rect 1616 35327 1684 35383
rect 1740 35327 1808 35383
rect 1864 35327 1874 35383
rect 1426 35259 1874 35327
rect 1426 35203 1436 35259
rect 1492 35203 1560 35259
rect 1616 35203 1684 35259
rect 1740 35203 1808 35259
rect 1864 35203 1874 35259
rect 1426 35135 1874 35203
rect 1426 35079 1436 35135
rect 1492 35079 1560 35135
rect 1616 35079 1684 35135
rect 1740 35079 1808 35135
rect 1864 35079 1874 35135
rect 1426 35011 1874 35079
rect 1426 34955 1436 35011
rect 1492 34955 1560 35011
rect 1616 34955 1684 35011
rect 1740 34955 1808 35011
rect 1864 34955 1874 35011
rect 1426 34887 1874 34955
rect 1426 34831 1436 34887
rect 1492 34831 1560 34887
rect 1616 34831 1684 34887
rect 1740 34831 1808 34887
rect 1864 34831 1874 34887
rect 1426 34763 1874 34831
rect 1426 34707 1436 34763
rect 1492 34707 1560 34763
rect 1616 34707 1684 34763
rect 1740 34707 1808 34763
rect 1864 34707 1874 34763
rect 1426 34639 1874 34707
rect 1426 34583 1436 34639
rect 1492 34583 1560 34639
rect 1616 34583 1684 34639
rect 1740 34583 1808 34639
rect 1864 34583 1874 34639
rect 1426 34515 1874 34583
rect 1426 34459 1436 34515
rect 1492 34459 1560 34515
rect 1616 34459 1684 34515
rect 1740 34459 1808 34515
rect 1864 34459 1874 34515
rect 1426 34391 1874 34459
rect 1426 34335 1436 34391
rect 1492 34335 1560 34391
rect 1616 34335 1684 34391
rect 1740 34335 1808 34391
rect 1864 34335 1874 34391
rect 1426 34267 1874 34335
rect 1426 34211 1436 34267
rect 1492 34211 1560 34267
rect 1616 34211 1684 34267
rect 1740 34211 1808 34267
rect 1864 34211 1874 34267
rect 1426 34143 1874 34211
rect 1426 34087 1436 34143
rect 1492 34087 1560 34143
rect 1616 34087 1684 34143
rect 1740 34087 1808 34143
rect 1864 34087 1874 34143
rect 1426 34019 1874 34087
rect 1426 33963 1436 34019
rect 1492 33963 1560 34019
rect 1616 33963 1684 34019
rect 1740 33963 1808 34019
rect 1864 33963 1874 34019
rect 1426 33895 1874 33963
rect 1426 33839 1436 33895
rect 1492 33839 1560 33895
rect 1616 33839 1684 33895
rect 1740 33839 1808 33895
rect 1864 33839 1874 33895
rect 1426 33771 1874 33839
rect 1426 33715 1436 33771
rect 1492 33715 1560 33771
rect 1616 33715 1684 33771
rect 1740 33715 1808 33771
rect 1864 33715 1874 33771
rect 1426 33647 1874 33715
rect 1426 33591 1436 33647
rect 1492 33591 1560 33647
rect 1616 33591 1684 33647
rect 1740 33591 1808 33647
rect 1864 33591 1874 33647
rect 1426 33523 1874 33591
rect 1426 33467 1436 33523
rect 1492 33467 1560 33523
rect 1616 33467 1684 33523
rect 1740 33467 1808 33523
rect 1864 33467 1874 33523
rect 1426 33399 1874 33467
rect 1426 33343 1436 33399
rect 1492 33343 1560 33399
rect 1616 33343 1684 33399
rect 1740 33343 1808 33399
rect 1864 33343 1874 33399
rect 1426 33333 1874 33343
rect 2562 36251 3010 36261
rect 2562 36195 2572 36251
rect 2628 36195 2696 36251
rect 2752 36195 2820 36251
rect 2876 36195 2944 36251
rect 3000 36195 3010 36251
rect 2562 36127 3010 36195
rect 2562 36071 2572 36127
rect 2628 36071 2696 36127
rect 2752 36071 2820 36127
rect 2876 36071 2944 36127
rect 3000 36071 3010 36127
rect 2562 36003 3010 36071
rect 2562 35947 2572 36003
rect 2628 35947 2696 36003
rect 2752 35947 2820 36003
rect 2876 35947 2944 36003
rect 3000 35947 3010 36003
rect 2562 35879 3010 35947
rect 2562 35823 2572 35879
rect 2628 35823 2696 35879
rect 2752 35823 2820 35879
rect 2876 35823 2944 35879
rect 3000 35823 3010 35879
rect 2562 35755 3010 35823
rect 2562 35699 2572 35755
rect 2628 35699 2696 35755
rect 2752 35699 2820 35755
rect 2876 35699 2944 35755
rect 3000 35699 3010 35755
rect 2562 35631 3010 35699
rect 2562 35575 2572 35631
rect 2628 35575 2696 35631
rect 2752 35575 2820 35631
rect 2876 35575 2944 35631
rect 3000 35575 3010 35631
rect 2562 35507 3010 35575
rect 2562 35451 2572 35507
rect 2628 35451 2696 35507
rect 2752 35451 2820 35507
rect 2876 35451 2944 35507
rect 3000 35451 3010 35507
rect 2562 35383 3010 35451
rect 2562 35327 2572 35383
rect 2628 35327 2696 35383
rect 2752 35327 2820 35383
rect 2876 35327 2944 35383
rect 3000 35327 3010 35383
rect 2562 35259 3010 35327
rect 2562 35203 2572 35259
rect 2628 35203 2696 35259
rect 2752 35203 2820 35259
rect 2876 35203 2944 35259
rect 3000 35203 3010 35259
rect 2562 35135 3010 35203
rect 2562 35079 2572 35135
rect 2628 35079 2696 35135
rect 2752 35079 2820 35135
rect 2876 35079 2944 35135
rect 3000 35079 3010 35135
rect 2562 35011 3010 35079
rect 2562 34955 2572 35011
rect 2628 34955 2696 35011
rect 2752 34955 2820 35011
rect 2876 34955 2944 35011
rect 3000 34955 3010 35011
rect 2562 34887 3010 34955
rect 2562 34831 2572 34887
rect 2628 34831 2696 34887
rect 2752 34831 2820 34887
rect 2876 34831 2944 34887
rect 3000 34831 3010 34887
rect 2562 34763 3010 34831
rect 2562 34707 2572 34763
rect 2628 34707 2696 34763
rect 2752 34707 2820 34763
rect 2876 34707 2944 34763
rect 3000 34707 3010 34763
rect 2562 34639 3010 34707
rect 2562 34583 2572 34639
rect 2628 34583 2696 34639
rect 2752 34583 2820 34639
rect 2876 34583 2944 34639
rect 3000 34583 3010 34639
rect 2562 34515 3010 34583
rect 2562 34459 2572 34515
rect 2628 34459 2696 34515
rect 2752 34459 2820 34515
rect 2876 34459 2944 34515
rect 3000 34459 3010 34515
rect 2562 34391 3010 34459
rect 2562 34335 2572 34391
rect 2628 34335 2696 34391
rect 2752 34335 2820 34391
rect 2876 34335 2944 34391
rect 3000 34335 3010 34391
rect 2562 34267 3010 34335
rect 2562 34211 2572 34267
rect 2628 34211 2696 34267
rect 2752 34211 2820 34267
rect 2876 34211 2944 34267
rect 3000 34211 3010 34267
rect 2562 34143 3010 34211
rect 2562 34087 2572 34143
rect 2628 34087 2696 34143
rect 2752 34087 2820 34143
rect 2876 34087 2944 34143
rect 3000 34087 3010 34143
rect 2562 34019 3010 34087
rect 2562 33963 2572 34019
rect 2628 33963 2696 34019
rect 2752 33963 2820 34019
rect 2876 33963 2944 34019
rect 3000 33963 3010 34019
rect 2562 33895 3010 33963
rect 2562 33839 2572 33895
rect 2628 33839 2696 33895
rect 2752 33839 2820 33895
rect 2876 33839 2944 33895
rect 3000 33839 3010 33895
rect 2562 33771 3010 33839
rect 2562 33715 2572 33771
rect 2628 33715 2696 33771
rect 2752 33715 2820 33771
rect 2876 33715 2944 33771
rect 3000 33715 3010 33771
rect 2562 33647 3010 33715
rect 2562 33591 2572 33647
rect 2628 33591 2696 33647
rect 2752 33591 2820 33647
rect 2876 33591 2944 33647
rect 3000 33591 3010 33647
rect 2562 33523 3010 33591
rect 2562 33467 2572 33523
rect 2628 33467 2696 33523
rect 2752 33467 2820 33523
rect 2876 33467 2944 33523
rect 3000 33467 3010 33523
rect 2562 33399 3010 33467
rect 2562 33343 2572 33399
rect 2628 33343 2696 33399
rect 2752 33343 2820 33399
rect 2876 33343 2944 33399
rect 3000 33343 3010 33399
rect 2562 33333 3010 33343
rect 4834 36251 5282 36261
rect 4834 36195 4844 36251
rect 4900 36195 4968 36251
rect 5024 36195 5092 36251
rect 5148 36195 5216 36251
rect 5272 36195 5282 36251
rect 4834 36127 5282 36195
rect 4834 36071 4844 36127
rect 4900 36071 4968 36127
rect 5024 36071 5092 36127
rect 5148 36071 5216 36127
rect 5272 36071 5282 36127
rect 4834 36003 5282 36071
rect 4834 35947 4844 36003
rect 4900 35947 4968 36003
rect 5024 35947 5092 36003
rect 5148 35947 5216 36003
rect 5272 35947 5282 36003
rect 4834 35879 5282 35947
rect 4834 35823 4844 35879
rect 4900 35823 4968 35879
rect 5024 35823 5092 35879
rect 5148 35823 5216 35879
rect 5272 35823 5282 35879
rect 4834 35755 5282 35823
rect 4834 35699 4844 35755
rect 4900 35699 4968 35755
rect 5024 35699 5092 35755
rect 5148 35699 5216 35755
rect 5272 35699 5282 35755
rect 4834 35631 5282 35699
rect 4834 35575 4844 35631
rect 4900 35575 4968 35631
rect 5024 35575 5092 35631
rect 5148 35575 5216 35631
rect 5272 35575 5282 35631
rect 4834 35507 5282 35575
rect 4834 35451 4844 35507
rect 4900 35451 4968 35507
rect 5024 35451 5092 35507
rect 5148 35451 5216 35507
rect 5272 35451 5282 35507
rect 4834 35383 5282 35451
rect 4834 35327 4844 35383
rect 4900 35327 4968 35383
rect 5024 35327 5092 35383
rect 5148 35327 5216 35383
rect 5272 35327 5282 35383
rect 4834 35259 5282 35327
rect 4834 35203 4844 35259
rect 4900 35203 4968 35259
rect 5024 35203 5092 35259
rect 5148 35203 5216 35259
rect 5272 35203 5282 35259
rect 4834 35135 5282 35203
rect 4834 35079 4844 35135
rect 4900 35079 4968 35135
rect 5024 35079 5092 35135
rect 5148 35079 5216 35135
rect 5272 35079 5282 35135
rect 4834 35011 5282 35079
rect 4834 34955 4844 35011
rect 4900 34955 4968 35011
rect 5024 34955 5092 35011
rect 5148 34955 5216 35011
rect 5272 34955 5282 35011
rect 4834 34887 5282 34955
rect 4834 34831 4844 34887
rect 4900 34831 4968 34887
rect 5024 34831 5092 34887
rect 5148 34831 5216 34887
rect 5272 34831 5282 34887
rect 4834 34763 5282 34831
rect 4834 34707 4844 34763
rect 4900 34707 4968 34763
rect 5024 34707 5092 34763
rect 5148 34707 5216 34763
rect 5272 34707 5282 34763
rect 4834 34639 5282 34707
rect 4834 34583 4844 34639
rect 4900 34583 4968 34639
rect 5024 34583 5092 34639
rect 5148 34583 5216 34639
rect 5272 34583 5282 34639
rect 4834 34515 5282 34583
rect 4834 34459 4844 34515
rect 4900 34459 4968 34515
rect 5024 34459 5092 34515
rect 5148 34459 5216 34515
rect 5272 34459 5282 34515
rect 4834 34391 5282 34459
rect 4834 34335 4844 34391
rect 4900 34335 4968 34391
rect 5024 34335 5092 34391
rect 5148 34335 5216 34391
rect 5272 34335 5282 34391
rect 4834 34267 5282 34335
rect 4834 34211 4844 34267
rect 4900 34211 4968 34267
rect 5024 34211 5092 34267
rect 5148 34211 5216 34267
rect 5272 34211 5282 34267
rect 4834 34143 5282 34211
rect 4834 34087 4844 34143
rect 4900 34087 4968 34143
rect 5024 34087 5092 34143
rect 5148 34087 5216 34143
rect 5272 34087 5282 34143
rect 4834 34019 5282 34087
rect 4834 33963 4844 34019
rect 4900 33963 4968 34019
rect 5024 33963 5092 34019
rect 5148 33963 5216 34019
rect 5272 33963 5282 34019
rect 4834 33895 5282 33963
rect 4834 33839 4844 33895
rect 4900 33839 4968 33895
rect 5024 33839 5092 33895
rect 5148 33839 5216 33895
rect 5272 33839 5282 33895
rect 4834 33771 5282 33839
rect 4834 33715 4844 33771
rect 4900 33715 4968 33771
rect 5024 33715 5092 33771
rect 5148 33715 5216 33771
rect 5272 33715 5282 33771
rect 4834 33647 5282 33715
rect 4834 33591 4844 33647
rect 4900 33591 4968 33647
rect 5024 33591 5092 33647
rect 5148 33591 5216 33647
rect 5272 33591 5282 33647
rect 4834 33523 5282 33591
rect 4834 33467 4844 33523
rect 4900 33467 4968 33523
rect 5024 33467 5092 33523
rect 5148 33467 5216 33523
rect 5272 33467 5282 33523
rect 4834 33399 5282 33467
rect 4834 33343 4844 33399
rect 4900 33343 4968 33399
rect 5024 33343 5092 33399
rect 5148 33343 5216 33399
rect 5272 33343 5282 33399
rect 4834 33333 5282 33343
rect 7127 36251 7451 36261
rect 7127 36195 7137 36251
rect 7193 36195 7261 36251
rect 7317 36195 7385 36251
rect 7441 36195 7451 36251
rect 7127 36127 7451 36195
rect 7127 36071 7137 36127
rect 7193 36071 7261 36127
rect 7317 36071 7385 36127
rect 7441 36071 7451 36127
rect 7127 36003 7451 36071
rect 7127 35947 7137 36003
rect 7193 35947 7261 36003
rect 7317 35947 7385 36003
rect 7441 35947 7451 36003
rect 7127 35879 7451 35947
rect 7127 35823 7137 35879
rect 7193 35823 7261 35879
rect 7317 35823 7385 35879
rect 7441 35823 7451 35879
rect 7127 35755 7451 35823
rect 7127 35699 7137 35755
rect 7193 35699 7261 35755
rect 7317 35699 7385 35755
rect 7441 35699 7451 35755
rect 7127 35631 7451 35699
rect 7127 35575 7137 35631
rect 7193 35575 7261 35631
rect 7317 35575 7385 35631
rect 7441 35575 7451 35631
rect 7127 35507 7451 35575
rect 7127 35451 7137 35507
rect 7193 35451 7261 35507
rect 7317 35451 7385 35507
rect 7441 35451 7451 35507
rect 7127 35383 7451 35451
rect 7127 35327 7137 35383
rect 7193 35327 7261 35383
rect 7317 35327 7385 35383
rect 7441 35327 7451 35383
rect 7127 35259 7451 35327
rect 7127 35203 7137 35259
rect 7193 35203 7261 35259
rect 7317 35203 7385 35259
rect 7441 35203 7451 35259
rect 7127 35135 7451 35203
rect 7127 35079 7137 35135
rect 7193 35079 7261 35135
rect 7317 35079 7385 35135
rect 7441 35079 7451 35135
rect 7127 35011 7451 35079
rect 7127 34955 7137 35011
rect 7193 34955 7261 35011
rect 7317 34955 7385 35011
rect 7441 34955 7451 35011
rect 7127 34887 7451 34955
rect 7127 34831 7137 34887
rect 7193 34831 7261 34887
rect 7317 34831 7385 34887
rect 7441 34831 7451 34887
rect 7127 34763 7451 34831
rect 7127 34707 7137 34763
rect 7193 34707 7261 34763
rect 7317 34707 7385 34763
rect 7441 34707 7451 34763
rect 7127 34639 7451 34707
rect 7127 34583 7137 34639
rect 7193 34583 7261 34639
rect 7317 34583 7385 34639
rect 7441 34583 7451 34639
rect 7127 34515 7451 34583
rect 7127 34459 7137 34515
rect 7193 34459 7261 34515
rect 7317 34459 7385 34515
rect 7441 34459 7451 34515
rect 7127 34391 7451 34459
rect 7127 34335 7137 34391
rect 7193 34335 7261 34391
rect 7317 34335 7385 34391
rect 7441 34335 7451 34391
rect 7127 34267 7451 34335
rect 7127 34211 7137 34267
rect 7193 34211 7261 34267
rect 7317 34211 7385 34267
rect 7441 34211 7451 34267
rect 7127 34143 7451 34211
rect 7127 34087 7137 34143
rect 7193 34087 7261 34143
rect 7317 34087 7385 34143
rect 7441 34087 7451 34143
rect 7127 34019 7451 34087
rect 7127 33963 7137 34019
rect 7193 33963 7261 34019
rect 7317 33963 7385 34019
rect 7441 33963 7451 34019
rect 7127 33895 7451 33963
rect 7127 33839 7137 33895
rect 7193 33839 7261 33895
rect 7317 33839 7385 33895
rect 7441 33839 7451 33895
rect 7127 33771 7451 33839
rect 7127 33715 7137 33771
rect 7193 33715 7261 33771
rect 7317 33715 7385 33771
rect 7441 33715 7451 33771
rect 7127 33647 7451 33715
rect 7127 33591 7137 33647
rect 7193 33591 7261 33647
rect 7317 33591 7385 33647
rect 7441 33591 7451 33647
rect 7127 33523 7451 33591
rect 7127 33467 7137 33523
rect 7193 33467 7261 33523
rect 7317 33467 7385 33523
rect 7441 33467 7451 33523
rect 7127 33399 7451 33467
rect 7127 33343 7137 33399
rect 7193 33343 7261 33399
rect 7317 33343 7385 33399
rect 7441 33343 7451 33399
rect 7127 33333 7451 33343
rect 7613 36251 7937 36261
rect 7613 36195 7623 36251
rect 7679 36195 7747 36251
rect 7803 36195 7871 36251
rect 7927 36195 7937 36251
rect 7613 36127 7937 36195
rect 7613 36071 7623 36127
rect 7679 36071 7747 36127
rect 7803 36071 7871 36127
rect 7927 36071 7937 36127
rect 7613 36003 7937 36071
rect 7613 35947 7623 36003
rect 7679 35947 7747 36003
rect 7803 35947 7871 36003
rect 7927 35947 7937 36003
rect 7613 35879 7937 35947
rect 7613 35823 7623 35879
rect 7679 35823 7747 35879
rect 7803 35823 7871 35879
rect 7927 35823 7937 35879
rect 7613 35755 7937 35823
rect 7613 35699 7623 35755
rect 7679 35699 7747 35755
rect 7803 35699 7871 35755
rect 7927 35699 7937 35755
rect 7613 35631 7937 35699
rect 7613 35575 7623 35631
rect 7679 35575 7747 35631
rect 7803 35575 7871 35631
rect 7927 35575 7937 35631
rect 7613 35507 7937 35575
rect 7613 35451 7623 35507
rect 7679 35451 7747 35507
rect 7803 35451 7871 35507
rect 7927 35451 7937 35507
rect 7613 35383 7937 35451
rect 7613 35327 7623 35383
rect 7679 35327 7747 35383
rect 7803 35327 7871 35383
rect 7927 35327 7937 35383
rect 7613 35259 7937 35327
rect 7613 35203 7623 35259
rect 7679 35203 7747 35259
rect 7803 35203 7871 35259
rect 7927 35203 7937 35259
rect 7613 35135 7937 35203
rect 7613 35079 7623 35135
rect 7679 35079 7747 35135
rect 7803 35079 7871 35135
rect 7927 35079 7937 35135
rect 7613 35011 7937 35079
rect 7613 34955 7623 35011
rect 7679 34955 7747 35011
rect 7803 34955 7871 35011
rect 7927 34955 7937 35011
rect 7613 34887 7937 34955
rect 7613 34831 7623 34887
rect 7679 34831 7747 34887
rect 7803 34831 7871 34887
rect 7927 34831 7937 34887
rect 7613 34763 7937 34831
rect 7613 34707 7623 34763
rect 7679 34707 7747 34763
rect 7803 34707 7871 34763
rect 7927 34707 7937 34763
rect 7613 34639 7937 34707
rect 7613 34583 7623 34639
rect 7679 34583 7747 34639
rect 7803 34583 7871 34639
rect 7927 34583 7937 34639
rect 7613 34515 7937 34583
rect 7613 34459 7623 34515
rect 7679 34459 7747 34515
rect 7803 34459 7871 34515
rect 7927 34459 7937 34515
rect 7613 34391 7937 34459
rect 7613 34335 7623 34391
rect 7679 34335 7747 34391
rect 7803 34335 7871 34391
rect 7927 34335 7937 34391
rect 7613 34267 7937 34335
rect 7613 34211 7623 34267
rect 7679 34211 7747 34267
rect 7803 34211 7871 34267
rect 7927 34211 7937 34267
rect 7613 34143 7937 34211
rect 7613 34087 7623 34143
rect 7679 34087 7747 34143
rect 7803 34087 7871 34143
rect 7927 34087 7937 34143
rect 7613 34019 7937 34087
rect 7613 33963 7623 34019
rect 7679 33963 7747 34019
rect 7803 33963 7871 34019
rect 7927 33963 7937 34019
rect 7613 33895 7937 33963
rect 7613 33839 7623 33895
rect 7679 33839 7747 33895
rect 7803 33839 7871 33895
rect 7927 33839 7937 33895
rect 7613 33771 7937 33839
rect 7613 33715 7623 33771
rect 7679 33715 7747 33771
rect 7803 33715 7871 33771
rect 7927 33715 7937 33771
rect 7613 33647 7937 33715
rect 7613 33591 7623 33647
rect 7679 33591 7747 33647
rect 7803 33591 7871 33647
rect 7927 33591 7937 33647
rect 7613 33523 7937 33591
rect 7613 33467 7623 33523
rect 7679 33467 7747 33523
rect 7803 33467 7871 33523
rect 7927 33467 7937 33523
rect 7613 33399 7937 33467
rect 7613 33343 7623 33399
rect 7679 33343 7747 33399
rect 7803 33343 7871 33399
rect 7927 33343 7937 33399
rect 7613 33333 7937 33343
rect 9782 36251 10230 36261
rect 9782 36195 9792 36251
rect 9848 36195 9916 36251
rect 9972 36195 10040 36251
rect 10096 36195 10164 36251
rect 10220 36195 10230 36251
rect 9782 36127 10230 36195
rect 9782 36071 9792 36127
rect 9848 36071 9916 36127
rect 9972 36071 10040 36127
rect 10096 36071 10164 36127
rect 10220 36071 10230 36127
rect 9782 36003 10230 36071
rect 9782 35947 9792 36003
rect 9848 35947 9916 36003
rect 9972 35947 10040 36003
rect 10096 35947 10164 36003
rect 10220 35947 10230 36003
rect 9782 35879 10230 35947
rect 9782 35823 9792 35879
rect 9848 35823 9916 35879
rect 9972 35823 10040 35879
rect 10096 35823 10164 35879
rect 10220 35823 10230 35879
rect 9782 35755 10230 35823
rect 9782 35699 9792 35755
rect 9848 35699 9916 35755
rect 9972 35699 10040 35755
rect 10096 35699 10164 35755
rect 10220 35699 10230 35755
rect 9782 35631 10230 35699
rect 9782 35575 9792 35631
rect 9848 35575 9916 35631
rect 9972 35575 10040 35631
rect 10096 35575 10164 35631
rect 10220 35575 10230 35631
rect 9782 35507 10230 35575
rect 9782 35451 9792 35507
rect 9848 35451 9916 35507
rect 9972 35451 10040 35507
rect 10096 35451 10164 35507
rect 10220 35451 10230 35507
rect 9782 35383 10230 35451
rect 9782 35327 9792 35383
rect 9848 35327 9916 35383
rect 9972 35327 10040 35383
rect 10096 35327 10164 35383
rect 10220 35327 10230 35383
rect 9782 35259 10230 35327
rect 9782 35203 9792 35259
rect 9848 35203 9916 35259
rect 9972 35203 10040 35259
rect 10096 35203 10164 35259
rect 10220 35203 10230 35259
rect 9782 35135 10230 35203
rect 9782 35079 9792 35135
rect 9848 35079 9916 35135
rect 9972 35079 10040 35135
rect 10096 35079 10164 35135
rect 10220 35079 10230 35135
rect 9782 35011 10230 35079
rect 9782 34955 9792 35011
rect 9848 34955 9916 35011
rect 9972 34955 10040 35011
rect 10096 34955 10164 35011
rect 10220 34955 10230 35011
rect 9782 34887 10230 34955
rect 9782 34831 9792 34887
rect 9848 34831 9916 34887
rect 9972 34831 10040 34887
rect 10096 34831 10164 34887
rect 10220 34831 10230 34887
rect 9782 34763 10230 34831
rect 9782 34707 9792 34763
rect 9848 34707 9916 34763
rect 9972 34707 10040 34763
rect 10096 34707 10164 34763
rect 10220 34707 10230 34763
rect 9782 34639 10230 34707
rect 9782 34583 9792 34639
rect 9848 34583 9916 34639
rect 9972 34583 10040 34639
rect 10096 34583 10164 34639
rect 10220 34583 10230 34639
rect 9782 34515 10230 34583
rect 9782 34459 9792 34515
rect 9848 34459 9916 34515
rect 9972 34459 10040 34515
rect 10096 34459 10164 34515
rect 10220 34459 10230 34515
rect 9782 34391 10230 34459
rect 9782 34335 9792 34391
rect 9848 34335 9916 34391
rect 9972 34335 10040 34391
rect 10096 34335 10164 34391
rect 10220 34335 10230 34391
rect 9782 34267 10230 34335
rect 9782 34211 9792 34267
rect 9848 34211 9916 34267
rect 9972 34211 10040 34267
rect 10096 34211 10164 34267
rect 10220 34211 10230 34267
rect 9782 34143 10230 34211
rect 9782 34087 9792 34143
rect 9848 34087 9916 34143
rect 9972 34087 10040 34143
rect 10096 34087 10164 34143
rect 10220 34087 10230 34143
rect 9782 34019 10230 34087
rect 9782 33963 9792 34019
rect 9848 33963 9916 34019
rect 9972 33963 10040 34019
rect 10096 33963 10164 34019
rect 10220 33963 10230 34019
rect 9782 33895 10230 33963
rect 9782 33839 9792 33895
rect 9848 33839 9916 33895
rect 9972 33839 10040 33895
rect 10096 33839 10164 33895
rect 10220 33839 10230 33895
rect 9782 33771 10230 33839
rect 9782 33715 9792 33771
rect 9848 33715 9916 33771
rect 9972 33715 10040 33771
rect 10096 33715 10164 33771
rect 10220 33715 10230 33771
rect 9782 33647 10230 33715
rect 9782 33591 9792 33647
rect 9848 33591 9916 33647
rect 9972 33591 10040 33647
rect 10096 33591 10164 33647
rect 10220 33591 10230 33647
rect 9782 33523 10230 33591
rect 9782 33467 9792 33523
rect 9848 33467 9916 33523
rect 9972 33467 10040 33523
rect 10096 33467 10164 33523
rect 10220 33467 10230 33523
rect 9782 33399 10230 33467
rect 9782 33343 9792 33399
rect 9848 33343 9916 33399
rect 9972 33343 10040 33399
rect 10096 33343 10164 33399
rect 10220 33343 10230 33399
rect 9782 33333 10230 33343
rect 12054 36251 12502 36261
rect 12054 36195 12064 36251
rect 12120 36195 12188 36251
rect 12244 36195 12312 36251
rect 12368 36195 12436 36251
rect 12492 36195 12502 36251
rect 12054 36127 12502 36195
rect 12054 36071 12064 36127
rect 12120 36071 12188 36127
rect 12244 36071 12312 36127
rect 12368 36071 12436 36127
rect 12492 36071 12502 36127
rect 12054 36003 12502 36071
rect 12054 35947 12064 36003
rect 12120 35947 12188 36003
rect 12244 35947 12312 36003
rect 12368 35947 12436 36003
rect 12492 35947 12502 36003
rect 12054 35879 12502 35947
rect 12054 35823 12064 35879
rect 12120 35823 12188 35879
rect 12244 35823 12312 35879
rect 12368 35823 12436 35879
rect 12492 35823 12502 35879
rect 12054 35755 12502 35823
rect 12054 35699 12064 35755
rect 12120 35699 12188 35755
rect 12244 35699 12312 35755
rect 12368 35699 12436 35755
rect 12492 35699 12502 35755
rect 12054 35631 12502 35699
rect 12054 35575 12064 35631
rect 12120 35575 12188 35631
rect 12244 35575 12312 35631
rect 12368 35575 12436 35631
rect 12492 35575 12502 35631
rect 12054 35507 12502 35575
rect 12054 35451 12064 35507
rect 12120 35451 12188 35507
rect 12244 35451 12312 35507
rect 12368 35451 12436 35507
rect 12492 35451 12502 35507
rect 12054 35383 12502 35451
rect 12054 35327 12064 35383
rect 12120 35327 12188 35383
rect 12244 35327 12312 35383
rect 12368 35327 12436 35383
rect 12492 35327 12502 35383
rect 12054 35259 12502 35327
rect 12054 35203 12064 35259
rect 12120 35203 12188 35259
rect 12244 35203 12312 35259
rect 12368 35203 12436 35259
rect 12492 35203 12502 35259
rect 12054 35135 12502 35203
rect 12054 35079 12064 35135
rect 12120 35079 12188 35135
rect 12244 35079 12312 35135
rect 12368 35079 12436 35135
rect 12492 35079 12502 35135
rect 12054 35011 12502 35079
rect 12054 34955 12064 35011
rect 12120 34955 12188 35011
rect 12244 34955 12312 35011
rect 12368 34955 12436 35011
rect 12492 34955 12502 35011
rect 12054 34887 12502 34955
rect 12054 34831 12064 34887
rect 12120 34831 12188 34887
rect 12244 34831 12312 34887
rect 12368 34831 12436 34887
rect 12492 34831 12502 34887
rect 12054 34763 12502 34831
rect 12054 34707 12064 34763
rect 12120 34707 12188 34763
rect 12244 34707 12312 34763
rect 12368 34707 12436 34763
rect 12492 34707 12502 34763
rect 12054 34639 12502 34707
rect 12054 34583 12064 34639
rect 12120 34583 12188 34639
rect 12244 34583 12312 34639
rect 12368 34583 12436 34639
rect 12492 34583 12502 34639
rect 12054 34515 12502 34583
rect 12054 34459 12064 34515
rect 12120 34459 12188 34515
rect 12244 34459 12312 34515
rect 12368 34459 12436 34515
rect 12492 34459 12502 34515
rect 12054 34391 12502 34459
rect 12054 34335 12064 34391
rect 12120 34335 12188 34391
rect 12244 34335 12312 34391
rect 12368 34335 12436 34391
rect 12492 34335 12502 34391
rect 12054 34267 12502 34335
rect 12054 34211 12064 34267
rect 12120 34211 12188 34267
rect 12244 34211 12312 34267
rect 12368 34211 12436 34267
rect 12492 34211 12502 34267
rect 12054 34143 12502 34211
rect 12054 34087 12064 34143
rect 12120 34087 12188 34143
rect 12244 34087 12312 34143
rect 12368 34087 12436 34143
rect 12492 34087 12502 34143
rect 12054 34019 12502 34087
rect 12054 33963 12064 34019
rect 12120 33963 12188 34019
rect 12244 33963 12312 34019
rect 12368 33963 12436 34019
rect 12492 33963 12502 34019
rect 12054 33895 12502 33963
rect 12054 33839 12064 33895
rect 12120 33839 12188 33895
rect 12244 33839 12312 33895
rect 12368 33839 12436 33895
rect 12492 33839 12502 33895
rect 12054 33771 12502 33839
rect 12054 33715 12064 33771
rect 12120 33715 12188 33771
rect 12244 33715 12312 33771
rect 12368 33715 12436 33771
rect 12492 33715 12502 33771
rect 12054 33647 12502 33715
rect 12054 33591 12064 33647
rect 12120 33591 12188 33647
rect 12244 33591 12312 33647
rect 12368 33591 12436 33647
rect 12492 33591 12502 33647
rect 12054 33523 12502 33591
rect 12054 33467 12064 33523
rect 12120 33467 12188 33523
rect 12244 33467 12312 33523
rect 12368 33467 12436 33523
rect 12492 33467 12502 33523
rect 12054 33399 12502 33467
rect 12054 33343 12064 33399
rect 12120 33343 12188 33399
rect 12244 33343 12312 33399
rect 12368 33343 12436 33399
rect 12492 33343 12502 33399
rect 12054 33333 12502 33343
rect 13190 36251 13638 36261
rect 13190 36195 13200 36251
rect 13256 36195 13324 36251
rect 13380 36195 13448 36251
rect 13504 36195 13572 36251
rect 13628 36195 13638 36251
rect 13190 36127 13638 36195
rect 13190 36071 13200 36127
rect 13256 36071 13324 36127
rect 13380 36071 13448 36127
rect 13504 36071 13572 36127
rect 13628 36071 13638 36127
rect 13190 36003 13638 36071
rect 13190 35947 13200 36003
rect 13256 35947 13324 36003
rect 13380 35947 13448 36003
rect 13504 35947 13572 36003
rect 13628 35947 13638 36003
rect 13190 35879 13638 35947
rect 13190 35823 13200 35879
rect 13256 35823 13324 35879
rect 13380 35823 13448 35879
rect 13504 35823 13572 35879
rect 13628 35823 13638 35879
rect 13190 35755 13638 35823
rect 13190 35699 13200 35755
rect 13256 35699 13324 35755
rect 13380 35699 13448 35755
rect 13504 35699 13572 35755
rect 13628 35699 13638 35755
rect 13190 35631 13638 35699
rect 13190 35575 13200 35631
rect 13256 35575 13324 35631
rect 13380 35575 13448 35631
rect 13504 35575 13572 35631
rect 13628 35575 13638 35631
rect 13190 35507 13638 35575
rect 13190 35451 13200 35507
rect 13256 35451 13324 35507
rect 13380 35451 13448 35507
rect 13504 35451 13572 35507
rect 13628 35451 13638 35507
rect 13190 35383 13638 35451
rect 13190 35327 13200 35383
rect 13256 35327 13324 35383
rect 13380 35327 13448 35383
rect 13504 35327 13572 35383
rect 13628 35327 13638 35383
rect 13190 35259 13638 35327
rect 13190 35203 13200 35259
rect 13256 35203 13324 35259
rect 13380 35203 13448 35259
rect 13504 35203 13572 35259
rect 13628 35203 13638 35259
rect 13190 35135 13638 35203
rect 13190 35079 13200 35135
rect 13256 35079 13324 35135
rect 13380 35079 13448 35135
rect 13504 35079 13572 35135
rect 13628 35079 13638 35135
rect 13190 35011 13638 35079
rect 13190 34955 13200 35011
rect 13256 34955 13324 35011
rect 13380 34955 13448 35011
rect 13504 34955 13572 35011
rect 13628 34955 13638 35011
rect 13190 34887 13638 34955
rect 13190 34831 13200 34887
rect 13256 34831 13324 34887
rect 13380 34831 13448 34887
rect 13504 34831 13572 34887
rect 13628 34831 13638 34887
rect 13190 34763 13638 34831
rect 13190 34707 13200 34763
rect 13256 34707 13324 34763
rect 13380 34707 13448 34763
rect 13504 34707 13572 34763
rect 13628 34707 13638 34763
rect 13190 34639 13638 34707
rect 13190 34583 13200 34639
rect 13256 34583 13324 34639
rect 13380 34583 13448 34639
rect 13504 34583 13572 34639
rect 13628 34583 13638 34639
rect 13190 34515 13638 34583
rect 13190 34459 13200 34515
rect 13256 34459 13324 34515
rect 13380 34459 13448 34515
rect 13504 34459 13572 34515
rect 13628 34459 13638 34515
rect 13190 34391 13638 34459
rect 13190 34335 13200 34391
rect 13256 34335 13324 34391
rect 13380 34335 13448 34391
rect 13504 34335 13572 34391
rect 13628 34335 13638 34391
rect 13190 34267 13638 34335
rect 13190 34211 13200 34267
rect 13256 34211 13324 34267
rect 13380 34211 13448 34267
rect 13504 34211 13572 34267
rect 13628 34211 13638 34267
rect 13190 34143 13638 34211
rect 13190 34087 13200 34143
rect 13256 34087 13324 34143
rect 13380 34087 13448 34143
rect 13504 34087 13572 34143
rect 13628 34087 13638 34143
rect 13190 34019 13638 34087
rect 13190 33963 13200 34019
rect 13256 33963 13324 34019
rect 13380 33963 13448 34019
rect 13504 33963 13572 34019
rect 13628 33963 13638 34019
rect 13190 33895 13638 33963
rect 13190 33839 13200 33895
rect 13256 33839 13324 33895
rect 13380 33839 13448 33895
rect 13504 33839 13572 33895
rect 13628 33839 13638 33895
rect 13190 33771 13638 33839
rect 13190 33715 13200 33771
rect 13256 33715 13324 33771
rect 13380 33715 13448 33771
rect 13504 33715 13572 33771
rect 13628 33715 13638 33771
rect 13190 33647 13638 33715
rect 13190 33591 13200 33647
rect 13256 33591 13324 33647
rect 13380 33591 13448 33647
rect 13504 33591 13572 33647
rect 13628 33591 13638 33647
rect 13190 33523 13638 33591
rect 13190 33467 13200 33523
rect 13256 33467 13324 33523
rect 13380 33467 13448 33523
rect 13504 33467 13572 33523
rect 13628 33467 13638 33523
rect 13190 33399 13638 33467
rect 13190 33343 13200 33399
rect 13256 33343 13324 33399
rect 13380 33343 13448 33399
rect 13504 33343 13572 33399
rect 13628 33343 13638 33399
rect 13190 33333 13638 33343
rect 14326 36251 14774 36261
rect 14326 36195 14336 36251
rect 14392 36195 14460 36251
rect 14516 36195 14584 36251
rect 14640 36195 14708 36251
rect 14764 36195 14774 36251
rect 14326 36127 14774 36195
rect 14326 36071 14336 36127
rect 14392 36071 14460 36127
rect 14516 36071 14584 36127
rect 14640 36071 14708 36127
rect 14764 36071 14774 36127
rect 14326 36003 14774 36071
rect 14326 35947 14336 36003
rect 14392 35947 14460 36003
rect 14516 35947 14584 36003
rect 14640 35947 14708 36003
rect 14764 35947 14774 36003
rect 14326 35879 14774 35947
rect 14326 35823 14336 35879
rect 14392 35823 14460 35879
rect 14516 35823 14584 35879
rect 14640 35823 14708 35879
rect 14764 35823 14774 35879
rect 14326 35755 14774 35823
rect 14326 35699 14336 35755
rect 14392 35699 14460 35755
rect 14516 35699 14584 35755
rect 14640 35699 14708 35755
rect 14764 35699 14774 35755
rect 14326 35631 14774 35699
rect 14326 35575 14336 35631
rect 14392 35575 14460 35631
rect 14516 35575 14584 35631
rect 14640 35575 14708 35631
rect 14764 35575 14774 35631
rect 14326 35507 14774 35575
rect 14326 35451 14336 35507
rect 14392 35451 14460 35507
rect 14516 35451 14584 35507
rect 14640 35451 14708 35507
rect 14764 35451 14774 35507
rect 14326 35383 14774 35451
rect 14326 35327 14336 35383
rect 14392 35327 14460 35383
rect 14516 35327 14584 35383
rect 14640 35327 14708 35383
rect 14764 35327 14774 35383
rect 14326 35259 14774 35327
rect 14326 35203 14336 35259
rect 14392 35203 14460 35259
rect 14516 35203 14584 35259
rect 14640 35203 14708 35259
rect 14764 35203 14774 35259
rect 14326 35135 14774 35203
rect 14326 35079 14336 35135
rect 14392 35079 14460 35135
rect 14516 35079 14584 35135
rect 14640 35079 14708 35135
rect 14764 35079 14774 35135
rect 14326 35011 14774 35079
rect 14326 34955 14336 35011
rect 14392 34955 14460 35011
rect 14516 34955 14584 35011
rect 14640 34955 14708 35011
rect 14764 34955 14774 35011
rect 14326 34887 14774 34955
rect 14326 34831 14336 34887
rect 14392 34831 14460 34887
rect 14516 34831 14584 34887
rect 14640 34831 14708 34887
rect 14764 34831 14774 34887
rect 14326 34763 14774 34831
rect 14326 34707 14336 34763
rect 14392 34707 14460 34763
rect 14516 34707 14584 34763
rect 14640 34707 14708 34763
rect 14764 34707 14774 34763
rect 14326 34639 14774 34707
rect 14326 34583 14336 34639
rect 14392 34583 14460 34639
rect 14516 34583 14584 34639
rect 14640 34583 14708 34639
rect 14764 34583 14774 34639
rect 14326 34515 14774 34583
rect 14326 34459 14336 34515
rect 14392 34459 14460 34515
rect 14516 34459 14584 34515
rect 14640 34459 14708 34515
rect 14764 34459 14774 34515
rect 14326 34391 14774 34459
rect 14326 34335 14336 34391
rect 14392 34335 14460 34391
rect 14516 34335 14584 34391
rect 14640 34335 14708 34391
rect 14764 34335 14774 34391
rect 14326 34267 14774 34335
rect 14326 34211 14336 34267
rect 14392 34211 14460 34267
rect 14516 34211 14584 34267
rect 14640 34211 14708 34267
rect 14764 34211 14774 34267
rect 14326 34143 14774 34211
rect 14326 34087 14336 34143
rect 14392 34087 14460 34143
rect 14516 34087 14584 34143
rect 14640 34087 14708 34143
rect 14764 34087 14774 34143
rect 14326 34019 14774 34087
rect 14326 33963 14336 34019
rect 14392 33963 14460 34019
rect 14516 33963 14584 34019
rect 14640 33963 14708 34019
rect 14764 33963 14774 34019
rect 14326 33895 14774 33963
rect 14326 33839 14336 33895
rect 14392 33839 14460 33895
rect 14516 33839 14584 33895
rect 14640 33839 14708 33895
rect 14764 33839 14774 33895
rect 14326 33771 14774 33839
rect 14326 33715 14336 33771
rect 14392 33715 14460 33771
rect 14516 33715 14584 33771
rect 14640 33715 14708 33771
rect 14764 33715 14774 33771
rect 14326 33647 14774 33715
rect 14326 33591 14336 33647
rect 14392 33591 14460 33647
rect 14516 33591 14584 33647
rect 14640 33591 14708 33647
rect 14764 33591 14774 33647
rect 14326 33523 14774 33591
rect 14326 33467 14336 33523
rect 14392 33467 14460 33523
rect 14516 33467 14584 33523
rect 14640 33467 14708 33523
rect 14764 33467 14774 33523
rect 14326 33399 14774 33467
rect 14326 33343 14336 33399
rect 14392 33343 14460 33399
rect 14516 33343 14584 33399
rect 14640 33343 14708 33399
rect 14764 33343 14774 33399
rect 14326 33333 14774 33343
rect 858 33051 1306 33061
rect 858 32995 868 33051
rect 924 32995 992 33051
rect 1048 32995 1116 33051
rect 1172 32995 1240 33051
rect 1296 32995 1306 33051
rect 858 32927 1306 32995
rect 858 32871 868 32927
rect 924 32871 992 32927
rect 1048 32871 1116 32927
rect 1172 32871 1240 32927
rect 1296 32871 1306 32927
rect 858 32803 1306 32871
rect 858 32747 868 32803
rect 924 32747 992 32803
rect 1048 32747 1116 32803
rect 1172 32747 1240 32803
rect 1296 32747 1306 32803
rect 858 32679 1306 32747
rect 858 32623 868 32679
rect 924 32623 992 32679
rect 1048 32623 1116 32679
rect 1172 32623 1240 32679
rect 1296 32623 1306 32679
rect 858 32555 1306 32623
rect 858 32499 868 32555
rect 924 32499 992 32555
rect 1048 32499 1116 32555
rect 1172 32499 1240 32555
rect 1296 32499 1306 32555
rect 858 32431 1306 32499
rect 858 32375 868 32431
rect 924 32375 992 32431
rect 1048 32375 1116 32431
rect 1172 32375 1240 32431
rect 1296 32375 1306 32431
rect 858 32307 1306 32375
rect 858 32251 868 32307
rect 924 32251 992 32307
rect 1048 32251 1116 32307
rect 1172 32251 1240 32307
rect 1296 32251 1306 32307
rect 858 32183 1306 32251
rect 858 32127 868 32183
rect 924 32127 992 32183
rect 1048 32127 1116 32183
rect 1172 32127 1240 32183
rect 1296 32127 1306 32183
rect 858 32059 1306 32127
rect 858 32003 868 32059
rect 924 32003 992 32059
rect 1048 32003 1116 32059
rect 1172 32003 1240 32059
rect 1296 32003 1306 32059
rect 858 31935 1306 32003
rect 858 31879 868 31935
rect 924 31879 992 31935
rect 1048 31879 1116 31935
rect 1172 31879 1240 31935
rect 1296 31879 1306 31935
rect 858 31811 1306 31879
rect 858 31755 868 31811
rect 924 31755 992 31811
rect 1048 31755 1116 31811
rect 1172 31755 1240 31811
rect 1296 31755 1306 31811
rect 858 31687 1306 31755
rect 858 31631 868 31687
rect 924 31631 992 31687
rect 1048 31631 1116 31687
rect 1172 31631 1240 31687
rect 1296 31631 1306 31687
rect 858 31563 1306 31631
rect 858 31507 868 31563
rect 924 31507 992 31563
rect 1048 31507 1116 31563
rect 1172 31507 1240 31563
rect 1296 31507 1306 31563
rect 858 31439 1306 31507
rect 858 31383 868 31439
rect 924 31383 992 31439
rect 1048 31383 1116 31439
rect 1172 31383 1240 31439
rect 1296 31383 1306 31439
rect 858 31315 1306 31383
rect 858 31259 868 31315
rect 924 31259 992 31315
rect 1048 31259 1116 31315
rect 1172 31259 1240 31315
rect 1296 31259 1306 31315
rect 858 31191 1306 31259
rect 858 31135 868 31191
rect 924 31135 992 31191
rect 1048 31135 1116 31191
rect 1172 31135 1240 31191
rect 1296 31135 1306 31191
rect 858 31067 1306 31135
rect 858 31011 868 31067
rect 924 31011 992 31067
rect 1048 31011 1116 31067
rect 1172 31011 1240 31067
rect 1296 31011 1306 31067
rect 858 30943 1306 31011
rect 858 30887 868 30943
rect 924 30887 992 30943
rect 1048 30887 1116 30943
rect 1172 30887 1240 30943
rect 1296 30887 1306 30943
rect 858 30819 1306 30887
rect 858 30763 868 30819
rect 924 30763 992 30819
rect 1048 30763 1116 30819
rect 1172 30763 1240 30819
rect 1296 30763 1306 30819
rect 858 30695 1306 30763
rect 858 30639 868 30695
rect 924 30639 992 30695
rect 1048 30639 1116 30695
rect 1172 30639 1240 30695
rect 1296 30639 1306 30695
rect 858 30571 1306 30639
rect 858 30515 868 30571
rect 924 30515 992 30571
rect 1048 30515 1116 30571
rect 1172 30515 1240 30571
rect 1296 30515 1306 30571
rect 858 30447 1306 30515
rect 858 30391 868 30447
rect 924 30391 992 30447
rect 1048 30391 1116 30447
rect 1172 30391 1240 30447
rect 1296 30391 1306 30447
rect 858 30323 1306 30391
rect 858 30267 868 30323
rect 924 30267 992 30323
rect 1048 30267 1116 30323
rect 1172 30267 1240 30323
rect 1296 30267 1306 30323
rect 858 30199 1306 30267
rect 858 30143 868 30199
rect 924 30143 992 30199
rect 1048 30143 1116 30199
rect 1172 30143 1240 30199
rect 1296 30143 1306 30199
rect 858 30133 1306 30143
rect 1994 33051 2442 33061
rect 1994 32995 2004 33051
rect 2060 32995 2128 33051
rect 2184 32995 2252 33051
rect 2308 32995 2376 33051
rect 2432 32995 2442 33051
rect 1994 32927 2442 32995
rect 1994 32871 2004 32927
rect 2060 32871 2128 32927
rect 2184 32871 2252 32927
rect 2308 32871 2376 32927
rect 2432 32871 2442 32927
rect 1994 32803 2442 32871
rect 1994 32747 2004 32803
rect 2060 32747 2128 32803
rect 2184 32747 2252 32803
rect 2308 32747 2376 32803
rect 2432 32747 2442 32803
rect 1994 32679 2442 32747
rect 1994 32623 2004 32679
rect 2060 32623 2128 32679
rect 2184 32623 2252 32679
rect 2308 32623 2376 32679
rect 2432 32623 2442 32679
rect 1994 32555 2442 32623
rect 1994 32499 2004 32555
rect 2060 32499 2128 32555
rect 2184 32499 2252 32555
rect 2308 32499 2376 32555
rect 2432 32499 2442 32555
rect 1994 32431 2442 32499
rect 1994 32375 2004 32431
rect 2060 32375 2128 32431
rect 2184 32375 2252 32431
rect 2308 32375 2376 32431
rect 2432 32375 2442 32431
rect 1994 32307 2442 32375
rect 1994 32251 2004 32307
rect 2060 32251 2128 32307
rect 2184 32251 2252 32307
rect 2308 32251 2376 32307
rect 2432 32251 2442 32307
rect 1994 32183 2442 32251
rect 1994 32127 2004 32183
rect 2060 32127 2128 32183
rect 2184 32127 2252 32183
rect 2308 32127 2376 32183
rect 2432 32127 2442 32183
rect 1994 32059 2442 32127
rect 1994 32003 2004 32059
rect 2060 32003 2128 32059
rect 2184 32003 2252 32059
rect 2308 32003 2376 32059
rect 2432 32003 2442 32059
rect 1994 31935 2442 32003
rect 1994 31879 2004 31935
rect 2060 31879 2128 31935
rect 2184 31879 2252 31935
rect 2308 31879 2376 31935
rect 2432 31879 2442 31935
rect 1994 31811 2442 31879
rect 1994 31755 2004 31811
rect 2060 31755 2128 31811
rect 2184 31755 2252 31811
rect 2308 31755 2376 31811
rect 2432 31755 2442 31811
rect 1994 31687 2442 31755
rect 1994 31631 2004 31687
rect 2060 31631 2128 31687
rect 2184 31631 2252 31687
rect 2308 31631 2376 31687
rect 2432 31631 2442 31687
rect 1994 31563 2442 31631
rect 1994 31507 2004 31563
rect 2060 31507 2128 31563
rect 2184 31507 2252 31563
rect 2308 31507 2376 31563
rect 2432 31507 2442 31563
rect 1994 31439 2442 31507
rect 1994 31383 2004 31439
rect 2060 31383 2128 31439
rect 2184 31383 2252 31439
rect 2308 31383 2376 31439
rect 2432 31383 2442 31439
rect 1994 31315 2442 31383
rect 1994 31259 2004 31315
rect 2060 31259 2128 31315
rect 2184 31259 2252 31315
rect 2308 31259 2376 31315
rect 2432 31259 2442 31315
rect 1994 31191 2442 31259
rect 1994 31135 2004 31191
rect 2060 31135 2128 31191
rect 2184 31135 2252 31191
rect 2308 31135 2376 31191
rect 2432 31135 2442 31191
rect 1994 31067 2442 31135
rect 1994 31011 2004 31067
rect 2060 31011 2128 31067
rect 2184 31011 2252 31067
rect 2308 31011 2376 31067
rect 2432 31011 2442 31067
rect 1994 30943 2442 31011
rect 1994 30887 2004 30943
rect 2060 30887 2128 30943
rect 2184 30887 2252 30943
rect 2308 30887 2376 30943
rect 2432 30887 2442 30943
rect 1994 30819 2442 30887
rect 1994 30763 2004 30819
rect 2060 30763 2128 30819
rect 2184 30763 2252 30819
rect 2308 30763 2376 30819
rect 2432 30763 2442 30819
rect 1994 30695 2442 30763
rect 1994 30639 2004 30695
rect 2060 30639 2128 30695
rect 2184 30639 2252 30695
rect 2308 30639 2376 30695
rect 2432 30639 2442 30695
rect 1994 30571 2442 30639
rect 1994 30515 2004 30571
rect 2060 30515 2128 30571
rect 2184 30515 2252 30571
rect 2308 30515 2376 30571
rect 2432 30515 2442 30571
rect 1994 30447 2442 30515
rect 1994 30391 2004 30447
rect 2060 30391 2128 30447
rect 2184 30391 2252 30447
rect 2308 30391 2376 30447
rect 2432 30391 2442 30447
rect 1994 30323 2442 30391
rect 1994 30267 2004 30323
rect 2060 30267 2128 30323
rect 2184 30267 2252 30323
rect 2308 30267 2376 30323
rect 2432 30267 2442 30323
rect 1994 30199 2442 30267
rect 1994 30143 2004 30199
rect 2060 30143 2128 30199
rect 2184 30143 2252 30199
rect 2308 30143 2376 30199
rect 2432 30143 2442 30199
rect 1994 30133 2442 30143
rect 3698 33051 4146 33061
rect 3698 32995 3708 33051
rect 3764 32995 3832 33051
rect 3888 32995 3956 33051
rect 4012 32995 4080 33051
rect 4136 32995 4146 33051
rect 3698 32927 4146 32995
rect 3698 32871 3708 32927
rect 3764 32871 3832 32927
rect 3888 32871 3956 32927
rect 4012 32871 4080 32927
rect 4136 32871 4146 32927
rect 3698 32803 4146 32871
rect 3698 32747 3708 32803
rect 3764 32747 3832 32803
rect 3888 32747 3956 32803
rect 4012 32747 4080 32803
rect 4136 32747 4146 32803
rect 3698 32679 4146 32747
rect 3698 32623 3708 32679
rect 3764 32623 3832 32679
rect 3888 32623 3956 32679
rect 4012 32623 4080 32679
rect 4136 32623 4146 32679
rect 3698 32555 4146 32623
rect 3698 32499 3708 32555
rect 3764 32499 3832 32555
rect 3888 32499 3956 32555
rect 4012 32499 4080 32555
rect 4136 32499 4146 32555
rect 3698 32431 4146 32499
rect 3698 32375 3708 32431
rect 3764 32375 3832 32431
rect 3888 32375 3956 32431
rect 4012 32375 4080 32431
rect 4136 32375 4146 32431
rect 3698 32307 4146 32375
rect 3698 32251 3708 32307
rect 3764 32251 3832 32307
rect 3888 32251 3956 32307
rect 4012 32251 4080 32307
rect 4136 32251 4146 32307
rect 3698 32183 4146 32251
rect 3698 32127 3708 32183
rect 3764 32127 3832 32183
rect 3888 32127 3956 32183
rect 4012 32127 4080 32183
rect 4136 32127 4146 32183
rect 3698 32059 4146 32127
rect 3698 32003 3708 32059
rect 3764 32003 3832 32059
rect 3888 32003 3956 32059
rect 4012 32003 4080 32059
rect 4136 32003 4146 32059
rect 3698 31935 4146 32003
rect 3698 31879 3708 31935
rect 3764 31879 3832 31935
rect 3888 31879 3956 31935
rect 4012 31879 4080 31935
rect 4136 31879 4146 31935
rect 3698 31811 4146 31879
rect 3698 31755 3708 31811
rect 3764 31755 3832 31811
rect 3888 31755 3956 31811
rect 4012 31755 4080 31811
rect 4136 31755 4146 31811
rect 3698 31687 4146 31755
rect 3698 31631 3708 31687
rect 3764 31631 3832 31687
rect 3888 31631 3956 31687
rect 4012 31631 4080 31687
rect 4136 31631 4146 31687
rect 3698 31563 4146 31631
rect 3698 31507 3708 31563
rect 3764 31507 3832 31563
rect 3888 31507 3956 31563
rect 4012 31507 4080 31563
rect 4136 31507 4146 31563
rect 3698 31439 4146 31507
rect 3698 31383 3708 31439
rect 3764 31383 3832 31439
rect 3888 31383 3956 31439
rect 4012 31383 4080 31439
rect 4136 31383 4146 31439
rect 3698 31315 4146 31383
rect 3698 31259 3708 31315
rect 3764 31259 3832 31315
rect 3888 31259 3956 31315
rect 4012 31259 4080 31315
rect 4136 31259 4146 31315
rect 3698 31191 4146 31259
rect 3698 31135 3708 31191
rect 3764 31135 3832 31191
rect 3888 31135 3956 31191
rect 4012 31135 4080 31191
rect 4136 31135 4146 31191
rect 3698 31067 4146 31135
rect 3698 31011 3708 31067
rect 3764 31011 3832 31067
rect 3888 31011 3956 31067
rect 4012 31011 4080 31067
rect 4136 31011 4146 31067
rect 3698 30943 4146 31011
rect 3698 30887 3708 30943
rect 3764 30887 3832 30943
rect 3888 30887 3956 30943
rect 4012 30887 4080 30943
rect 4136 30887 4146 30943
rect 3698 30819 4146 30887
rect 3698 30763 3708 30819
rect 3764 30763 3832 30819
rect 3888 30763 3956 30819
rect 4012 30763 4080 30819
rect 4136 30763 4146 30819
rect 3698 30695 4146 30763
rect 3698 30639 3708 30695
rect 3764 30639 3832 30695
rect 3888 30639 3956 30695
rect 4012 30639 4080 30695
rect 4136 30639 4146 30695
rect 3698 30571 4146 30639
rect 3698 30515 3708 30571
rect 3764 30515 3832 30571
rect 3888 30515 3956 30571
rect 4012 30515 4080 30571
rect 4136 30515 4146 30571
rect 3698 30447 4146 30515
rect 3698 30391 3708 30447
rect 3764 30391 3832 30447
rect 3888 30391 3956 30447
rect 4012 30391 4080 30447
rect 4136 30391 4146 30447
rect 3698 30323 4146 30391
rect 3698 30267 3708 30323
rect 3764 30267 3832 30323
rect 3888 30267 3956 30323
rect 4012 30267 4080 30323
rect 4136 30267 4146 30323
rect 3698 30199 4146 30267
rect 3698 30143 3708 30199
rect 3764 30143 3832 30199
rect 3888 30143 3956 30199
rect 4012 30143 4080 30199
rect 4136 30143 4146 30199
rect 3698 30133 4146 30143
rect 5970 33051 6418 33061
rect 5970 32995 5980 33051
rect 6036 32995 6104 33051
rect 6160 32995 6228 33051
rect 6284 32995 6352 33051
rect 6408 32995 6418 33051
rect 5970 32927 6418 32995
rect 5970 32871 5980 32927
rect 6036 32871 6104 32927
rect 6160 32871 6228 32927
rect 6284 32871 6352 32927
rect 6408 32871 6418 32927
rect 5970 32803 6418 32871
rect 5970 32747 5980 32803
rect 6036 32747 6104 32803
rect 6160 32747 6228 32803
rect 6284 32747 6352 32803
rect 6408 32747 6418 32803
rect 5970 32679 6418 32747
rect 5970 32623 5980 32679
rect 6036 32623 6104 32679
rect 6160 32623 6228 32679
rect 6284 32623 6352 32679
rect 6408 32623 6418 32679
rect 5970 32555 6418 32623
rect 5970 32499 5980 32555
rect 6036 32499 6104 32555
rect 6160 32499 6228 32555
rect 6284 32499 6352 32555
rect 6408 32499 6418 32555
rect 5970 32431 6418 32499
rect 5970 32375 5980 32431
rect 6036 32375 6104 32431
rect 6160 32375 6228 32431
rect 6284 32375 6352 32431
rect 6408 32375 6418 32431
rect 5970 32307 6418 32375
rect 5970 32251 5980 32307
rect 6036 32251 6104 32307
rect 6160 32251 6228 32307
rect 6284 32251 6352 32307
rect 6408 32251 6418 32307
rect 5970 32183 6418 32251
rect 5970 32127 5980 32183
rect 6036 32127 6104 32183
rect 6160 32127 6228 32183
rect 6284 32127 6352 32183
rect 6408 32127 6418 32183
rect 5970 32059 6418 32127
rect 5970 32003 5980 32059
rect 6036 32003 6104 32059
rect 6160 32003 6228 32059
rect 6284 32003 6352 32059
rect 6408 32003 6418 32059
rect 5970 31935 6418 32003
rect 5970 31879 5980 31935
rect 6036 31879 6104 31935
rect 6160 31879 6228 31935
rect 6284 31879 6352 31935
rect 6408 31879 6418 31935
rect 5970 31811 6418 31879
rect 5970 31755 5980 31811
rect 6036 31755 6104 31811
rect 6160 31755 6228 31811
rect 6284 31755 6352 31811
rect 6408 31755 6418 31811
rect 5970 31687 6418 31755
rect 5970 31631 5980 31687
rect 6036 31631 6104 31687
rect 6160 31631 6228 31687
rect 6284 31631 6352 31687
rect 6408 31631 6418 31687
rect 5970 31563 6418 31631
rect 5970 31507 5980 31563
rect 6036 31507 6104 31563
rect 6160 31507 6228 31563
rect 6284 31507 6352 31563
rect 6408 31507 6418 31563
rect 5970 31439 6418 31507
rect 5970 31383 5980 31439
rect 6036 31383 6104 31439
rect 6160 31383 6228 31439
rect 6284 31383 6352 31439
rect 6408 31383 6418 31439
rect 5970 31315 6418 31383
rect 5970 31259 5980 31315
rect 6036 31259 6104 31315
rect 6160 31259 6228 31315
rect 6284 31259 6352 31315
rect 6408 31259 6418 31315
rect 5970 31191 6418 31259
rect 5970 31135 5980 31191
rect 6036 31135 6104 31191
rect 6160 31135 6228 31191
rect 6284 31135 6352 31191
rect 6408 31135 6418 31191
rect 5970 31067 6418 31135
rect 5970 31011 5980 31067
rect 6036 31011 6104 31067
rect 6160 31011 6228 31067
rect 6284 31011 6352 31067
rect 6408 31011 6418 31067
rect 5970 30943 6418 31011
rect 5970 30887 5980 30943
rect 6036 30887 6104 30943
rect 6160 30887 6228 30943
rect 6284 30887 6352 30943
rect 6408 30887 6418 30943
rect 5970 30819 6418 30887
rect 5970 30763 5980 30819
rect 6036 30763 6104 30819
rect 6160 30763 6228 30819
rect 6284 30763 6352 30819
rect 6408 30763 6418 30819
rect 5970 30695 6418 30763
rect 5970 30639 5980 30695
rect 6036 30639 6104 30695
rect 6160 30639 6228 30695
rect 6284 30639 6352 30695
rect 6408 30639 6418 30695
rect 5970 30571 6418 30639
rect 5970 30515 5980 30571
rect 6036 30515 6104 30571
rect 6160 30515 6228 30571
rect 6284 30515 6352 30571
rect 6408 30515 6418 30571
rect 5970 30447 6418 30515
rect 5970 30391 5980 30447
rect 6036 30391 6104 30447
rect 6160 30391 6228 30447
rect 6284 30391 6352 30447
rect 6408 30391 6418 30447
rect 5970 30323 6418 30391
rect 5970 30267 5980 30323
rect 6036 30267 6104 30323
rect 6160 30267 6228 30323
rect 6284 30267 6352 30323
rect 6408 30267 6418 30323
rect 5970 30199 6418 30267
rect 5970 30143 5980 30199
rect 6036 30143 6104 30199
rect 6160 30143 6228 30199
rect 6284 30143 6352 30199
rect 6408 30143 6418 30199
rect 5970 30133 6418 30143
rect 8646 33051 9094 33061
rect 8646 32995 8656 33051
rect 8712 32995 8780 33051
rect 8836 32995 8904 33051
rect 8960 32995 9028 33051
rect 9084 32995 9094 33051
rect 8646 32927 9094 32995
rect 8646 32871 8656 32927
rect 8712 32871 8780 32927
rect 8836 32871 8904 32927
rect 8960 32871 9028 32927
rect 9084 32871 9094 32927
rect 8646 32803 9094 32871
rect 8646 32747 8656 32803
rect 8712 32747 8780 32803
rect 8836 32747 8904 32803
rect 8960 32747 9028 32803
rect 9084 32747 9094 32803
rect 8646 32679 9094 32747
rect 8646 32623 8656 32679
rect 8712 32623 8780 32679
rect 8836 32623 8904 32679
rect 8960 32623 9028 32679
rect 9084 32623 9094 32679
rect 8646 32555 9094 32623
rect 8646 32499 8656 32555
rect 8712 32499 8780 32555
rect 8836 32499 8904 32555
rect 8960 32499 9028 32555
rect 9084 32499 9094 32555
rect 8646 32431 9094 32499
rect 8646 32375 8656 32431
rect 8712 32375 8780 32431
rect 8836 32375 8904 32431
rect 8960 32375 9028 32431
rect 9084 32375 9094 32431
rect 8646 32307 9094 32375
rect 8646 32251 8656 32307
rect 8712 32251 8780 32307
rect 8836 32251 8904 32307
rect 8960 32251 9028 32307
rect 9084 32251 9094 32307
rect 8646 32183 9094 32251
rect 8646 32127 8656 32183
rect 8712 32127 8780 32183
rect 8836 32127 8904 32183
rect 8960 32127 9028 32183
rect 9084 32127 9094 32183
rect 8646 32059 9094 32127
rect 8646 32003 8656 32059
rect 8712 32003 8780 32059
rect 8836 32003 8904 32059
rect 8960 32003 9028 32059
rect 9084 32003 9094 32059
rect 8646 31935 9094 32003
rect 8646 31879 8656 31935
rect 8712 31879 8780 31935
rect 8836 31879 8904 31935
rect 8960 31879 9028 31935
rect 9084 31879 9094 31935
rect 8646 31811 9094 31879
rect 8646 31755 8656 31811
rect 8712 31755 8780 31811
rect 8836 31755 8904 31811
rect 8960 31755 9028 31811
rect 9084 31755 9094 31811
rect 8646 31687 9094 31755
rect 8646 31631 8656 31687
rect 8712 31631 8780 31687
rect 8836 31631 8904 31687
rect 8960 31631 9028 31687
rect 9084 31631 9094 31687
rect 8646 31563 9094 31631
rect 8646 31507 8656 31563
rect 8712 31507 8780 31563
rect 8836 31507 8904 31563
rect 8960 31507 9028 31563
rect 9084 31507 9094 31563
rect 8646 31439 9094 31507
rect 8646 31383 8656 31439
rect 8712 31383 8780 31439
rect 8836 31383 8904 31439
rect 8960 31383 9028 31439
rect 9084 31383 9094 31439
rect 8646 31315 9094 31383
rect 8646 31259 8656 31315
rect 8712 31259 8780 31315
rect 8836 31259 8904 31315
rect 8960 31259 9028 31315
rect 9084 31259 9094 31315
rect 8646 31191 9094 31259
rect 8646 31135 8656 31191
rect 8712 31135 8780 31191
rect 8836 31135 8904 31191
rect 8960 31135 9028 31191
rect 9084 31135 9094 31191
rect 8646 31067 9094 31135
rect 8646 31011 8656 31067
rect 8712 31011 8780 31067
rect 8836 31011 8904 31067
rect 8960 31011 9028 31067
rect 9084 31011 9094 31067
rect 8646 30943 9094 31011
rect 8646 30887 8656 30943
rect 8712 30887 8780 30943
rect 8836 30887 8904 30943
rect 8960 30887 9028 30943
rect 9084 30887 9094 30943
rect 8646 30819 9094 30887
rect 8646 30763 8656 30819
rect 8712 30763 8780 30819
rect 8836 30763 8904 30819
rect 8960 30763 9028 30819
rect 9084 30763 9094 30819
rect 8646 30695 9094 30763
rect 8646 30639 8656 30695
rect 8712 30639 8780 30695
rect 8836 30639 8904 30695
rect 8960 30639 9028 30695
rect 9084 30639 9094 30695
rect 8646 30571 9094 30639
rect 8646 30515 8656 30571
rect 8712 30515 8780 30571
rect 8836 30515 8904 30571
rect 8960 30515 9028 30571
rect 9084 30515 9094 30571
rect 8646 30447 9094 30515
rect 8646 30391 8656 30447
rect 8712 30391 8780 30447
rect 8836 30391 8904 30447
rect 8960 30391 9028 30447
rect 9084 30391 9094 30447
rect 8646 30323 9094 30391
rect 8646 30267 8656 30323
rect 8712 30267 8780 30323
rect 8836 30267 8904 30323
rect 8960 30267 9028 30323
rect 9084 30267 9094 30323
rect 8646 30199 9094 30267
rect 8646 30143 8656 30199
rect 8712 30143 8780 30199
rect 8836 30143 8904 30199
rect 8960 30143 9028 30199
rect 9084 30143 9094 30199
rect 8646 30133 9094 30143
rect 10918 33051 11366 33061
rect 10918 32995 10928 33051
rect 10984 32995 11052 33051
rect 11108 32995 11176 33051
rect 11232 32995 11300 33051
rect 11356 32995 11366 33051
rect 10918 32927 11366 32995
rect 10918 32871 10928 32927
rect 10984 32871 11052 32927
rect 11108 32871 11176 32927
rect 11232 32871 11300 32927
rect 11356 32871 11366 32927
rect 10918 32803 11366 32871
rect 10918 32747 10928 32803
rect 10984 32747 11052 32803
rect 11108 32747 11176 32803
rect 11232 32747 11300 32803
rect 11356 32747 11366 32803
rect 10918 32679 11366 32747
rect 10918 32623 10928 32679
rect 10984 32623 11052 32679
rect 11108 32623 11176 32679
rect 11232 32623 11300 32679
rect 11356 32623 11366 32679
rect 10918 32555 11366 32623
rect 10918 32499 10928 32555
rect 10984 32499 11052 32555
rect 11108 32499 11176 32555
rect 11232 32499 11300 32555
rect 11356 32499 11366 32555
rect 10918 32431 11366 32499
rect 10918 32375 10928 32431
rect 10984 32375 11052 32431
rect 11108 32375 11176 32431
rect 11232 32375 11300 32431
rect 11356 32375 11366 32431
rect 10918 32307 11366 32375
rect 10918 32251 10928 32307
rect 10984 32251 11052 32307
rect 11108 32251 11176 32307
rect 11232 32251 11300 32307
rect 11356 32251 11366 32307
rect 10918 32183 11366 32251
rect 10918 32127 10928 32183
rect 10984 32127 11052 32183
rect 11108 32127 11176 32183
rect 11232 32127 11300 32183
rect 11356 32127 11366 32183
rect 10918 32059 11366 32127
rect 10918 32003 10928 32059
rect 10984 32003 11052 32059
rect 11108 32003 11176 32059
rect 11232 32003 11300 32059
rect 11356 32003 11366 32059
rect 10918 31935 11366 32003
rect 10918 31879 10928 31935
rect 10984 31879 11052 31935
rect 11108 31879 11176 31935
rect 11232 31879 11300 31935
rect 11356 31879 11366 31935
rect 10918 31811 11366 31879
rect 10918 31755 10928 31811
rect 10984 31755 11052 31811
rect 11108 31755 11176 31811
rect 11232 31755 11300 31811
rect 11356 31755 11366 31811
rect 10918 31687 11366 31755
rect 10918 31631 10928 31687
rect 10984 31631 11052 31687
rect 11108 31631 11176 31687
rect 11232 31631 11300 31687
rect 11356 31631 11366 31687
rect 10918 31563 11366 31631
rect 10918 31507 10928 31563
rect 10984 31507 11052 31563
rect 11108 31507 11176 31563
rect 11232 31507 11300 31563
rect 11356 31507 11366 31563
rect 10918 31439 11366 31507
rect 10918 31383 10928 31439
rect 10984 31383 11052 31439
rect 11108 31383 11176 31439
rect 11232 31383 11300 31439
rect 11356 31383 11366 31439
rect 10918 31315 11366 31383
rect 10918 31259 10928 31315
rect 10984 31259 11052 31315
rect 11108 31259 11176 31315
rect 11232 31259 11300 31315
rect 11356 31259 11366 31315
rect 10918 31191 11366 31259
rect 10918 31135 10928 31191
rect 10984 31135 11052 31191
rect 11108 31135 11176 31191
rect 11232 31135 11300 31191
rect 11356 31135 11366 31191
rect 10918 31067 11366 31135
rect 10918 31011 10928 31067
rect 10984 31011 11052 31067
rect 11108 31011 11176 31067
rect 11232 31011 11300 31067
rect 11356 31011 11366 31067
rect 10918 30943 11366 31011
rect 10918 30887 10928 30943
rect 10984 30887 11052 30943
rect 11108 30887 11176 30943
rect 11232 30887 11300 30943
rect 11356 30887 11366 30943
rect 10918 30819 11366 30887
rect 10918 30763 10928 30819
rect 10984 30763 11052 30819
rect 11108 30763 11176 30819
rect 11232 30763 11300 30819
rect 11356 30763 11366 30819
rect 10918 30695 11366 30763
rect 10918 30639 10928 30695
rect 10984 30639 11052 30695
rect 11108 30639 11176 30695
rect 11232 30639 11300 30695
rect 11356 30639 11366 30695
rect 10918 30571 11366 30639
rect 10918 30515 10928 30571
rect 10984 30515 11052 30571
rect 11108 30515 11176 30571
rect 11232 30515 11300 30571
rect 11356 30515 11366 30571
rect 10918 30447 11366 30515
rect 10918 30391 10928 30447
rect 10984 30391 11052 30447
rect 11108 30391 11176 30447
rect 11232 30391 11300 30447
rect 11356 30391 11366 30447
rect 10918 30323 11366 30391
rect 10918 30267 10928 30323
rect 10984 30267 11052 30323
rect 11108 30267 11176 30323
rect 11232 30267 11300 30323
rect 11356 30267 11366 30323
rect 10918 30199 11366 30267
rect 10918 30143 10928 30199
rect 10984 30143 11052 30199
rect 11108 30143 11176 30199
rect 11232 30143 11300 30199
rect 11356 30143 11366 30199
rect 10918 30133 11366 30143
rect 12622 33051 13070 33061
rect 12622 32995 12632 33051
rect 12688 32995 12756 33051
rect 12812 32995 12880 33051
rect 12936 32995 13004 33051
rect 13060 32995 13070 33051
rect 12622 32927 13070 32995
rect 12622 32871 12632 32927
rect 12688 32871 12756 32927
rect 12812 32871 12880 32927
rect 12936 32871 13004 32927
rect 13060 32871 13070 32927
rect 12622 32803 13070 32871
rect 12622 32747 12632 32803
rect 12688 32747 12756 32803
rect 12812 32747 12880 32803
rect 12936 32747 13004 32803
rect 13060 32747 13070 32803
rect 12622 32679 13070 32747
rect 12622 32623 12632 32679
rect 12688 32623 12756 32679
rect 12812 32623 12880 32679
rect 12936 32623 13004 32679
rect 13060 32623 13070 32679
rect 12622 32555 13070 32623
rect 12622 32499 12632 32555
rect 12688 32499 12756 32555
rect 12812 32499 12880 32555
rect 12936 32499 13004 32555
rect 13060 32499 13070 32555
rect 12622 32431 13070 32499
rect 12622 32375 12632 32431
rect 12688 32375 12756 32431
rect 12812 32375 12880 32431
rect 12936 32375 13004 32431
rect 13060 32375 13070 32431
rect 12622 32307 13070 32375
rect 12622 32251 12632 32307
rect 12688 32251 12756 32307
rect 12812 32251 12880 32307
rect 12936 32251 13004 32307
rect 13060 32251 13070 32307
rect 12622 32183 13070 32251
rect 12622 32127 12632 32183
rect 12688 32127 12756 32183
rect 12812 32127 12880 32183
rect 12936 32127 13004 32183
rect 13060 32127 13070 32183
rect 12622 32059 13070 32127
rect 12622 32003 12632 32059
rect 12688 32003 12756 32059
rect 12812 32003 12880 32059
rect 12936 32003 13004 32059
rect 13060 32003 13070 32059
rect 12622 31935 13070 32003
rect 12622 31879 12632 31935
rect 12688 31879 12756 31935
rect 12812 31879 12880 31935
rect 12936 31879 13004 31935
rect 13060 31879 13070 31935
rect 12622 31811 13070 31879
rect 12622 31755 12632 31811
rect 12688 31755 12756 31811
rect 12812 31755 12880 31811
rect 12936 31755 13004 31811
rect 13060 31755 13070 31811
rect 12622 31687 13070 31755
rect 12622 31631 12632 31687
rect 12688 31631 12756 31687
rect 12812 31631 12880 31687
rect 12936 31631 13004 31687
rect 13060 31631 13070 31687
rect 12622 31563 13070 31631
rect 12622 31507 12632 31563
rect 12688 31507 12756 31563
rect 12812 31507 12880 31563
rect 12936 31507 13004 31563
rect 13060 31507 13070 31563
rect 12622 31439 13070 31507
rect 12622 31383 12632 31439
rect 12688 31383 12756 31439
rect 12812 31383 12880 31439
rect 12936 31383 13004 31439
rect 13060 31383 13070 31439
rect 12622 31315 13070 31383
rect 12622 31259 12632 31315
rect 12688 31259 12756 31315
rect 12812 31259 12880 31315
rect 12936 31259 13004 31315
rect 13060 31259 13070 31315
rect 12622 31191 13070 31259
rect 12622 31135 12632 31191
rect 12688 31135 12756 31191
rect 12812 31135 12880 31191
rect 12936 31135 13004 31191
rect 13060 31135 13070 31191
rect 12622 31067 13070 31135
rect 12622 31011 12632 31067
rect 12688 31011 12756 31067
rect 12812 31011 12880 31067
rect 12936 31011 13004 31067
rect 13060 31011 13070 31067
rect 12622 30943 13070 31011
rect 12622 30887 12632 30943
rect 12688 30887 12756 30943
rect 12812 30887 12880 30943
rect 12936 30887 13004 30943
rect 13060 30887 13070 30943
rect 12622 30819 13070 30887
rect 12622 30763 12632 30819
rect 12688 30763 12756 30819
rect 12812 30763 12880 30819
rect 12936 30763 13004 30819
rect 13060 30763 13070 30819
rect 12622 30695 13070 30763
rect 12622 30639 12632 30695
rect 12688 30639 12756 30695
rect 12812 30639 12880 30695
rect 12936 30639 13004 30695
rect 13060 30639 13070 30695
rect 12622 30571 13070 30639
rect 12622 30515 12632 30571
rect 12688 30515 12756 30571
rect 12812 30515 12880 30571
rect 12936 30515 13004 30571
rect 13060 30515 13070 30571
rect 12622 30447 13070 30515
rect 12622 30391 12632 30447
rect 12688 30391 12756 30447
rect 12812 30391 12880 30447
rect 12936 30391 13004 30447
rect 13060 30391 13070 30447
rect 12622 30323 13070 30391
rect 12622 30267 12632 30323
rect 12688 30267 12756 30323
rect 12812 30267 12880 30323
rect 12936 30267 13004 30323
rect 13060 30267 13070 30323
rect 12622 30199 13070 30267
rect 12622 30143 12632 30199
rect 12688 30143 12756 30199
rect 12812 30143 12880 30199
rect 12936 30143 13004 30199
rect 13060 30143 13070 30199
rect 12622 30133 13070 30143
rect 13758 33051 14206 33061
rect 13758 32995 13768 33051
rect 13824 32995 13892 33051
rect 13948 32995 14016 33051
rect 14072 32995 14140 33051
rect 14196 32995 14206 33051
rect 13758 32927 14206 32995
rect 13758 32871 13768 32927
rect 13824 32871 13892 32927
rect 13948 32871 14016 32927
rect 14072 32871 14140 32927
rect 14196 32871 14206 32927
rect 13758 32803 14206 32871
rect 13758 32747 13768 32803
rect 13824 32747 13892 32803
rect 13948 32747 14016 32803
rect 14072 32747 14140 32803
rect 14196 32747 14206 32803
rect 13758 32679 14206 32747
rect 13758 32623 13768 32679
rect 13824 32623 13892 32679
rect 13948 32623 14016 32679
rect 14072 32623 14140 32679
rect 14196 32623 14206 32679
rect 13758 32555 14206 32623
rect 13758 32499 13768 32555
rect 13824 32499 13892 32555
rect 13948 32499 14016 32555
rect 14072 32499 14140 32555
rect 14196 32499 14206 32555
rect 13758 32431 14206 32499
rect 13758 32375 13768 32431
rect 13824 32375 13892 32431
rect 13948 32375 14016 32431
rect 14072 32375 14140 32431
rect 14196 32375 14206 32431
rect 13758 32307 14206 32375
rect 13758 32251 13768 32307
rect 13824 32251 13892 32307
rect 13948 32251 14016 32307
rect 14072 32251 14140 32307
rect 14196 32251 14206 32307
rect 13758 32183 14206 32251
rect 13758 32127 13768 32183
rect 13824 32127 13892 32183
rect 13948 32127 14016 32183
rect 14072 32127 14140 32183
rect 14196 32127 14206 32183
rect 13758 32059 14206 32127
rect 13758 32003 13768 32059
rect 13824 32003 13892 32059
rect 13948 32003 14016 32059
rect 14072 32003 14140 32059
rect 14196 32003 14206 32059
rect 13758 31935 14206 32003
rect 13758 31879 13768 31935
rect 13824 31879 13892 31935
rect 13948 31879 14016 31935
rect 14072 31879 14140 31935
rect 14196 31879 14206 31935
rect 13758 31811 14206 31879
rect 13758 31755 13768 31811
rect 13824 31755 13892 31811
rect 13948 31755 14016 31811
rect 14072 31755 14140 31811
rect 14196 31755 14206 31811
rect 13758 31687 14206 31755
rect 13758 31631 13768 31687
rect 13824 31631 13892 31687
rect 13948 31631 14016 31687
rect 14072 31631 14140 31687
rect 14196 31631 14206 31687
rect 13758 31563 14206 31631
rect 13758 31507 13768 31563
rect 13824 31507 13892 31563
rect 13948 31507 14016 31563
rect 14072 31507 14140 31563
rect 14196 31507 14206 31563
rect 13758 31439 14206 31507
rect 13758 31383 13768 31439
rect 13824 31383 13892 31439
rect 13948 31383 14016 31439
rect 14072 31383 14140 31439
rect 14196 31383 14206 31439
rect 13758 31315 14206 31383
rect 13758 31259 13768 31315
rect 13824 31259 13892 31315
rect 13948 31259 14016 31315
rect 14072 31259 14140 31315
rect 14196 31259 14206 31315
rect 13758 31191 14206 31259
rect 13758 31135 13768 31191
rect 13824 31135 13892 31191
rect 13948 31135 14016 31191
rect 14072 31135 14140 31191
rect 14196 31135 14206 31191
rect 13758 31067 14206 31135
rect 13758 31011 13768 31067
rect 13824 31011 13892 31067
rect 13948 31011 14016 31067
rect 14072 31011 14140 31067
rect 14196 31011 14206 31067
rect 13758 30943 14206 31011
rect 13758 30887 13768 30943
rect 13824 30887 13892 30943
rect 13948 30887 14016 30943
rect 14072 30887 14140 30943
rect 14196 30887 14206 30943
rect 13758 30819 14206 30887
rect 13758 30763 13768 30819
rect 13824 30763 13892 30819
rect 13948 30763 14016 30819
rect 14072 30763 14140 30819
rect 14196 30763 14206 30819
rect 13758 30695 14206 30763
rect 13758 30639 13768 30695
rect 13824 30639 13892 30695
rect 13948 30639 14016 30695
rect 14072 30639 14140 30695
rect 14196 30639 14206 30695
rect 13758 30571 14206 30639
rect 13758 30515 13768 30571
rect 13824 30515 13892 30571
rect 13948 30515 14016 30571
rect 14072 30515 14140 30571
rect 14196 30515 14206 30571
rect 13758 30447 14206 30515
rect 13758 30391 13768 30447
rect 13824 30391 13892 30447
rect 13948 30391 14016 30447
rect 14072 30391 14140 30447
rect 14196 30391 14206 30447
rect 13758 30323 14206 30391
rect 13758 30267 13768 30323
rect 13824 30267 13892 30323
rect 13948 30267 14016 30323
rect 14072 30267 14140 30323
rect 14196 30267 14206 30323
rect 13758 30199 14206 30267
rect 13758 30143 13768 30199
rect 13824 30143 13892 30199
rect 13948 30143 14016 30199
rect 14072 30143 14140 30199
rect 14196 30143 14206 30199
rect 13758 30133 14206 30143
rect 858 29845 1306 29855
rect 858 29789 868 29845
rect 924 29789 992 29845
rect 1048 29789 1116 29845
rect 1172 29789 1240 29845
rect 1296 29789 1306 29845
rect 858 29721 1306 29789
rect 858 29665 868 29721
rect 924 29665 992 29721
rect 1048 29665 1116 29721
rect 1172 29665 1240 29721
rect 1296 29665 1306 29721
rect 858 29597 1306 29665
rect 858 29541 868 29597
rect 924 29541 992 29597
rect 1048 29541 1116 29597
rect 1172 29541 1240 29597
rect 1296 29541 1306 29597
rect 858 29473 1306 29541
rect 858 29417 868 29473
rect 924 29417 992 29473
rect 1048 29417 1116 29473
rect 1172 29417 1240 29473
rect 1296 29417 1306 29473
rect 858 29349 1306 29417
rect 858 29293 868 29349
rect 924 29293 992 29349
rect 1048 29293 1116 29349
rect 1172 29293 1240 29349
rect 1296 29293 1306 29349
rect 858 29225 1306 29293
rect 858 29169 868 29225
rect 924 29169 992 29225
rect 1048 29169 1116 29225
rect 1172 29169 1240 29225
rect 1296 29169 1306 29225
rect 858 29101 1306 29169
rect 858 29045 868 29101
rect 924 29045 992 29101
rect 1048 29045 1116 29101
rect 1172 29045 1240 29101
rect 1296 29045 1306 29101
rect 858 28977 1306 29045
rect 858 28921 868 28977
rect 924 28921 992 28977
rect 1048 28921 1116 28977
rect 1172 28921 1240 28977
rect 1296 28921 1306 28977
rect 858 28853 1306 28921
rect 858 28797 868 28853
rect 924 28797 992 28853
rect 1048 28797 1116 28853
rect 1172 28797 1240 28853
rect 1296 28797 1306 28853
rect 858 28729 1306 28797
rect 858 28673 868 28729
rect 924 28673 992 28729
rect 1048 28673 1116 28729
rect 1172 28673 1240 28729
rect 1296 28673 1306 28729
rect 858 28605 1306 28673
rect 858 28549 868 28605
rect 924 28549 992 28605
rect 1048 28549 1116 28605
rect 1172 28549 1240 28605
rect 1296 28549 1306 28605
rect 858 28539 1306 28549
rect 1994 29845 2442 29855
rect 1994 29789 2004 29845
rect 2060 29789 2128 29845
rect 2184 29789 2252 29845
rect 2308 29789 2376 29845
rect 2432 29789 2442 29845
rect 1994 29721 2442 29789
rect 1994 29665 2004 29721
rect 2060 29665 2128 29721
rect 2184 29665 2252 29721
rect 2308 29665 2376 29721
rect 2432 29665 2442 29721
rect 1994 29597 2442 29665
rect 1994 29541 2004 29597
rect 2060 29541 2128 29597
rect 2184 29541 2252 29597
rect 2308 29541 2376 29597
rect 2432 29541 2442 29597
rect 1994 29473 2442 29541
rect 1994 29417 2004 29473
rect 2060 29417 2128 29473
rect 2184 29417 2252 29473
rect 2308 29417 2376 29473
rect 2432 29417 2442 29473
rect 1994 29349 2442 29417
rect 1994 29293 2004 29349
rect 2060 29293 2128 29349
rect 2184 29293 2252 29349
rect 2308 29293 2376 29349
rect 2432 29293 2442 29349
rect 1994 29225 2442 29293
rect 1994 29169 2004 29225
rect 2060 29169 2128 29225
rect 2184 29169 2252 29225
rect 2308 29169 2376 29225
rect 2432 29169 2442 29225
rect 1994 29101 2442 29169
rect 1994 29045 2004 29101
rect 2060 29045 2128 29101
rect 2184 29045 2252 29101
rect 2308 29045 2376 29101
rect 2432 29045 2442 29101
rect 1994 28977 2442 29045
rect 1994 28921 2004 28977
rect 2060 28921 2128 28977
rect 2184 28921 2252 28977
rect 2308 28921 2376 28977
rect 2432 28921 2442 28977
rect 1994 28853 2442 28921
rect 1994 28797 2004 28853
rect 2060 28797 2128 28853
rect 2184 28797 2252 28853
rect 2308 28797 2376 28853
rect 2432 28797 2442 28853
rect 1994 28729 2442 28797
rect 1994 28673 2004 28729
rect 2060 28673 2128 28729
rect 2184 28673 2252 28729
rect 2308 28673 2376 28729
rect 2432 28673 2442 28729
rect 1994 28605 2442 28673
rect 1994 28549 2004 28605
rect 2060 28549 2128 28605
rect 2184 28549 2252 28605
rect 2308 28549 2376 28605
rect 2432 28549 2442 28605
rect 1994 28539 2442 28549
rect 3698 29845 4146 29855
rect 3698 29789 3708 29845
rect 3764 29789 3832 29845
rect 3888 29789 3956 29845
rect 4012 29789 4080 29845
rect 4136 29789 4146 29845
rect 3698 29721 4146 29789
rect 3698 29665 3708 29721
rect 3764 29665 3832 29721
rect 3888 29665 3956 29721
rect 4012 29665 4080 29721
rect 4136 29665 4146 29721
rect 3698 29597 4146 29665
rect 3698 29541 3708 29597
rect 3764 29541 3832 29597
rect 3888 29541 3956 29597
rect 4012 29541 4080 29597
rect 4136 29541 4146 29597
rect 3698 29473 4146 29541
rect 3698 29417 3708 29473
rect 3764 29417 3832 29473
rect 3888 29417 3956 29473
rect 4012 29417 4080 29473
rect 4136 29417 4146 29473
rect 3698 29349 4146 29417
rect 3698 29293 3708 29349
rect 3764 29293 3832 29349
rect 3888 29293 3956 29349
rect 4012 29293 4080 29349
rect 4136 29293 4146 29349
rect 3698 29225 4146 29293
rect 3698 29169 3708 29225
rect 3764 29169 3832 29225
rect 3888 29169 3956 29225
rect 4012 29169 4080 29225
rect 4136 29169 4146 29225
rect 3698 29101 4146 29169
rect 3698 29045 3708 29101
rect 3764 29045 3832 29101
rect 3888 29045 3956 29101
rect 4012 29045 4080 29101
rect 4136 29045 4146 29101
rect 3698 28977 4146 29045
rect 3698 28921 3708 28977
rect 3764 28921 3832 28977
rect 3888 28921 3956 28977
rect 4012 28921 4080 28977
rect 4136 28921 4146 28977
rect 3698 28853 4146 28921
rect 3698 28797 3708 28853
rect 3764 28797 3832 28853
rect 3888 28797 3956 28853
rect 4012 28797 4080 28853
rect 4136 28797 4146 28853
rect 3698 28729 4146 28797
rect 3698 28673 3708 28729
rect 3764 28673 3832 28729
rect 3888 28673 3956 28729
rect 4012 28673 4080 28729
rect 4136 28673 4146 28729
rect 3698 28605 4146 28673
rect 3698 28549 3708 28605
rect 3764 28549 3832 28605
rect 3888 28549 3956 28605
rect 4012 28549 4080 28605
rect 4136 28549 4146 28605
rect 3698 28539 4146 28549
rect 5970 29845 6418 29855
rect 5970 29789 5980 29845
rect 6036 29789 6104 29845
rect 6160 29789 6228 29845
rect 6284 29789 6352 29845
rect 6408 29789 6418 29845
rect 5970 29721 6418 29789
rect 5970 29665 5980 29721
rect 6036 29665 6104 29721
rect 6160 29665 6228 29721
rect 6284 29665 6352 29721
rect 6408 29665 6418 29721
rect 5970 29597 6418 29665
rect 5970 29541 5980 29597
rect 6036 29541 6104 29597
rect 6160 29541 6228 29597
rect 6284 29541 6352 29597
rect 6408 29541 6418 29597
rect 5970 29473 6418 29541
rect 5970 29417 5980 29473
rect 6036 29417 6104 29473
rect 6160 29417 6228 29473
rect 6284 29417 6352 29473
rect 6408 29417 6418 29473
rect 5970 29349 6418 29417
rect 5970 29293 5980 29349
rect 6036 29293 6104 29349
rect 6160 29293 6228 29349
rect 6284 29293 6352 29349
rect 6408 29293 6418 29349
rect 5970 29225 6418 29293
rect 5970 29169 5980 29225
rect 6036 29169 6104 29225
rect 6160 29169 6228 29225
rect 6284 29169 6352 29225
rect 6408 29169 6418 29225
rect 5970 29101 6418 29169
rect 5970 29045 5980 29101
rect 6036 29045 6104 29101
rect 6160 29045 6228 29101
rect 6284 29045 6352 29101
rect 6408 29045 6418 29101
rect 5970 28977 6418 29045
rect 5970 28921 5980 28977
rect 6036 28921 6104 28977
rect 6160 28921 6228 28977
rect 6284 28921 6352 28977
rect 6408 28921 6418 28977
rect 5970 28853 6418 28921
rect 5970 28797 5980 28853
rect 6036 28797 6104 28853
rect 6160 28797 6228 28853
rect 6284 28797 6352 28853
rect 6408 28797 6418 28853
rect 5970 28729 6418 28797
rect 5970 28673 5980 28729
rect 6036 28673 6104 28729
rect 6160 28673 6228 28729
rect 6284 28673 6352 28729
rect 6408 28673 6418 28729
rect 5970 28605 6418 28673
rect 5970 28549 5980 28605
rect 6036 28549 6104 28605
rect 6160 28549 6228 28605
rect 6284 28549 6352 28605
rect 6408 28549 6418 28605
rect 5970 28539 6418 28549
rect 8646 29845 9094 29855
rect 8646 29789 8656 29845
rect 8712 29789 8780 29845
rect 8836 29789 8904 29845
rect 8960 29789 9028 29845
rect 9084 29789 9094 29845
rect 8646 29721 9094 29789
rect 8646 29665 8656 29721
rect 8712 29665 8780 29721
rect 8836 29665 8904 29721
rect 8960 29665 9028 29721
rect 9084 29665 9094 29721
rect 8646 29597 9094 29665
rect 8646 29541 8656 29597
rect 8712 29541 8780 29597
rect 8836 29541 8904 29597
rect 8960 29541 9028 29597
rect 9084 29541 9094 29597
rect 8646 29473 9094 29541
rect 8646 29417 8656 29473
rect 8712 29417 8780 29473
rect 8836 29417 8904 29473
rect 8960 29417 9028 29473
rect 9084 29417 9094 29473
rect 8646 29349 9094 29417
rect 8646 29293 8656 29349
rect 8712 29293 8780 29349
rect 8836 29293 8904 29349
rect 8960 29293 9028 29349
rect 9084 29293 9094 29349
rect 8646 29225 9094 29293
rect 8646 29169 8656 29225
rect 8712 29169 8780 29225
rect 8836 29169 8904 29225
rect 8960 29169 9028 29225
rect 9084 29169 9094 29225
rect 8646 29101 9094 29169
rect 8646 29045 8656 29101
rect 8712 29045 8780 29101
rect 8836 29045 8904 29101
rect 8960 29045 9028 29101
rect 9084 29045 9094 29101
rect 8646 28977 9094 29045
rect 8646 28921 8656 28977
rect 8712 28921 8780 28977
rect 8836 28921 8904 28977
rect 8960 28921 9028 28977
rect 9084 28921 9094 28977
rect 8646 28853 9094 28921
rect 8646 28797 8656 28853
rect 8712 28797 8780 28853
rect 8836 28797 8904 28853
rect 8960 28797 9028 28853
rect 9084 28797 9094 28853
rect 8646 28729 9094 28797
rect 8646 28673 8656 28729
rect 8712 28673 8780 28729
rect 8836 28673 8904 28729
rect 8960 28673 9028 28729
rect 9084 28673 9094 28729
rect 8646 28605 9094 28673
rect 8646 28549 8656 28605
rect 8712 28549 8780 28605
rect 8836 28549 8904 28605
rect 8960 28549 9028 28605
rect 9084 28549 9094 28605
rect 8646 28539 9094 28549
rect 10918 29845 11366 29855
rect 10918 29789 10928 29845
rect 10984 29789 11052 29845
rect 11108 29789 11176 29845
rect 11232 29789 11300 29845
rect 11356 29789 11366 29845
rect 10918 29721 11366 29789
rect 10918 29665 10928 29721
rect 10984 29665 11052 29721
rect 11108 29665 11176 29721
rect 11232 29665 11300 29721
rect 11356 29665 11366 29721
rect 10918 29597 11366 29665
rect 10918 29541 10928 29597
rect 10984 29541 11052 29597
rect 11108 29541 11176 29597
rect 11232 29541 11300 29597
rect 11356 29541 11366 29597
rect 10918 29473 11366 29541
rect 10918 29417 10928 29473
rect 10984 29417 11052 29473
rect 11108 29417 11176 29473
rect 11232 29417 11300 29473
rect 11356 29417 11366 29473
rect 10918 29349 11366 29417
rect 10918 29293 10928 29349
rect 10984 29293 11052 29349
rect 11108 29293 11176 29349
rect 11232 29293 11300 29349
rect 11356 29293 11366 29349
rect 10918 29225 11366 29293
rect 10918 29169 10928 29225
rect 10984 29169 11052 29225
rect 11108 29169 11176 29225
rect 11232 29169 11300 29225
rect 11356 29169 11366 29225
rect 10918 29101 11366 29169
rect 10918 29045 10928 29101
rect 10984 29045 11052 29101
rect 11108 29045 11176 29101
rect 11232 29045 11300 29101
rect 11356 29045 11366 29101
rect 10918 28977 11366 29045
rect 10918 28921 10928 28977
rect 10984 28921 11052 28977
rect 11108 28921 11176 28977
rect 11232 28921 11300 28977
rect 11356 28921 11366 28977
rect 10918 28853 11366 28921
rect 10918 28797 10928 28853
rect 10984 28797 11052 28853
rect 11108 28797 11176 28853
rect 11232 28797 11300 28853
rect 11356 28797 11366 28853
rect 10918 28729 11366 28797
rect 10918 28673 10928 28729
rect 10984 28673 11052 28729
rect 11108 28673 11176 28729
rect 11232 28673 11300 28729
rect 11356 28673 11366 28729
rect 10918 28605 11366 28673
rect 10918 28549 10928 28605
rect 10984 28549 11052 28605
rect 11108 28549 11176 28605
rect 11232 28549 11300 28605
rect 11356 28549 11366 28605
rect 10918 28539 11366 28549
rect 12622 29845 13070 29855
rect 12622 29789 12632 29845
rect 12688 29789 12756 29845
rect 12812 29789 12880 29845
rect 12936 29789 13004 29845
rect 13060 29789 13070 29845
rect 12622 29721 13070 29789
rect 12622 29665 12632 29721
rect 12688 29665 12756 29721
rect 12812 29665 12880 29721
rect 12936 29665 13004 29721
rect 13060 29665 13070 29721
rect 12622 29597 13070 29665
rect 12622 29541 12632 29597
rect 12688 29541 12756 29597
rect 12812 29541 12880 29597
rect 12936 29541 13004 29597
rect 13060 29541 13070 29597
rect 12622 29473 13070 29541
rect 12622 29417 12632 29473
rect 12688 29417 12756 29473
rect 12812 29417 12880 29473
rect 12936 29417 13004 29473
rect 13060 29417 13070 29473
rect 12622 29349 13070 29417
rect 12622 29293 12632 29349
rect 12688 29293 12756 29349
rect 12812 29293 12880 29349
rect 12936 29293 13004 29349
rect 13060 29293 13070 29349
rect 12622 29225 13070 29293
rect 12622 29169 12632 29225
rect 12688 29169 12756 29225
rect 12812 29169 12880 29225
rect 12936 29169 13004 29225
rect 13060 29169 13070 29225
rect 12622 29101 13070 29169
rect 12622 29045 12632 29101
rect 12688 29045 12756 29101
rect 12812 29045 12880 29101
rect 12936 29045 13004 29101
rect 13060 29045 13070 29101
rect 12622 28977 13070 29045
rect 12622 28921 12632 28977
rect 12688 28921 12756 28977
rect 12812 28921 12880 28977
rect 12936 28921 13004 28977
rect 13060 28921 13070 28977
rect 12622 28853 13070 28921
rect 12622 28797 12632 28853
rect 12688 28797 12756 28853
rect 12812 28797 12880 28853
rect 12936 28797 13004 28853
rect 13060 28797 13070 28853
rect 12622 28729 13070 28797
rect 12622 28673 12632 28729
rect 12688 28673 12756 28729
rect 12812 28673 12880 28729
rect 12936 28673 13004 28729
rect 13060 28673 13070 28729
rect 12622 28605 13070 28673
rect 12622 28549 12632 28605
rect 12688 28549 12756 28605
rect 12812 28549 12880 28605
rect 12936 28549 13004 28605
rect 13060 28549 13070 28605
rect 12622 28539 13070 28549
rect 13758 29845 14206 29855
rect 13758 29789 13768 29845
rect 13824 29789 13892 29845
rect 13948 29789 14016 29845
rect 14072 29789 14140 29845
rect 14196 29789 14206 29845
rect 13758 29721 14206 29789
rect 13758 29665 13768 29721
rect 13824 29665 13892 29721
rect 13948 29665 14016 29721
rect 14072 29665 14140 29721
rect 14196 29665 14206 29721
rect 13758 29597 14206 29665
rect 13758 29541 13768 29597
rect 13824 29541 13892 29597
rect 13948 29541 14016 29597
rect 14072 29541 14140 29597
rect 14196 29541 14206 29597
rect 13758 29473 14206 29541
rect 13758 29417 13768 29473
rect 13824 29417 13892 29473
rect 13948 29417 14016 29473
rect 14072 29417 14140 29473
rect 14196 29417 14206 29473
rect 13758 29349 14206 29417
rect 13758 29293 13768 29349
rect 13824 29293 13892 29349
rect 13948 29293 14016 29349
rect 14072 29293 14140 29349
rect 14196 29293 14206 29349
rect 13758 29225 14206 29293
rect 13758 29169 13768 29225
rect 13824 29169 13892 29225
rect 13948 29169 14016 29225
rect 14072 29169 14140 29225
rect 14196 29169 14206 29225
rect 13758 29101 14206 29169
rect 13758 29045 13768 29101
rect 13824 29045 13892 29101
rect 13948 29045 14016 29101
rect 14072 29045 14140 29101
rect 14196 29045 14206 29101
rect 13758 28977 14206 29045
rect 13758 28921 13768 28977
rect 13824 28921 13892 28977
rect 13948 28921 14016 28977
rect 14072 28921 14140 28977
rect 14196 28921 14206 28977
rect 13758 28853 14206 28921
rect 13758 28797 13768 28853
rect 13824 28797 13892 28853
rect 13948 28797 14016 28853
rect 14072 28797 14140 28853
rect 14196 28797 14206 28853
rect 13758 28729 14206 28797
rect 13758 28673 13768 28729
rect 13824 28673 13892 28729
rect 13948 28673 14016 28729
rect 14072 28673 14140 28729
rect 14196 28673 14206 28729
rect 13758 28605 14206 28673
rect 13758 28549 13768 28605
rect 13824 28549 13892 28605
rect 13948 28549 14016 28605
rect 14072 28549 14140 28605
rect 14196 28549 14206 28605
rect 13758 28539 14206 28549
rect 290 28245 738 28255
rect 290 28189 300 28245
rect 356 28189 424 28245
rect 480 28189 548 28245
rect 604 28189 672 28245
rect 728 28189 738 28245
rect 290 28121 738 28189
rect 290 28065 300 28121
rect 356 28065 424 28121
rect 480 28065 548 28121
rect 604 28065 672 28121
rect 728 28065 738 28121
rect 290 27997 738 28065
rect 290 27941 300 27997
rect 356 27941 424 27997
rect 480 27941 548 27997
rect 604 27941 672 27997
rect 728 27941 738 27997
rect 290 27873 738 27941
rect 290 27817 300 27873
rect 356 27817 424 27873
rect 480 27817 548 27873
rect 604 27817 672 27873
rect 728 27817 738 27873
rect 290 27749 738 27817
rect 290 27693 300 27749
rect 356 27693 424 27749
rect 480 27693 548 27749
rect 604 27693 672 27749
rect 728 27693 738 27749
rect 290 27625 738 27693
rect 290 27569 300 27625
rect 356 27569 424 27625
rect 480 27569 548 27625
rect 604 27569 672 27625
rect 728 27569 738 27625
rect 290 27501 738 27569
rect 290 27445 300 27501
rect 356 27445 424 27501
rect 480 27445 548 27501
rect 604 27445 672 27501
rect 728 27445 738 27501
rect 290 27377 738 27445
rect 290 27321 300 27377
rect 356 27321 424 27377
rect 480 27321 548 27377
rect 604 27321 672 27377
rect 728 27321 738 27377
rect 290 27253 738 27321
rect 290 27197 300 27253
rect 356 27197 424 27253
rect 480 27197 548 27253
rect 604 27197 672 27253
rect 728 27197 738 27253
rect 290 27129 738 27197
rect 290 27073 300 27129
rect 356 27073 424 27129
rect 480 27073 548 27129
rect 604 27073 672 27129
rect 728 27073 738 27129
rect 290 27005 738 27073
rect 290 26949 300 27005
rect 356 26949 424 27005
rect 480 26949 548 27005
rect 604 26949 672 27005
rect 728 26949 738 27005
rect 290 26939 738 26949
rect 1426 28245 1874 28255
rect 1426 28189 1436 28245
rect 1492 28189 1560 28245
rect 1616 28189 1684 28245
rect 1740 28189 1808 28245
rect 1864 28189 1874 28245
rect 1426 28121 1874 28189
rect 1426 28065 1436 28121
rect 1492 28065 1560 28121
rect 1616 28065 1684 28121
rect 1740 28065 1808 28121
rect 1864 28065 1874 28121
rect 1426 27997 1874 28065
rect 1426 27941 1436 27997
rect 1492 27941 1560 27997
rect 1616 27941 1684 27997
rect 1740 27941 1808 27997
rect 1864 27941 1874 27997
rect 1426 27873 1874 27941
rect 1426 27817 1436 27873
rect 1492 27817 1560 27873
rect 1616 27817 1684 27873
rect 1740 27817 1808 27873
rect 1864 27817 1874 27873
rect 1426 27749 1874 27817
rect 1426 27693 1436 27749
rect 1492 27693 1560 27749
rect 1616 27693 1684 27749
rect 1740 27693 1808 27749
rect 1864 27693 1874 27749
rect 1426 27625 1874 27693
rect 1426 27569 1436 27625
rect 1492 27569 1560 27625
rect 1616 27569 1684 27625
rect 1740 27569 1808 27625
rect 1864 27569 1874 27625
rect 1426 27501 1874 27569
rect 1426 27445 1436 27501
rect 1492 27445 1560 27501
rect 1616 27445 1684 27501
rect 1740 27445 1808 27501
rect 1864 27445 1874 27501
rect 1426 27377 1874 27445
rect 1426 27321 1436 27377
rect 1492 27321 1560 27377
rect 1616 27321 1684 27377
rect 1740 27321 1808 27377
rect 1864 27321 1874 27377
rect 1426 27253 1874 27321
rect 1426 27197 1436 27253
rect 1492 27197 1560 27253
rect 1616 27197 1684 27253
rect 1740 27197 1808 27253
rect 1864 27197 1874 27253
rect 1426 27129 1874 27197
rect 1426 27073 1436 27129
rect 1492 27073 1560 27129
rect 1616 27073 1684 27129
rect 1740 27073 1808 27129
rect 1864 27073 1874 27129
rect 1426 27005 1874 27073
rect 1426 26949 1436 27005
rect 1492 26949 1560 27005
rect 1616 26949 1684 27005
rect 1740 26949 1808 27005
rect 1864 26949 1874 27005
rect 1426 26939 1874 26949
rect 2562 28245 3010 28255
rect 2562 28189 2572 28245
rect 2628 28189 2696 28245
rect 2752 28189 2820 28245
rect 2876 28189 2944 28245
rect 3000 28189 3010 28245
rect 2562 28121 3010 28189
rect 2562 28065 2572 28121
rect 2628 28065 2696 28121
rect 2752 28065 2820 28121
rect 2876 28065 2944 28121
rect 3000 28065 3010 28121
rect 2562 27997 3010 28065
rect 2562 27941 2572 27997
rect 2628 27941 2696 27997
rect 2752 27941 2820 27997
rect 2876 27941 2944 27997
rect 3000 27941 3010 27997
rect 2562 27873 3010 27941
rect 2562 27817 2572 27873
rect 2628 27817 2696 27873
rect 2752 27817 2820 27873
rect 2876 27817 2944 27873
rect 3000 27817 3010 27873
rect 2562 27749 3010 27817
rect 2562 27693 2572 27749
rect 2628 27693 2696 27749
rect 2752 27693 2820 27749
rect 2876 27693 2944 27749
rect 3000 27693 3010 27749
rect 2562 27625 3010 27693
rect 2562 27569 2572 27625
rect 2628 27569 2696 27625
rect 2752 27569 2820 27625
rect 2876 27569 2944 27625
rect 3000 27569 3010 27625
rect 2562 27501 3010 27569
rect 2562 27445 2572 27501
rect 2628 27445 2696 27501
rect 2752 27445 2820 27501
rect 2876 27445 2944 27501
rect 3000 27445 3010 27501
rect 2562 27377 3010 27445
rect 2562 27321 2572 27377
rect 2628 27321 2696 27377
rect 2752 27321 2820 27377
rect 2876 27321 2944 27377
rect 3000 27321 3010 27377
rect 2562 27253 3010 27321
rect 2562 27197 2572 27253
rect 2628 27197 2696 27253
rect 2752 27197 2820 27253
rect 2876 27197 2944 27253
rect 3000 27197 3010 27253
rect 2562 27129 3010 27197
rect 2562 27073 2572 27129
rect 2628 27073 2696 27129
rect 2752 27073 2820 27129
rect 2876 27073 2944 27129
rect 3000 27073 3010 27129
rect 2562 27005 3010 27073
rect 2562 26949 2572 27005
rect 2628 26949 2696 27005
rect 2752 26949 2820 27005
rect 2876 26949 2944 27005
rect 3000 26949 3010 27005
rect 2562 26939 3010 26949
rect 4834 28245 5282 28255
rect 4834 28189 4844 28245
rect 4900 28189 4968 28245
rect 5024 28189 5092 28245
rect 5148 28189 5216 28245
rect 5272 28189 5282 28245
rect 4834 28121 5282 28189
rect 4834 28065 4844 28121
rect 4900 28065 4968 28121
rect 5024 28065 5092 28121
rect 5148 28065 5216 28121
rect 5272 28065 5282 28121
rect 4834 27997 5282 28065
rect 4834 27941 4844 27997
rect 4900 27941 4968 27997
rect 5024 27941 5092 27997
rect 5148 27941 5216 27997
rect 5272 27941 5282 27997
rect 4834 27873 5282 27941
rect 4834 27817 4844 27873
rect 4900 27817 4968 27873
rect 5024 27817 5092 27873
rect 5148 27817 5216 27873
rect 5272 27817 5282 27873
rect 4834 27749 5282 27817
rect 4834 27693 4844 27749
rect 4900 27693 4968 27749
rect 5024 27693 5092 27749
rect 5148 27693 5216 27749
rect 5272 27693 5282 27749
rect 4834 27625 5282 27693
rect 4834 27569 4844 27625
rect 4900 27569 4968 27625
rect 5024 27569 5092 27625
rect 5148 27569 5216 27625
rect 5272 27569 5282 27625
rect 4834 27501 5282 27569
rect 4834 27445 4844 27501
rect 4900 27445 4968 27501
rect 5024 27445 5092 27501
rect 5148 27445 5216 27501
rect 5272 27445 5282 27501
rect 4834 27377 5282 27445
rect 4834 27321 4844 27377
rect 4900 27321 4968 27377
rect 5024 27321 5092 27377
rect 5148 27321 5216 27377
rect 5272 27321 5282 27377
rect 4834 27253 5282 27321
rect 4834 27197 4844 27253
rect 4900 27197 4968 27253
rect 5024 27197 5092 27253
rect 5148 27197 5216 27253
rect 5272 27197 5282 27253
rect 4834 27129 5282 27197
rect 4834 27073 4844 27129
rect 4900 27073 4968 27129
rect 5024 27073 5092 27129
rect 5148 27073 5216 27129
rect 5272 27073 5282 27129
rect 4834 27005 5282 27073
rect 4834 26949 4844 27005
rect 4900 26949 4968 27005
rect 5024 26949 5092 27005
rect 5148 26949 5216 27005
rect 5272 26949 5282 27005
rect 4834 26939 5282 26949
rect 7127 28245 7451 28255
rect 7127 28189 7137 28245
rect 7193 28189 7261 28245
rect 7317 28189 7385 28245
rect 7441 28189 7451 28245
rect 7127 28121 7451 28189
rect 7127 28065 7137 28121
rect 7193 28065 7261 28121
rect 7317 28065 7385 28121
rect 7441 28065 7451 28121
rect 7127 27997 7451 28065
rect 7127 27941 7137 27997
rect 7193 27941 7261 27997
rect 7317 27941 7385 27997
rect 7441 27941 7451 27997
rect 7127 27873 7451 27941
rect 7127 27817 7137 27873
rect 7193 27817 7261 27873
rect 7317 27817 7385 27873
rect 7441 27817 7451 27873
rect 7127 27749 7451 27817
rect 7127 27693 7137 27749
rect 7193 27693 7261 27749
rect 7317 27693 7385 27749
rect 7441 27693 7451 27749
rect 7127 27625 7451 27693
rect 7127 27569 7137 27625
rect 7193 27569 7261 27625
rect 7317 27569 7385 27625
rect 7441 27569 7451 27625
rect 7127 27501 7451 27569
rect 7127 27445 7137 27501
rect 7193 27445 7261 27501
rect 7317 27445 7385 27501
rect 7441 27445 7451 27501
rect 7127 27377 7451 27445
rect 7127 27321 7137 27377
rect 7193 27321 7261 27377
rect 7317 27321 7385 27377
rect 7441 27321 7451 27377
rect 7127 27253 7451 27321
rect 7127 27197 7137 27253
rect 7193 27197 7261 27253
rect 7317 27197 7385 27253
rect 7441 27197 7451 27253
rect 7127 27129 7451 27197
rect 7127 27073 7137 27129
rect 7193 27073 7261 27129
rect 7317 27073 7385 27129
rect 7441 27073 7451 27129
rect 7127 27005 7451 27073
rect 7127 26949 7137 27005
rect 7193 26949 7261 27005
rect 7317 26949 7385 27005
rect 7441 26949 7451 27005
rect 7127 26939 7451 26949
rect 7613 28245 7937 28255
rect 7613 28189 7623 28245
rect 7679 28189 7747 28245
rect 7803 28189 7871 28245
rect 7927 28189 7937 28245
rect 7613 28121 7937 28189
rect 7613 28065 7623 28121
rect 7679 28065 7747 28121
rect 7803 28065 7871 28121
rect 7927 28065 7937 28121
rect 7613 27997 7937 28065
rect 7613 27941 7623 27997
rect 7679 27941 7747 27997
rect 7803 27941 7871 27997
rect 7927 27941 7937 27997
rect 7613 27873 7937 27941
rect 7613 27817 7623 27873
rect 7679 27817 7747 27873
rect 7803 27817 7871 27873
rect 7927 27817 7937 27873
rect 7613 27749 7937 27817
rect 7613 27693 7623 27749
rect 7679 27693 7747 27749
rect 7803 27693 7871 27749
rect 7927 27693 7937 27749
rect 7613 27625 7937 27693
rect 7613 27569 7623 27625
rect 7679 27569 7747 27625
rect 7803 27569 7871 27625
rect 7927 27569 7937 27625
rect 7613 27501 7937 27569
rect 7613 27445 7623 27501
rect 7679 27445 7747 27501
rect 7803 27445 7871 27501
rect 7927 27445 7937 27501
rect 7613 27377 7937 27445
rect 7613 27321 7623 27377
rect 7679 27321 7747 27377
rect 7803 27321 7871 27377
rect 7927 27321 7937 27377
rect 7613 27253 7937 27321
rect 7613 27197 7623 27253
rect 7679 27197 7747 27253
rect 7803 27197 7871 27253
rect 7927 27197 7937 27253
rect 7613 27129 7937 27197
rect 7613 27073 7623 27129
rect 7679 27073 7747 27129
rect 7803 27073 7871 27129
rect 7927 27073 7937 27129
rect 7613 27005 7937 27073
rect 7613 26949 7623 27005
rect 7679 26949 7747 27005
rect 7803 26949 7871 27005
rect 7927 26949 7937 27005
rect 7613 26939 7937 26949
rect 9782 28245 10230 28255
rect 9782 28189 9792 28245
rect 9848 28189 9916 28245
rect 9972 28189 10040 28245
rect 10096 28189 10164 28245
rect 10220 28189 10230 28245
rect 9782 28121 10230 28189
rect 9782 28065 9792 28121
rect 9848 28065 9916 28121
rect 9972 28065 10040 28121
rect 10096 28065 10164 28121
rect 10220 28065 10230 28121
rect 9782 27997 10230 28065
rect 9782 27941 9792 27997
rect 9848 27941 9916 27997
rect 9972 27941 10040 27997
rect 10096 27941 10164 27997
rect 10220 27941 10230 27997
rect 9782 27873 10230 27941
rect 9782 27817 9792 27873
rect 9848 27817 9916 27873
rect 9972 27817 10040 27873
rect 10096 27817 10164 27873
rect 10220 27817 10230 27873
rect 9782 27749 10230 27817
rect 9782 27693 9792 27749
rect 9848 27693 9916 27749
rect 9972 27693 10040 27749
rect 10096 27693 10164 27749
rect 10220 27693 10230 27749
rect 9782 27625 10230 27693
rect 9782 27569 9792 27625
rect 9848 27569 9916 27625
rect 9972 27569 10040 27625
rect 10096 27569 10164 27625
rect 10220 27569 10230 27625
rect 9782 27501 10230 27569
rect 9782 27445 9792 27501
rect 9848 27445 9916 27501
rect 9972 27445 10040 27501
rect 10096 27445 10164 27501
rect 10220 27445 10230 27501
rect 9782 27377 10230 27445
rect 9782 27321 9792 27377
rect 9848 27321 9916 27377
rect 9972 27321 10040 27377
rect 10096 27321 10164 27377
rect 10220 27321 10230 27377
rect 9782 27253 10230 27321
rect 9782 27197 9792 27253
rect 9848 27197 9916 27253
rect 9972 27197 10040 27253
rect 10096 27197 10164 27253
rect 10220 27197 10230 27253
rect 9782 27129 10230 27197
rect 9782 27073 9792 27129
rect 9848 27073 9916 27129
rect 9972 27073 10040 27129
rect 10096 27073 10164 27129
rect 10220 27073 10230 27129
rect 9782 27005 10230 27073
rect 9782 26949 9792 27005
rect 9848 26949 9916 27005
rect 9972 26949 10040 27005
rect 10096 26949 10164 27005
rect 10220 26949 10230 27005
rect 9782 26939 10230 26949
rect 12054 28245 12502 28255
rect 12054 28189 12064 28245
rect 12120 28189 12188 28245
rect 12244 28189 12312 28245
rect 12368 28189 12436 28245
rect 12492 28189 12502 28245
rect 12054 28121 12502 28189
rect 12054 28065 12064 28121
rect 12120 28065 12188 28121
rect 12244 28065 12312 28121
rect 12368 28065 12436 28121
rect 12492 28065 12502 28121
rect 12054 27997 12502 28065
rect 12054 27941 12064 27997
rect 12120 27941 12188 27997
rect 12244 27941 12312 27997
rect 12368 27941 12436 27997
rect 12492 27941 12502 27997
rect 12054 27873 12502 27941
rect 12054 27817 12064 27873
rect 12120 27817 12188 27873
rect 12244 27817 12312 27873
rect 12368 27817 12436 27873
rect 12492 27817 12502 27873
rect 12054 27749 12502 27817
rect 12054 27693 12064 27749
rect 12120 27693 12188 27749
rect 12244 27693 12312 27749
rect 12368 27693 12436 27749
rect 12492 27693 12502 27749
rect 12054 27625 12502 27693
rect 12054 27569 12064 27625
rect 12120 27569 12188 27625
rect 12244 27569 12312 27625
rect 12368 27569 12436 27625
rect 12492 27569 12502 27625
rect 12054 27501 12502 27569
rect 12054 27445 12064 27501
rect 12120 27445 12188 27501
rect 12244 27445 12312 27501
rect 12368 27445 12436 27501
rect 12492 27445 12502 27501
rect 12054 27377 12502 27445
rect 12054 27321 12064 27377
rect 12120 27321 12188 27377
rect 12244 27321 12312 27377
rect 12368 27321 12436 27377
rect 12492 27321 12502 27377
rect 12054 27253 12502 27321
rect 12054 27197 12064 27253
rect 12120 27197 12188 27253
rect 12244 27197 12312 27253
rect 12368 27197 12436 27253
rect 12492 27197 12502 27253
rect 12054 27129 12502 27197
rect 12054 27073 12064 27129
rect 12120 27073 12188 27129
rect 12244 27073 12312 27129
rect 12368 27073 12436 27129
rect 12492 27073 12502 27129
rect 12054 27005 12502 27073
rect 12054 26949 12064 27005
rect 12120 26949 12188 27005
rect 12244 26949 12312 27005
rect 12368 26949 12436 27005
rect 12492 26949 12502 27005
rect 12054 26939 12502 26949
rect 13190 28245 13638 28255
rect 13190 28189 13200 28245
rect 13256 28189 13324 28245
rect 13380 28189 13448 28245
rect 13504 28189 13572 28245
rect 13628 28189 13638 28245
rect 13190 28121 13638 28189
rect 13190 28065 13200 28121
rect 13256 28065 13324 28121
rect 13380 28065 13448 28121
rect 13504 28065 13572 28121
rect 13628 28065 13638 28121
rect 13190 27997 13638 28065
rect 13190 27941 13200 27997
rect 13256 27941 13324 27997
rect 13380 27941 13448 27997
rect 13504 27941 13572 27997
rect 13628 27941 13638 27997
rect 13190 27873 13638 27941
rect 13190 27817 13200 27873
rect 13256 27817 13324 27873
rect 13380 27817 13448 27873
rect 13504 27817 13572 27873
rect 13628 27817 13638 27873
rect 13190 27749 13638 27817
rect 13190 27693 13200 27749
rect 13256 27693 13324 27749
rect 13380 27693 13448 27749
rect 13504 27693 13572 27749
rect 13628 27693 13638 27749
rect 13190 27625 13638 27693
rect 13190 27569 13200 27625
rect 13256 27569 13324 27625
rect 13380 27569 13448 27625
rect 13504 27569 13572 27625
rect 13628 27569 13638 27625
rect 13190 27501 13638 27569
rect 13190 27445 13200 27501
rect 13256 27445 13324 27501
rect 13380 27445 13448 27501
rect 13504 27445 13572 27501
rect 13628 27445 13638 27501
rect 13190 27377 13638 27445
rect 13190 27321 13200 27377
rect 13256 27321 13324 27377
rect 13380 27321 13448 27377
rect 13504 27321 13572 27377
rect 13628 27321 13638 27377
rect 13190 27253 13638 27321
rect 13190 27197 13200 27253
rect 13256 27197 13324 27253
rect 13380 27197 13448 27253
rect 13504 27197 13572 27253
rect 13628 27197 13638 27253
rect 13190 27129 13638 27197
rect 13190 27073 13200 27129
rect 13256 27073 13324 27129
rect 13380 27073 13448 27129
rect 13504 27073 13572 27129
rect 13628 27073 13638 27129
rect 13190 27005 13638 27073
rect 13190 26949 13200 27005
rect 13256 26949 13324 27005
rect 13380 26949 13448 27005
rect 13504 26949 13572 27005
rect 13628 26949 13638 27005
rect 13190 26939 13638 26949
rect 14326 28245 14774 28255
rect 14326 28189 14336 28245
rect 14392 28189 14460 28245
rect 14516 28189 14584 28245
rect 14640 28189 14708 28245
rect 14764 28189 14774 28245
rect 14326 28121 14774 28189
rect 14326 28065 14336 28121
rect 14392 28065 14460 28121
rect 14516 28065 14584 28121
rect 14640 28065 14708 28121
rect 14764 28065 14774 28121
rect 14326 27997 14774 28065
rect 14326 27941 14336 27997
rect 14392 27941 14460 27997
rect 14516 27941 14584 27997
rect 14640 27941 14708 27997
rect 14764 27941 14774 27997
rect 14326 27873 14774 27941
rect 14326 27817 14336 27873
rect 14392 27817 14460 27873
rect 14516 27817 14584 27873
rect 14640 27817 14708 27873
rect 14764 27817 14774 27873
rect 14326 27749 14774 27817
rect 14326 27693 14336 27749
rect 14392 27693 14460 27749
rect 14516 27693 14584 27749
rect 14640 27693 14708 27749
rect 14764 27693 14774 27749
rect 14326 27625 14774 27693
rect 14326 27569 14336 27625
rect 14392 27569 14460 27625
rect 14516 27569 14584 27625
rect 14640 27569 14708 27625
rect 14764 27569 14774 27625
rect 14326 27501 14774 27569
rect 14326 27445 14336 27501
rect 14392 27445 14460 27501
rect 14516 27445 14584 27501
rect 14640 27445 14708 27501
rect 14764 27445 14774 27501
rect 14326 27377 14774 27445
rect 14326 27321 14336 27377
rect 14392 27321 14460 27377
rect 14516 27321 14584 27377
rect 14640 27321 14708 27377
rect 14764 27321 14774 27377
rect 14326 27253 14774 27321
rect 14326 27197 14336 27253
rect 14392 27197 14460 27253
rect 14516 27197 14584 27253
rect 14640 27197 14708 27253
rect 14764 27197 14774 27253
rect 14326 27129 14774 27197
rect 14326 27073 14336 27129
rect 14392 27073 14460 27129
rect 14516 27073 14584 27129
rect 14640 27073 14708 27129
rect 14764 27073 14774 27129
rect 14326 27005 14774 27073
rect 14326 26949 14336 27005
rect 14392 26949 14460 27005
rect 14516 26949 14584 27005
rect 14640 26949 14708 27005
rect 14764 26949 14774 27005
rect 14326 26939 14774 26949
rect 858 26651 1306 26661
rect 858 26595 868 26651
rect 924 26595 992 26651
rect 1048 26595 1116 26651
rect 1172 26595 1240 26651
rect 1296 26595 1306 26651
rect 858 26527 1306 26595
rect 858 26471 868 26527
rect 924 26471 992 26527
rect 1048 26471 1116 26527
rect 1172 26471 1240 26527
rect 1296 26471 1306 26527
rect 858 26403 1306 26471
rect 858 26347 868 26403
rect 924 26347 992 26403
rect 1048 26347 1116 26403
rect 1172 26347 1240 26403
rect 1296 26347 1306 26403
rect 858 26279 1306 26347
rect 858 26223 868 26279
rect 924 26223 992 26279
rect 1048 26223 1116 26279
rect 1172 26223 1240 26279
rect 1296 26223 1306 26279
rect 858 26155 1306 26223
rect 858 26099 868 26155
rect 924 26099 992 26155
rect 1048 26099 1116 26155
rect 1172 26099 1240 26155
rect 1296 26099 1306 26155
rect 858 26031 1306 26099
rect 858 25975 868 26031
rect 924 25975 992 26031
rect 1048 25975 1116 26031
rect 1172 25975 1240 26031
rect 1296 25975 1306 26031
rect 858 25907 1306 25975
rect 858 25851 868 25907
rect 924 25851 992 25907
rect 1048 25851 1116 25907
rect 1172 25851 1240 25907
rect 1296 25851 1306 25907
rect 858 25783 1306 25851
rect 858 25727 868 25783
rect 924 25727 992 25783
rect 1048 25727 1116 25783
rect 1172 25727 1240 25783
rect 1296 25727 1306 25783
rect 858 25659 1306 25727
rect 858 25603 868 25659
rect 924 25603 992 25659
rect 1048 25603 1116 25659
rect 1172 25603 1240 25659
rect 1296 25603 1306 25659
rect 858 25535 1306 25603
rect 858 25479 868 25535
rect 924 25479 992 25535
rect 1048 25479 1116 25535
rect 1172 25479 1240 25535
rect 1296 25479 1306 25535
rect 858 25411 1306 25479
rect 858 25355 868 25411
rect 924 25355 992 25411
rect 1048 25355 1116 25411
rect 1172 25355 1240 25411
rect 1296 25355 1306 25411
rect 858 25287 1306 25355
rect 858 25231 868 25287
rect 924 25231 992 25287
rect 1048 25231 1116 25287
rect 1172 25231 1240 25287
rect 1296 25231 1306 25287
rect 858 25163 1306 25231
rect 858 25107 868 25163
rect 924 25107 992 25163
rect 1048 25107 1116 25163
rect 1172 25107 1240 25163
rect 1296 25107 1306 25163
rect 858 25039 1306 25107
rect 858 24983 868 25039
rect 924 24983 992 25039
rect 1048 24983 1116 25039
rect 1172 24983 1240 25039
rect 1296 24983 1306 25039
rect 858 24915 1306 24983
rect 858 24859 868 24915
rect 924 24859 992 24915
rect 1048 24859 1116 24915
rect 1172 24859 1240 24915
rect 1296 24859 1306 24915
rect 858 24791 1306 24859
rect 858 24735 868 24791
rect 924 24735 992 24791
rect 1048 24735 1116 24791
rect 1172 24735 1240 24791
rect 1296 24735 1306 24791
rect 858 24667 1306 24735
rect 858 24611 868 24667
rect 924 24611 992 24667
rect 1048 24611 1116 24667
rect 1172 24611 1240 24667
rect 1296 24611 1306 24667
rect 858 24543 1306 24611
rect 858 24487 868 24543
rect 924 24487 992 24543
rect 1048 24487 1116 24543
rect 1172 24487 1240 24543
rect 1296 24487 1306 24543
rect 858 24419 1306 24487
rect 858 24363 868 24419
rect 924 24363 992 24419
rect 1048 24363 1116 24419
rect 1172 24363 1240 24419
rect 1296 24363 1306 24419
rect 858 24295 1306 24363
rect 858 24239 868 24295
rect 924 24239 992 24295
rect 1048 24239 1116 24295
rect 1172 24239 1240 24295
rect 1296 24239 1306 24295
rect 858 24171 1306 24239
rect 858 24115 868 24171
rect 924 24115 992 24171
rect 1048 24115 1116 24171
rect 1172 24115 1240 24171
rect 1296 24115 1306 24171
rect 858 24047 1306 24115
rect 858 23991 868 24047
rect 924 23991 992 24047
rect 1048 23991 1116 24047
rect 1172 23991 1240 24047
rect 1296 23991 1306 24047
rect 858 23923 1306 23991
rect 858 23867 868 23923
rect 924 23867 992 23923
rect 1048 23867 1116 23923
rect 1172 23867 1240 23923
rect 1296 23867 1306 23923
rect 858 23799 1306 23867
rect 858 23743 868 23799
rect 924 23743 992 23799
rect 1048 23743 1116 23799
rect 1172 23743 1240 23799
rect 1296 23743 1306 23799
rect 858 23733 1306 23743
rect 1994 26651 2442 26661
rect 1994 26595 2004 26651
rect 2060 26595 2128 26651
rect 2184 26595 2252 26651
rect 2308 26595 2376 26651
rect 2432 26595 2442 26651
rect 1994 26527 2442 26595
rect 1994 26471 2004 26527
rect 2060 26471 2128 26527
rect 2184 26471 2252 26527
rect 2308 26471 2376 26527
rect 2432 26471 2442 26527
rect 1994 26403 2442 26471
rect 1994 26347 2004 26403
rect 2060 26347 2128 26403
rect 2184 26347 2252 26403
rect 2308 26347 2376 26403
rect 2432 26347 2442 26403
rect 1994 26279 2442 26347
rect 1994 26223 2004 26279
rect 2060 26223 2128 26279
rect 2184 26223 2252 26279
rect 2308 26223 2376 26279
rect 2432 26223 2442 26279
rect 1994 26155 2442 26223
rect 1994 26099 2004 26155
rect 2060 26099 2128 26155
rect 2184 26099 2252 26155
rect 2308 26099 2376 26155
rect 2432 26099 2442 26155
rect 1994 26031 2442 26099
rect 1994 25975 2004 26031
rect 2060 25975 2128 26031
rect 2184 25975 2252 26031
rect 2308 25975 2376 26031
rect 2432 25975 2442 26031
rect 1994 25907 2442 25975
rect 1994 25851 2004 25907
rect 2060 25851 2128 25907
rect 2184 25851 2252 25907
rect 2308 25851 2376 25907
rect 2432 25851 2442 25907
rect 1994 25783 2442 25851
rect 1994 25727 2004 25783
rect 2060 25727 2128 25783
rect 2184 25727 2252 25783
rect 2308 25727 2376 25783
rect 2432 25727 2442 25783
rect 1994 25659 2442 25727
rect 1994 25603 2004 25659
rect 2060 25603 2128 25659
rect 2184 25603 2252 25659
rect 2308 25603 2376 25659
rect 2432 25603 2442 25659
rect 1994 25535 2442 25603
rect 1994 25479 2004 25535
rect 2060 25479 2128 25535
rect 2184 25479 2252 25535
rect 2308 25479 2376 25535
rect 2432 25479 2442 25535
rect 1994 25411 2442 25479
rect 1994 25355 2004 25411
rect 2060 25355 2128 25411
rect 2184 25355 2252 25411
rect 2308 25355 2376 25411
rect 2432 25355 2442 25411
rect 1994 25287 2442 25355
rect 1994 25231 2004 25287
rect 2060 25231 2128 25287
rect 2184 25231 2252 25287
rect 2308 25231 2376 25287
rect 2432 25231 2442 25287
rect 1994 25163 2442 25231
rect 1994 25107 2004 25163
rect 2060 25107 2128 25163
rect 2184 25107 2252 25163
rect 2308 25107 2376 25163
rect 2432 25107 2442 25163
rect 1994 25039 2442 25107
rect 1994 24983 2004 25039
rect 2060 24983 2128 25039
rect 2184 24983 2252 25039
rect 2308 24983 2376 25039
rect 2432 24983 2442 25039
rect 1994 24915 2442 24983
rect 1994 24859 2004 24915
rect 2060 24859 2128 24915
rect 2184 24859 2252 24915
rect 2308 24859 2376 24915
rect 2432 24859 2442 24915
rect 1994 24791 2442 24859
rect 1994 24735 2004 24791
rect 2060 24735 2128 24791
rect 2184 24735 2252 24791
rect 2308 24735 2376 24791
rect 2432 24735 2442 24791
rect 1994 24667 2442 24735
rect 1994 24611 2004 24667
rect 2060 24611 2128 24667
rect 2184 24611 2252 24667
rect 2308 24611 2376 24667
rect 2432 24611 2442 24667
rect 1994 24543 2442 24611
rect 1994 24487 2004 24543
rect 2060 24487 2128 24543
rect 2184 24487 2252 24543
rect 2308 24487 2376 24543
rect 2432 24487 2442 24543
rect 1994 24419 2442 24487
rect 1994 24363 2004 24419
rect 2060 24363 2128 24419
rect 2184 24363 2252 24419
rect 2308 24363 2376 24419
rect 2432 24363 2442 24419
rect 1994 24295 2442 24363
rect 1994 24239 2004 24295
rect 2060 24239 2128 24295
rect 2184 24239 2252 24295
rect 2308 24239 2376 24295
rect 2432 24239 2442 24295
rect 1994 24171 2442 24239
rect 1994 24115 2004 24171
rect 2060 24115 2128 24171
rect 2184 24115 2252 24171
rect 2308 24115 2376 24171
rect 2432 24115 2442 24171
rect 1994 24047 2442 24115
rect 1994 23991 2004 24047
rect 2060 23991 2128 24047
rect 2184 23991 2252 24047
rect 2308 23991 2376 24047
rect 2432 23991 2442 24047
rect 1994 23923 2442 23991
rect 1994 23867 2004 23923
rect 2060 23867 2128 23923
rect 2184 23867 2252 23923
rect 2308 23867 2376 23923
rect 2432 23867 2442 23923
rect 1994 23799 2442 23867
rect 1994 23743 2004 23799
rect 2060 23743 2128 23799
rect 2184 23743 2252 23799
rect 2308 23743 2376 23799
rect 2432 23743 2442 23799
rect 1994 23733 2442 23743
rect 3698 26651 4146 26661
rect 3698 26595 3708 26651
rect 3764 26595 3832 26651
rect 3888 26595 3956 26651
rect 4012 26595 4080 26651
rect 4136 26595 4146 26651
rect 3698 26527 4146 26595
rect 3698 26471 3708 26527
rect 3764 26471 3832 26527
rect 3888 26471 3956 26527
rect 4012 26471 4080 26527
rect 4136 26471 4146 26527
rect 3698 26403 4146 26471
rect 3698 26347 3708 26403
rect 3764 26347 3832 26403
rect 3888 26347 3956 26403
rect 4012 26347 4080 26403
rect 4136 26347 4146 26403
rect 3698 26279 4146 26347
rect 3698 26223 3708 26279
rect 3764 26223 3832 26279
rect 3888 26223 3956 26279
rect 4012 26223 4080 26279
rect 4136 26223 4146 26279
rect 3698 26155 4146 26223
rect 3698 26099 3708 26155
rect 3764 26099 3832 26155
rect 3888 26099 3956 26155
rect 4012 26099 4080 26155
rect 4136 26099 4146 26155
rect 3698 26031 4146 26099
rect 3698 25975 3708 26031
rect 3764 25975 3832 26031
rect 3888 25975 3956 26031
rect 4012 25975 4080 26031
rect 4136 25975 4146 26031
rect 3698 25907 4146 25975
rect 3698 25851 3708 25907
rect 3764 25851 3832 25907
rect 3888 25851 3956 25907
rect 4012 25851 4080 25907
rect 4136 25851 4146 25907
rect 3698 25783 4146 25851
rect 3698 25727 3708 25783
rect 3764 25727 3832 25783
rect 3888 25727 3956 25783
rect 4012 25727 4080 25783
rect 4136 25727 4146 25783
rect 3698 25659 4146 25727
rect 3698 25603 3708 25659
rect 3764 25603 3832 25659
rect 3888 25603 3956 25659
rect 4012 25603 4080 25659
rect 4136 25603 4146 25659
rect 3698 25535 4146 25603
rect 3698 25479 3708 25535
rect 3764 25479 3832 25535
rect 3888 25479 3956 25535
rect 4012 25479 4080 25535
rect 4136 25479 4146 25535
rect 3698 25411 4146 25479
rect 3698 25355 3708 25411
rect 3764 25355 3832 25411
rect 3888 25355 3956 25411
rect 4012 25355 4080 25411
rect 4136 25355 4146 25411
rect 3698 25287 4146 25355
rect 3698 25231 3708 25287
rect 3764 25231 3832 25287
rect 3888 25231 3956 25287
rect 4012 25231 4080 25287
rect 4136 25231 4146 25287
rect 3698 25163 4146 25231
rect 3698 25107 3708 25163
rect 3764 25107 3832 25163
rect 3888 25107 3956 25163
rect 4012 25107 4080 25163
rect 4136 25107 4146 25163
rect 3698 25039 4146 25107
rect 3698 24983 3708 25039
rect 3764 24983 3832 25039
rect 3888 24983 3956 25039
rect 4012 24983 4080 25039
rect 4136 24983 4146 25039
rect 3698 24915 4146 24983
rect 3698 24859 3708 24915
rect 3764 24859 3832 24915
rect 3888 24859 3956 24915
rect 4012 24859 4080 24915
rect 4136 24859 4146 24915
rect 3698 24791 4146 24859
rect 3698 24735 3708 24791
rect 3764 24735 3832 24791
rect 3888 24735 3956 24791
rect 4012 24735 4080 24791
rect 4136 24735 4146 24791
rect 3698 24667 4146 24735
rect 3698 24611 3708 24667
rect 3764 24611 3832 24667
rect 3888 24611 3956 24667
rect 4012 24611 4080 24667
rect 4136 24611 4146 24667
rect 3698 24543 4146 24611
rect 3698 24487 3708 24543
rect 3764 24487 3832 24543
rect 3888 24487 3956 24543
rect 4012 24487 4080 24543
rect 4136 24487 4146 24543
rect 3698 24419 4146 24487
rect 3698 24363 3708 24419
rect 3764 24363 3832 24419
rect 3888 24363 3956 24419
rect 4012 24363 4080 24419
rect 4136 24363 4146 24419
rect 3698 24295 4146 24363
rect 3698 24239 3708 24295
rect 3764 24239 3832 24295
rect 3888 24239 3956 24295
rect 4012 24239 4080 24295
rect 4136 24239 4146 24295
rect 3698 24171 4146 24239
rect 3698 24115 3708 24171
rect 3764 24115 3832 24171
rect 3888 24115 3956 24171
rect 4012 24115 4080 24171
rect 4136 24115 4146 24171
rect 3698 24047 4146 24115
rect 3698 23991 3708 24047
rect 3764 23991 3832 24047
rect 3888 23991 3956 24047
rect 4012 23991 4080 24047
rect 4136 23991 4146 24047
rect 3698 23923 4146 23991
rect 3698 23867 3708 23923
rect 3764 23867 3832 23923
rect 3888 23867 3956 23923
rect 4012 23867 4080 23923
rect 4136 23867 4146 23923
rect 3698 23799 4146 23867
rect 3698 23743 3708 23799
rect 3764 23743 3832 23799
rect 3888 23743 3956 23799
rect 4012 23743 4080 23799
rect 4136 23743 4146 23799
rect 3698 23733 4146 23743
rect 5970 26651 6418 26661
rect 5970 26595 5980 26651
rect 6036 26595 6104 26651
rect 6160 26595 6228 26651
rect 6284 26595 6352 26651
rect 6408 26595 6418 26651
rect 5970 26527 6418 26595
rect 5970 26471 5980 26527
rect 6036 26471 6104 26527
rect 6160 26471 6228 26527
rect 6284 26471 6352 26527
rect 6408 26471 6418 26527
rect 5970 26403 6418 26471
rect 5970 26347 5980 26403
rect 6036 26347 6104 26403
rect 6160 26347 6228 26403
rect 6284 26347 6352 26403
rect 6408 26347 6418 26403
rect 5970 26279 6418 26347
rect 5970 26223 5980 26279
rect 6036 26223 6104 26279
rect 6160 26223 6228 26279
rect 6284 26223 6352 26279
rect 6408 26223 6418 26279
rect 5970 26155 6418 26223
rect 5970 26099 5980 26155
rect 6036 26099 6104 26155
rect 6160 26099 6228 26155
rect 6284 26099 6352 26155
rect 6408 26099 6418 26155
rect 5970 26031 6418 26099
rect 5970 25975 5980 26031
rect 6036 25975 6104 26031
rect 6160 25975 6228 26031
rect 6284 25975 6352 26031
rect 6408 25975 6418 26031
rect 5970 25907 6418 25975
rect 5970 25851 5980 25907
rect 6036 25851 6104 25907
rect 6160 25851 6228 25907
rect 6284 25851 6352 25907
rect 6408 25851 6418 25907
rect 5970 25783 6418 25851
rect 5970 25727 5980 25783
rect 6036 25727 6104 25783
rect 6160 25727 6228 25783
rect 6284 25727 6352 25783
rect 6408 25727 6418 25783
rect 5970 25659 6418 25727
rect 5970 25603 5980 25659
rect 6036 25603 6104 25659
rect 6160 25603 6228 25659
rect 6284 25603 6352 25659
rect 6408 25603 6418 25659
rect 5970 25535 6418 25603
rect 5970 25479 5980 25535
rect 6036 25479 6104 25535
rect 6160 25479 6228 25535
rect 6284 25479 6352 25535
rect 6408 25479 6418 25535
rect 5970 25411 6418 25479
rect 5970 25355 5980 25411
rect 6036 25355 6104 25411
rect 6160 25355 6228 25411
rect 6284 25355 6352 25411
rect 6408 25355 6418 25411
rect 5970 25287 6418 25355
rect 5970 25231 5980 25287
rect 6036 25231 6104 25287
rect 6160 25231 6228 25287
rect 6284 25231 6352 25287
rect 6408 25231 6418 25287
rect 5970 25163 6418 25231
rect 5970 25107 5980 25163
rect 6036 25107 6104 25163
rect 6160 25107 6228 25163
rect 6284 25107 6352 25163
rect 6408 25107 6418 25163
rect 5970 25039 6418 25107
rect 5970 24983 5980 25039
rect 6036 24983 6104 25039
rect 6160 24983 6228 25039
rect 6284 24983 6352 25039
rect 6408 24983 6418 25039
rect 5970 24915 6418 24983
rect 5970 24859 5980 24915
rect 6036 24859 6104 24915
rect 6160 24859 6228 24915
rect 6284 24859 6352 24915
rect 6408 24859 6418 24915
rect 5970 24791 6418 24859
rect 5970 24735 5980 24791
rect 6036 24735 6104 24791
rect 6160 24735 6228 24791
rect 6284 24735 6352 24791
rect 6408 24735 6418 24791
rect 5970 24667 6418 24735
rect 5970 24611 5980 24667
rect 6036 24611 6104 24667
rect 6160 24611 6228 24667
rect 6284 24611 6352 24667
rect 6408 24611 6418 24667
rect 5970 24543 6418 24611
rect 5970 24487 5980 24543
rect 6036 24487 6104 24543
rect 6160 24487 6228 24543
rect 6284 24487 6352 24543
rect 6408 24487 6418 24543
rect 5970 24419 6418 24487
rect 5970 24363 5980 24419
rect 6036 24363 6104 24419
rect 6160 24363 6228 24419
rect 6284 24363 6352 24419
rect 6408 24363 6418 24419
rect 5970 24295 6418 24363
rect 5970 24239 5980 24295
rect 6036 24239 6104 24295
rect 6160 24239 6228 24295
rect 6284 24239 6352 24295
rect 6408 24239 6418 24295
rect 5970 24171 6418 24239
rect 5970 24115 5980 24171
rect 6036 24115 6104 24171
rect 6160 24115 6228 24171
rect 6284 24115 6352 24171
rect 6408 24115 6418 24171
rect 5970 24047 6418 24115
rect 5970 23991 5980 24047
rect 6036 23991 6104 24047
rect 6160 23991 6228 24047
rect 6284 23991 6352 24047
rect 6408 23991 6418 24047
rect 5970 23923 6418 23991
rect 5970 23867 5980 23923
rect 6036 23867 6104 23923
rect 6160 23867 6228 23923
rect 6284 23867 6352 23923
rect 6408 23867 6418 23923
rect 5970 23799 6418 23867
rect 5970 23743 5980 23799
rect 6036 23743 6104 23799
rect 6160 23743 6228 23799
rect 6284 23743 6352 23799
rect 6408 23743 6418 23799
rect 5970 23733 6418 23743
rect 8646 26651 9094 26661
rect 8646 26595 8656 26651
rect 8712 26595 8780 26651
rect 8836 26595 8904 26651
rect 8960 26595 9028 26651
rect 9084 26595 9094 26651
rect 8646 26527 9094 26595
rect 8646 26471 8656 26527
rect 8712 26471 8780 26527
rect 8836 26471 8904 26527
rect 8960 26471 9028 26527
rect 9084 26471 9094 26527
rect 8646 26403 9094 26471
rect 8646 26347 8656 26403
rect 8712 26347 8780 26403
rect 8836 26347 8904 26403
rect 8960 26347 9028 26403
rect 9084 26347 9094 26403
rect 8646 26279 9094 26347
rect 8646 26223 8656 26279
rect 8712 26223 8780 26279
rect 8836 26223 8904 26279
rect 8960 26223 9028 26279
rect 9084 26223 9094 26279
rect 8646 26155 9094 26223
rect 8646 26099 8656 26155
rect 8712 26099 8780 26155
rect 8836 26099 8904 26155
rect 8960 26099 9028 26155
rect 9084 26099 9094 26155
rect 8646 26031 9094 26099
rect 8646 25975 8656 26031
rect 8712 25975 8780 26031
rect 8836 25975 8904 26031
rect 8960 25975 9028 26031
rect 9084 25975 9094 26031
rect 8646 25907 9094 25975
rect 8646 25851 8656 25907
rect 8712 25851 8780 25907
rect 8836 25851 8904 25907
rect 8960 25851 9028 25907
rect 9084 25851 9094 25907
rect 8646 25783 9094 25851
rect 8646 25727 8656 25783
rect 8712 25727 8780 25783
rect 8836 25727 8904 25783
rect 8960 25727 9028 25783
rect 9084 25727 9094 25783
rect 8646 25659 9094 25727
rect 8646 25603 8656 25659
rect 8712 25603 8780 25659
rect 8836 25603 8904 25659
rect 8960 25603 9028 25659
rect 9084 25603 9094 25659
rect 8646 25535 9094 25603
rect 8646 25479 8656 25535
rect 8712 25479 8780 25535
rect 8836 25479 8904 25535
rect 8960 25479 9028 25535
rect 9084 25479 9094 25535
rect 8646 25411 9094 25479
rect 8646 25355 8656 25411
rect 8712 25355 8780 25411
rect 8836 25355 8904 25411
rect 8960 25355 9028 25411
rect 9084 25355 9094 25411
rect 8646 25287 9094 25355
rect 8646 25231 8656 25287
rect 8712 25231 8780 25287
rect 8836 25231 8904 25287
rect 8960 25231 9028 25287
rect 9084 25231 9094 25287
rect 8646 25163 9094 25231
rect 8646 25107 8656 25163
rect 8712 25107 8780 25163
rect 8836 25107 8904 25163
rect 8960 25107 9028 25163
rect 9084 25107 9094 25163
rect 8646 25039 9094 25107
rect 8646 24983 8656 25039
rect 8712 24983 8780 25039
rect 8836 24983 8904 25039
rect 8960 24983 9028 25039
rect 9084 24983 9094 25039
rect 8646 24915 9094 24983
rect 8646 24859 8656 24915
rect 8712 24859 8780 24915
rect 8836 24859 8904 24915
rect 8960 24859 9028 24915
rect 9084 24859 9094 24915
rect 8646 24791 9094 24859
rect 8646 24735 8656 24791
rect 8712 24735 8780 24791
rect 8836 24735 8904 24791
rect 8960 24735 9028 24791
rect 9084 24735 9094 24791
rect 8646 24667 9094 24735
rect 8646 24611 8656 24667
rect 8712 24611 8780 24667
rect 8836 24611 8904 24667
rect 8960 24611 9028 24667
rect 9084 24611 9094 24667
rect 8646 24543 9094 24611
rect 8646 24487 8656 24543
rect 8712 24487 8780 24543
rect 8836 24487 8904 24543
rect 8960 24487 9028 24543
rect 9084 24487 9094 24543
rect 8646 24419 9094 24487
rect 8646 24363 8656 24419
rect 8712 24363 8780 24419
rect 8836 24363 8904 24419
rect 8960 24363 9028 24419
rect 9084 24363 9094 24419
rect 8646 24295 9094 24363
rect 8646 24239 8656 24295
rect 8712 24239 8780 24295
rect 8836 24239 8904 24295
rect 8960 24239 9028 24295
rect 9084 24239 9094 24295
rect 8646 24171 9094 24239
rect 8646 24115 8656 24171
rect 8712 24115 8780 24171
rect 8836 24115 8904 24171
rect 8960 24115 9028 24171
rect 9084 24115 9094 24171
rect 8646 24047 9094 24115
rect 8646 23991 8656 24047
rect 8712 23991 8780 24047
rect 8836 23991 8904 24047
rect 8960 23991 9028 24047
rect 9084 23991 9094 24047
rect 8646 23923 9094 23991
rect 8646 23867 8656 23923
rect 8712 23867 8780 23923
rect 8836 23867 8904 23923
rect 8960 23867 9028 23923
rect 9084 23867 9094 23923
rect 8646 23799 9094 23867
rect 8646 23743 8656 23799
rect 8712 23743 8780 23799
rect 8836 23743 8904 23799
rect 8960 23743 9028 23799
rect 9084 23743 9094 23799
rect 8646 23733 9094 23743
rect 10918 26651 11366 26661
rect 10918 26595 10928 26651
rect 10984 26595 11052 26651
rect 11108 26595 11176 26651
rect 11232 26595 11300 26651
rect 11356 26595 11366 26651
rect 10918 26527 11366 26595
rect 10918 26471 10928 26527
rect 10984 26471 11052 26527
rect 11108 26471 11176 26527
rect 11232 26471 11300 26527
rect 11356 26471 11366 26527
rect 10918 26403 11366 26471
rect 10918 26347 10928 26403
rect 10984 26347 11052 26403
rect 11108 26347 11176 26403
rect 11232 26347 11300 26403
rect 11356 26347 11366 26403
rect 10918 26279 11366 26347
rect 10918 26223 10928 26279
rect 10984 26223 11052 26279
rect 11108 26223 11176 26279
rect 11232 26223 11300 26279
rect 11356 26223 11366 26279
rect 10918 26155 11366 26223
rect 10918 26099 10928 26155
rect 10984 26099 11052 26155
rect 11108 26099 11176 26155
rect 11232 26099 11300 26155
rect 11356 26099 11366 26155
rect 10918 26031 11366 26099
rect 10918 25975 10928 26031
rect 10984 25975 11052 26031
rect 11108 25975 11176 26031
rect 11232 25975 11300 26031
rect 11356 25975 11366 26031
rect 10918 25907 11366 25975
rect 10918 25851 10928 25907
rect 10984 25851 11052 25907
rect 11108 25851 11176 25907
rect 11232 25851 11300 25907
rect 11356 25851 11366 25907
rect 10918 25783 11366 25851
rect 10918 25727 10928 25783
rect 10984 25727 11052 25783
rect 11108 25727 11176 25783
rect 11232 25727 11300 25783
rect 11356 25727 11366 25783
rect 10918 25659 11366 25727
rect 10918 25603 10928 25659
rect 10984 25603 11052 25659
rect 11108 25603 11176 25659
rect 11232 25603 11300 25659
rect 11356 25603 11366 25659
rect 10918 25535 11366 25603
rect 10918 25479 10928 25535
rect 10984 25479 11052 25535
rect 11108 25479 11176 25535
rect 11232 25479 11300 25535
rect 11356 25479 11366 25535
rect 10918 25411 11366 25479
rect 10918 25355 10928 25411
rect 10984 25355 11052 25411
rect 11108 25355 11176 25411
rect 11232 25355 11300 25411
rect 11356 25355 11366 25411
rect 10918 25287 11366 25355
rect 10918 25231 10928 25287
rect 10984 25231 11052 25287
rect 11108 25231 11176 25287
rect 11232 25231 11300 25287
rect 11356 25231 11366 25287
rect 10918 25163 11366 25231
rect 10918 25107 10928 25163
rect 10984 25107 11052 25163
rect 11108 25107 11176 25163
rect 11232 25107 11300 25163
rect 11356 25107 11366 25163
rect 10918 25039 11366 25107
rect 10918 24983 10928 25039
rect 10984 24983 11052 25039
rect 11108 24983 11176 25039
rect 11232 24983 11300 25039
rect 11356 24983 11366 25039
rect 10918 24915 11366 24983
rect 10918 24859 10928 24915
rect 10984 24859 11052 24915
rect 11108 24859 11176 24915
rect 11232 24859 11300 24915
rect 11356 24859 11366 24915
rect 10918 24791 11366 24859
rect 10918 24735 10928 24791
rect 10984 24735 11052 24791
rect 11108 24735 11176 24791
rect 11232 24735 11300 24791
rect 11356 24735 11366 24791
rect 10918 24667 11366 24735
rect 10918 24611 10928 24667
rect 10984 24611 11052 24667
rect 11108 24611 11176 24667
rect 11232 24611 11300 24667
rect 11356 24611 11366 24667
rect 10918 24543 11366 24611
rect 10918 24487 10928 24543
rect 10984 24487 11052 24543
rect 11108 24487 11176 24543
rect 11232 24487 11300 24543
rect 11356 24487 11366 24543
rect 10918 24419 11366 24487
rect 10918 24363 10928 24419
rect 10984 24363 11052 24419
rect 11108 24363 11176 24419
rect 11232 24363 11300 24419
rect 11356 24363 11366 24419
rect 10918 24295 11366 24363
rect 10918 24239 10928 24295
rect 10984 24239 11052 24295
rect 11108 24239 11176 24295
rect 11232 24239 11300 24295
rect 11356 24239 11366 24295
rect 10918 24171 11366 24239
rect 10918 24115 10928 24171
rect 10984 24115 11052 24171
rect 11108 24115 11176 24171
rect 11232 24115 11300 24171
rect 11356 24115 11366 24171
rect 10918 24047 11366 24115
rect 10918 23991 10928 24047
rect 10984 23991 11052 24047
rect 11108 23991 11176 24047
rect 11232 23991 11300 24047
rect 11356 23991 11366 24047
rect 10918 23923 11366 23991
rect 10918 23867 10928 23923
rect 10984 23867 11052 23923
rect 11108 23867 11176 23923
rect 11232 23867 11300 23923
rect 11356 23867 11366 23923
rect 10918 23799 11366 23867
rect 10918 23743 10928 23799
rect 10984 23743 11052 23799
rect 11108 23743 11176 23799
rect 11232 23743 11300 23799
rect 11356 23743 11366 23799
rect 10918 23733 11366 23743
rect 12622 26651 13070 26661
rect 12622 26595 12632 26651
rect 12688 26595 12756 26651
rect 12812 26595 12880 26651
rect 12936 26595 13004 26651
rect 13060 26595 13070 26651
rect 12622 26527 13070 26595
rect 12622 26471 12632 26527
rect 12688 26471 12756 26527
rect 12812 26471 12880 26527
rect 12936 26471 13004 26527
rect 13060 26471 13070 26527
rect 12622 26403 13070 26471
rect 12622 26347 12632 26403
rect 12688 26347 12756 26403
rect 12812 26347 12880 26403
rect 12936 26347 13004 26403
rect 13060 26347 13070 26403
rect 12622 26279 13070 26347
rect 12622 26223 12632 26279
rect 12688 26223 12756 26279
rect 12812 26223 12880 26279
rect 12936 26223 13004 26279
rect 13060 26223 13070 26279
rect 12622 26155 13070 26223
rect 12622 26099 12632 26155
rect 12688 26099 12756 26155
rect 12812 26099 12880 26155
rect 12936 26099 13004 26155
rect 13060 26099 13070 26155
rect 12622 26031 13070 26099
rect 12622 25975 12632 26031
rect 12688 25975 12756 26031
rect 12812 25975 12880 26031
rect 12936 25975 13004 26031
rect 13060 25975 13070 26031
rect 12622 25907 13070 25975
rect 12622 25851 12632 25907
rect 12688 25851 12756 25907
rect 12812 25851 12880 25907
rect 12936 25851 13004 25907
rect 13060 25851 13070 25907
rect 12622 25783 13070 25851
rect 12622 25727 12632 25783
rect 12688 25727 12756 25783
rect 12812 25727 12880 25783
rect 12936 25727 13004 25783
rect 13060 25727 13070 25783
rect 12622 25659 13070 25727
rect 12622 25603 12632 25659
rect 12688 25603 12756 25659
rect 12812 25603 12880 25659
rect 12936 25603 13004 25659
rect 13060 25603 13070 25659
rect 12622 25535 13070 25603
rect 12622 25479 12632 25535
rect 12688 25479 12756 25535
rect 12812 25479 12880 25535
rect 12936 25479 13004 25535
rect 13060 25479 13070 25535
rect 12622 25411 13070 25479
rect 12622 25355 12632 25411
rect 12688 25355 12756 25411
rect 12812 25355 12880 25411
rect 12936 25355 13004 25411
rect 13060 25355 13070 25411
rect 12622 25287 13070 25355
rect 12622 25231 12632 25287
rect 12688 25231 12756 25287
rect 12812 25231 12880 25287
rect 12936 25231 13004 25287
rect 13060 25231 13070 25287
rect 12622 25163 13070 25231
rect 12622 25107 12632 25163
rect 12688 25107 12756 25163
rect 12812 25107 12880 25163
rect 12936 25107 13004 25163
rect 13060 25107 13070 25163
rect 12622 25039 13070 25107
rect 12622 24983 12632 25039
rect 12688 24983 12756 25039
rect 12812 24983 12880 25039
rect 12936 24983 13004 25039
rect 13060 24983 13070 25039
rect 12622 24915 13070 24983
rect 12622 24859 12632 24915
rect 12688 24859 12756 24915
rect 12812 24859 12880 24915
rect 12936 24859 13004 24915
rect 13060 24859 13070 24915
rect 12622 24791 13070 24859
rect 12622 24735 12632 24791
rect 12688 24735 12756 24791
rect 12812 24735 12880 24791
rect 12936 24735 13004 24791
rect 13060 24735 13070 24791
rect 12622 24667 13070 24735
rect 12622 24611 12632 24667
rect 12688 24611 12756 24667
rect 12812 24611 12880 24667
rect 12936 24611 13004 24667
rect 13060 24611 13070 24667
rect 12622 24543 13070 24611
rect 12622 24487 12632 24543
rect 12688 24487 12756 24543
rect 12812 24487 12880 24543
rect 12936 24487 13004 24543
rect 13060 24487 13070 24543
rect 12622 24419 13070 24487
rect 12622 24363 12632 24419
rect 12688 24363 12756 24419
rect 12812 24363 12880 24419
rect 12936 24363 13004 24419
rect 13060 24363 13070 24419
rect 12622 24295 13070 24363
rect 12622 24239 12632 24295
rect 12688 24239 12756 24295
rect 12812 24239 12880 24295
rect 12936 24239 13004 24295
rect 13060 24239 13070 24295
rect 12622 24171 13070 24239
rect 12622 24115 12632 24171
rect 12688 24115 12756 24171
rect 12812 24115 12880 24171
rect 12936 24115 13004 24171
rect 13060 24115 13070 24171
rect 12622 24047 13070 24115
rect 12622 23991 12632 24047
rect 12688 23991 12756 24047
rect 12812 23991 12880 24047
rect 12936 23991 13004 24047
rect 13060 23991 13070 24047
rect 12622 23923 13070 23991
rect 12622 23867 12632 23923
rect 12688 23867 12756 23923
rect 12812 23867 12880 23923
rect 12936 23867 13004 23923
rect 13060 23867 13070 23923
rect 12622 23799 13070 23867
rect 12622 23743 12632 23799
rect 12688 23743 12756 23799
rect 12812 23743 12880 23799
rect 12936 23743 13004 23799
rect 13060 23743 13070 23799
rect 12622 23733 13070 23743
rect 13758 26651 14206 26661
rect 13758 26595 13768 26651
rect 13824 26595 13892 26651
rect 13948 26595 14016 26651
rect 14072 26595 14140 26651
rect 14196 26595 14206 26651
rect 13758 26527 14206 26595
rect 13758 26471 13768 26527
rect 13824 26471 13892 26527
rect 13948 26471 14016 26527
rect 14072 26471 14140 26527
rect 14196 26471 14206 26527
rect 13758 26403 14206 26471
rect 13758 26347 13768 26403
rect 13824 26347 13892 26403
rect 13948 26347 14016 26403
rect 14072 26347 14140 26403
rect 14196 26347 14206 26403
rect 13758 26279 14206 26347
rect 13758 26223 13768 26279
rect 13824 26223 13892 26279
rect 13948 26223 14016 26279
rect 14072 26223 14140 26279
rect 14196 26223 14206 26279
rect 13758 26155 14206 26223
rect 13758 26099 13768 26155
rect 13824 26099 13892 26155
rect 13948 26099 14016 26155
rect 14072 26099 14140 26155
rect 14196 26099 14206 26155
rect 13758 26031 14206 26099
rect 13758 25975 13768 26031
rect 13824 25975 13892 26031
rect 13948 25975 14016 26031
rect 14072 25975 14140 26031
rect 14196 25975 14206 26031
rect 13758 25907 14206 25975
rect 13758 25851 13768 25907
rect 13824 25851 13892 25907
rect 13948 25851 14016 25907
rect 14072 25851 14140 25907
rect 14196 25851 14206 25907
rect 13758 25783 14206 25851
rect 13758 25727 13768 25783
rect 13824 25727 13892 25783
rect 13948 25727 14016 25783
rect 14072 25727 14140 25783
rect 14196 25727 14206 25783
rect 13758 25659 14206 25727
rect 13758 25603 13768 25659
rect 13824 25603 13892 25659
rect 13948 25603 14016 25659
rect 14072 25603 14140 25659
rect 14196 25603 14206 25659
rect 13758 25535 14206 25603
rect 13758 25479 13768 25535
rect 13824 25479 13892 25535
rect 13948 25479 14016 25535
rect 14072 25479 14140 25535
rect 14196 25479 14206 25535
rect 13758 25411 14206 25479
rect 13758 25355 13768 25411
rect 13824 25355 13892 25411
rect 13948 25355 14016 25411
rect 14072 25355 14140 25411
rect 14196 25355 14206 25411
rect 13758 25287 14206 25355
rect 13758 25231 13768 25287
rect 13824 25231 13892 25287
rect 13948 25231 14016 25287
rect 14072 25231 14140 25287
rect 14196 25231 14206 25287
rect 13758 25163 14206 25231
rect 13758 25107 13768 25163
rect 13824 25107 13892 25163
rect 13948 25107 14016 25163
rect 14072 25107 14140 25163
rect 14196 25107 14206 25163
rect 13758 25039 14206 25107
rect 13758 24983 13768 25039
rect 13824 24983 13892 25039
rect 13948 24983 14016 25039
rect 14072 24983 14140 25039
rect 14196 24983 14206 25039
rect 13758 24915 14206 24983
rect 13758 24859 13768 24915
rect 13824 24859 13892 24915
rect 13948 24859 14016 24915
rect 14072 24859 14140 24915
rect 14196 24859 14206 24915
rect 13758 24791 14206 24859
rect 13758 24735 13768 24791
rect 13824 24735 13892 24791
rect 13948 24735 14016 24791
rect 14072 24735 14140 24791
rect 14196 24735 14206 24791
rect 13758 24667 14206 24735
rect 13758 24611 13768 24667
rect 13824 24611 13892 24667
rect 13948 24611 14016 24667
rect 14072 24611 14140 24667
rect 14196 24611 14206 24667
rect 13758 24543 14206 24611
rect 13758 24487 13768 24543
rect 13824 24487 13892 24543
rect 13948 24487 14016 24543
rect 14072 24487 14140 24543
rect 14196 24487 14206 24543
rect 13758 24419 14206 24487
rect 13758 24363 13768 24419
rect 13824 24363 13892 24419
rect 13948 24363 14016 24419
rect 14072 24363 14140 24419
rect 14196 24363 14206 24419
rect 13758 24295 14206 24363
rect 13758 24239 13768 24295
rect 13824 24239 13892 24295
rect 13948 24239 14016 24295
rect 14072 24239 14140 24295
rect 14196 24239 14206 24295
rect 13758 24171 14206 24239
rect 13758 24115 13768 24171
rect 13824 24115 13892 24171
rect 13948 24115 14016 24171
rect 14072 24115 14140 24171
rect 14196 24115 14206 24171
rect 13758 24047 14206 24115
rect 13758 23991 13768 24047
rect 13824 23991 13892 24047
rect 13948 23991 14016 24047
rect 14072 23991 14140 24047
rect 14196 23991 14206 24047
rect 13758 23923 14206 23991
rect 13758 23867 13768 23923
rect 13824 23867 13892 23923
rect 13948 23867 14016 23923
rect 14072 23867 14140 23923
rect 14196 23867 14206 23923
rect 13758 23799 14206 23867
rect 13758 23743 13768 23799
rect 13824 23743 13892 23799
rect 13948 23743 14016 23799
rect 14072 23743 14140 23799
rect 14196 23743 14206 23799
rect 13758 23733 14206 23743
rect 858 23451 1306 23461
rect 858 23395 868 23451
rect 924 23395 992 23451
rect 1048 23395 1116 23451
rect 1172 23395 1240 23451
rect 1296 23395 1306 23451
rect 858 23327 1306 23395
rect 858 23271 868 23327
rect 924 23271 992 23327
rect 1048 23271 1116 23327
rect 1172 23271 1240 23327
rect 1296 23271 1306 23327
rect 858 23203 1306 23271
rect 858 23147 868 23203
rect 924 23147 992 23203
rect 1048 23147 1116 23203
rect 1172 23147 1240 23203
rect 1296 23147 1306 23203
rect 858 23079 1306 23147
rect 858 23023 868 23079
rect 924 23023 992 23079
rect 1048 23023 1116 23079
rect 1172 23023 1240 23079
rect 1296 23023 1306 23079
rect 858 22955 1306 23023
rect 858 22899 868 22955
rect 924 22899 992 22955
rect 1048 22899 1116 22955
rect 1172 22899 1240 22955
rect 1296 22899 1306 22955
rect 858 22831 1306 22899
rect 858 22775 868 22831
rect 924 22775 992 22831
rect 1048 22775 1116 22831
rect 1172 22775 1240 22831
rect 1296 22775 1306 22831
rect 858 22707 1306 22775
rect 858 22651 868 22707
rect 924 22651 992 22707
rect 1048 22651 1116 22707
rect 1172 22651 1240 22707
rect 1296 22651 1306 22707
rect 858 22583 1306 22651
rect 858 22527 868 22583
rect 924 22527 992 22583
rect 1048 22527 1116 22583
rect 1172 22527 1240 22583
rect 1296 22527 1306 22583
rect 858 22459 1306 22527
rect 858 22403 868 22459
rect 924 22403 992 22459
rect 1048 22403 1116 22459
rect 1172 22403 1240 22459
rect 1296 22403 1306 22459
rect 858 22335 1306 22403
rect 858 22279 868 22335
rect 924 22279 992 22335
rect 1048 22279 1116 22335
rect 1172 22279 1240 22335
rect 1296 22279 1306 22335
rect 858 22211 1306 22279
rect 858 22155 868 22211
rect 924 22155 992 22211
rect 1048 22155 1116 22211
rect 1172 22155 1240 22211
rect 1296 22155 1306 22211
rect 858 22087 1306 22155
rect 858 22031 868 22087
rect 924 22031 992 22087
rect 1048 22031 1116 22087
rect 1172 22031 1240 22087
rect 1296 22031 1306 22087
rect 858 21963 1306 22031
rect 858 21907 868 21963
rect 924 21907 992 21963
rect 1048 21907 1116 21963
rect 1172 21907 1240 21963
rect 1296 21907 1306 21963
rect 858 21839 1306 21907
rect 858 21783 868 21839
rect 924 21783 992 21839
rect 1048 21783 1116 21839
rect 1172 21783 1240 21839
rect 1296 21783 1306 21839
rect 858 21715 1306 21783
rect 858 21659 868 21715
rect 924 21659 992 21715
rect 1048 21659 1116 21715
rect 1172 21659 1240 21715
rect 1296 21659 1306 21715
rect 858 21591 1306 21659
rect 858 21535 868 21591
rect 924 21535 992 21591
rect 1048 21535 1116 21591
rect 1172 21535 1240 21591
rect 1296 21535 1306 21591
rect 858 21467 1306 21535
rect 858 21411 868 21467
rect 924 21411 992 21467
rect 1048 21411 1116 21467
rect 1172 21411 1240 21467
rect 1296 21411 1306 21467
rect 858 21343 1306 21411
rect 858 21287 868 21343
rect 924 21287 992 21343
rect 1048 21287 1116 21343
rect 1172 21287 1240 21343
rect 1296 21287 1306 21343
rect 858 21219 1306 21287
rect 858 21163 868 21219
rect 924 21163 992 21219
rect 1048 21163 1116 21219
rect 1172 21163 1240 21219
rect 1296 21163 1306 21219
rect 858 21095 1306 21163
rect 858 21039 868 21095
rect 924 21039 992 21095
rect 1048 21039 1116 21095
rect 1172 21039 1240 21095
rect 1296 21039 1306 21095
rect 858 20971 1306 21039
rect 858 20915 868 20971
rect 924 20915 992 20971
rect 1048 20915 1116 20971
rect 1172 20915 1240 20971
rect 1296 20915 1306 20971
rect 858 20847 1306 20915
rect 858 20791 868 20847
rect 924 20791 992 20847
rect 1048 20791 1116 20847
rect 1172 20791 1240 20847
rect 1296 20791 1306 20847
rect 858 20723 1306 20791
rect 858 20667 868 20723
rect 924 20667 992 20723
rect 1048 20667 1116 20723
rect 1172 20667 1240 20723
rect 1296 20667 1306 20723
rect 858 20599 1306 20667
rect 858 20543 868 20599
rect 924 20543 992 20599
rect 1048 20543 1116 20599
rect 1172 20543 1240 20599
rect 1296 20543 1306 20599
rect 858 20533 1306 20543
rect 1994 23451 2442 23461
rect 1994 23395 2004 23451
rect 2060 23395 2128 23451
rect 2184 23395 2252 23451
rect 2308 23395 2376 23451
rect 2432 23395 2442 23451
rect 1994 23327 2442 23395
rect 1994 23271 2004 23327
rect 2060 23271 2128 23327
rect 2184 23271 2252 23327
rect 2308 23271 2376 23327
rect 2432 23271 2442 23327
rect 1994 23203 2442 23271
rect 1994 23147 2004 23203
rect 2060 23147 2128 23203
rect 2184 23147 2252 23203
rect 2308 23147 2376 23203
rect 2432 23147 2442 23203
rect 1994 23079 2442 23147
rect 1994 23023 2004 23079
rect 2060 23023 2128 23079
rect 2184 23023 2252 23079
rect 2308 23023 2376 23079
rect 2432 23023 2442 23079
rect 1994 22955 2442 23023
rect 1994 22899 2004 22955
rect 2060 22899 2128 22955
rect 2184 22899 2252 22955
rect 2308 22899 2376 22955
rect 2432 22899 2442 22955
rect 1994 22831 2442 22899
rect 1994 22775 2004 22831
rect 2060 22775 2128 22831
rect 2184 22775 2252 22831
rect 2308 22775 2376 22831
rect 2432 22775 2442 22831
rect 1994 22707 2442 22775
rect 1994 22651 2004 22707
rect 2060 22651 2128 22707
rect 2184 22651 2252 22707
rect 2308 22651 2376 22707
rect 2432 22651 2442 22707
rect 1994 22583 2442 22651
rect 1994 22527 2004 22583
rect 2060 22527 2128 22583
rect 2184 22527 2252 22583
rect 2308 22527 2376 22583
rect 2432 22527 2442 22583
rect 1994 22459 2442 22527
rect 1994 22403 2004 22459
rect 2060 22403 2128 22459
rect 2184 22403 2252 22459
rect 2308 22403 2376 22459
rect 2432 22403 2442 22459
rect 1994 22335 2442 22403
rect 1994 22279 2004 22335
rect 2060 22279 2128 22335
rect 2184 22279 2252 22335
rect 2308 22279 2376 22335
rect 2432 22279 2442 22335
rect 1994 22211 2442 22279
rect 1994 22155 2004 22211
rect 2060 22155 2128 22211
rect 2184 22155 2252 22211
rect 2308 22155 2376 22211
rect 2432 22155 2442 22211
rect 1994 22087 2442 22155
rect 1994 22031 2004 22087
rect 2060 22031 2128 22087
rect 2184 22031 2252 22087
rect 2308 22031 2376 22087
rect 2432 22031 2442 22087
rect 1994 21963 2442 22031
rect 1994 21907 2004 21963
rect 2060 21907 2128 21963
rect 2184 21907 2252 21963
rect 2308 21907 2376 21963
rect 2432 21907 2442 21963
rect 1994 21839 2442 21907
rect 1994 21783 2004 21839
rect 2060 21783 2128 21839
rect 2184 21783 2252 21839
rect 2308 21783 2376 21839
rect 2432 21783 2442 21839
rect 1994 21715 2442 21783
rect 1994 21659 2004 21715
rect 2060 21659 2128 21715
rect 2184 21659 2252 21715
rect 2308 21659 2376 21715
rect 2432 21659 2442 21715
rect 1994 21591 2442 21659
rect 1994 21535 2004 21591
rect 2060 21535 2128 21591
rect 2184 21535 2252 21591
rect 2308 21535 2376 21591
rect 2432 21535 2442 21591
rect 1994 21467 2442 21535
rect 1994 21411 2004 21467
rect 2060 21411 2128 21467
rect 2184 21411 2252 21467
rect 2308 21411 2376 21467
rect 2432 21411 2442 21467
rect 1994 21343 2442 21411
rect 1994 21287 2004 21343
rect 2060 21287 2128 21343
rect 2184 21287 2252 21343
rect 2308 21287 2376 21343
rect 2432 21287 2442 21343
rect 1994 21219 2442 21287
rect 1994 21163 2004 21219
rect 2060 21163 2128 21219
rect 2184 21163 2252 21219
rect 2308 21163 2376 21219
rect 2432 21163 2442 21219
rect 1994 21095 2442 21163
rect 1994 21039 2004 21095
rect 2060 21039 2128 21095
rect 2184 21039 2252 21095
rect 2308 21039 2376 21095
rect 2432 21039 2442 21095
rect 1994 20971 2442 21039
rect 1994 20915 2004 20971
rect 2060 20915 2128 20971
rect 2184 20915 2252 20971
rect 2308 20915 2376 20971
rect 2432 20915 2442 20971
rect 1994 20847 2442 20915
rect 1994 20791 2004 20847
rect 2060 20791 2128 20847
rect 2184 20791 2252 20847
rect 2308 20791 2376 20847
rect 2432 20791 2442 20847
rect 1994 20723 2442 20791
rect 1994 20667 2004 20723
rect 2060 20667 2128 20723
rect 2184 20667 2252 20723
rect 2308 20667 2376 20723
rect 2432 20667 2442 20723
rect 1994 20599 2442 20667
rect 1994 20543 2004 20599
rect 2060 20543 2128 20599
rect 2184 20543 2252 20599
rect 2308 20543 2376 20599
rect 2432 20543 2442 20599
rect 1994 20533 2442 20543
rect 3698 23451 4146 23461
rect 3698 23395 3708 23451
rect 3764 23395 3832 23451
rect 3888 23395 3956 23451
rect 4012 23395 4080 23451
rect 4136 23395 4146 23451
rect 3698 23327 4146 23395
rect 3698 23271 3708 23327
rect 3764 23271 3832 23327
rect 3888 23271 3956 23327
rect 4012 23271 4080 23327
rect 4136 23271 4146 23327
rect 3698 23203 4146 23271
rect 3698 23147 3708 23203
rect 3764 23147 3832 23203
rect 3888 23147 3956 23203
rect 4012 23147 4080 23203
rect 4136 23147 4146 23203
rect 3698 23079 4146 23147
rect 3698 23023 3708 23079
rect 3764 23023 3832 23079
rect 3888 23023 3956 23079
rect 4012 23023 4080 23079
rect 4136 23023 4146 23079
rect 3698 22955 4146 23023
rect 3698 22899 3708 22955
rect 3764 22899 3832 22955
rect 3888 22899 3956 22955
rect 4012 22899 4080 22955
rect 4136 22899 4146 22955
rect 3698 22831 4146 22899
rect 3698 22775 3708 22831
rect 3764 22775 3832 22831
rect 3888 22775 3956 22831
rect 4012 22775 4080 22831
rect 4136 22775 4146 22831
rect 3698 22707 4146 22775
rect 3698 22651 3708 22707
rect 3764 22651 3832 22707
rect 3888 22651 3956 22707
rect 4012 22651 4080 22707
rect 4136 22651 4146 22707
rect 3698 22583 4146 22651
rect 3698 22527 3708 22583
rect 3764 22527 3832 22583
rect 3888 22527 3956 22583
rect 4012 22527 4080 22583
rect 4136 22527 4146 22583
rect 3698 22459 4146 22527
rect 3698 22403 3708 22459
rect 3764 22403 3832 22459
rect 3888 22403 3956 22459
rect 4012 22403 4080 22459
rect 4136 22403 4146 22459
rect 3698 22335 4146 22403
rect 3698 22279 3708 22335
rect 3764 22279 3832 22335
rect 3888 22279 3956 22335
rect 4012 22279 4080 22335
rect 4136 22279 4146 22335
rect 3698 22211 4146 22279
rect 3698 22155 3708 22211
rect 3764 22155 3832 22211
rect 3888 22155 3956 22211
rect 4012 22155 4080 22211
rect 4136 22155 4146 22211
rect 3698 22087 4146 22155
rect 3698 22031 3708 22087
rect 3764 22031 3832 22087
rect 3888 22031 3956 22087
rect 4012 22031 4080 22087
rect 4136 22031 4146 22087
rect 3698 21963 4146 22031
rect 3698 21907 3708 21963
rect 3764 21907 3832 21963
rect 3888 21907 3956 21963
rect 4012 21907 4080 21963
rect 4136 21907 4146 21963
rect 3698 21839 4146 21907
rect 3698 21783 3708 21839
rect 3764 21783 3832 21839
rect 3888 21783 3956 21839
rect 4012 21783 4080 21839
rect 4136 21783 4146 21839
rect 3698 21715 4146 21783
rect 3698 21659 3708 21715
rect 3764 21659 3832 21715
rect 3888 21659 3956 21715
rect 4012 21659 4080 21715
rect 4136 21659 4146 21715
rect 3698 21591 4146 21659
rect 3698 21535 3708 21591
rect 3764 21535 3832 21591
rect 3888 21535 3956 21591
rect 4012 21535 4080 21591
rect 4136 21535 4146 21591
rect 3698 21467 4146 21535
rect 3698 21411 3708 21467
rect 3764 21411 3832 21467
rect 3888 21411 3956 21467
rect 4012 21411 4080 21467
rect 4136 21411 4146 21467
rect 3698 21343 4146 21411
rect 3698 21287 3708 21343
rect 3764 21287 3832 21343
rect 3888 21287 3956 21343
rect 4012 21287 4080 21343
rect 4136 21287 4146 21343
rect 3698 21219 4146 21287
rect 3698 21163 3708 21219
rect 3764 21163 3832 21219
rect 3888 21163 3956 21219
rect 4012 21163 4080 21219
rect 4136 21163 4146 21219
rect 3698 21095 4146 21163
rect 3698 21039 3708 21095
rect 3764 21039 3832 21095
rect 3888 21039 3956 21095
rect 4012 21039 4080 21095
rect 4136 21039 4146 21095
rect 3698 20971 4146 21039
rect 3698 20915 3708 20971
rect 3764 20915 3832 20971
rect 3888 20915 3956 20971
rect 4012 20915 4080 20971
rect 4136 20915 4146 20971
rect 3698 20847 4146 20915
rect 3698 20791 3708 20847
rect 3764 20791 3832 20847
rect 3888 20791 3956 20847
rect 4012 20791 4080 20847
rect 4136 20791 4146 20847
rect 3698 20723 4146 20791
rect 3698 20667 3708 20723
rect 3764 20667 3832 20723
rect 3888 20667 3956 20723
rect 4012 20667 4080 20723
rect 4136 20667 4146 20723
rect 3698 20599 4146 20667
rect 3698 20543 3708 20599
rect 3764 20543 3832 20599
rect 3888 20543 3956 20599
rect 4012 20543 4080 20599
rect 4136 20543 4146 20599
rect 3698 20533 4146 20543
rect 5970 23451 6418 23461
rect 5970 23395 5980 23451
rect 6036 23395 6104 23451
rect 6160 23395 6228 23451
rect 6284 23395 6352 23451
rect 6408 23395 6418 23451
rect 5970 23327 6418 23395
rect 5970 23271 5980 23327
rect 6036 23271 6104 23327
rect 6160 23271 6228 23327
rect 6284 23271 6352 23327
rect 6408 23271 6418 23327
rect 5970 23203 6418 23271
rect 5970 23147 5980 23203
rect 6036 23147 6104 23203
rect 6160 23147 6228 23203
rect 6284 23147 6352 23203
rect 6408 23147 6418 23203
rect 5970 23079 6418 23147
rect 5970 23023 5980 23079
rect 6036 23023 6104 23079
rect 6160 23023 6228 23079
rect 6284 23023 6352 23079
rect 6408 23023 6418 23079
rect 5970 22955 6418 23023
rect 5970 22899 5980 22955
rect 6036 22899 6104 22955
rect 6160 22899 6228 22955
rect 6284 22899 6352 22955
rect 6408 22899 6418 22955
rect 5970 22831 6418 22899
rect 5970 22775 5980 22831
rect 6036 22775 6104 22831
rect 6160 22775 6228 22831
rect 6284 22775 6352 22831
rect 6408 22775 6418 22831
rect 5970 22707 6418 22775
rect 5970 22651 5980 22707
rect 6036 22651 6104 22707
rect 6160 22651 6228 22707
rect 6284 22651 6352 22707
rect 6408 22651 6418 22707
rect 5970 22583 6418 22651
rect 5970 22527 5980 22583
rect 6036 22527 6104 22583
rect 6160 22527 6228 22583
rect 6284 22527 6352 22583
rect 6408 22527 6418 22583
rect 5970 22459 6418 22527
rect 5970 22403 5980 22459
rect 6036 22403 6104 22459
rect 6160 22403 6228 22459
rect 6284 22403 6352 22459
rect 6408 22403 6418 22459
rect 5970 22335 6418 22403
rect 5970 22279 5980 22335
rect 6036 22279 6104 22335
rect 6160 22279 6228 22335
rect 6284 22279 6352 22335
rect 6408 22279 6418 22335
rect 5970 22211 6418 22279
rect 5970 22155 5980 22211
rect 6036 22155 6104 22211
rect 6160 22155 6228 22211
rect 6284 22155 6352 22211
rect 6408 22155 6418 22211
rect 5970 22087 6418 22155
rect 5970 22031 5980 22087
rect 6036 22031 6104 22087
rect 6160 22031 6228 22087
rect 6284 22031 6352 22087
rect 6408 22031 6418 22087
rect 5970 21963 6418 22031
rect 5970 21907 5980 21963
rect 6036 21907 6104 21963
rect 6160 21907 6228 21963
rect 6284 21907 6352 21963
rect 6408 21907 6418 21963
rect 5970 21839 6418 21907
rect 5970 21783 5980 21839
rect 6036 21783 6104 21839
rect 6160 21783 6228 21839
rect 6284 21783 6352 21839
rect 6408 21783 6418 21839
rect 5970 21715 6418 21783
rect 5970 21659 5980 21715
rect 6036 21659 6104 21715
rect 6160 21659 6228 21715
rect 6284 21659 6352 21715
rect 6408 21659 6418 21715
rect 5970 21591 6418 21659
rect 5970 21535 5980 21591
rect 6036 21535 6104 21591
rect 6160 21535 6228 21591
rect 6284 21535 6352 21591
rect 6408 21535 6418 21591
rect 5970 21467 6418 21535
rect 5970 21411 5980 21467
rect 6036 21411 6104 21467
rect 6160 21411 6228 21467
rect 6284 21411 6352 21467
rect 6408 21411 6418 21467
rect 5970 21343 6418 21411
rect 5970 21287 5980 21343
rect 6036 21287 6104 21343
rect 6160 21287 6228 21343
rect 6284 21287 6352 21343
rect 6408 21287 6418 21343
rect 5970 21219 6418 21287
rect 5970 21163 5980 21219
rect 6036 21163 6104 21219
rect 6160 21163 6228 21219
rect 6284 21163 6352 21219
rect 6408 21163 6418 21219
rect 5970 21095 6418 21163
rect 5970 21039 5980 21095
rect 6036 21039 6104 21095
rect 6160 21039 6228 21095
rect 6284 21039 6352 21095
rect 6408 21039 6418 21095
rect 5970 20971 6418 21039
rect 5970 20915 5980 20971
rect 6036 20915 6104 20971
rect 6160 20915 6228 20971
rect 6284 20915 6352 20971
rect 6408 20915 6418 20971
rect 5970 20847 6418 20915
rect 5970 20791 5980 20847
rect 6036 20791 6104 20847
rect 6160 20791 6228 20847
rect 6284 20791 6352 20847
rect 6408 20791 6418 20847
rect 5970 20723 6418 20791
rect 5970 20667 5980 20723
rect 6036 20667 6104 20723
rect 6160 20667 6228 20723
rect 6284 20667 6352 20723
rect 6408 20667 6418 20723
rect 5970 20599 6418 20667
rect 5970 20543 5980 20599
rect 6036 20543 6104 20599
rect 6160 20543 6228 20599
rect 6284 20543 6352 20599
rect 6408 20543 6418 20599
rect 5970 20533 6418 20543
rect 8646 23451 9094 23461
rect 8646 23395 8656 23451
rect 8712 23395 8780 23451
rect 8836 23395 8904 23451
rect 8960 23395 9028 23451
rect 9084 23395 9094 23451
rect 8646 23327 9094 23395
rect 8646 23271 8656 23327
rect 8712 23271 8780 23327
rect 8836 23271 8904 23327
rect 8960 23271 9028 23327
rect 9084 23271 9094 23327
rect 8646 23203 9094 23271
rect 8646 23147 8656 23203
rect 8712 23147 8780 23203
rect 8836 23147 8904 23203
rect 8960 23147 9028 23203
rect 9084 23147 9094 23203
rect 8646 23079 9094 23147
rect 8646 23023 8656 23079
rect 8712 23023 8780 23079
rect 8836 23023 8904 23079
rect 8960 23023 9028 23079
rect 9084 23023 9094 23079
rect 8646 22955 9094 23023
rect 8646 22899 8656 22955
rect 8712 22899 8780 22955
rect 8836 22899 8904 22955
rect 8960 22899 9028 22955
rect 9084 22899 9094 22955
rect 8646 22831 9094 22899
rect 8646 22775 8656 22831
rect 8712 22775 8780 22831
rect 8836 22775 8904 22831
rect 8960 22775 9028 22831
rect 9084 22775 9094 22831
rect 8646 22707 9094 22775
rect 8646 22651 8656 22707
rect 8712 22651 8780 22707
rect 8836 22651 8904 22707
rect 8960 22651 9028 22707
rect 9084 22651 9094 22707
rect 8646 22583 9094 22651
rect 8646 22527 8656 22583
rect 8712 22527 8780 22583
rect 8836 22527 8904 22583
rect 8960 22527 9028 22583
rect 9084 22527 9094 22583
rect 8646 22459 9094 22527
rect 8646 22403 8656 22459
rect 8712 22403 8780 22459
rect 8836 22403 8904 22459
rect 8960 22403 9028 22459
rect 9084 22403 9094 22459
rect 8646 22335 9094 22403
rect 8646 22279 8656 22335
rect 8712 22279 8780 22335
rect 8836 22279 8904 22335
rect 8960 22279 9028 22335
rect 9084 22279 9094 22335
rect 8646 22211 9094 22279
rect 8646 22155 8656 22211
rect 8712 22155 8780 22211
rect 8836 22155 8904 22211
rect 8960 22155 9028 22211
rect 9084 22155 9094 22211
rect 8646 22087 9094 22155
rect 8646 22031 8656 22087
rect 8712 22031 8780 22087
rect 8836 22031 8904 22087
rect 8960 22031 9028 22087
rect 9084 22031 9094 22087
rect 8646 21963 9094 22031
rect 8646 21907 8656 21963
rect 8712 21907 8780 21963
rect 8836 21907 8904 21963
rect 8960 21907 9028 21963
rect 9084 21907 9094 21963
rect 8646 21839 9094 21907
rect 8646 21783 8656 21839
rect 8712 21783 8780 21839
rect 8836 21783 8904 21839
rect 8960 21783 9028 21839
rect 9084 21783 9094 21839
rect 8646 21715 9094 21783
rect 8646 21659 8656 21715
rect 8712 21659 8780 21715
rect 8836 21659 8904 21715
rect 8960 21659 9028 21715
rect 9084 21659 9094 21715
rect 8646 21591 9094 21659
rect 8646 21535 8656 21591
rect 8712 21535 8780 21591
rect 8836 21535 8904 21591
rect 8960 21535 9028 21591
rect 9084 21535 9094 21591
rect 8646 21467 9094 21535
rect 8646 21411 8656 21467
rect 8712 21411 8780 21467
rect 8836 21411 8904 21467
rect 8960 21411 9028 21467
rect 9084 21411 9094 21467
rect 8646 21343 9094 21411
rect 8646 21287 8656 21343
rect 8712 21287 8780 21343
rect 8836 21287 8904 21343
rect 8960 21287 9028 21343
rect 9084 21287 9094 21343
rect 8646 21219 9094 21287
rect 8646 21163 8656 21219
rect 8712 21163 8780 21219
rect 8836 21163 8904 21219
rect 8960 21163 9028 21219
rect 9084 21163 9094 21219
rect 8646 21095 9094 21163
rect 8646 21039 8656 21095
rect 8712 21039 8780 21095
rect 8836 21039 8904 21095
rect 8960 21039 9028 21095
rect 9084 21039 9094 21095
rect 8646 20971 9094 21039
rect 8646 20915 8656 20971
rect 8712 20915 8780 20971
rect 8836 20915 8904 20971
rect 8960 20915 9028 20971
rect 9084 20915 9094 20971
rect 8646 20847 9094 20915
rect 8646 20791 8656 20847
rect 8712 20791 8780 20847
rect 8836 20791 8904 20847
rect 8960 20791 9028 20847
rect 9084 20791 9094 20847
rect 8646 20723 9094 20791
rect 8646 20667 8656 20723
rect 8712 20667 8780 20723
rect 8836 20667 8904 20723
rect 8960 20667 9028 20723
rect 9084 20667 9094 20723
rect 8646 20599 9094 20667
rect 8646 20543 8656 20599
rect 8712 20543 8780 20599
rect 8836 20543 8904 20599
rect 8960 20543 9028 20599
rect 9084 20543 9094 20599
rect 8646 20533 9094 20543
rect 10918 23451 11366 23461
rect 10918 23395 10928 23451
rect 10984 23395 11052 23451
rect 11108 23395 11176 23451
rect 11232 23395 11300 23451
rect 11356 23395 11366 23451
rect 10918 23327 11366 23395
rect 10918 23271 10928 23327
rect 10984 23271 11052 23327
rect 11108 23271 11176 23327
rect 11232 23271 11300 23327
rect 11356 23271 11366 23327
rect 10918 23203 11366 23271
rect 10918 23147 10928 23203
rect 10984 23147 11052 23203
rect 11108 23147 11176 23203
rect 11232 23147 11300 23203
rect 11356 23147 11366 23203
rect 10918 23079 11366 23147
rect 10918 23023 10928 23079
rect 10984 23023 11052 23079
rect 11108 23023 11176 23079
rect 11232 23023 11300 23079
rect 11356 23023 11366 23079
rect 10918 22955 11366 23023
rect 10918 22899 10928 22955
rect 10984 22899 11052 22955
rect 11108 22899 11176 22955
rect 11232 22899 11300 22955
rect 11356 22899 11366 22955
rect 10918 22831 11366 22899
rect 10918 22775 10928 22831
rect 10984 22775 11052 22831
rect 11108 22775 11176 22831
rect 11232 22775 11300 22831
rect 11356 22775 11366 22831
rect 10918 22707 11366 22775
rect 10918 22651 10928 22707
rect 10984 22651 11052 22707
rect 11108 22651 11176 22707
rect 11232 22651 11300 22707
rect 11356 22651 11366 22707
rect 10918 22583 11366 22651
rect 10918 22527 10928 22583
rect 10984 22527 11052 22583
rect 11108 22527 11176 22583
rect 11232 22527 11300 22583
rect 11356 22527 11366 22583
rect 10918 22459 11366 22527
rect 10918 22403 10928 22459
rect 10984 22403 11052 22459
rect 11108 22403 11176 22459
rect 11232 22403 11300 22459
rect 11356 22403 11366 22459
rect 10918 22335 11366 22403
rect 10918 22279 10928 22335
rect 10984 22279 11052 22335
rect 11108 22279 11176 22335
rect 11232 22279 11300 22335
rect 11356 22279 11366 22335
rect 10918 22211 11366 22279
rect 10918 22155 10928 22211
rect 10984 22155 11052 22211
rect 11108 22155 11176 22211
rect 11232 22155 11300 22211
rect 11356 22155 11366 22211
rect 10918 22087 11366 22155
rect 10918 22031 10928 22087
rect 10984 22031 11052 22087
rect 11108 22031 11176 22087
rect 11232 22031 11300 22087
rect 11356 22031 11366 22087
rect 10918 21963 11366 22031
rect 10918 21907 10928 21963
rect 10984 21907 11052 21963
rect 11108 21907 11176 21963
rect 11232 21907 11300 21963
rect 11356 21907 11366 21963
rect 10918 21839 11366 21907
rect 10918 21783 10928 21839
rect 10984 21783 11052 21839
rect 11108 21783 11176 21839
rect 11232 21783 11300 21839
rect 11356 21783 11366 21839
rect 10918 21715 11366 21783
rect 10918 21659 10928 21715
rect 10984 21659 11052 21715
rect 11108 21659 11176 21715
rect 11232 21659 11300 21715
rect 11356 21659 11366 21715
rect 10918 21591 11366 21659
rect 10918 21535 10928 21591
rect 10984 21535 11052 21591
rect 11108 21535 11176 21591
rect 11232 21535 11300 21591
rect 11356 21535 11366 21591
rect 10918 21467 11366 21535
rect 10918 21411 10928 21467
rect 10984 21411 11052 21467
rect 11108 21411 11176 21467
rect 11232 21411 11300 21467
rect 11356 21411 11366 21467
rect 10918 21343 11366 21411
rect 10918 21287 10928 21343
rect 10984 21287 11052 21343
rect 11108 21287 11176 21343
rect 11232 21287 11300 21343
rect 11356 21287 11366 21343
rect 10918 21219 11366 21287
rect 10918 21163 10928 21219
rect 10984 21163 11052 21219
rect 11108 21163 11176 21219
rect 11232 21163 11300 21219
rect 11356 21163 11366 21219
rect 10918 21095 11366 21163
rect 10918 21039 10928 21095
rect 10984 21039 11052 21095
rect 11108 21039 11176 21095
rect 11232 21039 11300 21095
rect 11356 21039 11366 21095
rect 10918 20971 11366 21039
rect 10918 20915 10928 20971
rect 10984 20915 11052 20971
rect 11108 20915 11176 20971
rect 11232 20915 11300 20971
rect 11356 20915 11366 20971
rect 10918 20847 11366 20915
rect 10918 20791 10928 20847
rect 10984 20791 11052 20847
rect 11108 20791 11176 20847
rect 11232 20791 11300 20847
rect 11356 20791 11366 20847
rect 10918 20723 11366 20791
rect 10918 20667 10928 20723
rect 10984 20667 11052 20723
rect 11108 20667 11176 20723
rect 11232 20667 11300 20723
rect 11356 20667 11366 20723
rect 10918 20599 11366 20667
rect 10918 20543 10928 20599
rect 10984 20543 11052 20599
rect 11108 20543 11176 20599
rect 11232 20543 11300 20599
rect 11356 20543 11366 20599
rect 10918 20533 11366 20543
rect 12622 23451 13070 23461
rect 12622 23395 12632 23451
rect 12688 23395 12756 23451
rect 12812 23395 12880 23451
rect 12936 23395 13004 23451
rect 13060 23395 13070 23451
rect 12622 23327 13070 23395
rect 12622 23271 12632 23327
rect 12688 23271 12756 23327
rect 12812 23271 12880 23327
rect 12936 23271 13004 23327
rect 13060 23271 13070 23327
rect 12622 23203 13070 23271
rect 12622 23147 12632 23203
rect 12688 23147 12756 23203
rect 12812 23147 12880 23203
rect 12936 23147 13004 23203
rect 13060 23147 13070 23203
rect 12622 23079 13070 23147
rect 12622 23023 12632 23079
rect 12688 23023 12756 23079
rect 12812 23023 12880 23079
rect 12936 23023 13004 23079
rect 13060 23023 13070 23079
rect 12622 22955 13070 23023
rect 12622 22899 12632 22955
rect 12688 22899 12756 22955
rect 12812 22899 12880 22955
rect 12936 22899 13004 22955
rect 13060 22899 13070 22955
rect 12622 22831 13070 22899
rect 12622 22775 12632 22831
rect 12688 22775 12756 22831
rect 12812 22775 12880 22831
rect 12936 22775 13004 22831
rect 13060 22775 13070 22831
rect 12622 22707 13070 22775
rect 12622 22651 12632 22707
rect 12688 22651 12756 22707
rect 12812 22651 12880 22707
rect 12936 22651 13004 22707
rect 13060 22651 13070 22707
rect 12622 22583 13070 22651
rect 12622 22527 12632 22583
rect 12688 22527 12756 22583
rect 12812 22527 12880 22583
rect 12936 22527 13004 22583
rect 13060 22527 13070 22583
rect 12622 22459 13070 22527
rect 12622 22403 12632 22459
rect 12688 22403 12756 22459
rect 12812 22403 12880 22459
rect 12936 22403 13004 22459
rect 13060 22403 13070 22459
rect 12622 22335 13070 22403
rect 12622 22279 12632 22335
rect 12688 22279 12756 22335
rect 12812 22279 12880 22335
rect 12936 22279 13004 22335
rect 13060 22279 13070 22335
rect 12622 22211 13070 22279
rect 12622 22155 12632 22211
rect 12688 22155 12756 22211
rect 12812 22155 12880 22211
rect 12936 22155 13004 22211
rect 13060 22155 13070 22211
rect 12622 22087 13070 22155
rect 12622 22031 12632 22087
rect 12688 22031 12756 22087
rect 12812 22031 12880 22087
rect 12936 22031 13004 22087
rect 13060 22031 13070 22087
rect 12622 21963 13070 22031
rect 12622 21907 12632 21963
rect 12688 21907 12756 21963
rect 12812 21907 12880 21963
rect 12936 21907 13004 21963
rect 13060 21907 13070 21963
rect 12622 21839 13070 21907
rect 12622 21783 12632 21839
rect 12688 21783 12756 21839
rect 12812 21783 12880 21839
rect 12936 21783 13004 21839
rect 13060 21783 13070 21839
rect 12622 21715 13070 21783
rect 12622 21659 12632 21715
rect 12688 21659 12756 21715
rect 12812 21659 12880 21715
rect 12936 21659 13004 21715
rect 13060 21659 13070 21715
rect 12622 21591 13070 21659
rect 12622 21535 12632 21591
rect 12688 21535 12756 21591
rect 12812 21535 12880 21591
rect 12936 21535 13004 21591
rect 13060 21535 13070 21591
rect 12622 21467 13070 21535
rect 12622 21411 12632 21467
rect 12688 21411 12756 21467
rect 12812 21411 12880 21467
rect 12936 21411 13004 21467
rect 13060 21411 13070 21467
rect 12622 21343 13070 21411
rect 12622 21287 12632 21343
rect 12688 21287 12756 21343
rect 12812 21287 12880 21343
rect 12936 21287 13004 21343
rect 13060 21287 13070 21343
rect 12622 21219 13070 21287
rect 12622 21163 12632 21219
rect 12688 21163 12756 21219
rect 12812 21163 12880 21219
rect 12936 21163 13004 21219
rect 13060 21163 13070 21219
rect 12622 21095 13070 21163
rect 12622 21039 12632 21095
rect 12688 21039 12756 21095
rect 12812 21039 12880 21095
rect 12936 21039 13004 21095
rect 13060 21039 13070 21095
rect 12622 20971 13070 21039
rect 12622 20915 12632 20971
rect 12688 20915 12756 20971
rect 12812 20915 12880 20971
rect 12936 20915 13004 20971
rect 13060 20915 13070 20971
rect 12622 20847 13070 20915
rect 12622 20791 12632 20847
rect 12688 20791 12756 20847
rect 12812 20791 12880 20847
rect 12936 20791 13004 20847
rect 13060 20791 13070 20847
rect 12622 20723 13070 20791
rect 12622 20667 12632 20723
rect 12688 20667 12756 20723
rect 12812 20667 12880 20723
rect 12936 20667 13004 20723
rect 13060 20667 13070 20723
rect 12622 20599 13070 20667
rect 12622 20543 12632 20599
rect 12688 20543 12756 20599
rect 12812 20543 12880 20599
rect 12936 20543 13004 20599
rect 13060 20543 13070 20599
rect 12622 20533 13070 20543
rect 13758 23451 14206 23461
rect 13758 23395 13768 23451
rect 13824 23395 13892 23451
rect 13948 23395 14016 23451
rect 14072 23395 14140 23451
rect 14196 23395 14206 23451
rect 13758 23327 14206 23395
rect 13758 23271 13768 23327
rect 13824 23271 13892 23327
rect 13948 23271 14016 23327
rect 14072 23271 14140 23327
rect 14196 23271 14206 23327
rect 13758 23203 14206 23271
rect 13758 23147 13768 23203
rect 13824 23147 13892 23203
rect 13948 23147 14016 23203
rect 14072 23147 14140 23203
rect 14196 23147 14206 23203
rect 13758 23079 14206 23147
rect 13758 23023 13768 23079
rect 13824 23023 13892 23079
rect 13948 23023 14016 23079
rect 14072 23023 14140 23079
rect 14196 23023 14206 23079
rect 13758 22955 14206 23023
rect 13758 22899 13768 22955
rect 13824 22899 13892 22955
rect 13948 22899 14016 22955
rect 14072 22899 14140 22955
rect 14196 22899 14206 22955
rect 13758 22831 14206 22899
rect 13758 22775 13768 22831
rect 13824 22775 13892 22831
rect 13948 22775 14016 22831
rect 14072 22775 14140 22831
rect 14196 22775 14206 22831
rect 13758 22707 14206 22775
rect 13758 22651 13768 22707
rect 13824 22651 13892 22707
rect 13948 22651 14016 22707
rect 14072 22651 14140 22707
rect 14196 22651 14206 22707
rect 13758 22583 14206 22651
rect 13758 22527 13768 22583
rect 13824 22527 13892 22583
rect 13948 22527 14016 22583
rect 14072 22527 14140 22583
rect 14196 22527 14206 22583
rect 13758 22459 14206 22527
rect 13758 22403 13768 22459
rect 13824 22403 13892 22459
rect 13948 22403 14016 22459
rect 14072 22403 14140 22459
rect 14196 22403 14206 22459
rect 13758 22335 14206 22403
rect 13758 22279 13768 22335
rect 13824 22279 13892 22335
rect 13948 22279 14016 22335
rect 14072 22279 14140 22335
rect 14196 22279 14206 22335
rect 13758 22211 14206 22279
rect 13758 22155 13768 22211
rect 13824 22155 13892 22211
rect 13948 22155 14016 22211
rect 14072 22155 14140 22211
rect 14196 22155 14206 22211
rect 13758 22087 14206 22155
rect 13758 22031 13768 22087
rect 13824 22031 13892 22087
rect 13948 22031 14016 22087
rect 14072 22031 14140 22087
rect 14196 22031 14206 22087
rect 13758 21963 14206 22031
rect 13758 21907 13768 21963
rect 13824 21907 13892 21963
rect 13948 21907 14016 21963
rect 14072 21907 14140 21963
rect 14196 21907 14206 21963
rect 13758 21839 14206 21907
rect 13758 21783 13768 21839
rect 13824 21783 13892 21839
rect 13948 21783 14016 21839
rect 14072 21783 14140 21839
rect 14196 21783 14206 21839
rect 13758 21715 14206 21783
rect 13758 21659 13768 21715
rect 13824 21659 13892 21715
rect 13948 21659 14016 21715
rect 14072 21659 14140 21715
rect 14196 21659 14206 21715
rect 13758 21591 14206 21659
rect 13758 21535 13768 21591
rect 13824 21535 13892 21591
rect 13948 21535 14016 21591
rect 14072 21535 14140 21591
rect 14196 21535 14206 21591
rect 13758 21467 14206 21535
rect 13758 21411 13768 21467
rect 13824 21411 13892 21467
rect 13948 21411 14016 21467
rect 14072 21411 14140 21467
rect 14196 21411 14206 21467
rect 13758 21343 14206 21411
rect 13758 21287 13768 21343
rect 13824 21287 13892 21343
rect 13948 21287 14016 21343
rect 14072 21287 14140 21343
rect 14196 21287 14206 21343
rect 13758 21219 14206 21287
rect 13758 21163 13768 21219
rect 13824 21163 13892 21219
rect 13948 21163 14016 21219
rect 14072 21163 14140 21219
rect 14196 21163 14206 21219
rect 13758 21095 14206 21163
rect 13758 21039 13768 21095
rect 13824 21039 13892 21095
rect 13948 21039 14016 21095
rect 14072 21039 14140 21095
rect 14196 21039 14206 21095
rect 13758 20971 14206 21039
rect 13758 20915 13768 20971
rect 13824 20915 13892 20971
rect 13948 20915 14016 20971
rect 14072 20915 14140 20971
rect 14196 20915 14206 20971
rect 13758 20847 14206 20915
rect 13758 20791 13768 20847
rect 13824 20791 13892 20847
rect 13948 20791 14016 20847
rect 14072 20791 14140 20847
rect 14196 20791 14206 20847
rect 13758 20723 14206 20791
rect 13758 20667 13768 20723
rect 13824 20667 13892 20723
rect 13948 20667 14016 20723
rect 14072 20667 14140 20723
rect 14196 20667 14206 20723
rect 13758 20599 14206 20667
rect 13758 20543 13768 20599
rect 13824 20543 13892 20599
rect 13948 20543 14016 20599
rect 14072 20543 14140 20599
rect 14196 20543 14206 20599
rect 13758 20533 14206 20543
rect 858 20251 1306 20261
rect 858 20195 868 20251
rect 924 20195 992 20251
rect 1048 20195 1116 20251
rect 1172 20195 1240 20251
rect 1296 20195 1306 20251
rect 858 20127 1306 20195
rect 858 20071 868 20127
rect 924 20071 992 20127
rect 1048 20071 1116 20127
rect 1172 20071 1240 20127
rect 1296 20071 1306 20127
rect 858 20003 1306 20071
rect 858 19947 868 20003
rect 924 19947 992 20003
rect 1048 19947 1116 20003
rect 1172 19947 1240 20003
rect 1296 19947 1306 20003
rect 858 19879 1306 19947
rect 858 19823 868 19879
rect 924 19823 992 19879
rect 1048 19823 1116 19879
rect 1172 19823 1240 19879
rect 1296 19823 1306 19879
rect 858 19755 1306 19823
rect 858 19699 868 19755
rect 924 19699 992 19755
rect 1048 19699 1116 19755
rect 1172 19699 1240 19755
rect 1296 19699 1306 19755
rect 858 19631 1306 19699
rect 858 19575 868 19631
rect 924 19575 992 19631
rect 1048 19575 1116 19631
rect 1172 19575 1240 19631
rect 1296 19575 1306 19631
rect 858 19507 1306 19575
rect 858 19451 868 19507
rect 924 19451 992 19507
rect 1048 19451 1116 19507
rect 1172 19451 1240 19507
rect 1296 19451 1306 19507
rect 858 19383 1306 19451
rect 858 19327 868 19383
rect 924 19327 992 19383
rect 1048 19327 1116 19383
rect 1172 19327 1240 19383
rect 1296 19327 1306 19383
rect 858 19259 1306 19327
rect 858 19203 868 19259
rect 924 19203 992 19259
rect 1048 19203 1116 19259
rect 1172 19203 1240 19259
rect 1296 19203 1306 19259
rect 858 19135 1306 19203
rect 858 19079 868 19135
rect 924 19079 992 19135
rect 1048 19079 1116 19135
rect 1172 19079 1240 19135
rect 1296 19079 1306 19135
rect 858 19011 1306 19079
rect 858 18955 868 19011
rect 924 18955 992 19011
rect 1048 18955 1116 19011
rect 1172 18955 1240 19011
rect 1296 18955 1306 19011
rect 858 18887 1306 18955
rect 858 18831 868 18887
rect 924 18831 992 18887
rect 1048 18831 1116 18887
rect 1172 18831 1240 18887
rect 1296 18831 1306 18887
rect 858 18763 1306 18831
rect 858 18707 868 18763
rect 924 18707 992 18763
rect 1048 18707 1116 18763
rect 1172 18707 1240 18763
rect 1296 18707 1306 18763
rect 858 18639 1306 18707
rect 858 18583 868 18639
rect 924 18583 992 18639
rect 1048 18583 1116 18639
rect 1172 18583 1240 18639
rect 1296 18583 1306 18639
rect 858 18515 1306 18583
rect 858 18459 868 18515
rect 924 18459 992 18515
rect 1048 18459 1116 18515
rect 1172 18459 1240 18515
rect 1296 18459 1306 18515
rect 858 18391 1306 18459
rect 858 18335 868 18391
rect 924 18335 992 18391
rect 1048 18335 1116 18391
rect 1172 18335 1240 18391
rect 1296 18335 1306 18391
rect 858 18267 1306 18335
rect 858 18211 868 18267
rect 924 18211 992 18267
rect 1048 18211 1116 18267
rect 1172 18211 1240 18267
rect 1296 18211 1306 18267
rect 858 18143 1306 18211
rect 858 18087 868 18143
rect 924 18087 992 18143
rect 1048 18087 1116 18143
rect 1172 18087 1240 18143
rect 1296 18087 1306 18143
rect 858 18019 1306 18087
rect 858 17963 868 18019
rect 924 17963 992 18019
rect 1048 17963 1116 18019
rect 1172 17963 1240 18019
rect 1296 17963 1306 18019
rect 858 17895 1306 17963
rect 858 17839 868 17895
rect 924 17839 992 17895
rect 1048 17839 1116 17895
rect 1172 17839 1240 17895
rect 1296 17839 1306 17895
rect 858 17771 1306 17839
rect 858 17715 868 17771
rect 924 17715 992 17771
rect 1048 17715 1116 17771
rect 1172 17715 1240 17771
rect 1296 17715 1306 17771
rect 858 17647 1306 17715
rect 858 17591 868 17647
rect 924 17591 992 17647
rect 1048 17591 1116 17647
rect 1172 17591 1240 17647
rect 1296 17591 1306 17647
rect 858 17523 1306 17591
rect 858 17467 868 17523
rect 924 17467 992 17523
rect 1048 17467 1116 17523
rect 1172 17467 1240 17523
rect 1296 17467 1306 17523
rect 858 17399 1306 17467
rect 858 17343 868 17399
rect 924 17343 992 17399
rect 1048 17343 1116 17399
rect 1172 17343 1240 17399
rect 1296 17343 1306 17399
rect 858 17333 1306 17343
rect 1994 20251 2442 20261
rect 1994 20195 2004 20251
rect 2060 20195 2128 20251
rect 2184 20195 2252 20251
rect 2308 20195 2376 20251
rect 2432 20195 2442 20251
rect 1994 20127 2442 20195
rect 1994 20071 2004 20127
rect 2060 20071 2128 20127
rect 2184 20071 2252 20127
rect 2308 20071 2376 20127
rect 2432 20071 2442 20127
rect 1994 20003 2442 20071
rect 1994 19947 2004 20003
rect 2060 19947 2128 20003
rect 2184 19947 2252 20003
rect 2308 19947 2376 20003
rect 2432 19947 2442 20003
rect 1994 19879 2442 19947
rect 1994 19823 2004 19879
rect 2060 19823 2128 19879
rect 2184 19823 2252 19879
rect 2308 19823 2376 19879
rect 2432 19823 2442 19879
rect 1994 19755 2442 19823
rect 1994 19699 2004 19755
rect 2060 19699 2128 19755
rect 2184 19699 2252 19755
rect 2308 19699 2376 19755
rect 2432 19699 2442 19755
rect 1994 19631 2442 19699
rect 1994 19575 2004 19631
rect 2060 19575 2128 19631
rect 2184 19575 2252 19631
rect 2308 19575 2376 19631
rect 2432 19575 2442 19631
rect 1994 19507 2442 19575
rect 1994 19451 2004 19507
rect 2060 19451 2128 19507
rect 2184 19451 2252 19507
rect 2308 19451 2376 19507
rect 2432 19451 2442 19507
rect 1994 19383 2442 19451
rect 1994 19327 2004 19383
rect 2060 19327 2128 19383
rect 2184 19327 2252 19383
rect 2308 19327 2376 19383
rect 2432 19327 2442 19383
rect 1994 19259 2442 19327
rect 1994 19203 2004 19259
rect 2060 19203 2128 19259
rect 2184 19203 2252 19259
rect 2308 19203 2376 19259
rect 2432 19203 2442 19259
rect 1994 19135 2442 19203
rect 1994 19079 2004 19135
rect 2060 19079 2128 19135
rect 2184 19079 2252 19135
rect 2308 19079 2376 19135
rect 2432 19079 2442 19135
rect 1994 19011 2442 19079
rect 1994 18955 2004 19011
rect 2060 18955 2128 19011
rect 2184 18955 2252 19011
rect 2308 18955 2376 19011
rect 2432 18955 2442 19011
rect 1994 18887 2442 18955
rect 1994 18831 2004 18887
rect 2060 18831 2128 18887
rect 2184 18831 2252 18887
rect 2308 18831 2376 18887
rect 2432 18831 2442 18887
rect 1994 18763 2442 18831
rect 1994 18707 2004 18763
rect 2060 18707 2128 18763
rect 2184 18707 2252 18763
rect 2308 18707 2376 18763
rect 2432 18707 2442 18763
rect 1994 18639 2442 18707
rect 1994 18583 2004 18639
rect 2060 18583 2128 18639
rect 2184 18583 2252 18639
rect 2308 18583 2376 18639
rect 2432 18583 2442 18639
rect 1994 18515 2442 18583
rect 1994 18459 2004 18515
rect 2060 18459 2128 18515
rect 2184 18459 2252 18515
rect 2308 18459 2376 18515
rect 2432 18459 2442 18515
rect 1994 18391 2442 18459
rect 1994 18335 2004 18391
rect 2060 18335 2128 18391
rect 2184 18335 2252 18391
rect 2308 18335 2376 18391
rect 2432 18335 2442 18391
rect 1994 18267 2442 18335
rect 1994 18211 2004 18267
rect 2060 18211 2128 18267
rect 2184 18211 2252 18267
rect 2308 18211 2376 18267
rect 2432 18211 2442 18267
rect 1994 18143 2442 18211
rect 1994 18087 2004 18143
rect 2060 18087 2128 18143
rect 2184 18087 2252 18143
rect 2308 18087 2376 18143
rect 2432 18087 2442 18143
rect 1994 18019 2442 18087
rect 1994 17963 2004 18019
rect 2060 17963 2128 18019
rect 2184 17963 2252 18019
rect 2308 17963 2376 18019
rect 2432 17963 2442 18019
rect 1994 17895 2442 17963
rect 1994 17839 2004 17895
rect 2060 17839 2128 17895
rect 2184 17839 2252 17895
rect 2308 17839 2376 17895
rect 2432 17839 2442 17895
rect 1994 17771 2442 17839
rect 1994 17715 2004 17771
rect 2060 17715 2128 17771
rect 2184 17715 2252 17771
rect 2308 17715 2376 17771
rect 2432 17715 2442 17771
rect 1994 17647 2442 17715
rect 1994 17591 2004 17647
rect 2060 17591 2128 17647
rect 2184 17591 2252 17647
rect 2308 17591 2376 17647
rect 2432 17591 2442 17647
rect 1994 17523 2442 17591
rect 1994 17467 2004 17523
rect 2060 17467 2128 17523
rect 2184 17467 2252 17523
rect 2308 17467 2376 17523
rect 2432 17467 2442 17523
rect 1994 17399 2442 17467
rect 1994 17343 2004 17399
rect 2060 17343 2128 17399
rect 2184 17343 2252 17399
rect 2308 17343 2376 17399
rect 2432 17343 2442 17399
rect 1994 17333 2442 17343
rect 3698 20251 4146 20261
rect 3698 20195 3708 20251
rect 3764 20195 3832 20251
rect 3888 20195 3956 20251
rect 4012 20195 4080 20251
rect 4136 20195 4146 20251
rect 3698 20127 4146 20195
rect 3698 20071 3708 20127
rect 3764 20071 3832 20127
rect 3888 20071 3956 20127
rect 4012 20071 4080 20127
rect 4136 20071 4146 20127
rect 3698 20003 4146 20071
rect 3698 19947 3708 20003
rect 3764 19947 3832 20003
rect 3888 19947 3956 20003
rect 4012 19947 4080 20003
rect 4136 19947 4146 20003
rect 3698 19879 4146 19947
rect 3698 19823 3708 19879
rect 3764 19823 3832 19879
rect 3888 19823 3956 19879
rect 4012 19823 4080 19879
rect 4136 19823 4146 19879
rect 3698 19755 4146 19823
rect 3698 19699 3708 19755
rect 3764 19699 3832 19755
rect 3888 19699 3956 19755
rect 4012 19699 4080 19755
rect 4136 19699 4146 19755
rect 3698 19631 4146 19699
rect 3698 19575 3708 19631
rect 3764 19575 3832 19631
rect 3888 19575 3956 19631
rect 4012 19575 4080 19631
rect 4136 19575 4146 19631
rect 3698 19507 4146 19575
rect 3698 19451 3708 19507
rect 3764 19451 3832 19507
rect 3888 19451 3956 19507
rect 4012 19451 4080 19507
rect 4136 19451 4146 19507
rect 3698 19383 4146 19451
rect 3698 19327 3708 19383
rect 3764 19327 3832 19383
rect 3888 19327 3956 19383
rect 4012 19327 4080 19383
rect 4136 19327 4146 19383
rect 3698 19259 4146 19327
rect 3698 19203 3708 19259
rect 3764 19203 3832 19259
rect 3888 19203 3956 19259
rect 4012 19203 4080 19259
rect 4136 19203 4146 19259
rect 3698 19135 4146 19203
rect 3698 19079 3708 19135
rect 3764 19079 3832 19135
rect 3888 19079 3956 19135
rect 4012 19079 4080 19135
rect 4136 19079 4146 19135
rect 3698 19011 4146 19079
rect 3698 18955 3708 19011
rect 3764 18955 3832 19011
rect 3888 18955 3956 19011
rect 4012 18955 4080 19011
rect 4136 18955 4146 19011
rect 3698 18887 4146 18955
rect 3698 18831 3708 18887
rect 3764 18831 3832 18887
rect 3888 18831 3956 18887
rect 4012 18831 4080 18887
rect 4136 18831 4146 18887
rect 3698 18763 4146 18831
rect 3698 18707 3708 18763
rect 3764 18707 3832 18763
rect 3888 18707 3956 18763
rect 4012 18707 4080 18763
rect 4136 18707 4146 18763
rect 3698 18639 4146 18707
rect 3698 18583 3708 18639
rect 3764 18583 3832 18639
rect 3888 18583 3956 18639
rect 4012 18583 4080 18639
rect 4136 18583 4146 18639
rect 3698 18515 4146 18583
rect 3698 18459 3708 18515
rect 3764 18459 3832 18515
rect 3888 18459 3956 18515
rect 4012 18459 4080 18515
rect 4136 18459 4146 18515
rect 3698 18391 4146 18459
rect 3698 18335 3708 18391
rect 3764 18335 3832 18391
rect 3888 18335 3956 18391
rect 4012 18335 4080 18391
rect 4136 18335 4146 18391
rect 3698 18267 4146 18335
rect 3698 18211 3708 18267
rect 3764 18211 3832 18267
rect 3888 18211 3956 18267
rect 4012 18211 4080 18267
rect 4136 18211 4146 18267
rect 3698 18143 4146 18211
rect 3698 18087 3708 18143
rect 3764 18087 3832 18143
rect 3888 18087 3956 18143
rect 4012 18087 4080 18143
rect 4136 18087 4146 18143
rect 3698 18019 4146 18087
rect 3698 17963 3708 18019
rect 3764 17963 3832 18019
rect 3888 17963 3956 18019
rect 4012 17963 4080 18019
rect 4136 17963 4146 18019
rect 3698 17895 4146 17963
rect 3698 17839 3708 17895
rect 3764 17839 3832 17895
rect 3888 17839 3956 17895
rect 4012 17839 4080 17895
rect 4136 17839 4146 17895
rect 3698 17771 4146 17839
rect 3698 17715 3708 17771
rect 3764 17715 3832 17771
rect 3888 17715 3956 17771
rect 4012 17715 4080 17771
rect 4136 17715 4146 17771
rect 3698 17647 4146 17715
rect 3698 17591 3708 17647
rect 3764 17591 3832 17647
rect 3888 17591 3956 17647
rect 4012 17591 4080 17647
rect 4136 17591 4146 17647
rect 3698 17523 4146 17591
rect 3698 17467 3708 17523
rect 3764 17467 3832 17523
rect 3888 17467 3956 17523
rect 4012 17467 4080 17523
rect 4136 17467 4146 17523
rect 3698 17399 4146 17467
rect 3698 17343 3708 17399
rect 3764 17343 3832 17399
rect 3888 17343 3956 17399
rect 4012 17343 4080 17399
rect 4136 17343 4146 17399
rect 3698 17333 4146 17343
rect 5970 20251 6418 20261
rect 5970 20195 5980 20251
rect 6036 20195 6104 20251
rect 6160 20195 6228 20251
rect 6284 20195 6352 20251
rect 6408 20195 6418 20251
rect 5970 20127 6418 20195
rect 5970 20071 5980 20127
rect 6036 20071 6104 20127
rect 6160 20071 6228 20127
rect 6284 20071 6352 20127
rect 6408 20071 6418 20127
rect 5970 20003 6418 20071
rect 5970 19947 5980 20003
rect 6036 19947 6104 20003
rect 6160 19947 6228 20003
rect 6284 19947 6352 20003
rect 6408 19947 6418 20003
rect 5970 19879 6418 19947
rect 5970 19823 5980 19879
rect 6036 19823 6104 19879
rect 6160 19823 6228 19879
rect 6284 19823 6352 19879
rect 6408 19823 6418 19879
rect 5970 19755 6418 19823
rect 5970 19699 5980 19755
rect 6036 19699 6104 19755
rect 6160 19699 6228 19755
rect 6284 19699 6352 19755
rect 6408 19699 6418 19755
rect 5970 19631 6418 19699
rect 5970 19575 5980 19631
rect 6036 19575 6104 19631
rect 6160 19575 6228 19631
rect 6284 19575 6352 19631
rect 6408 19575 6418 19631
rect 5970 19507 6418 19575
rect 5970 19451 5980 19507
rect 6036 19451 6104 19507
rect 6160 19451 6228 19507
rect 6284 19451 6352 19507
rect 6408 19451 6418 19507
rect 5970 19383 6418 19451
rect 5970 19327 5980 19383
rect 6036 19327 6104 19383
rect 6160 19327 6228 19383
rect 6284 19327 6352 19383
rect 6408 19327 6418 19383
rect 5970 19259 6418 19327
rect 5970 19203 5980 19259
rect 6036 19203 6104 19259
rect 6160 19203 6228 19259
rect 6284 19203 6352 19259
rect 6408 19203 6418 19259
rect 5970 19135 6418 19203
rect 5970 19079 5980 19135
rect 6036 19079 6104 19135
rect 6160 19079 6228 19135
rect 6284 19079 6352 19135
rect 6408 19079 6418 19135
rect 5970 19011 6418 19079
rect 5970 18955 5980 19011
rect 6036 18955 6104 19011
rect 6160 18955 6228 19011
rect 6284 18955 6352 19011
rect 6408 18955 6418 19011
rect 5970 18887 6418 18955
rect 5970 18831 5980 18887
rect 6036 18831 6104 18887
rect 6160 18831 6228 18887
rect 6284 18831 6352 18887
rect 6408 18831 6418 18887
rect 5970 18763 6418 18831
rect 5970 18707 5980 18763
rect 6036 18707 6104 18763
rect 6160 18707 6228 18763
rect 6284 18707 6352 18763
rect 6408 18707 6418 18763
rect 5970 18639 6418 18707
rect 5970 18583 5980 18639
rect 6036 18583 6104 18639
rect 6160 18583 6228 18639
rect 6284 18583 6352 18639
rect 6408 18583 6418 18639
rect 5970 18515 6418 18583
rect 5970 18459 5980 18515
rect 6036 18459 6104 18515
rect 6160 18459 6228 18515
rect 6284 18459 6352 18515
rect 6408 18459 6418 18515
rect 5970 18391 6418 18459
rect 5970 18335 5980 18391
rect 6036 18335 6104 18391
rect 6160 18335 6228 18391
rect 6284 18335 6352 18391
rect 6408 18335 6418 18391
rect 5970 18267 6418 18335
rect 5970 18211 5980 18267
rect 6036 18211 6104 18267
rect 6160 18211 6228 18267
rect 6284 18211 6352 18267
rect 6408 18211 6418 18267
rect 5970 18143 6418 18211
rect 5970 18087 5980 18143
rect 6036 18087 6104 18143
rect 6160 18087 6228 18143
rect 6284 18087 6352 18143
rect 6408 18087 6418 18143
rect 5970 18019 6418 18087
rect 5970 17963 5980 18019
rect 6036 17963 6104 18019
rect 6160 17963 6228 18019
rect 6284 17963 6352 18019
rect 6408 17963 6418 18019
rect 5970 17895 6418 17963
rect 5970 17839 5980 17895
rect 6036 17839 6104 17895
rect 6160 17839 6228 17895
rect 6284 17839 6352 17895
rect 6408 17839 6418 17895
rect 5970 17771 6418 17839
rect 5970 17715 5980 17771
rect 6036 17715 6104 17771
rect 6160 17715 6228 17771
rect 6284 17715 6352 17771
rect 6408 17715 6418 17771
rect 5970 17647 6418 17715
rect 5970 17591 5980 17647
rect 6036 17591 6104 17647
rect 6160 17591 6228 17647
rect 6284 17591 6352 17647
rect 6408 17591 6418 17647
rect 5970 17523 6418 17591
rect 5970 17467 5980 17523
rect 6036 17467 6104 17523
rect 6160 17467 6228 17523
rect 6284 17467 6352 17523
rect 6408 17467 6418 17523
rect 5970 17399 6418 17467
rect 5970 17343 5980 17399
rect 6036 17343 6104 17399
rect 6160 17343 6228 17399
rect 6284 17343 6352 17399
rect 6408 17343 6418 17399
rect 5970 17333 6418 17343
rect 8646 20251 9094 20261
rect 8646 20195 8656 20251
rect 8712 20195 8780 20251
rect 8836 20195 8904 20251
rect 8960 20195 9028 20251
rect 9084 20195 9094 20251
rect 8646 20127 9094 20195
rect 8646 20071 8656 20127
rect 8712 20071 8780 20127
rect 8836 20071 8904 20127
rect 8960 20071 9028 20127
rect 9084 20071 9094 20127
rect 8646 20003 9094 20071
rect 8646 19947 8656 20003
rect 8712 19947 8780 20003
rect 8836 19947 8904 20003
rect 8960 19947 9028 20003
rect 9084 19947 9094 20003
rect 8646 19879 9094 19947
rect 8646 19823 8656 19879
rect 8712 19823 8780 19879
rect 8836 19823 8904 19879
rect 8960 19823 9028 19879
rect 9084 19823 9094 19879
rect 8646 19755 9094 19823
rect 8646 19699 8656 19755
rect 8712 19699 8780 19755
rect 8836 19699 8904 19755
rect 8960 19699 9028 19755
rect 9084 19699 9094 19755
rect 8646 19631 9094 19699
rect 8646 19575 8656 19631
rect 8712 19575 8780 19631
rect 8836 19575 8904 19631
rect 8960 19575 9028 19631
rect 9084 19575 9094 19631
rect 8646 19507 9094 19575
rect 8646 19451 8656 19507
rect 8712 19451 8780 19507
rect 8836 19451 8904 19507
rect 8960 19451 9028 19507
rect 9084 19451 9094 19507
rect 8646 19383 9094 19451
rect 8646 19327 8656 19383
rect 8712 19327 8780 19383
rect 8836 19327 8904 19383
rect 8960 19327 9028 19383
rect 9084 19327 9094 19383
rect 8646 19259 9094 19327
rect 8646 19203 8656 19259
rect 8712 19203 8780 19259
rect 8836 19203 8904 19259
rect 8960 19203 9028 19259
rect 9084 19203 9094 19259
rect 8646 19135 9094 19203
rect 8646 19079 8656 19135
rect 8712 19079 8780 19135
rect 8836 19079 8904 19135
rect 8960 19079 9028 19135
rect 9084 19079 9094 19135
rect 8646 19011 9094 19079
rect 8646 18955 8656 19011
rect 8712 18955 8780 19011
rect 8836 18955 8904 19011
rect 8960 18955 9028 19011
rect 9084 18955 9094 19011
rect 8646 18887 9094 18955
rect 8646 18831 8656 18887
rect 8712 18831 8780 18887
rect 8836 18831 8904 18887
rect 8960 18831 9028 18887
rect 9084 18831 9094 18887
rect 8646 18763 9094 18831
rect 8646 18707 8656 18763
rect 8712 18707 8780 18763
rect 8836 18707 8904 18763
rect 8960 18707 9028 18763
rect 9084 18707 9094 18763
rect 8646 18639 9094 18707
rect 8646 18583 8656 18639
rect 8712 18583 8780 18639
rect 8836 18583 8904 18639
rect 8960 18583 9028 18639
rect 9084 18583 9094 18639
rect 8646 18515 9094 18583
rect 8646 18459 8656 18515
rect 8712 18459 8780 18515
rect 8836 18459 8904 18515
rect 8960 18459 9028 18515
rect 9084 18459 9094 18515
rect 8646 18391 9094 18459
rect 8646 18335 8656 18391
rect 8712 18335 8780 18391
rect 8836 18335 8904 18391
rect 8960 18335 9028 18391
rect 9084 18335 9094 18391
rect 8646 18267 9094 18335
rect 8646 18211 8656 18267
rect 8712 18211 8780 18267
rect 8836 18211 8904 18267
rect 8960 18211 9028 18267
rect 9084 18211 9094 18267
rect 8646 18143 9094 18211
rect 8646 18087 8656 18143
rect 8712 18087 8780 18143
rect 8836 18087 8904 18143
rect 8960 18087 9028 18143
rect 9084 18087 9094 18143
rect 8646 18019 9094 18087
rect 8646 17963 8656 18019
rect 8712 17963 8780 18019
rect 8836 17963 8904 18019
rect 8960 17963 9028 18019
rect 9084 17963 9094 18019
rect 8646 17895 9094 17963
rect 8646 17839 8656 17895
rect 8712 17839 8780 17895
rect 8836 17839 8904 17895
rect 8960 17839 9028 17895
rect 9084 17839 9094 17895
rect 8646 17771 9094 17839
rect 8646 17715 8656 17771
rect 8712 17715 8780 17771
rect 8836 17715 8904 17771
rect 8960 17715 9028 17771
rect 9084 17715 9094 17771
rect 8646 17647 9094 17715
rect 8646 17591 8656 17647
rect 8712 17591 8780 17647
rect 8836 17591 8904 17647
rect 8960 17591 9028 17647
rect 9084 17591 9094 17647
rect 8646 17523 9094 17591
rect 8646 17467 8656 17523
rect 8712 17467 8780 17523
rect 8836 17467 8904 17523
rect 8960 17467 9028 17523
rect 9084 17467 9094 17523
rect 8646 17399 9094 17467
rect 8646 17343 8656 17399
rect 8712 17343 8780 17399
rect 8836 17343 8904 17399
rect 8960 17343 9028 17399
rect 9084 17343 9094 17399
rect 8646 17333 9094 17343
rect 10918 20251 11366 20261
rect 10918 20195 10928 20251
rect 10984 20195 11052 20251
rect 11108 20195 11176 20251
rect 11232 20195 11300 20251
rect 11356 20195 11366 20251
rect 10918 20127 11366 20195
rect 10918 20071 10928 20127
rect 10984 20071 11052 20127
rect 11108 20071 11176 20127
rect 11232 20071 11300 20127
rect 11356 20071 11366 20127
rect 10918 20003 11366 20071
rect 10918 19947 10928 20003
rect 10984 19947 11052 20003
rect 11108 19947 11176 20003
rect 11232 19947 11300 20003
rect 11356 19947 11366 20003
rect 10918 19879 11366 19947
rect 10918 19823 10928 19879
rect 10984 19823 11052 19879
rect 11108 19823 11176 19879
rect 11232 19823 11300 19879
rect 11356 19823 11366 19879
rect 10918 19755 11366 19823
rect 10918 19699 10928 19755
rect 10984 19699 11052 19755
rect 11108 19699 11176 19755
rect 11232 19699 11300 19755
rect 11356 19699 11366 19755
rect 10918 19631 11366 19699
rect 10918 19575 10928 19631
rect 10984 19575 11052 19631
rect 11108 19575 11176 19631
rect 11232 19575 11300 19631
rect 11356 19575 11366 19631
rect 10918 19507 11366 19575
rect 10918 19451 10928 19507
rect 10984 19451 11052 19507
rect 11108 19451 11176 19507
rect 11232 19451 11300 19507
rect 11356 19451 11366 19507
rect 10918 19383 11366 19451
rect 10918 19327 10928 19383
rect 10984 19327 11052 19383
rect 11108 19327 11176 19383
rect 11232 19327 11300 19383
rect 11356 19327 11366 19383
rect 10918 19259 11366 19327
rect 10918 19203 10928 19259
rect 10984 19203 11052 19259
rect 11108 19203 11176 19259
rect 11232 19203 11300 19259
rect 11356 19203 11366 19259
rect 10918 19135 11366 19203
rect 10918 19079 10928 19135
rect 10984 19079 11052 19135
rect 11108 19079 11176 19135
rect 11232 19079 11300 19135
rect 11356 19079 11366 19135
rect 10918 19011 11366 19079
rect 10918 18955 10928 19011
rect 10984 18955 11052 19011
rect 11108 18955 11176 19011
rect 11232 18955 11300 19011
rect 11356 18955 11366 19011
rect 10918 18887 11366 18955
rect 10918 18831 10928 18887
rect 10984 18831 11052 18887
rect 11108 18831 11176 18887
rect 11232 18831 11300 18887
rect 11356 18831 11366 18887
rect 10918 18763 11366 18831
rect 10918 18707 10928 18763
rect 10984 18707 11052 18763
rect 11108 18707 11176 18763
rect 11232 18707 11300 18763
rect 11356 18707 11366 18763
rect 10918 18639 11366 18707
rect 10918 18583 10928 18639
rect 10984 18583 11052 18639
rect 11108 18583 11176 18639
rect 11232 18583 11300 18639
rect 11356 18583 11366 18639
rect 10918 18515 11366 18583
rect 10918 18459 10928 18515
rect 10984 18459 11052 18515
rect 11108 18459 11176 18515
rect 11232 18459 11300 18515
rect 11356 18459 11366 18515
rect 10918 18391 11366 18459
rect 10918 18335 10928 18391
rect 10984 18335 11052 18391
rect 11108 18335 11176 18391
rect 11232 18335 11300 18391
rect 11356 18335 11366 18391
rect 10918 18267 11366 18335
rect 10918 18211 10928 18267
rect 10984 18211 11052 18267
rect 11108 18211 11176 18267
rect 11232 18211 11300 18267
rect 11356 18211 11366 18267
rect 10918 18143 11366 18211
rect 10918 18087 10928 18143
rect 10984 18087 11052 18143
rect 11108 18087 11176 18143
rect 11232 18087 11300 18143
rect 11356 18087 11366 18143
rect 10918 18019 11366 18087
rect 10918 17963 10928 18019
rect 10984 17963 11052 18019
rect 11108 17963 11176 18019
rect 11232 17963 11300 18019
rect 11356 17963 11366 18019
rect 10918 17895 11366 17963
rect 10918 17839 10928 17895
rect 10984 17839 11052 17895
rect 11108 17839 11176 17895
rect 11232 17839 11300 17895
rect 11356 17839 11366 17895
rect 10918 17771 11366 17839
rect 10918 17715 10928 17771
rect 10984 17715 11052 17771
rect 11108 17715 11176 17771
rect 11232 17715 11300 17771
rect 11356 17715 11366 17771
rect 10918 17647 11366 17715
rect 10918 17591 10928 17647
rect 10984 17591 11052 17647
rect 11108 17591 11176 17647
rect 11232 17591 11300 17647
rect 11356 17591 11366 17647
rect 10918 17523 11366 17591
rect 10918 17467 10928 17523
rect 10984 17467 11052 17523
rect 11108 17467 11176 17523
rect 11232 17467 11300 17523
rect 11356 17467 11366 17523
rect 10918 17399 11366 17467
rect 10918 17343 10928 17399
rect 10984 17343 11052 17399
rect 11108 17343 11176 17399
rect 11232 17343 11300 17399
rect 11356 17343 11366 17399
rect 10918 17333 11366 17343
rect 12622 20251 13070 20261
rect 12622 20195 12632 20251
rect 12688 20195 12756 20251
rect 12812 20195 12880 20251
rect 12936 20195 13004 20251
rect 13060 20195 13070 20251
rect 12622 20127 13070 20195
rect 12622 20071 12632 20127
rect 12688 20071 12756 20127
rect 12812 20071 12880 20127
rect 12936 20071 13004 20127
rect 13060 20071 13070 20127
rect 12622 20003 13070 20071
rect 12622 19947 12632 20003
rect 12688 19947 12756 20003
rect 12812 19947 12880 20003
rect 12936 19947 13004 20003
rect 13060 19947 13070 20003
rect 12622 19879 13070 19947
rect 12622 19823 12632 19879
rect 12688 19823 12756 19879
rect 12812 19823 12880 19879
rect 12936 19823 13004 19879
rect 13060 19823 13070 19879
rect 12622 19755 13070 19823
rect 12622 19699 12632 19755
rect 12688 19699 12756 19755
rect 12812 19699 12880 19755
rect 12936 19699 13004 19755
rect 13060 19699 13070 19755
rect 12622 19631 13070 19699
rect 12622 19575 12632 19631
rect 12688 19575 12756 19631
rect 12812 19575 12880 19631
rect 12936 19575 13004 19631
rect 13060 19575 13070 19631
rect 12622 19507 13070 19575
rect 12622 19451 12632 19507
rect 12688 19451 12756 19507
rect 12812 19451 12880 19507
rect 12936 19451 13004 19507
rect 13060 19451 13070 19507
rect 12622 19383 13070 19451
rect 12622 19327 12632 19383
rect 12688 19327 12756 19383
rect 12812 19327 12880 19383
rect 12936 19327 13004 19383
rect 13060 19327 13070 19383
rect 12622 19259 13070 19327
rect 12622 19203 12632 19259
rect 12688 19203 12756 19259
rect 12812 19203 12880 19259
rect 12936 19203 13004 19259
rect 13060 19203 13070 19259
rect 12622 19135 13070 19203
rect 12622 19079 12632 19135
rect 12688 19079 12756 19135
rect 12812 19079 12880 19135
rect 12936 19079 13004 19135
rect 13060 19079 13070 19135
rect 12622 19011 13070 19079
rect 12622 18955 12632 19011
rect 12688 18955 12756 19011
rect 12812 18955 12880 19011
rect 12936 18955 13004 19011
rect 13060 18955 13070 19011
rect 12622 18887 13070 18955
rect 12622 18831 12632 18887
rect 12688 18831 12756 18887
rect 12812 18831 12880 18887
rect 12936 18831 13004 18887
rect 13060 18831 13070 18887
rect 12622 18763 13070 18831
rect 12622 18707 12632 18763
rect 12688 18707 12756 18763
rect 12812 18707 12880 18763
rect 12936 18707 13004 18763
rect 13060 18707 13070 18763
rect 12622 18639 13070 18707
rect 12622 18583 12632 18639
rect 12688 18583 12756 18639
rect 12812 18583 12880 18639
rect 12936 18583 13004 18639
rect 13060 18583 13070 18639
rect 12622 18515 13070 18583
rect 12622 18459 12632 18515
rect 12688 18459 12756 18515
rect 12812 18459 12880 18515
rect 12936 18459 13004 18515
rect 13060 18459 13070 18515
rect 12622 18391 13070 18459
rect 12622 18335 12632 18391
rect 12688 18335 12756 18391
rect 12812 18335 12880 18391
rect 12936 18335 13004 18391
rect 13060 18335 13070 18391
rect 12622 18267 13070 18335
rect 12622 18211 12632 18267
rect 12688 18211 12756 18267
rect 12812 18211 12880 18267
rect 12936 18211 13004 18267
rect 13060 18211 13070 18267
rect 12622 18143 13070 18211
rect 12622 18087 12632 18143
rect 12688 18087 12756 18143
rect 12812 18087 12880 18143
rect 12936 18087 13004 18143
rect 13060 18087 13070 18143
rect 12622 18019 13070 18087
rect 12622 17963 12632 18019
rect 12688 17963 12756 18019
rect 12812 17963 12880 18019
rect 12936 17963 13004 18019
rect 13060 17963 13070 18019
rect 12622 17895 13070 17963
rect 12622 17839 12632 17895
rect 12688 17839 12756 17895
rect 12812 17839 12880 17895
rect 12936 17839 13004 17895
rect 13060 17839 13070 17895
rect 12622 17771 13070 17839
rect 12622 17715 12632 17771
rect 12688 17715 12756 17771
rect 12812 17715 12880 17771
rect 12936 17715 13004 17771
rect 13060 17715 13070 17771
rect 12622 17647 13070 17715
rect 12622 17591 12632 17647
rect 12688 17591 12756 17647
rect 12812 17591 12880 17647
rect 12936 17591 13004 17647
rect 13060 17591 13070 17647
rect 12622 17523 13070 17591
rect 12622 17467 12632 17523
rect 12688 17467 12756 17523
rect 12812 17467 12880 17523
rect 12936 17467 13004 17523
rect 13060 17467 13070 17523
rect 12622 17399 13070 17467
rect 12622 17343 12632 17399
rect 12688 17343 12756 17399
rect 12812 17343 12880 17399
rect 12936 17343 13004 17399
rect 13060 17343 13070 17399
rect 12622 17333 13070 17343
rect 13758 20251 14206 20261
rect 13758 20195 13768 20251
rect 13824 20195 13892 20251
rect 13948 20195 14016 20251
rect 14072 20195 14140 20251
rect 14196 20195 14206 20251
rect 13758 20127 14206 20195
rect 13758 20071 13768 20127
rect 13824 20071 13892 20127
rect 13948 20071 14016 20127
rect 14072 20071 14140 20127
rect 14196 20071 14206 20127
rect 13758 20003 14206 20071
rect 13758 19947 13768 20003
rect 13824 19947 13892 20003
rect 13948 19947 14016 20003
rect 14072 19947 14140 20003
rect 14196 19947 14206 20003
rect 13758 19879 14206 19947
rect 13758 19823 13768 19879
rect 13824 19823 13892 19879
rect 13948 19823 14016 19879
rect 14072 19823 14140 19879
rect 14196 19823 14206 19879
rect 13758 19755 14206 19823
rect 13758 19699 13768 19755
rect 13824 19699 13892 19755
rect 13948 19699 14016 19755
rect 14072 19699 14140 19755
rect 14196 19699 14206 19755
rect 13758 19631 14206 19699
rect 13758 19575 13768 19631
rect 13824 19575 13892 19631
rect 13948 19575 14016 19631
rect 14072 19575 14140 19631
rect 14196 19575 14206 19631
rect 13758 19507 14206 19575
rect 13758 19451 13768 19507
rect 13824 19451 13892 19507
rect 13948 19451 14016 19507
rect 14072 19451 14140 19507
rect 14196 19451 14206 19507
rect 13758 19383 14206 19451
rect 13758 19327 13768 19383
rect 13824 19327 13892 19383
rect 13948 19327 14016 19383
rect 14072 19327 14140 19383
rect 14196 19327 14206 19383
rect 13758 19259 14206 19327
rect 13758 19203 13768 19259
rect 13824 19203 13892 19259
rect 13948 19203 14016 19259
rect 14072 19203 14140 19259
rect 14196 19203 14206 19259
rect 13758 19135 14206 19203
rect 13758 19079 13768 19135
rect 13824 19079 13892 19135
rect 13948 19079 14016 19135
rect 14072 19079 14140 19135
rect 14196 19079 14206 19135
rect 13758 19011 14206 19079
rect 13758 18955 13768 19011
rect 13824 18955 13892 19011
rect 13948 18955 14016 19011
rect 14072 18955 14140 19011
rect 14196 18955 14206 19011
rect 13758 18887 14206 18955
rect 13758 18831 13768 18887
rect 13824 18831 13892 18887
rect 13948 18831 14016 18887
rect 14072 18831 14140 18887
rect 14196 18831 14206 18887
rect 13758 18763 14206 18831
rect 13758 18707 13768 18763
rect 13824 18707 13892 18763
rect 13948 18707 14016 18763
rect 14072 18707 14140 18763
rect 14196 18707 14206 18763
rect 13758 18639 14206 18707
rect 13758 18583 13768 18639
rect 13824 18583 13892 18639
rect 13948 18583 14016 18639
rect 14072 18583 14140 18639
rect 14196 18583 14206 18639
rect 13758 18515 14206 18583
rect 13758 18459 13768 18515
rect 13824 18459 13892 18515
rect 13948 18459 14016 18515
rect 14072 18459 14140 18515
rect 14196 18459 14206 18515
rect 13758 18391 14206 18459
rect 13758 18335 13768 18391
rect 13824 18335 13892 18391
rect 13948 18335 14016 18391
rect 14072 18335 14140 18391
rect 14196 18335 14206 18391
rect 13758 18267 14206 18335
rect 13758 18211 13768 18267
rect 13824 18211 13892 18267
rect 13948 18211 14016 18267
rect 14072 18211 14140 18267
rect 14196 18211 14206 18267
rect 13758 18143 14206 18211
rect 13758 18087 13768 18143
rect 13824 18087 13892 18143
rect 13948 18087 14016 18143
rect 14072 18087 14140 18143
rect 14196 18087 14206 18143
rect 13758 18019 14206 18087
rect 13758 17963 13768 18019
rect 13824 17963 13892 18019
rect 13948 17963 14016 18019
rect 14072 17963 14140 18019
rect 14196 17963 14206 18019
rect 13758 17895 14206 17963
rect 13758 17839 13768 17895
rect 13824 17839 13892 17895
rect 13948 17839 14016 17895
rect 14072 17839 14140 17895
rect 14196 17839 14206 17895
rect 13758 17771 14206 17839
rect 13758 17715 13768 17771
rect 13824 17715 13892 17771
rect 13948 17715 14016 17771
rect 14072 17715 14140 17771
rect 14196 17715 14206 17771
rect 13758 17647 14206 17715
rect 13758 17591 13768 17647
rect 13824 17591 13892 17647
rect 13948 17591 14016 17647
rect 14072 17591 14140 17647
rect 14196 17591 14206 17647
rect 13758 17523 14206 17591
rect 13758 17467 13768 17523
rect 13824 17467 13892 17523
rect 13948 17467 14016 17523
rect 14072 17467 14140 17523
rect 14196 17467 14206 17523
rect 13758 17399 14206 17467
rect 13758 17343 13768 17399
rect 13824 17343 13892 17399
rect 13948 17343 14016 17399
rect 14072 17343 14140 17399
rect 14196 17343 14206 17399
rect 13758 17333 14206 17343
rect 858 17051 1306 17061
rect 858 16995 868 17051
rect 924 16995 992 17051
rect 1048 16995 1116 17051
rect 1172 16995 1240 17051
rect 1296 16995 1306 17051
rect 858 16927 1306 16995
rect 858 16871 868 16927
rect 924 16871 992 16927
rect 1048 16871 1116 16927
rect 1172 16871 1240 16927
rect 1296 16871 1306 16927
rect 858 16803 1306 16871
rect 858 16747 868 16803
rect 924 16747 992 16803
rect 1048 16747 1116 16803
rect 1172 16747 1240 16803
rect 1296 16747 1306 16803
rect 858 16679 1306 16747
rect 858 16623 868 16679
rect 924 16623 992 16679
rect 1048 16623 1116 16679
rect 1172 16623 1240 16679
rect 1296 16623 1306 16679
rect 858 16555 1306 16623
rect 858 16499 868 16555
rect 924 16499 992 16555
rect 1048 16499 1116 16555
rect 1172 16499 1240 16555
rect 1296 16499 1306 16555
rect 858 16431 1306 16499
rect 858 16375 868 16431
rect 924 16375 992 16431
rect 1048 16375 1116 16431
rect 1172 16375 1240 16431
rect 1296 16375 1306 16431
rect 858 16307 1306 16375
rect 858 16251 868 16307
rect 924 16251 992 16307
rect 1048 16251 1116 16307
rect 1172 16251 1240 16307
rect 1296 16251 1306 16307
rect 858 16183 1306 16251
rect 858 16127 868 16183
rect 924 16127 992 16183
rect 1048 16127 1116 16183
rect 1172 16127 1240 16183
rect 1296 16127 1306 16183
rect 858 16059 1306 16127
rect 858 16003 868 16059
rect 924 16003 992 16059
rect 1048 16003 1116 16059
rect 1172 16003 1240 16059
rect 1296 16003 1306 16059
rect 858 15935 1306 16003
rect 858 15879 868 15935
rect 924 15879 992 15935
rect 1048 15879 1116 15935
rect 1172 15879 1240 15935
rect 1296 15879 1306 15935
rect 858 15811 1306 15879
rect 858 15755 868 15811
rect 924 15755 992 15811
rect 1048 15755 1116 15811
rect 1172 15755 1240 15811
rect 1296 15755 1306 15811
rect 858 15687 1306 15755
rect 858 15631 868 15687
rect 924 15631 992 15687
rect 1048 15631 1116 15687
rect 1172 15631 1240 15687
rect 1296 15631 1306 15687
rect 858 15563 1306 15631
rect 858 15507 868 15563
rect 924 15507 992 15563
rect 1048 15507 1116 15563
rect 1172 15507 1240 15563
rect 1296 15507 1306 15563
rect 858 15439 1306 15507
rect 858 15383 868 15439
rect 924 15383 992 15439
rect 1048 15383 1116 15439
rect 1172 15383 1240 15439
rect 1296 15383 1306 15439
rect 858 15315 1306 15383
rect 858 15259 868 15315
rect 924 15259 992 15315
rect 1048 15259 1116 15315
rect 1172 15259 1240 15315
rect 1296 15259 1306 15315
rect 858 15191 1306 15259
rect 858 15135 868 15191
rect 924 15135 992 15191
rect 1048 15135 1116 15191
rect 1172 15135 1240 15191
rect 1296 15135 1306 15191
rect 858 15067 1306 15135
rect 858 15011 868 15067
rect 924 15011 992 15067
rect 1048 15011 1116 15067
rect 1172 15011 1240 15067
rect 1296 15011 1306 15067
rect 858 14943 1306 15011
rect 858 14887 868 14943
rect 924 14887 992 14943
rect 1048 14887 1116 14943
rect 1172 14887 1240 14943
rect 1296 14887 1306 14943
rect 858 14819 1306 14887
rect 858 14763 868 14819
rect 924 14763 992 14819
rect 1048 14763 1116 14819
rect 1172 14763 1240 14819
rect 1296 14763 1306 14819
rect 858 14695 1306 14763
rect 858 14639 868 14695
rect 924 14639 992 14695
rect 1048 14639 1116 14695
rect 1172 14639 1240 14695
rect 1296 14639 1306 14695
rect 858 14571 1306 14639
rect 858 14515 868 14571
rect 924 14515 992 14571
rect 1048 14515 1116 14571
rect 1172 14515 1240 14571
rect 1296 14515 1306 14571
rect 858 14447 1306 14515
rect 858 14391 868 14447
rect 924 14391 992 14447
rect 1048 14391 1116 14447
rect 1172 14391 1240 14447
rect 1296 14391 1306 14447
rect 858 14323 1306 14391
rect 858 14267 868 14323
rect 924 14267 992 14323
rect 1048 14267 1116 14323
rect 1172 14267 1240 14323
rect 1296 14267 1306 14323
rect 858 14199 1306 14267
rect 858 14143 868 14199
rect 924 14143 992 14199
rect 1048 14143 1116 14199
rect 1172 14143 1240 14199
rect 1296 14143 1306 14199
rect 858 14133 1306 14143
rect 1994 17051 2442 17061
rect 1994 16995 2004 17051
rect 2060 16995 2128 17051
rect 2184 16995 2252 17051
rect 2308 16995 2376 17051
rect 2432 16995 2442 17051
rect 1994 16927 2442 16995
rect 1994 16871 2004 16927
rect 2060 16871 2128 16927
rect 2184 16871 2252 16927
rect 2308 16871 2376 16927
rect 2432 16871 2442 16927
rect 1994 16803 2442 16871
rect 1994 16747 2004 16803
rect 2060 16747 2128 16803
rect 2184 16747 2252 16803
rect 2308 16747 2376 16803
rect 2432 16747 2442 16803
rect 1994 16679 2442 16747
rect 1994 16623 2004 16679
rect 2060 16623 2128 16679
rect 2184 16623 2252 16679
rect 2308 16623 2376 16679
rect 2432 16623 2442 16679
rect 1994 16555 2442 16623
rect 1994 16499 2004 16555
rect 2060 16499 2128 16555
rect 2184 16499 2252 16555
rect 2308 16499 2376 16555
rect 2432 16499 2442 16555
rect 1994 16431 2442 16499
rect 1994 16375 2004 16431
rect 2060 16375 2128 16431
rect 2184 16375 2252 16431
rect 2308 16375 2376 16431
rect 2432 16375 2442 16431
rect 1994 16307 2442 16375
rect 1994 16251 2004 16307
rect 2060 16251 2128 16307
rect 2184 16251 2252 16307
rect 2308 16251 2376 16307
rect 2432 16251 2442 16307
rect 1994 16183 2442 16251
rect 1994 16127 2004 16183
rect 2060 16127 2128 16183
rect 2184 16127 2252 16183
rect 2308 16127 2376 16183
rect 2432 16127 2442 16183
rect 1994 16059 2442 16127
rect 1994 16003 2004 16059
rect 2060 16003 2128 16059
rect 2184 16003 2252 16059
rect 2308 16003 2376 16059
rect 2432 16003 2442 16059
rect 1994 15935 2442 16003
rect 1994 15879 2004 15935
rect 2060 15879 2128 15935
rect 2184 15879 2252 15935
rect 2308 15879 2376 15935
rect 2432 15879 2442 15935
rect 1994 15811 2442 15879
rect 1994 15755 2004 15811
rect 2060 15755 2128 15811
rect 2184 15755 2252 15811
rect 2308 15755 2376 15811
rect 2432 15755 2442 15811
rect 1994 15687 2442 15755
rect 1994 15631 2004 15687
rect 2060 15631 2128 15687
rect 2184 15631 2252 15687
rect 2308 15631 2376 15687
rect 2432 15631 2442 15687
rect 1994 15563 2442 15631
rect 1994 15507 2004 15563
rect 2060 15507 2128 15563
rect 2184 15507 2252 15563
rect 2308 15507 2376 15563
rect 2432 15507 2442 15563
rect 1994 15439 2442 15507
rect 1994 15383 2004 15439
rect 2060 15383 2128 15439
rect 2184 15383 2252 15439
rect 2308 15383 2376 15439
rect 2432 15383 2442 15439
rect 1994 15315 2442 15383
rect 1994 15259 2004 15315
rect 2060 15259 2128 15315
rect 2184 15259 2252 15315
rect 2308 15259 2376 15315
rect 2432 15259 2442 15315
rect 1994 15191 2442 15259
rect 1994 15135 2004 15191
rect 2060 15135 2128 15191
rect 2184 15135 2252 15191
rect 2308 15135 2376 15191
rect 2432 15135 2442 15191
rect 1994 15067 2442 15135
rect 1994 15011 2004 15067
rect 2060 15011 2128 15067
rect 2184 15011 2252 15067
rect 2308 15011 2376 15067
rect 2432 15011 2442 15067
rect 1994 14943 2442 15011
rect 1994 14887 2004 14943
rect 2060 14887 2128 14943
rect 2184 14887 2252 14943
rect 2308 14887 2376 14943
rect 2432 14887 2442 14943
rect 1994 14819 2442 14887
rect 1994 14763 2004 14819
rect 2060 14763 2128 14819
rect 2184 14763 2252 14819
rect 2308 14763 2376 14819
rect 2432 14763 2442 14819
rect 1994 14695 2442 14763
rect 1994 14639 2004 14695
rect 2060 14639 2128 14695
rect 2184 14639 2252 14695
rect 2308 14639 2376 14695
rect 2432 14639 2442 14695
rect 1994 14571 2442 14639
rect 1994 14515 2004 14571
rect 2060 14515 2128 14571
rect 2184 14515 2252 14571
rect 2308 14515 2376 14571
rect 2432 14515 2442 14571
rect 1994 14447 2442 14515
rect 1994 14391 2004 14447
rect 2060 14391 2128 14447
rect 2184 14391 2252 14447
rect 2308 14391 2376 14447
rect 2432 14391 2442 14447
rect 1994 14323 2442 14391
rect 1994 14267 2004 14323
rect 2060 14267 2128 14323
rect 2184 14267 2252 14323
rect 2308 14267 2376 14323
rect 2432 14267 2442 14323
rect 1994 14199 2442 14267
rect 1994 14143 2004 14199
rect 2060 14143 2128 14199
rect 2184 14143 2252 14199
rect 2308 14143 2376 14199
rect 2432 14143 2442 14199
rect 1994 14133 2442 14143
rect 3698 17051 4146 17061
rect 3698 16995 3708 17051
rect 3764 16995 3832 17051
rect 3888 16995 3956 17051
rect 4012 16995 4080 17051
rect 4136 16995 4146 17051
rect 3698 16927 4146 16995
rect 3698 16871 3708 16927
rect 3764 16871 3832 16927
rect 3888 16871 3956 16927
rect 4012 16871 4080 16927
rect 4136 16871 4146 16927
rect 3698 16803 4146 16871
rect 3698 16747 3708 16803
rect 3764 16747 3832 16803
rect 3888 16747 3956 16803
rect 4012 16747 4080 16803
rect 4136 16747 4146 16803
rect 3698 16679 4146 16747
rect 3698 16623 3708 16679
rect 3764 16623 3832 16679
rect 3888 16623 3956 16679
rect 4012 16623 4080 16679
rect 4136 16623 4146 16679
rect 3698 16555 4146 16623
rect 3698 16499 3708 16555
rect 3764 16499 3832 16555
rect 3888 16499 3956 16555
rect 4012 16499 4080 16555
rect 4136 16499 4146 16555
rect 3698 16431 4146 16499
rect 3698 16375 3708 16431
rect 3764 16375 3832 16431
rect 3888 16375 3956 16431
rect 4012 16375 4080 16431
rect 4136 16375 4146 16431
rect 3698 16307 4146 16375
rect 3698 16251 3708 16307
rect 3764 16251 3832 16307
rect 3888 16251 3956 16307
rect 4012 16251 4080 16307
rect 4136 16251 4146 16307
rect 3698 16183 4146 16251
rect 3698 16127 3708 16183
rect 3764 16127 3832 16183
rect 3888 16127 3956 16183
rect 4012 16127 4080 16183
rect 4136 16127 4146 16183
rect 3698 16059 4146 16127
rect 3698 16003 3708 16059
rect 3764 16003 3832 16059
rect 3888 16003 3956 16059
rect 4012 16003 4080 16059
rect 4136 16003 4146 16059
rect 3698 15935 4146 16003
rect 3698 15879 3708 15935
rect 3764 15879 3832 15935
rect 3888 15879 3956 15935
rect 4012 15879 4080 15935
rect 4136 15879 4146 15935
rect 3698 15811 4146 15879
rect 3698 15755 3708 15811
rect 3764 15755 3832 15811
rect 3888 15755 3956 15811
rect 4012 15755 4080 15811
rect 4136 15755 4146 15811
rect 3698 15687 4146 15755
rect 3698 15631 3708 15687
rect 3764 15631 3832 15687
rect 3888 15631 3956 15687
rect 4012 15631 4080 15687
rect 4136 15631 4146 15687
rect 3698 15563 4146 15631
rect 3698 15507 3708 15563
rect 3764 15507 3832 15563
rect 3888 15507 3956 15563
rect 4012 15507 4080 15563
rect 4136 15507 4146 15563
rect 3698 15439 4146 15507
rect 3698 15383 3708 15439
rect 3764 15383 3832 15439
rect 3888 15383 3956 15439
rect 4012 15383 4080 15439
rect 4136 15383 4146 15439
rect 3698 15315 4146 15383
rect 3698 15259 3708 15315
rect 3764 15259 3832 15315
rect 3888 15259 3956 15315
rect 4012 15259 4080 15315
rect 4136 15259 4146 15315
rect 3698 15191 4146 15259
rect 3698 15135 3708 15191
rect 3764 15135 3832 15191
rect 3888 15135 3956 15191
rect 4012 15135 4080 15191
rect 4136 15135 4146 15191
rect 3698 15067 4146 15135
rect 3698 15011 3708 15067
rect 3764 15011 3832 15067
rect 3888 15011 3956 15067
rect 4012 15011 4080 15067
rect 4136 15011 4146 15067
rect 3698 14943 4146 15011
rect 3698 14887 3708 14943
rect 3764 14887 3832 14943
rect 3888 14887 3956 14943
rect 4012 14887 4080 14943
rect 4136 14887 4146 14943
rect 3698 14819 4146 14887
rect 3698 14763 3708 14819
rect 3764 14763 3832 14819
rect 3888 14763 3956 14819
rect 4012 14763 4080 14819
rect 4136 14763 4146 14819
rect 3698 14695 4146 14763
rect 3698 14639 3708 14695
rect 3764 14639 3832 14695
rect 3888 14639 3956 14695
rect 4012 14639 4080 14695
rect 4136 14639 4146 14695
rect 3698 14571 4146 14639
rect 3698 14515 3708 14571
rect 3764 14515 3832 14571
rect 3888 14515 3956 14571
rect 4012 14515 4080 14571
rect 4136 14515 4146 14571
rect 3698 14447 4146 14515
rect 3698 14391 3708 14447
rect 3764 14391 3832 14447
rect 3888 14391 3956 14447
rect 4012 14391 4080 14447
rect 4136 14391 4146 14447
rect 3698 14323 4146 14391
rect 3698 14267 3708 14323
rect 3764 14267 3832 14323
rect 3888 14267 3956 14323
rect 4012 14267 4080 14323
rect 4136 14267 4146 14323
rect 3698 14199 4146 14267
rect 3698 14143 3708 14199
rect 3764 14143 3832 14199
rect 3888 14143 3956 14199
rect 4012 14143 4080 14199
rect 4136 14143 4146 14199
rect 3698 14133 4146 14143
rect 5970 17051 6418 17061
rect 5970 16995 5980 17051
rect 6036 16995 6104 17051
rect 6160 16995 6228 17051
rect 6284 16995 6352 17051
rect 6408 16995 6418 17051
rect 5970 16927 6418 16995
rect 5970 16871 5980 16927
rect 6036 16871 6104 16927
rect 6160 16871 6228 16927
rect 6284 16871 6352 16927
rect 6408 16871 6418 16927
rect 5970 16803 6418 16871
rect 5970 16747 5980 16803
rect 6036 16747 6104 16803
rect 6160 16747 6228 16803
rect 6284 16747 6352 16803
rect 6408 16747 6418 16803
rect 5970 16679 6418 16747
rect 5970 16623 5980 16679
rect 6036 16623 6104 16679
rect 6160 16623 6228 16679
rect 6284 16623 6352 16679
rect 6408 16623 6418 16679
rect 5970 16555 6418 16623
rect 5970 16499 5980 16555
rect 6036 16499 6104 16555
rect 6160 16499 6228 16555
rect 6284 16499 6352 16555
rect 6408 16499 6418 16555
rect 5970 16431 6418 16499
rect 5970 16375 5980 16431
rect 6036 16375 6104 16431
rect 6160 16375 6228 16431
rect 6284 16375 6352 16431
rect 6408 16375 6418 16431
rect 5970 16307 6418 16375
rect 5970 16251 5980 16307
rect 6036 16251 6104 16307
rect 6160 16251 6228 16307
rect 6284 16251 6352 16307
rect 6408 16251 6418 16307
rect 5970 16183 6418 16251
rect 5970 16127 5980 16183
rect 6036 16127 6104 16183
rect 6160 16127 6228 16183
rect 6284 16127 6352 16183
rect 6408 16127 6418 16183
rect 5970 16059 6418 16127
rect 5970 16003 5980 16059
rect 6036 16003 6104 16059
rect 6160 16003 6228 16059
rect 6284 16003 6352 16059
rect 6408 16003 6418 16059
rect 5970 15935 6418 16003
rect 5970 15879 5980 15935
rect 6036 15879 6104 15935
rect 6160 15879 6228 15935
rect 6284 15879 6352 15935
rect 6408 15879 6418 15935
rect 5970 15811 6418 15879
rect 5970 15755 5980 15811
rect 6036 15755 6104 15811
rect 6160 15755 6228 15811
rect 6284 15755 6352 15811
rect 6408 15755 6418 15811
rect 5970 15687 6418 15755
rect 5970 15631 5980 15687
rect 6036 15631 6104 15687
rect 6160 15631 6228 15687
rect 6284 15631 6352 15687
rect 6408 15631 6418 15687
rect 5970 15563 6418 15631
rect 5970 15507 5980 15563
rect 6036 15507 6104 15563
rect 6160 15507 6228 15563
rect 6284 15507 6352 15563
rect 6408 15507 6418 15563
rect 5970 15439 6418 15507
rect 5970 15383 5980 15439
rect 6036 15383 6104 15439
rect 6160 15383 6228 15439
rect 6284 15383 6352 15439
rect 6408 15383 6418 15439
rect 5970 15315 6418 15383
rect 5970 15259 5980 15315
rect 6036 15259 6104 15315
rect 6160 15259 6228 15315
rect 6284 15259 6352 15315
rect 6408 15259 6418 15315
rect 5970 15191 6418 15259
rect 5970 15135 5980 15191
rect 6036 15135 6104 15191
rect 6160 15135 6228 15191
rect 6284 15135 6352 15191
rect 6408 15135 6418 15191
rect 5970 15067 6418 15135
rect 5970 15011 5980 15067
rect 6036 15011 6104 15067
rect 6160 15011 6228 15067
rect 6284 15011 6352 15067
rect 6408 15011 6418 15067
rect 5970 14943 6418 15011
rect 5970 14887 5980 14943
rect 6036 14887 6104 14943
rect 6160 14887 6228 14943
rect 6284 14887 6352 14943
rect 6408 14887 6418 14943
rect 5970 14819 6418 14887
rect 5970 14763 5980 14819
rect 6036 14763 6104 14819
rect 6160 14763 6228 14819
rect 6284 14763 6352 14819
rect 6408 14763 6418 14819
rect 5970 14695 6418 14763
rect 5970 14639 5980 14695
rect 6036 14639 6104 14695
rect 6160 14639 6228 14695
rect 6284 14639 6352 14695
rect 6408 14639 6418 14695
rect 5970 14571 6418 14639
rect 5970 14515 5980 14571
rect 6036 14515 6104 14571
rect 6160 14515 6228 14571
rect 6284 14515 6352 14571
rect 6408 14515 6418 14571
rect 5970 14447 6418 14515
rect 5970 14391 5980 14447
rect 6036 14391 6104 14447
rect 6160 14391 6228 14447
rect 6284 14391 6352 14447
rect 6408 14391 6418 14447
rect 5970 14323 6418 14391
rect 5970 14267 5980 14323
rect 6036 14267 6104 14323
rect 6160 14267 6228 14323
rect 6284 14267 6352 14323
rect 6408 14267 6418 14323
rect 5970 14199 6418 14267
rect 5970 14143 5980 14199
rect 6036 14143 6104 14199
rect 6160 14143 6228 14199
rect 6284 14143 6352 14199
rect 6408 14143 6418 14199
rect 5970 14133 6418 14143
rect 8646 17051 9094 17061
rect 8646 16995 8656 17051
rect 8712 16995 8780 17051
rect 8836 16995 8904 17051
rect 8960 16995 9028 17051
rect 9084 16995 9094 17051
rect 8646 16927 9094 16995
rect 8646 16871 8656 16927
rect 8712 16871 8780 16927
rect 8836 16871 8904 16927
rect 8960 16871 9028 16927
rect 9084 16871 9094 16927
rect 8646 16803 9094 16871
rect 8646 16747 8656 16803
rect 8712 16747 8780 16803
rect 8836 16747 8904 16803
rect 8960 16747 9028 16803
rect 9084 16747 9094 16803
rect 8646 16679 9094 16747
rect 8646 16623 8656 16679
rect 8712 16623 8780 16679
rect 8836 16623 8904 16679
rect 8960 16623 9028 16679
rect 9084 16623 9094 16679
rect 8646 16555 9094 16623
rect 8646 16499 8656 16555
rect 8712 16499 8780 16555
rect 8836 16499 8904 16555
rect 8960 16499 9028 16555
rect 9084 16499 9094 16555
rect 8646 16431 9094 16499
rect 8646 16375 8656 16431
rect 8712 16375 8780 16431
rect 8836 16375 8904 16431
rect 8960 16375 9028 16431
rect 9084 16375 9094 16431
rect 8646 16307 9094 16375
rect 8646 16251 8656 16307
rect 8712 16251 8780 16307
rect 8836 16251 8904 16307
rect 8960 16251 9028 16307
rect 9084 16251 9094 16307
rect 8646 16183 9094 16251
rect 8646 16127 8656 16183
rect 8712 16127 8780 16183
rect 8836 16127 8904 16183
rect 8960 16127 9028 16183
rect 9084 16127 9094 16183
rect 8646 16059 9094 16127
rect 8646 16003 8656 16059
rect 8712 16003 8780 16059
rect 8836 16003 8904 16059
rect 8960 16003 9028 16059
rect 9084 16003 9094 16059
rect 8646 15935 9094 16003
rect 8646 15879 8656 15935
rect 8712 15879 8780 15935
rect 8836 15879 8904 15935
rect 8960 15879 9028 15935
rect 9084 15879 9094 15935
rect 8646 15811 9094 15879
rect 8646 15755 8656 15811
rect 8712 15755 8780 15811
rect 8836 15755 8904 15811
rect 8960 15755 9028 15811
rect 9084 15755 9094 15811
rect 8646 15687 9094 15755
rect 8646 15631 8656 15687
rect 8712 15631 8780 15687
rect 8836 15631 8904 15687
rect 8960 15631 9028 15687
rect 9084 15631 9094 15687
rect 8646 15563 9094 15631
rect 8646 15507 8656 15563
rect 8712 15507 8780 15563
rect 8836 15507 8904 15563
rect 8960 15507 9028 15563
rect 9084 15507 9094 15563
rect 8646 15439 9094 15507
rect 8646 15383 8656 15439
rect 8712 15383 8780 15439
rect 8836 15383 8904 15439
rect 8960 15383 9028 15439
rect 9084 15383 9094 15439
rect 8646 15315 9094 15383
rect 8646 15259 8656 15315
rect 8712 15259 8780 15315
rect 8836 15259 8904 15315
rect 8960 15259 9028 15315
rect 9084 15259 9094 15315
rect 8646 15191 9094 15259
rect 8646 15135 8656 15191
rect 8712 15135 8780 15191
rect 8836 15135 8904 15191
rect 8960 15135 9028 15191
rect 9084 15135 9094 15191
rect 8646 15067 9094 15135
rect 8646 15011 8656 15067
rect 8712 15011 8780 15067
rect 8836 15011 8904 15067
rect 8960 15011 9028 15067
rect 9084 15011 9094 15067
rect 8646 14943 9094 15011
rect 8646 14887 8656 14943
rect 8712 14887 8780 14943
rect 8836 14887 8904 14943
rect 8960 14887 9028 14943
rect 9084 14887 9094 14943
rect 8646 14819 9094 14887
rect 8646 14763 8656 14819
rect 8712 14763 8780 14819
rect 8836 14763 8904 14819
rect 8960 14763 9028 14819
rect 9084 14763 9094 14819
rect 8646 14695 9094 14763
rect 8646 14639 8656 14695
rect 8712 14639 8780 14695
rect 8836 14639 8904 14695
rect 8960 14639 9028 14695
rect 9084 14639 9094 14695
rect 8646 14571 9094 14639
rect 8646 14515 8656 14571
rect 8712 14515 8780 14571
rect 8836 14515 8904 14571
rect 8960 14515 9028 14571
rect 9084 14515 9094 14571
rect 8646 14447 9094 14515
rect 8646 14391 8656 14447
rect 8712 14391 8780 14447
rect 8836 14391 8904 14447
rect 8960 14391 9028 14447
rect 9084 14391 9094 14447
rect 8646 14323 9094 14391
rect 8646 14267 8656 14323
rect 8712 14267 8780 14323
rect 8836 14267 8904 14323
rect 8960 14267 9028 14323
rect 9084 14267 9094 14323
rect 8646 14199 9094 14267
rect 8646 14143 8656 14199
rect 8712 14143 8780 14199
rect 8836 14143 8904 14199
rect 8960 14143 9028 14199
rect 9084 14143 9094 14199
rect 8646 14133 9094 14143
rect 10918 17051 11366 17061
rect 10918 16995 10928 17051
rect 10984 16995 11052 17051
rect 11108 16995 11176 17051
rect 11232 16995 11300 17051
rect 11356 16995 11366 17051
rect 10918 16927 11366 16995
rect 10918 16871 10928 16927
rect 10984 16871 11052 16927
rect 11108 16871 11176 16927
rect 11232 16871 11300 16927
rect 11356 16871 11366 16927
rect 10918 16803 11366 16871
rect 10918 16747 10928 16803
rect 10984 16747 11052 16803
rect 11108 16747 11176 16803
rect 11232 16747 11300 16803
rect 11356 16747 11366 16803
rect 10918 16679 11366 16747
rect 10918 16623 10928 16679
rect 10984 16623 11052 16679
rect 11108 16623 11176 16679
rect 11232 16623 11300 16679
rect 11356 16623 11366 16679
rect 10918 16555 11366 16623
rect 10918 16499 10928 16555
rect 10984 16499 11052 16555
rect 11108 16499 11176 16555
rect 11232 16499 11300 16555
rect 11356 16499 11366 16555
rect 10918 16431 11366 16499
rect 10918 16375 10928 16431
rect 10984 16375 11052 16431
rect 11108 16375 11176 16431
rect 11232 16375 11300 16431
rect 11356 16375 11366 16431
rect 10918 16307 11366 16375
rect 10918 16251 10928 16307
rect 10984 16251 11052 16307
rect 11108 16251 11176 16307
rect 11232 16251 11300 16307
rect 11356 16251 11366 16307
rect 10918 16183 11366 16251
rect 10918 16127 10928 16183
rect 10984 16127 11052 16183
rect 11108 16127 11176 16183
rect 11232 16127 11300 16183
rect 11356 16127 11366 16183
rect 10918 16059 11366 16127
rect 10918 16003 10928 16059
rect 10984 16003 11052 16059
rect 11108 16003 11176 16059
rect 11232 16003 11300 16059
rect 11356 16003 11366 16059
rect 10918 15935 11366 16003
rect 10918 15879 10928 15935
rect 10984 15879 11052 15935
rect 11108 15879 11176 15935
rect 11232 15879 11300 15935
rect 11356 15879 11366 15935
rect 10918 15811 11366 15879
rect 10918 15755 10928 15811
rect 10984 15755 11052 15811
rect 11108 15755 11176 15811
rect 11232 15755 11300 15811
rect 11356 15755 11366 15811
rect 10918 15687 11366 15755
rect 10918 15631 10928 15687
rect 10984 15631 11052 15687
rect 11108 15631 11176 15687
rect 11232 15631 11300 15687
rect 11356 15631 11366 15687
rect 10918 15563 11366 15631
rect 10918 15507 10928 15563
rect 10984 15507 11052 15563
rect 11108 15507 11176 15563
rect 11232 15507 11300 15563
rect 11356 15507 11366 15563
rect 10918 15439 11366 15507
rect 10918 15383 10928 15439
rect 10984 15383 11052 15439
rect 11108 15383 11176 15439
rect 11232 15383 11300 15439
rect 11356 15383 11366 15439
rect 10918 15315 11366 15383
rect 10918 15259 10928 15315
rect 10984 15259 11052 15315
rect 11108 15259 11176 15315
rect 11232 15259 11300 15315
rect 11356 15259 11366 15315
rect 10918 15191 11366 15259
rect 10918 15135 10928 15191
rect 10984 15135 11052 15191
rect 11108 15135 11176 15191
rect 11232 15135 11300 15191
rect 11356 15135 11366 15191
rect 10918 15067 11366 15135
rect 10918 15011 10928 15067
rect 10984 15011 11052 15067
rect 11108 15011 11176 15067
rect 11232 15011 11300 15067
rect 11356 15011 11366 15067
rect 10918 14943 11366 15011
rect 10918 14887 10928 14943
rect 10984 14887 11052 14943
rect 11108 14887 11176 14943
rect 11232 14887 11300 14943
rect 11356 14887 11366 14943
rect 10918 14819 11366 14887
rect 10918 14763 10928 14819
rect 10984 14763 11052 14819
rect 11108 14763 11176 14819
rect 11232 14763 11300 14819
rect 11356 14763 11366 14819
rect 10918 14695 11366 14763
rect 10918 14639 10928 14695
rect 10984 14639 11052 14695
rect 11108 14639 11176 14695
rect 11232 14639 11300 14695
rect 11356 14639 11366 14695
rect 10918 14571 11366 14639
rect 10918 14515 10928 14571
rect 10984 14515 11052 14571
rect 11108 14515 11176 14571
rect 11232 14515 11300 14571
rect 11356 14515 11366 14571
rect 10918 14447 11366 14515
rect 10918 14391 10928 14447
rect 10984 14391 11052 14447
rect 11108 14391 11176 14447
rect 11232 14391 11300 14447
rect 11356 14391 11366 14447
rect 10918 14323 11366 14391
rect 10918 14267 10928 14323
rect 10984 14267 11052 14323
rect 11108 14267 11176 14323
rect 11232 14267 11300 14323
rect 11356 14267 11366 14323
rect 10918 14199 11366 14267
rect 10918 14143 10928 14199
rect 10984 14143 11052 14199
rect 11108 14143 11176 14199
rect 11232 14143 11300 14199
rect 11356 14143 11366 14199
rect 10918 14133 11366 14143
rect 12622 17051 13070 17061
rect 12622 16995 12632 17051
rect 12688 16995 12756 17051
rect 12812 16995 12880 17051
rect 12936 16995 13004 17051
rect 13060 16995 13070 17051
rect 12622 16927 13070 16995
rect 12622 16871 12632 16927
rect 12688 16871 12756 16927
rect 12812 16871 12880 16927
rect 12936 16871 13004 16927
rect 13060 16871 13070 16927
rect 12622 16803 13070 16871
rect 12622 16747 12632 16803
rect 12688 16747 12756 16803
rect 12812 16747 12880 16803
rect 12936 16747 13004 16803
rect 13060 16747 13070 16803
rect 12622 16679 13070 16747
rect 12622 16623 12632 16679
rect 12688 16623 12756 16679
rect 12812 16623 12880 16679
rect 12936 16623 13004 16679
rect 13060 16623 13070 16679
rect 12622 16555 13070 16623
rect 12622 16499 12632 16555
rect 12688 16499 12756 16555
rect 12812 16499 12880 16555
rect 12936 16499 13004 16555
rect 13060 16499 13070 16555
rect 12622 16431 13070 16499
rect 12622 16375 12632 16431
rect 12688 16375 12756 16431
rect 12812 16375 12880 16431
rect 12936 16375 13004 16431
rect 13060 16375 13070 16431
rect 12622 16307 13070 16375
rect 12622 16251 12632 16307
rect 12688 16251 12756 16307
rect 12812 16251 12880 16307
rect 12936 16251 13004 16307
rect 13060 16251 13070 16307
rect 12622 16183 13070 16251
rect 12622 16127 12632 16183
rect 12688 16127 12756 16183
rect 12812 16127 12880 16183
rect 12936 16127 13004 16183
rect 13060 16127 13070 16183
rect 12622 16059 13070 16127
rect 12622 16003 12632 16059
rect 12688 16003 12756 16059
rect 12812 16003 12880 16059
rect 12936 16003 13004 16059
rect 13060 16003 13070 16059
rect 12622 15935 13070 16003
rect 12622 15879 12632 15935
rect 12688 15879 12756 15935
rect 12812 15879 12880 15935
rect 12936 15879 13004 15935
rect 13060 15879 13070 15935
rect 12622 15811 13070 15879
rect 12622 15755 12632 15811
rect 12688 15755 12756 15811
rect 12812 15755 12880 15811
rect 12936 15755 13004 15811
rect 13060 15755 13070 15811
rect 12622 15687 13070 15755
rect 12622 15631 12632 15687
rect 12688 15631 12756 15687
rect 12812 15631 12880 15687
rect 12936 15631 13004 15687
rect 13060 15631 13070 15687
rect 12622 15563 13070 15631
rect 12622 15507 12632 15563
rect 12688 15507 12756 15563
rect 12812 15507 12880 15563
rect 12936 15507 13004 15563
rect 13060 15507 13070 15563
rect 12622 15439 13070 15507
rect 12622 15383 12632 15439
rect 12688 15383 12756 15439
rect 12812 15383 12880 15439
rect 12936 15383 13004 15439
rect 13060 15383 13070 15439
rect 12622 15315 13070 15383
rect 12622 15259 12632 15315
rect 12688 15259 12756 15315
rect 12812 15259 12880 15315
rect 12936 15259 13004 15315
rect 13060 15259 13070 15315
rect 12622 15191 13070 15259
rect 12622 15135 12632 15191
rect 12688 15135 12756 15191
rect 12812 15135 12880 15191
rect 12936 15135 13004 15191
rect 13060 15135 13070 15191
rect 12622 15067 13070 15135
rect 12622 15011 12632 15067
rect 12688 15011 12756 15067
rect 12812 15011 12880 15067
rect 12936 15011 13004 15067
rect 13060 15011 13070 15067
rect 12622 14943 13070 15011
rect 12622 14887 12632 14943
rect 12688 14887 12756 14943
rect 12812 14887 12880 14943
rect 12936 14887 13004 14943
rect 13060 14887 13070 14943
rect 12622 14819 13070 14887
rect 12622 14763 12632 14819
rect 12688 14763 12756 14819
rect 12812 14763 12880 14819
rect 12936 14763 13004 14819
rect 13060 14763 13070 14819
rect 12622 14695 13070 14763
rect 12622 14639 12632 14695
rect 12688 14639 12756 14695
rect 12812 14639 12880 14695
rect 12936 14639 13004 14695
rect 13060 14639 13070 14695
rect 12622 14571 13070 14639
rect 12622 14515 12632 14571
rect 12688 14515 12756 14571
rect 12812 14515 12880 14571
rect 12936 14515 13004 14571
rect 13060 14515 13070 14571
rect 12622 14447 13070 14515
rect 12622 14391 12632 14447
rect 12688 14391 12756 14447
rect 12812 14391 12880 14447
rect 12936 14391 13004 14447
rect 13060 14391 13070 14447
rect 12622 14323 13070 14391
rect 12622 14267 12632 14323
rect 12688 14267 12756 14323
rect 12812 14267 12880 14323
rect 12936 14267 13004 14323
rect 13060 14267 13070 14323
rect 12622 14199 13070 14267
rect 12622 14143 12632 14199
rect 12688 14143 12756 14199
rect 12812 14143 12880 14199
rect 12936 14143 13004 14199
rect 13060 14143 13070 14199
rect 12622 14133 13070 14143
rect 13758 17051 14206 17061
rect 13758 16995 13768 17051
rect 13824 16995 13892 17051
rect 13948 16995 14016 17051
rect 14072 16995 14140 17051
rect 14196 16995 14206 17051
rect 13758 16927 14206 16995
rect 13758 16871 13768 16927
rect 13824 16871 13892 16927
rect 13948 16871 14016 16927
rect 14072 16871 14140 16927
rect 14196 16871 14206 16927
rect 13758 16803 14206 16871
rect 13758 16747 13768 16803
rect 13824 16747 13892 16803
rect 13948 16747 14016 16803
rect 14072 16747 14140 16803
rect 14196 16747 14206 16803
rect 13758 16679 14206 16747
rect 13758 16623 13768 16679
rect 13824 16623 13892 16679
rect 13948 16623 14016 16679
rect 14072 16623 14140 16679
rect 14196 16623 14206 16679
rect 13758 16555 14206 16623
rect 13758 16499 13768 16555
rect 13824 16499 13892 16555
rect 13948 16499 14016 16555
rect 14072 16499 14140 16555
rect 14196 16499 14206 16555
rect 13758 16431 14206 16499
rect 13758 16375 13768 16431
rect 13824 16375 13892 16431
rect 13948 16375 14016 16431
rect 14072 16375 14140 16431
rect 14196 16375 14206 16431
rect 13758 16307 14206 16375
rect 13758 16251 13768 16307
rect 13824 16251 13892 16307
rect 13948 16251 14016 16307
rect 14072 16251 14140 16307
rect 14196 16251 14206 16307
rect 13758 16183 14206 16251
rect 13758 16127 13768 16183
rect 13824 16127 13892 16183
rect 13948 16127 14016 16183
rect 14072 16127 14140 16183
rect 14196 16127 14206 16183
rect 13758 16059 14206 16127
rect 13758 16003 13768 16059
rect 13824 16003 13892 16059
rect 13948 16003 14016 16059
rect 14072 16003 14140 16059
rect 14196 16003 14206 16059
rect 13758 15935 14206 16003
rect 13758 15879 13768 15935
rect 13824 15879 13892 15935
rect 13948 15879 14016 15935
rect 14072 15879 14140 15935
rect 14196 15879 14206 15935
rect 13758 15811 14206 15879
rect 13758 15755 13768 15811
rect 13824 15755 13892 15811
rect 13948 15755 14016 15811
rect 14072 15755 14140 15811
rect 14196 15755 14206 15811
rect 13758 15687 14206 15755
rect 13758 15631 13768 15687
rect 13824 15631 13892 15687
rect 13948 15631 14016 15687
rect 14072 15631 14140 15687
rect 14196 15631 14206 15687
rect 13758 15563 14206 15631
rect 13758 15507 13768 15563
rect 13824 15507 13892 15563
rect 13948 15507 14016 15563
rect 14072 15507 14140 15563
rect 14196 15507 14206 15563
rect 13758 15439 14206 15507
rect 13758 15383 13768 15439
rect 13824 15383 13892 15439
rect 13948 15383 14016 15439
rect 14072 15383 14140 15439
rect 14196 15383 14206 15439
rect 13758 15315 14206 15383
rect 13758 15259 13768 15315
rect 13824 15259 13892 15315
rect 13948 15259 14016 15315
rect 14072 15259 14140 15315
rect 14196 15259 14206 15315
rect 13758 15191 14206 15259
rect 13758 15135 13768 15191
rect 13824 15135 13892 15191
rect 13948 15135 14016 15191
rect 14072 15135 14140 15191
rect 14196 15135 14206 15191
rect 13758 15067 14206 15135
rect 13758 15011 13768 15067
rect 13824 15011 13892 15067
rect 13948 15011 14016 15067
rect 14072 15011 14140 15067
rect 14196 15011 14206 15067
rect 13758 14943 14206 15011
rect 13758 14887 13768 14943
rect 13824 14887 13892 14943
rect 13948 14887 14016 14943
rect 14072 14887 14140 14943
rect 14196 14887 14206 14943
rect 13758 14819 14206 14887
rect 13758 14763 13768 14819
rect 13824 14763 13892 14819
rect 13948 14763 14016 14819
rect 14072 14763 14140 14819
rect 14196 14763 14206 14819
rect 13758 14695 14206 14763
rect 13758 14639 13768 14695
rect 13824 14639 13892 14695
rect 13948 14639 14016 14695
rect 14072 14639 14140 14695
rect 14196 14639 14206 14695
rect 13758 14571 14206 14639
rect 13758 14515 13768 14571
rect 13824 14515 13892 14571
rect 13948 14515 14016 14571
rect 14072 14515 14140 14571
rect 14196 14515 14206 14571
rect 13758 14447 14206 14515
rect 13758 14391 13768 14447
rect 13824 14391 13892 14447
rect 13948 14391 14016 14447
rect 14072 14391 14140 14447
rect 14196 14391 14206 14447
rect 13758 14323 14206 14391
rect 13758 14267 13768 14323
rect 13824 14267 13892 14323
rect 13948 14267 14016 14323
rect 14072 14267 14140 14323
rect 14196 14267 14206 14323
rect 13758 14199 14206 14267
rect 13758 14143 13768 14199
rect 13824 14143 13892 14199
rect 13948 14143 14016 14199
rect 14072 14143 14140 14199
rect 14196 14143 14206 14199
rect 13758 14133 14206 14143
rect 290 13845 738 13855
rect 290 13789 300 13845
rect 356 13789 424 13845
rect 480 13789 548 13845
rect 604 13789 672 13845
rect 728 13789 738 13845
rect 290 13721 738 13789
rect 290 13665 300 13721
rect 356 13665 424 13721
rect 480 13665 548 13721
rect 604 13665 672 13721
rect 728 13665 738 13721
rect 290 13597 738 13665
rect 290 13541 300 13597
rect 356 13541 424 13597
rect 480 13541 548 13597
rect 604 13541 672 13597
rect 728 13541 738 13597
rect 290 13473 738 13541
rect 290 13417 300 13473
rect 356 13417 424 13473
rect 480 13417 548 13473
rect 604 13417 672 13473
rect 728 13417 738 13473
rect 290 13349 738 13417
rect 290 13293 300 13349
rect 356 13293 424 13349
rect 480 13293 548 13349
rect 604 13293 672 13349
rect 728 13293 738 13349
rect 290 13225 738 13293
rect 290 13169 300 13225
rect 356 13169 424 13225
rect 480 13169 548 13225
rect 604 13169 672 13225
rect 728 13169 738 13225
rect 290 13101 738 13169
rect 290 13045 300 13101
rect 356 13045 424 13101
rect 480 13045 548 13101
rect 604 13045 672 13101
rect 728 13045 738 13101
rect 290 12977 738 13045
rect 290 12921 300 12977
rect 356 12921 424 12977
rect 480 12921 548 12977
rect 604 12921 672 12977
rect 728 12921 738 12977
rect 290 12853 738 12921
rect 290 12797 300 12853
rect 356 12797 424 12853
rect 480 12797 548 12853
rect 604 12797 672 12853
rect 728 12797 738 12853
rect 290 12729 738 12797
rect 290 12673 300 12729
rect 356 12673 424 12729
rect 480 12673 548 12729
rect 604 12673 672 12729
rect 728 12673 738 12729
rect 290 12605 738 12673
rect 290 12549 300 12605
rect 356 12549 424 12605
rect 480 12549 548 12605
rect 604 12549 672 12605
rect 728 12549 738 12605
rect 290 12539 738 12549
rect 1426 13845 1874 13855
rect 1426 13789 1436 13845
rect 1492 13789 1560 13845
rect 1616 13789 1684 13845
rect 1740 13789 1808 13845
rect 1864 13789 1874 13845
rect 1426 13721 1874 13789
rect 1426 13665 1436 13721
rect 1492 13665 1560 13721
rect 1616 13665 1684 13721
rect 1740 13665 1808 13721
rect 1864 13665 1874 13721
rect 1426 13597 1874 13665
rect 1426 13541 1436 13597
rect 1492 13541 1560 13597
rect 1616 13541 1684 13597
rect 1740 13541 1808 13597
rect 1864 13541 1874 13597
rect 1426 13473 1874 13541
rect 1426 13417 1436 13473
rect 1492 13417 1560 13473
rect 1616 13417 1684 13473
rect 1740 13417 1808 13473
rect 1864 13417 1874 13473
rect 1426 13349 1874 13417
rect 1426 13293 1436 13349
rect 1492 13293 1560 13349
rect 1616 13293 1684 13349
rect 1740 13293 1808 13349
rect 1864 13293 1874 13349
rect 1426 13225 1874 13293
rect 1426 13169 1436 13225
rect 1492 13169 1560 13225
rect 1616 13169 1684 13225
rect 1740 13169 1808 13225
rect 1864 13169 1874 13225
rect 1426 13101 1874 13169
rect 1426 13045 1436 13101
rect 1492 13045 1560 13101
rect 1616 13045 1684 13101
rect 1740 13045 1808 13101
rect 1864 13045 1874 13101
rect 1426 12977 1874 13045
rect 1426 12921 1436 12977
rect 1492 12921 1560 12977
rect 1616 12921 1684 12977
rect 1740 12921 1808 12977
rect 1864 12921 1874 12977
rect 1426 12853 1874 12921
rect 1426 12797 1436 12853
rect 1492 12797 1560 12853
rect 1616 12797 1684 12853
rect 1740 12797 1808 12853
rect 1864 12797 1874 12853
rect 1426 12729 1874 12797
rect 1426 12673 1436 12729
rect 1492 12673 1560 12729
rect 1616 12673 1684 12729
rect 1740 12673 1808 12729
rect 1864 12673 1874 12729
rect 1426 12605 1874 12673
rect 1426 12549 1436 12605
rect 1492 12549 1560 12605
rect 1616 12549 1684 12605
rect 1740 12549 1808 12605
rect 1864 12549 1874 12605
rect 1426 12539 1874 12549
rect 2562 13845 3010 13855
rect 2562 13789 2572 13845
rect 2628 13789 2696 13845
rect 2752 13789 2820 13845
rect 2876 13789 2944 13845
rect 3000 13789 3010 13845
rect 2562 13721 3010 13789
rect 2562 13665 2572 13721
rect 2628 13665 2696 13721
rect 2752 13665 2820 13721
rect 2876 13665 2944 13721
rect 3000 13665 3010 13721
rect 2562 13597 3010 13665
rect 2562 13541 2572 13597
rect 2628 13541 2696 13597
rect 2752 13541 2820 13597
rect 2876 13541 2944 13597
rect 3000 13541 3010 13597
rect 2562 13473 3010 13541
rect 2562 13417 2572 13473
rect 2628 13417 2696 13473
rect 2752 13417 2820 13473
rect 2876 13417 2944 13473
rect 3000 13417 3010 13473
rect 2562 13349 3010 13417
rect 2562 13293 2572 13349
rect 2628 13293 2696 13349
rect 2752 13293 2820 13349
rect 2876 13293 2944 13349
rect 3000 13293 3010 13349
rect 2562 13225 3010 13293
rect 2562 13169 2572 13225
rect 2628 13169 2696 13225
rect 2752 13169 2820 13225
rect 2876 13169 2944 13225
rect 3000 13169 3010 13225
rect 2562 13101 3010 13169
rect 2562 13045 2572 13101
rect 2628 13045 2696 13101
rect 2752 13045 2820 13101
rect 2876 13045 2944 13101
rect 3000 13045 3010 13101
rect 2562 12977 3010 13045
rect 2562 12921 2572 12977
rect 2628 12921 2696 12977
rect 2752 12921 2820 12977
rect 2876 12921 2944 12977
rect 3000 12921 3010 12977
rect 2562 12853 3010 12921
rect 2562 12797 2572 12853
rect 2628 12797 2696 12853
rect 2752 12797 2820 12853
rect 2876 12797 2944 12853
rect 3000 12797 3010 12853
rect 2562 12729 3010 12797
rect 2562 12673 2572 12729
rect 2628 12673 2696 12729
rect 2752 12673 2820 12729
rect 2876 12673 2944 12729
rect 3000 12673 3010 12729
rect 2562 12605 3010 12673
rect 2562 12549 2572 12605
rect 2628 12549 2696 12605
rect 2752 12549 2820 12605
rect 2876 12549 2944 12605
rect 3000 12549 3010 12605
rect 2562 12539 3010 12549
rect 4834 13845 5282 13855
rect 4834 13789 4844 13845
rect 4900 13789 4968 13845
rect 5024 13789 5092 13845
rect 5148 13789 5216 13845
rect 5272 13789 5282 13845
rect 4834 13721 5282 13789
rect 4834 13665 4844 13721
rect 4900 13665 4968 13721
rect 5024 13665 5092 13721
rect 5148 13665 5216 13721
rect 5272 13665 5282 13721
rect 4834 13597 5282 13665
rect 4834 13541 4844 13597
rect 4900 13541 4968 13597
rect 5024 13541 5092 13597
rect 5148 13541 5216 13597
rect 5272 13541 5282 13597
rect 4834 13473 5282 13541
rect 4834 13417 4844 13473
rect 4900 13417 4968 13473
rect 5024 13417 5092 13473
rect 5148 13417 5216 13473
rect 5272 13417 5282 13473
rect 4834 13349 5282 13417
rect 4834 13293 4844 13349
rect 4900 13293 4968 13349
rect 5024 13293 5092 13349
rect 5148 13293 5216 13349
rect 5272 13293 5282 13349
rect 4834 13225 5282 13293
rect 4834 13169 4844 13225
rect 4900 13169 4968 13225
rect 5024 13169 5092 13225
rect 5148 13169 5216 13225
rect 5272 13169 5282 13225
rect 4834 13101 5282 13169
rect 4834 13045 4844 13101
rect 4900 13045 4968 13101
rect 5024 13045 5092 13101
rect 5148 13045 5216 13101
rect 5272 13045 5282 13101
rect 4834 12977 5282 13045
rect 4834 12921 4844 12977
rect 4900 12921 4968 12977
rect 5024 12921 5092 12977
rect 5148 12921 5216 12977
rect 5272 12921 5282 12977
rect 4834 12853 5282 12921
rect 4834 12797 4844 12853
rect 4900 12797 4968 12853
rect 5024 12797 5092 12853
rect 5148 12797 5216 12853
rect 5272 12797 5282 12853
rect 4834 12729 5282 12797
rect 4834 12673 4844 12729
rect 4900 12673 4968 12729
rect 5024 12673 5092 12729
rect 5148 12673 5216 12729
rect 5272 12673 5282 12729
rect 4834 12605 5282 12673
rect 4834 12549 4844 12605
rect 4900 12549 4968 12605
rect 5024 12549 5092 12605
rect 5148 12549 5216 12605
rect 5272 12549 5282 12605
rect 4834 12539 5282 12549
rect 7127 13845 7451 13855
rect 7127 13789 7137 13845
rect 7193 13789 7261 13845
rect 7317 13789 7385 13845
rect 7441 13789 7451 13845
rect 7127 13721 7451 13789
rect 7127 13665 7137 13721
rect 7193 13665 7261 13721
rect 7317 13665 7385 13721
rect 7441 13665 7451 13721
rect 7127 13597 7451 13665
rect 7127 13541 7137 13597
rect 7193 13541 7261 13597
rect 7317 13541 7385 13597
rect 7441 13541 7451 13597
rect 7127 13473 7451 13541
rect 7127 13417 7137 13473
rect 7193 13417 7261 13473
rect 7317 13417 7385 13473
rect 7441 13417 7451 13473
rect 7127 13349 7451 13417
rect 7127 13293 7137 13349
rect 7193 13293 7261 13349
rect 7317 13293 7385 13349
rect 7441 13293 7451 13349
rect 7127 13225 7451 13293
rect 7127 13169 7137 13225
rect 7193 13169 7261 13225
rect 7317 13169 7385 13225
rect 7441 13169 7451 13225
rect 7127 13101 7451 13169
rect 7127 13045 7137 13101
rect 7193 13045 7261 13101
rect 7317 13045 7385 13101
rect 7441 13045 7451 13101
rect 7127 12977 7451 13045
rect 7127 12921 7137 12977
rect 7193 12921 7261 12977
rect 7317 12921 7385 12977
rect 7441 12921 7451 12977
rect 7127 12853 7451 12921
rect 7127 12797 7137 12853
rect 7193 12797 7261 12853
rect 7317 12797 7385 12853
rect 7441 12797 7451 12853
rect 7127 12729 7451 12797
rect 7127 12673 7137 12729
rect 7193 12673 7261 12729
rect 7317 12673 7385 12729
rect 7441 12673 7451 12729
rect 7127 12605 7451 12673
rect 7127 12549 7137 12605
rect 7193 12549 7261 12605
rect 7317 12549 7385 12605
rect 7441 12549 7451 12605
rect 7127 12539 7451 12549
rect 7613 13845 7937 13855
rect 7613 13789 7623 13845
rect 7679 13789 7747 13845
rect 7803 13789 7871 13845
rect 7927 13789 7937 13845
rect 7613 13721 7937 13789
rect 7613 13665 7623 13721
rect 7679 13665 7747 13721
rect 7803 13665 7871 13721
rect 7927 13665 7937 13721
rect 7613 13597 7937 13665
rect 7613 13541 7623 13597
rect 7679 13541 7747 13597
rect 7803 13541 7871 13597
rect 7927 13541 7937 13597
rect 7613 13473 7937 13541
rect 7613 13417 7623 13473
rect 7679 13417 7747 13473
rect 7803 13417 7871 13473
rect 7927 13417 7937 13473
rect 7613 13349 7937 13417
rect 7613 13293 7623 13349
rect 7679 13293 7747 13349
rect 7803 13293 7871 13349
rect 7927 13293 7937 13349
rect 7613 13225 7937 13293
rect 7613 13169 7623 13225
rect 7679 13169 7747 13225
rect 7803 13169 7871 13225
rect 7927 13169 7937 13225
rect 7613 13101 7937 13169
rect 7613 13045 7623 13101
rect 7679 13045 7747 13101
rect 7803 13045 7871 13101
rect 7927 13045 7937 13101
rect 7613 12977 7937 13045
rect 7613 12921 7623 12977
rect 7679 12921 7747 12977
rect 7803 12921 7871 12977
rect 7927 12921 7937 12977
rect 7613 12853 7937 12921
rect 7613 12797 7623 12853
rect 7679 12797 7747 12853
rect 7803 12797 7871 12853
rect 7927 12797 7937 12853
rect 7613 12729 7937 12797
rect 7613 12673 7623 12729
rect 7679 12673 7747 12729
rect 7803 12673 7871 12729
rect 7927 12673 7937 12729
rect 7613 12605 7937 12673
rect 7613 12549 7623 12605
rect 7679 12549 7747 12605
rect 7803 12549 7871 12605
rect 7927 12549 7937 12605
rect 7613 12539 7937 12549
rect 9782 13845 10230 13855
rect 9782 13789 9792 13845
rect 9848 13789 9916 13845
rect 9972 13789 10040 13845
rect 10096 13789 10164 13845
rect 10220 13789 10230 13845
rect 9782 13721 10230 13789
rect 9782 13665 9792 13721
rect 9848 13665 9916 13721
rect 9972 13665 10040 13721
rect 10096 13665 10164 13721
rect 10220 13665 10230 13721
rect 9782 13597 10230 13665
rect 9782 13541 9792 13597
rect 9848 13541 9916 13597
rect 9972 13541 10040 13597
rect 10096 13541 10164 13597
rect 10220 13541 10230 13597
rect 9782 13473 10230 13541
rect 9782 13417 9792 13473
rect 9848 13417 9916 13473
rect 9972 13417 10040 13473
rect 10096 13417 10164 13473
rect 10220 13417 10230 13473
rect 9782 13349 10230 13417
rect 9782 13293 9792 13349
rect 9848 13293 9916 13349
rect 9972 13293 10040 13349
rect 10096 13293 10164 13349
rect 10220 13293 10230 13349
rect 9782 13225 10230 13293
rect 9782 13169 9792 13225
rect 9848 13169 9916 13225
rect 9972 13169 10040 13225
rect 10096 13169 10164 13225
rect 10220 13169 10230 13225
rect 9782 13101 10230 13169
rect 9782 13045 9792 13101
rect 9848 13045 9916 13101
rect 9972 13045 10040 13101
rect 10096 13045 10164 13101
rect 10220 13045 10230 13101
rect 9782 12977 10230 13045
rect 9782 12921 9792 12977
rect 9848 12921 9916 12977
rect 9972 12921 10040 12977
rect 10096 12921 10164 12977
rect 10220 12921 10230 12977
rect 9782 12853 10230 12921
rect 9782 12797 9792 12853
rect 9848 12797 9916 12853
rect 9972 12797 10040 12853
rect 10096 12797 10164 12853
rect 10220 12797 10230 12853
rect 9782 12729 10230 12797
rect 9782 12673 9792 12729
rect 9848 12673 9916 12729
rect 9972 12673 10040 12729
rect 10096 12673 10164 12729
rect 10220 12673 10230 12729
rect 9782 12605 10230 12673
rect 9782 12549 9792 12605
rect 9848 12549 9916 12605
rect 9972 12549 10040 12605
rect 10096 12549 10164 12605
rect 10220 12549 10230 12605
rect 9782 12539 10230 12549
rect 12054 13845 12502 13855
rect 12054 13789 12064 13845
rect 12120 13789 12188 13845
rect 12244 13789 12312 13845
rect 12368 13789 12436 13845
rect 12492 13789 12502 13845
rect 12054 13721 12502 13789
rect 12054 13665 12064 13721
rect 12120 13665 12188 13721
rect 12244 13665 12312 13721
rect 12368 13665 12436 13721
rect 12492 13665 12502 13721
rect 12054 13597 12502 13665
rect 12054 13541 12064 13597
rect 12120 13541 12188 13597
rect 12244 13541 12312 13597
rect 12368 13541 12436 13597
rect 12492 13541 12502 13597
rect 12054 13473 12502 13541
rect 12054 13417 12064 13473
rect 12120 13417 12188 13473
rect 12244 13417 12312 13473
rect 12368 13417 12436 13473
rect 12492 13417 12502 13473
rect 12054 13349 12502 13417
rect 12054 13293 12064 13349
rect 12120 13293 12188 13349
rect 12244 13293 12312 13349
rect 12368 13293 12436 13349
rect 12492 13293 12502 13349
rect 12054 13225 12502 13293
rect 12054 13169 12064 13225
rect 12120 13169 12188 13225
rect 12244 13169 12312 13225
rect 12368 13169 12436 13225
rect 12492 13169 12502 13225
rect 12054 13101 12502 13169
rect 12054 13045 12064 13101
rect 12120 13045 12188 13101
rect 12244 13045 12312 13101
rect 12368 13045 12436 13101
rect 12492 13045 12502 13101
rect 12054 12977 12502 13045
rect 12054 12921 12064 12977
rect 12120 12921 12188 12977
rect 12244 12921 12312 12977
rect 12368 12921 12436 12977
rect 12492 12921 12502 12977
rect 12054 12853 12502 12921
rect 12054 12797 12064 12853
rect 12120 12797 12188 12853
rect 12244 12797 12312 12853
rect 12368 12797 12436 12853
rect 12492 12797 12502 12853
rect 12054 12729 12502 12797
rect 12054 12673 12064 12729
rect 12120 12673 12188 12729
rect 12244 12673 12312 12729
rect 12368 12673 12436 12729
rect 12492 12673 12502 12729
rect 12054 12605 12502 12673
rect 12054 12549 12064 12605
rect 12120 12549 12188 12605
rect 12244 12549 12312 12605
rect 12368 12549 12436 12605
rect 12492 12549 12502 12605
rect 12054 12539 12502 12549
rect 13190 13845 13638 13855
rect 13190 13789 13200 13845
rect 13256 13789 13324 13845
rect 13380 13789 13448 13845
rect 13504 13789 13572 13845
rect 13628 13789 13638 13845
rect 13190 13721 13638 13789
rect 13190 13665 13200 13721
rect 13256 13665 13324 13721
rect 13380 13665 13448 13721
rect 13504 13665 13572 13721
rect 13628 13665 13638 13721
rect 13190 13597 13638 13665
rect 13190 13541 13200 13597
rect 13256 13541 13324 13597
rect 13380 13541 13448 13597
rect 13504 13541 13572 13597
rect 13628 13541 13638 13597
rect 13190 13473 13638 13541
rect 13190 13417 13200 13473
rect 13256 13417 13324 13473
rect 13380 13417 13448 13473
rect 13504 13417 13572 13473
rect 13628 13417 13638 13473
rect 13190 13349 13638 13417
rect 13190 13293 13200 13349
rect 13256 13293 13324 13349
rect 13380 13293 13448 13349
rect 13504 13293 13572 13349
rect 13628 13293 13638 13349
rect 13190 13225 13638 13293
rect 13190 13169 13200 13225
rect 13256 13169 13324 13225
rect 13380 13169 13448 13225
rect 13504 13169 13572 13225
rect 13628 13169 13638 13225
rect 13190 13101 13638 13169
rect 13190 13045 13200 13101
rect 13256 13045 13324 13101
rect 13380 13045 13448 13101
rect 13504 13045 13572 13101
rect 13628 13045 13638 13101
rect 13190 12977 13638 13045
rect 13190 12921 13200 12977
rect 13256 12921 13324 12977
rect 13380 12921 13448 12977
rect 13504 12921 13572 12977
rect 13628 12921 13638 12977
rect 13190 12853 13638 12921
rect 13190 12797 13200 12853
rect 13256 12797 13324 12853
rect 13380 12797 13448 12853
rect 13504 12797 13572 12853
rect 13628 12797 13638 12853
rect 13190 12729 13638 12797
rect 13190 12673 13200 12729
rect 13256 12673 13324 12729
rect 13380 12673 13448 12729
rect 13504 12673 13572 12729
rect 13628 12673 13638 12729
rect 13190 12605 13638 12673
rect 13190 12549 13200 12605
rect 13256 12549 13324 12605
rect 13380 12549 13448 12605
rect 13504 12549 13572 12605
rect 13628 12549 13638 12605
rect 13190 12539 13638 12549
rect 14326 13845 14774 13855
rect 14326 13789 14336 13845
rect 14392 13789 14460 13845
rect 14516 13789 14584 13845
rect 14640 13789 14708 13845
rect 14764 13789 14774 13845
rect 14326 13721 14774 13789
rect 14326 13665 14336 13721
rect 14392 13665 14460 13721
rect 14516 13665 14584 13721
rect 14640 13665 14708 13721
rect 14764 13665 14774 13721
rect 14326 13597 14774 13665
rect 14326 13541 14336 13597
rect 14392 13541 14460 13597
rect 14516 13541 14584 13597
rect 14640 13541 14708 13597
rect 14764 13541 14774 13597
rect 14326 13473 14774 13541
rect 14326 13417 14336 13473
rect 14392 13417 14460 13473
rect 14516 13417 14584 13473
rect 14640 13417 14708 13473
rect 14764 13417 14774 13473
rect 14326 13349 14774 13417
rect 14326 13293 14336 13349
rect 14392 13293 14460 13349
rect 14516 13293 14584 13349
rect 14640 13293 14708 13349
rect 14764 13293 14774 13349
rect 14326 13225 14774 13293
rect 14326 13169 14336 13225
rect 14392 13169 14460 13225
rect 14516 13169 14584 13225
rect 14640 13169 14708 13225
rect 14764 13169 14774 13225
rect 14326 13101 14774 13169
rect 14326 13045 14336 13101
rect 14392 13045 14460 13101
rect 14516 13045 14584 13101
rect 14640 13045 14708 13101
rect 14764 13045 14774 13101
rect 14326 12977 14774 13045
rect 14326 12921 14336 12977
rect 14392 12921 14460 12977
rect 14516 12921 14584 12977
rect 14640 12921 14708 12977
rect 14764 12921 14774 12977
rect 14326 12853 14774 12921
rect 14326 12797 14336 12853
rect 14392 12797 14460 12853
rect 14516 12797 14584 12853
rect 14640 12797 14708 12853
rect 14764 12797 14774 12853
rect 14326 12729 14774 12797
rect 14326 12673 14336 12729
rect 14392 12673 14460 12729
rect 14516 12673 14584 12729
rect 14640 12673 14708 12729
rect 14764 12673 14774 12729
rect 14326 12605 14774 12673
rect 14326 12549 14336 12605
rect 14392 12549 14460 12605
rect 14516 12549 14584 12605
rect 14640 12549 14708 12605
rect 14764 12549 14774 12605
rect 14326 12539 14774 12549
rect 858 12245 1306 12255
rect 858 12189 868 12245
rect 924 12189 992 12245
rect 1048 12189 1116 12245
rect 1172 12189 1240 12245
rect 1296 12189 1306 12245
rect 858 12121 1306 12189
rect 858 12065 868 12121
rect 924 12065 992 12121
rect 1048 12065 1116 12121
rect 1172 12065 1240 12121
rect 1296 12065 1306 12121
rect 858 11997 1306 12065
rect 858 11941 868 11997
rect 924 11941 992 11997
rect 1048 11941 1116 11997
rect 1172 11941 1240 11997
rect 1296 11941 1306 11997
rect 858 11873 1306 11941
rect 858 11817 868 11873
rect 924 11817 992 11873
rect 1048 11817 1116 11873
rect 1172 11817 1240 11873
rect 1296 11817 1306 11873
rect 858 11749 1306 11817
rect 858 11693 868 11749
rect 924 11693 992 11749
rect 1048 11693 1116 11749
rect 1172 11693 1240 11749
rect 1296 11693 1306 11749
rect 858 11625 1306 11693
rect 858 11569 868 11625
rect 924 11569 992 11625
rect 1048 11569 1116 11625
rect 1172 11569 1240 11625
rect 1296 11569 1306 11625
rect 858 11501 1306 11569
rect 858 11445 868 11501
rect 924 11445 992 11501
rect 1048 11445 1116 11501
rect 1172 11445 1240 11501
rect 1296 11445 1306 11501
rect 858 11377 1306 11445
rect 858 11321 868 11377
rect 924 11321 992 11377
rect 1048 11321 1116 11377
rect 1172 11321 1240 11377
rect 1296 11321 1306 11377
rect 858 11253 1306 11321
rect 858 11197 868 11253
rect 924 11197 992 11253
rect 1048 11197 1116 11253
rect 1172 11197 1240 11253
rect 1296 11197 1306 11253
rect 858 11129 1306 11197
rect 858 11073 868 11129
rect 924 11073 992 11129
rect 1048 11073 1116 11129
rect 1172 11073 1240 11129
rect 1296 11073 1306 11129
rect 858 11005 1306 11073
rect 858 10949 868 11005
rect 924 10949 992 11005
rect 1048 10949 1116 11005
rect 1172 10949 1240 11005
rect 1296 10949 1306 11005
rect 858 10939 1306 10949
rect 1994 12245 2442 12255
rect 1994 12189 2004 12245
rect 2060 12189 2128 12245
rect 2184 12189 2252 12245
rect 2308 12189 2376 12245
rect 2432 12189 2442 12245
rect 1994 12121 2442 12189
rect 1994 12065 2004 12121
rect 2060 12065 2128 12121
rect 2184 12065 2252 12121
rect 2308 12065 2376 12121
rect 2432 12065 2442 12121
rect 1994 11997 2442 12065
rect 1994 11941 2004 11997
rect 2060 11941 2128 11997
rect 2184 11941 2252 11997
rect 2308 11941 2376 11997
rect 2432 11941 2442 11997
rect 1994 11873 2442 11941
rect 1994 11817 2004 11873
rect 2060 11817 2128 11873
rect 2184 11817 2252 11873
rect 2308 11817 2376 11873
rect 2432 11817 2442 11873
rect 1994 11749 2442 11817
rect 1994 11693 2004 11749
rect 2060 11693 2128 11749
rect 2184 11693 2252 11749
rect 2308 11693 2376 11749
rect 2432 11693 2442 11749
rect 1994 11625 2442 11693
rect 1994 11569 2004 11625
rect 2060 11569 2128 11625
rect 2184 11569 2252 11625
rect 2308 11569 2376 11625
rect 2432 11569 2442 11625
rect 1994 11501 2442 11569
rect 1994 11445 2004 11501
rect 2060 11445 2128 11501
rect 2184 11445 2252 11501
rect 2308 11445 2376 11501
rect 2432 11445 2442 11501
rect 1994 11377 2442 11445
rect 1994 11321 2004 11377
rect 2060 11321 2128 11377
rect 2184 11321 2252 11377
rect 2308 11321 2376 11377
rect 2432 11321 2442 11377
rect 1994 11253 2442 11321
rect 1994 11197 2004 11253
rect 2060 11197 2128 11253
rect 2184 11197 2252 11253
rect 2308 11197 2376 11253
rect 2432 11197 2442 11253
rect 1994 11129 2442 11197
rect 1994 11073 2004 11129
rect 2060 11073 2128 11129
rect 2184 11073 2252 11129
rect 2308 11073 2376 11129
rect 2432 11073 2442 11129
rect 1994 11005 2442 11073
rect 1994 10949 2004 11005
rect 2060 10949 2128 11005
rect 2184 10949 2252 11005
rect 2308 10949 2376 11005
rect 2432 10949 2442 11005
rect 1994 10939 2442 10949
rect 3698 12245 4146 12255
rect 3698 12189 3708 12245
rect 3764 12189 3832 12245
rect 3888 12189 3956 12245
rect 4012 12189 4080 12245
rect 4136 12189 4146 12245
rect 3698 12121 4146 12189
rect 3698 12065 3708 12121
rect 3764 12065 3832 12121
rect 3888 12065 3956 12121
rect 4012 12065 4080 12121
rect 4136 12065 4146 12121
rect 3698 11997 4146 12065
rect 3698 11941 3708 11997
rect 3764 11941 3832 11997
rect 3888 11941 3956 11997
rect 4012 11941 4080 11997
rect 4136 11941 4146 11997
rect 3698 11873 4146 11941
rect 3698 11817 3708 11873
rect 3764 11817 3832 11873
rect 3888 11817 3956 11873
rect 4012 11817 4080 11873
rect 4136 11817 4146 11873
rect 3698 11749 4146 11817
rect 3698 11693 3708 11749
rect 3764 11693 3832 11749
rect 3888 11693 3956 11749
rect 4012 11693 4080 11749
rect 4136 11693 4146 11749
rect 3698 11625 4146 11693
rect 3698 11569 3708 11625
rect 3764 11569 3832 11625
rect 3888 11569 3956 11625
rect 4012 11569 4080 11625
rect 4136 11569 4146 11625
rect 3698 11501 4146 11569
rect 3698 11445 3708 11501
rect 3764 11445 3832 11501
rect 3888 11445 3956 11501
rect 4012 11445 4080 11501
rect 4136 11445 4146 11501
rect 3698 11377 4146 11445
rect 3698 11321 3708 11377
rect 3764 11321 3832 11377
rect 3888 11321 3956 11377
rect 4012 11321 4080 11377
rect 4136 11321 4146 11377
rect 3698 11253 4146 11321
rect 3698 11197 3708 11253
rect 3764 11197 3832 11253
rect 3888 11197 3956 11253
rect 4012 11197 4080 11253
rect 4136 11197 4146 11253
rect 3698 11129 4146 11197
rect 3698 11073 3708 11129
rect 3764 11073 3832 11129
rect 3888 11073 3956 11129
rect 4012 11073 4080 11129
rect 4136 11073 4146 11129
rect 3698 11005 4146 11073
rect 3698 10949 3708 11005
rect 3764 10949 3832 11005
rect 3888 10949 3956 11005
rect 4012 10949 4080 11005
rect 4136 10949 4146 11005
rect 3698 10939 4146 10949
rect 5970 12245 6418 12255
rect 5970 12189 5980 12245
rect 6036 12189 6104 12245
rect 6160 12189 6228 12245
rect 6284 12189 6352 12245
rect 6408 12189 6418 12245
rect 5970 12121 6418 12189
rect 5970 12065 5980 12121
rect 6036 12065 6104 12121
rect 6160 12065 6228 12121
rect 6284 12065 6352 12121
rect 6408 12065 6418 12121
rect 5970 11997 6418 12065
rect 5970 11941 5980 11997
rect 6036 11941 6104 11997
rect 6160 11941 6228 11997
rect 6284 11941 6352 11997
rect 6408 11941 6418 11997
rect 5970 11873 6418 11941
rect 5970 11817 5980 11873
rect 6036 11817 6104 11873
rect 6160 11817 6228 11873
rect 6284 11817 6352 11873
rect 6408 11817 6418 11873
rect 5970 11749 6418 11817
rect 5970 11693 5980 11749
rect 6036 11693 6104 11749
rect 6160 11693 6228 11749
rect 6284 11693 6352 11749
rect 6408 11693 6418 11749
rect 5970 11625 6418 11693
rect 5970 11569 5980 11625
rect 6036 11569 6104 11625
rect 6160 11569 6228 11625
rect 6284 11569 6352 11625
rect 6408 11569 6418 11625
rect 5970 11501 6418 11569
rect 5970 11445 5980 11501
rect 6036 11445 6104 11501
rect 6160 11445 6228 11501
rect 6284 11445 6352 11501
rect 6408 11445 6418 11501
rect 5970 11377 6418 11445
rect 5970 11321 5980 11377
rect 6036 11321 6104 11377
rect 6160 11321 6228 11377
rect 6284 11321 6352 11377
rect 6408 11321 6418 11377
rect 5970 11253 6418 11321
rect 5970 11197 5980 11253
rect 6036 11197 6104 11253
rect 6160 11197 6228 11253
rect 6284 11197 6352 11253
rect 6408 11197 6418 11253
rect 5970 11129 6418 11197
rect 5970 11073 5980 11129
rect 6036 11073 6104 11129
rect 6160 11073 6228 11129
rect 6284 11073 6352 11129
rect 6408 11073 6418 11129
rect 5970 11005 6418 11073
rect 5970 10949 5980 11005
rect 6036 10949 6104 11005
rect 6160 10949 6228 11005
rect 6284 10949 6352 11005
rect 6408 10949 6418 11005
rect 5970 10939 6418 10949
rect 8646 12245 9094 12255
rect 8646 12189 8656 12245
rect 8712 12189 8780 12245
rect 8836 12189 8904 12245
rect 8960 12189 9028 12245
rect 9084 12189 9094 12245
rect 8646 12121 9094 12189
rect 8646 12065 8656 12121
rect 8712 12065 8780 12121
rect 8836 12065 8904 12121
rect 8960 12065 9028 12121
rect 9084 12065 9094 12121
rect 8646 11997 9094 12065
rect 8646 11941 8656 11997
rect 8712 11941 8780 11997
rect 8836 11941 8904 11997
rect 8960 11941 9028 11997
rect 9084 11941 9094 11997
rect 8646 11873 9094 11941
rect 8646 11817 8656 11873
rect 8712 11817 8780 11873
rect 8836 11817 8904 11873
rect 8960 11817 9028 11873
rect 9084 11817 9094 11873
rect 8646 11749 9094 11817
rect 8646 11693 8656 11749
rect 8712 11693 8780 11749
rect 8836 11693 8904 11749
rect 8960 11693 9028 11749
rect 9084 11693 9094 11749
rect 8646 11625 9094 11693
rect 8646 11569 8656 11625
rect 8712 11569 8780 11625
rect 8836 11569 8904 11625
rect 8960 11569 9028 11625
rect 9084 11569 9094 11625
rect 8646 11501 9094 11569
rect 8646 11445 8656 11501
rect 8712 11445 8780 11501
rect 8836 11445 8904 11501
rect 8960 11445 9028 11501
rect 9084 11445 9094 11501
rect 8646 11377 9094 11445
rect 8646 11321 8656 11377
rect 8712 11321 8780 11377
rect 8836 11321 8904 11377
rect 8960 11321 9028 11377
rect 9084 11321 9094 11377
rect 8646 11253 9094 11321
rect 8646 11197 8656 11253
rect 8712 11197 8780 11253
rect 8836 11197 8904 11253
rect 8960 11197 9028 11253
rect 9084 11197 9094 11253
rect 8646 11129 9094 11197
rect 8646 11073 8656 11129
rect 8712 11073 8780 11129
rect 8836 11073 8904 11129
rect 8960 11073 9028 11129
rect 9084 11073 9094 11129
rect 8646 11005 9094 11073
rect 8646 10949 8656 11005
rect 8712 10949 8780 11005
rect 8836 10949 8904 11005
rect 8960 10949 9028 11005
rect 9084 10949 9094 11005
rect 8646 10939 9094 10949
rect 10918 12245 11366 12255
rect 10918 12189 10928 12245
rect 10984 12189 11052 12245
rect 11108 12189 11176 12245
rect 11232 12189 11300 12245
rect 11356 12189 11366 12245
rect 10918 12121 11366 12189
rect 10918 12065 10928 12121
rect 10984 12065 11052 12121
rect 11108 12065 11176 12121
rect 11232 12065 11300 12121
rect 11356 12065 11366 12121
rect 10918 11997 11366 12065
rect 10918 11941 10928 11997
rect 10984 11941 11052 11997
rect 11108 11941 11176 11997
rect 11232 11941 11300 11997
rect 11356 11941 11366 11997
rect 10918 11873 11366 11941
rect 10918 11817 10928 11873
rect 10984 11817 11052 11873
rect 11108 11817 11176 11873
rect 11232 11817 11300 11873
rect 11356 11817 11366 11873
rect 10918 11749 11366 11817
rect 10918 11693 10928 11749
rect 10984 11693 11052 11749
rect 11108 11693 11176 11749
rect 11232 11693 11300 11749
rect 11356 11693 11366 11749
rect 10918 11625 11366 11693
rect 10918 11569 10928 11625
rect 10984 11569 11052 11625
rect 11108 11569 11176 11625
rect 11232 11569 11300 11625
rect 11356 11569 11366 11625
rect 10918 11501 11366 11569
rect 10918 11445 10928 11501
rect 10984 11445 11052 11501
rect 11108 11445 11176 11501
rect 11232 11445 11300 11501
rect 11356 11445 11366 11501
rect 10918 11377 11366 11445
rect 10918 11321 10928 11377
rect 10984 11321 11052 11377
rect 11108 11321 11176 11377
rect 11232 11321 11300 11377
rect 11356 11321 11366 11377
rect 10918 11253 11366 11321
rect 10918 11197 10928 11253
rect 10984 11197 11052 11253
rect 11108 11197 11176 11253
rect 11232 11197 11300 11253
rect 11356 11197 11366 11253
rect 10918 11129 11366 11197
rect 10918 11073 10928 11129
rect 10984 11073 11052 11129
rect 11108 11073 11176 11129
rect 11232 11073 11300 11129
rect 11356 11073 11366 11129
rect 10918 11005 11366 11073
rect 10918 10949 10928 11005
rect 10984 10949 11052 11005
rect 11108 10949 11176 11005
rect 11232 10949 11300 11005
rect 11356 10949 11366 11005
rect 10918 10939 11366 10949
rect 12622 12245 13070 12255
rect 12622 12189 12632 12245
rect 12688 12189 12756 12245
rect 12812 12189 12880 12245
rect 12936 12189 13004 12245
rect 13060 12189 13070 12245
rect 12622 12121 13070 12189
rect 12622 12065 12632 12121
rect 12688 12065 12756 12121
rect 12812 12065 12880 12121
rect 12936 12065 13004 12121
rect 13060 12065 13070 12121
rect 12622 11997 13070 12065
rect 12622 11941 12632 11997
rect 12688 11941 12756 11997
rect 12812 11941 12880 11997
rect 12936 11941 13004 11997
rect 13060 11941 13070 11997
rect 12622 11873 13070 11941
rect 12622 11817 12632 11873
rect 12688 11817 12756 11873
rect 12812 11817 12880 11873
rect 12936 11817 13004 11873
rect 13060 11817 13070 11873
rect 12622 11749 13070 11817
rect 12622 11693 12632 11749
rect 12688 11693 12756 11749
rect 12812 11693 12880 11749
rect 12936 11693 13004 11749
rect 13060 11693 13070 11749
rect 12622 11625 13070 11693
rect 12622 11569 12632 11625
rect 12688 11569 12756 11625
rect 12812 11569 12880 11625
rect 12936 11569 13004 11625
rect 13060 11569 13070 11625
rect 12622 11501 13070 11569
rect 12622 11445 12632 11501
rect 12688 11445 12756 11501
rect 12812 11445 12880 11501
rect 12936 11445 13004 11501
rect 13060 11445 13070 11501
rect 12622 11377 13070 11445
rect 12622 11321 12632 11377
rect 12688 11321 12756 11377
rect 12812 11321 12880 11377
rect 12936 11321 13004 11377
rect 13060 11321 13070 11377
rect 12622 11253 13070 11321
rect 12622 11197 12632 11253
rect 12688 11197 12756 11253
rect 12812 11197 12880 11253
rect 12936 11197 13004 11253
rect 13060 11197 13070 11253
rect 12622 11129 13070 11197
rect 12622 11073 12632 11129
rect 12688 11073 12756 11129
rect 12812 11073 12880 11129
rect 12936 11073 13004 11129
rect 13060 11073 13070 11129
rect 12622 11005 13070 11073
rect 12622 10949 12632 11005
rect 12688 10949 12756 11005
rect 12812 10949 12880 11005
rect 12936 10949 13004 11005
rect 13060 10949 13070 11005
rect 12622 10939 13070 10949
rect 13758 12245 14206 12255
rect 13758 12189 13768 12245
rect 13824 12189 13892 12245
rect 13948 12189 14016 12245
rect 14072 12189 14140 12245
rect 14196 12189 14206 12245
rect 13758 12121 14206 12189
rect 13758 12065 13768 12121
rect 13824 12065 13892 12121
rect 13948 12065 14016 12121
rect 14072 12065 14140 12121
rect 14196 12065 14206 12121
rect 13758 11997 14206 12065
rect 13758 11941 13768 11997
rect 13824 11941 13892 11997
rect 13948 11941 14016 11997
rect 14072 11941 14140 11997
rect 14196 11941 14206 11997
rect 13758 11873 14206 11941
rect 13758 11817 13768 11873
rect 13824 11817 13892 11873
rect 13948 11817 14016 11873
rect 14072 11817 14140 11873
rect 14196 11817 14206 11873
rect 13758 11749 14206 11817
rect 13758 11693 13768 11749
rect 13824 11693 13892 11749
rect 13948 11693 14016 11749
rect 14072 11693 14140 11749
rect 14196 11693 14206 11749
rect 13758 11625 14206 11693
rect 13758 11569 13768 11625
rect 13824 11569 13892 11625
rect 13948 11569 14016 11625
rect 14072 11569 14140 11625
rect 14196 11569 14206 11625
rect 13758 11501 14206 11569
rect 13758 11445 13768 11501
rect 13824 11445 13892 11501
rect 13948 11445 14016 11501
rect 14072 11445 14140 11501
rect 14196 11445 14206 11501
rect 13758 11377 14206 11445
rect 13758 11321 13768 11377
rect 13824 11321 13892 11377
rect 13948 11321 14016 11377
rect 14072 11321 14140 11377
rect 14196 11321 14206 11377
rect 13758 11253 14206 11321
rect 13758 11197 13768 11253
rect 13824 11197 13892 11253
rect 13948 11197 14016 11253
rect 14072 11197 14140 11253
rect 14196 11197 14206 11253
rect 13758 11129 14206 11197
rect 13758 11073 13768 11129
rect 13824 11073 13892 11129
rect 13948 11073 14016 11129
rect 14072 11073 14140 11129
rect 14196 11073 14206 11129
rect 13758 11005 14206 11073
rect 13758 10949 13768 11005
rect 13824 10949 13892 11005
rect 13948 10949 14016 11005
rect 14072 10949 14140 11005
rect 14196 10949 14206 11005
rect 13758 10939 14206 10949
rect 290 10651 738 10661
rect 290 10595 300 10651
rect 356 10595 424 10651
rect 480 10595 548 10651
rect 604 10595 672 10651
rect 728 10595 738 10651
rect 290 10527 738 10595
rect 290 10471 300 10527
rect 356 10471 424 10527
rect 480 10471 548 10527
rect 604 10471 672 10527
rect 728 10471 738 10527
rect 290 10403 738 10471
rect 290 10347 300 10403
rect 356 10347 424 10403
rect 480 10347 548 10403
rect 604 10347 672 10403
rect 728 10347 738 10403
rect 290 10279 738 10347
rect 290 10223 300 10279
rect 356 10223 424 10279
rect 480 10223 548 10279
rect 604 10223 672 10279
rect 728 10223 738 10279
rect 290 10155 738 10223
rect 290 10099 300 10155
rect 356 10099 424 10155
rect 480 10099 548 10155
rect 604 10099 672 10155
rect 728 10099 738 10155
rect 290 10031 738 10099
rect 290 9975 300 10031
rect 356 9975 424 10031
rect 480 9975 548 10031
rect 604 9975 672 10031
rect 728 9975 738 10031
rect 290 9907 738 9975
rect 290 9851 300 9907
rect 356 9851 424 9907
rect 480 9851 548 9907
rect 604 9851 672 9907
rect 728 9851 738 9907
rect 290 9783 738 9851
rect 290 9727 300 9783
rect 356 9727 424 9783
rect 480 9727 548 9783
rect 604 9727 672 9783
rect 728 9727 738 9783
rect 290 9659 738 9727
rect 290 9603 300 9659
rect 356 9603 424 9659
rect 480 9603 548 9659
rect 604 9603 672 9659
rect 728 9603 738 9659
rect 290 9535 738 9603
rect 290 9479 300 9535
rect 356 9479 424 9535
rect 480 9479 548 9535
rect 604 9479 672 9535
rect 728 9479 738 9535
rect 290 9411 738 9479
rect 290 9355 300 9411
rect 356 9355 424 9411
rect 480 9355 548 9411
rect 604 9355 672 9411
rect 728 9355 738 9411
rect 290 9287 738 9355
rect 290 9231 300 9287
rect 356 9231 424 9287
rect 480 9231 548 9287
rect 604 9231 672 9287
rect 728 9231 738 9287
rect 290 9163 738 9231
rect 290 9107 300 9163
rect 356 9107 424 9163
rect 480 9107 548 9163
rect 604 9107 672 9163
rect 728 9107 738 9163
rect 290 9039 738 9107
rect 290 8983 300 9039
rect 356 8983 424 9039
rect 480 8983 548 9039
rect 604 8983 672 9039
rect 728 8983 738 9039
rect 290 8915 738 8983
rect 290 8859 300 8915
rect 356 8859 424 8915
rect 480 8859 548 8915
rect 604 8859 672 8915
rect 728 8859 738 8915
rect 290 8791 738 8859
rect 290 8735 300 8791
rect 356 8735 424 8791
rect 480 8735 548 8791
rect 604 8735 672 8791
rect 728 8735 738 8791
rect 290 8667 738 8735
rect 290 8611 300 8667
rect 356 8611 424 8667
rect 480 8611 548 8667
rect 604 8611 672 8667
rect 728 8611 738 8667
rect 290 8543 738 8611
rect 290 8487 300 8543
rect 356 8487 424 8543
rect 480 8487 548 8543
rect 604 8487 672 8543
rect 728 8487 738 8543
rect 290 8419 738 8487
rect 290 8363 300 8419
rect 356 8363 424 8419
rect 480 8363 548 8419
rect 604 8363 672 8419
rect 728 8363 738 8419
rect 290 8295 738 8363
rect 290 8239 300 8295
rect 356 8239 424 8295
rect 480 8239 548 8295
rect 604 8239 672 8295
rect 728 8239 738 8295
rect 290 8171 738 8239
rect 290 8115 300 8171
rect 356 8115 424 8171
rect 480 8115 548 8171
rect 604 8115 672 8171
rect 728 8115 738 8171
rect 290 8047 738 8115
rect 290 7991 300 8047
rect 356 7991 424 8047
rect 480 7991 548 8047
rect 604 7991 672 8047
rect 728 7991 738 8047
rect 290 7923 738 7991
rect 290 7867 300 7923
rect 356 7867 424 7923
rect 480 7867 548 7923
rect 604 7867 672 7923
rect 728 7867 738 7923
rect 290 7799 738 7867
rect 290 7743 300 7799
rect 356 7743 424 7799
rect 480 7743 548 7799
rect 604 7743 672 7799
rect 728 7743 738 7799
rect 290 7733 738 7743
rect 1426 10651 1874 10661
rect 1426 10595 1436 10651
rect 1492 10595 1560 10651
rect 1616 10595 1684 10651
rect 1740 10595 1808 10651
rect 1864 10595 1874 10651
rect 1426 10527 1874 10595
rect 1426 10471 1436 10527
rect 1492 10471 1560 10527
rect 1616 10471 1684 10527
rect 1740 10471 1808 10527
rect 1864 10471 1874 10527
rect 1426 10403 1874 10471
rect 1426 10347 1436 10403
rect 1492 10347 1560 10403
rect 1616 10347 1684 10403
rect 1740 10347 1808 10403
rect 1864 10347 1874 10403
rect 1426 10279 1874 10347
rect 1426 10223 1436 10279
rect 1492 10223 1560 10279
rect 1616 10223 1684 10279
rect 1740 10223 1808 10279
rect 1864 10223 1874 10279
rect 1426 10155 1874 10223
rect 1426 10099 1436 10155
rect 1492 10099 1560 10155
rect 1616 10099 1684 10155
rect 1740 10099 1808 10155
rect 1864 10099 1874 10155
rect 1426 10031 1874 10099
rect 1426 9975 1436 10031
rect 1492 9975 1560 10031
rect 1616 9975 1684 10031
rect 1740 9975 1808 10031
rect 1864 9975 1874 10031
rect 1426 9907 1874 9975
rect 1426 9851 1436 9907
rect 1492 9851 1560 9907
rect 1616 9851 1684 9907
rect 1740 9851 1808 9907
rect 1864 9851 1874 9907
rect 1426 9783 1874 9851
rect 1426 9727 1436 9783
rect 1492 9727 1560 9783
rect 1616 9727 1684 9783
rect 1740 9727 1808 9783
rect 1864 9727 1874 9783
rect 1426 9659 1874 9727
rect 1426 9603 1436 9659
rect 1492 9603 1560 9659
rect 1616 9603 1684 9659
rect 1740 9603 1808 9659
rect 1864 9603 1874 9659
rect 1426 9535 1874 9603
rect 1426 9479 1436 9535
rect 1492 9479 1560 9535
rect 1616 9479 1684 9535
rect 1740 9479 1808 9535
rect 1864 9479 1874 9535
rect 1426 9411 1874 9479
rect 1426 9355 1436 9411
rect 1492 9355 1560 9411
rect 1616 9355 1684 9411
rect 1740 9355 1808 9411
rect 1864 9355 1874 9411
rect 1426 9287 1874 9355
rect 1426 9231 1436 9287
rect 1492 9231 1560 9287
rect 1616 9231 1684 9287
rect 1740 9231 1808 9287
rect 1864 9231 1874 9287
rect 1426 9163 1874 9231
rect 1426 9107 1436 9163
rect 1492 9107 1560 9163
rect 1616 9107 1684 9163
rect 1740 9107 1808 9163
rect 1864 9107 1874 9163
rect 1426 9039 1874 9107
rect 1426 8983 1436 9039
rect 1492 8983 1560 9039
rect 1616 8983 1684 9039
rect 1740 8983 1808 9039
rect 1864 8983 1874 9039
rect 1426 8915 1874 8983
rect 1426 8859 1436 8915
rect 1492 8859 1560 8915
rect 1616 8859 1684 8915
rect 1740 8859 1808 8915
rect 1864 8859 1874 8915
rect 1426 8791 1874 8859
rect 1426 8735 1436 8791
rect 1492 8735 1560 8791
rect 1616 8735 1684 8791
rect 1740 8735 1808 8791
rect 1864 8735 1874 8791
rect 1426 8667 1874 8735
rect 1426 8611 1436 8667
rect 1492 8611 1560 8667
rect 1616 8611 1684 8667
rect 1740 8611 1808 8667
rect 1864 8611 1874 8667
rect 1426 8543 1874 8611
rect 1426 8487 1436 8543
rect 1492 8487 1560 8543
rect 1616 8487 1684 8543
rect 1740 8487 1808 8543
rect 1864 8487 1874 8543
rect 1426 8419 1874 8487
rect 1426 8363 1436 8419
rect 1492 8363 1560 8419
rect 1616 8363 1684 8419
rect 1740 8363 1808 8419
rect 1864 8363 1874 8419
rect 1426 8295 1874 8363
rect 1426 8239 1436 8295
rect 1492 8239 1560 8295
rect 1616 8239 1684 8295
rect 1740 8239 1808 8295
rect 1864 8239 1874 8295
rect 1426 8171 1874 8239
rect 1426 8115 1436 8171
rect 1492 8115 1560 8171
rect 1616 8115 1684 8171
rect 1740 8115 1808 8171
rect 1864 8115 1874 8171
rect 1426 8047 1874 8115
rect 1426 7991 1436 8047
rect 1492 7991 1560 8047
rect 1616 7991 1684 8047
rect 1740 7991 1808 8047
rect 1864 7991 1874 8047
rect 1426 7923 1874 7991
rect 1426 7867 1436 7923
rect 1492 7867 1560 7923
rect 1616 7867 1684 7923
rect 1740 7867 1808 7923
rect 1864 7867 1874 7923
rect 1426 7799 1874 7867
rect 1426 7743 1436 7799
rect 1492 7743 1560 7799
rect 1616 7743 1684 7799
rect 1740 7743 1808 7799
rect 1864 7743 1874 7799
rect 1426 7733 1874 7743
rect 2562 10651 3010 10661
rect 2562 10595 2572 10651
rect 2628 10595 2696 10651
rect 2752 10595 2820 10651
rect 2876 10595 2944 10651
rect 3000 10595 3010 10651
rect 2562 10527 3010 10595
rect 2562 10471 2572 10527
rect 2628 10471 2696 10527
rect 2752 10471 2820 10527
rect 2876 10471 2944 10527
rect 3000 10471 3010 10527
rect 2562 10403 3010 10471
rect 2562 10347 2572 10403
rect 2628 10347 2696 10403
rect 2752 10347 2820 10403
rect 2876 10347 2944 10403
rect 3000 10347 3010 10403
rect 2562 10279 3010 10347
rect 2562 10223 2572 10279
rect 2628 10223 2696 10279
rect 2752 10223 2820 10279
rect 2876 10223 2944 10279
rect 3000 10223 3010 10279
rect 2562 10155 3010 10223
rect 2562 10099 2572 10155
rect 2628 10099 2696 10155
rect 2752 10099 2820 10155
rect 2876 10099 2944 10155
rect 3000 10099 3010 10155
rect 2562 10031 3010 10099
rect 2562 9975 2572 10031
rect 2628 9975 2696 10031
rect 2752 9975 2820 10031
rect 2876 9975 2944 10031
rect 3000 9975 3010 10031
rect 2562 9907 3010 9975
rect 2562 9851 2572 9907
rect 2628 9851 2696 9907
rect 2752 9851 2820 9907
rect 2876 9851 2944 9907
rect 3000 9851 3010 9907
rect 2562 9783 3010 9851
rect 2562 9727 2572 9783
rect 2628 9727 2696 9783
rect 2752 9727 2820 9783
rect 2876 9727 2944 9783
rect 3000 9727 3010 9783
rect 2562 9659 3010 9727
rect 2562 9603 2572 9659
rect 2628 9603 2696 9659
rect 2752 9603 2820 9659
rect 2876 9603 2944 9659
rect 3000 9603 3010 9659
rect 2562 9535 3010 9603
rect 2562 9479 2572 9535
rect 2628 9479 2696 9535
rect 2752 9479 2820 9535
rect 2876 9479 2944 9535
rect 3000 9479 3010 9535
rect 2562 9411 3010 9479
rect 2562 9355 2572 9411
rect 2628 9355 2696 9411
rect 2752 9355 2820 9411
rect 2876 9355 2944 9411
rect 3000 9355 3010 9411
rect 2562 9287 3010 9355
rect 2562 9231 2572 9287
rect 2628 9231 2696 9287
rect 2752 9231 2820 9287
rect 2876 9231 2944 9287
rect 3000 9231 3010 9287
rect 2562 9163 3010 9231
rect 2562 9107 2572 9163
rect 2628 9107 2696 9163
rect 2752 9107 2820 9163
rect 2876 9107 2944 9163
rect 3000 9107 3010 9163
rect 2562 9039 3010 9107
rect 2562 8983 2572 9039
rect 2628 8983 2696 9039
rect 2752 8983 2820 9039
rect 2876 8983 2944 9039
rect 3000 8983 3010 9039
rect 2562 8915 3010 8983
rect 2562 8859 2572 8915
rect 2628 8859 2696 8915
rect 2752 8859 2820 8915
rect 2876 8859 2944 8915
rect 3000 8859 3010 8915
rect 2562 8791 3010 8859
rect 2562 8735 2572 8791
rect 2628 8735 2696 8791
rect 2752 8735 2820 8791
rect 2876 8735 2944 8791
rect 3000 8735 3010 8791
rect 2562 8667 3010 8735
rect 2562 8611 2572 8667
rect 2628 8611 2696 8667
rect 2752 8611 2820 8667
rect 2876 8611 2944 8667
rect 3000 8611 3010 8667
rect 2562 8543 3010 8611
rect 2562 8487 2572 8543
rect 2628 8487 2696 8543
rect 2752 8487 2820 8543
rect 2876 8487 2944 8543
rect 3000 8487 3010 8543
rect 2562 8419 3010 8487
rect 2562 8363 2572 8419
rect 2628 8363 2696 8419
rect 2752 8363 2820 8419
rect 2876 8363 2944 8419
rect 3000 8363 3010 8419
rect 2562 8295 3010 8363
rect 2562 8239 2572 8295
rect 2628 8239 2696 8295
rect 2752 8239 2820 8295
rect 2876 8239 2944 8295
rect 3000 8239 3010 8295
rect 2562 8171 3010 8239
rect 2562 8115 2572 8171
rect 2628 8115 2696 8171
rect 2752 8115 2820 8171
rect 2876 8115 2944 8171
rect 3000 8115 3010 8171
rect 2562 8047 3010 8115
rect 2562 7991 2572 8047
rect 2628 7991 2696 8047
rect 2752 7991 2820 8047
rect 2876 7991 2944 8047
rect 3000 7991 3010 8047
rect 2562 7923 3010 7991
rect 2562 7867 2572 7923
rect 2628 7867 2696 7923
rect 2752 7867 2820 7923
rect 2876 7867 2944 7923
rect 3000 7867 3010 7923
rect 2562 7799 3010 7867
rect 2562 7743 2572 7799
rect 2628 7743 2696 7799
rect 2752 7743 2820 7799
rect 2876 7743 2944 7799
rect 3000 7743 3010 7799
rect 2562 7733 3010 7743
rect 4834 10651 5282 10661
rect 4834 10595 4844 10651
rect 4900 10595 4968 10651
rect 5024 10595 5092 10651
rect 5148 10595 5216 10651
rect 5272 10595 5282 10651
rect 4834 10527 5282 10595
rect 4834 10471 4844 10527
rect 4900 10471 4968 10527
rect 5024 10471 5092 10527
rect 5148 10471 5216 10527
rect 5272 10471 5282 10527
rect 4834 10403 5282 10471
rect 4834 10347 4844 10403
rect 4900 10347 4968 10403
rect 5024 10347 5092 10403
rect 5148 10347 5216 10403
rect 5272 10347 5282 10403
rect 4834 10279 5282 10347
rect 4834 10223 4844 10279
rect 4900 10223 4968 10279
rect 5024 10223 5092 10279
rect 5148 10223 5216 10279
rect 5272 10223 5282 10279
rect 4834 10155 5282 10223
rect 4834 10099 4844 10155
rect 4900 10099 4968 10155
rect 5024 10099 5092 10155
rect 5148 10099 5216 10155
rect 5272 10099 5282 10155
rect 4834 10031 5282 10099
rect 4834 9975 4844 10031
rect 4900 9975 4968 10031
rect 5024 9975 5092 10031
rect 5148 9975 5216 10031
rect 5272 9975 5282 10031
rect 4834 9907 5282 9975
rect 4834 9851 4844 9907
rect 4900 9851 4968 9907
rect 5024 9851 5092 9907
rect 5148 9851 5216 9907
rect 5272 9851 5282 9907
rect 4834 9783 5282 9851
rect 4834 9727 4844 9783
rect 4900 9727 4968 9783
rect 5024 9727 5092 9783
rect 5148 9727 5216 9783
rect 5272 9727 5282 9783
rect 4834 9659 5282 9727
rect 4834 9603 4844 9659
rect 4900 9603 4968 9659
rect 5024 9603 5092 9659
rect 5148 9603 5216 9659
rect 5272 9603 5282 9659
rect 4834 9535 5282 9603
rect 4834 9479 4844 9535
rect 4900 9479 4968 9535
rect 5024 9479 5092 9535
rect 5148 9479 5216 9535
rect 5272 9479 5282 9535
rect 4834 9411 5282 9479
rect 4834 9355 4844 9411
rect 4900 9355 4968 9411
rect 5024 9355 5092 9411
rect 5148 9355 5216 9411
rect 5272 9355 5282 9411
rect 4834 9287 5282 9355
rect 4834 9231 4844 9287
rect 4900 9231 4968 9287
rect 5024 9231 5092 9287
rect 5148 9231 5216 9287
rect 5272 9231 5282 9287
rect 4834 9163 5282 9231
rect 4834 9107 4844 9163
rect 4900 9107 4968 9163
rect 5024 9107 5092 9163
rect 5148 9107 5216 9163
rect 5272 9107 5282 9163
rect 4834 9039 5282 9107
rect 4834 8983 4844 9039
rect 4900 8983 4968 9039
rect 5024 8983 5092 9039
rect 5148 8983 5216 9039
rect 5272 8983 5282 9039
rect 4834 8915 5282 8983
rect 4834 8859 4844 8915
rect 4900 8859 4968 8915
rect 5024 8859 5092 8915
rect 5148 8859 5216 8915
rect 5272 8859 5282 8915
rect 4834 8791 5282 8859
rect 4834 8735 4844 8791
rect 4900 8735 4968 8791
rect 5024 8735 5092 8791
rect 5148 8735 5216 8791
rect 5272 8735 5282 8791
rect 4834 8667 5282 8735
rect 4834 8611 4844 8667
rect 4900 8611 4968 8667
rect 5024 8611 5092 8667
rect 5148 8611 5216 8667
rect 5272 8611 5282 8667
rect 4834 8543 5282 8611
rect 4834 8487 4844 8543
rect 4900 8487 4968 8543
rect 5024 8487 5092 8543
rect 5148 8487 5216 8543
rect 5272 8487 5282 8543
rect 4834 8419 5282 8487
rect 4834 8363 4844 8419
rect 4900 8363 4968 8419
rect 5024 8363 5092 8419
rect 5148 8363 5216 8419
rect 5272 8363 5282 8419
rect 4834 8295 5282 8363
rect 4834 8239 4844 8295
rect 4900 8239 4968 8295
rect 5024 8239 5092 8295
rect 5148 8239 5216 8295
rect 5272 8239 5282 8295
rect 4834 8171 5282 8239
rect 4834 8115 4844 8171
rect 4900 8115 4968 8171
rect 5024 8115 5092 8171
rect 5148 8115 5216 8171
rect 5272 8115 5282 8171
rect 4834 8047 5282 8115
rect 4834 7991 4844 8047
rect 4900 7991 4968 8047
rect 5024 7991 5092 8047
rect 5148 7991 5216 8047
rect 5272 7991 5282 8047
rect 4834 7923 5282 7991
rect 4834 7867 4844 7923
rect 4900 7867 4968 7923
rect 5024 7867 5092 7923
rect 5148 7867 5216 7923
rect 5272 7867 5282 7923
rect 4834 7799 5282 7867
rect 4834 7743 4844 7799
rect 4900 7743 4968 7799
rect 5024 7743 5092 7799
rect 5148 7743 5216 7799
rect 5272 7743 5282 7799
rect 4834 7733 5282 7743
rect 7127 10651 7451 10661
rect 7127 10595 7137 10651
rect 7193 10595 7261 10651
rect 7317 10595 7385 10651
rect 7441 10595 7451 10651
rect 7127 10527 7451 10595
rect 7127 10471 7137 10527
rect 7193 10471 7261 10527
rect 7317 10471 7385 10527
rect 7441 10471 7451 10527
rect 7127 10403 7451 10471
rect 7127 10347 7137 10403
rect 7193 10347 7261 10403
rect 7317 10347 7385 10403
rect 7441 10347 7451 10403
rect 7127 10279 7451 10347
rect 7127 10223 7137 10279
rect 7193 10223 7261 10279
rect 7317 10223 7385 10279
rect 7441 10223 7451 10279
rect 7127 10155 7451 10223
rect 7127 10099 7137 10155
rect 7193 10099 7261 10155
rect 7317 10099 7385 10155
rect 7441 10099 7451 10155
rect 7127 10031 7451 10099
rect 7127 9975 7137 10031
rect 7193 9975 7261 10031
rect 7317 9975 7385 10031
rect 7441 9975 7451 10031
rect 7127 9907 7451 9975
rect 7127 9851 7137 9907
rect 7193 9851 7261 9907
rect 7317 9851 7385 9907
rect 7441 9851 7451 9907
rect 7127 9783 7451 9851
rect 7127 9727 7137 9783
rect 7193 9727 7261 9783
rect 7317 9727 7385 9783
rect 7441 9727 7451 9783
rect 7127 9659 7451 9727
rect 7127 9603 7137 9659
rect 7193 9603 7261 9659
rect 7317 9603 7385 9659
rect 7441 9603 7451 9659
rect 7127 9535 7451 9603
rect 7127 9479 7137 9535
rect 7193 9479 7261 9535
rect 7317 9479 7385 9535
rect 7441 9479 7451 9535
rect 7127 9411 7451 9479
rect 7127 9355 7137 9411
rect 7193 9355 7261 9411
rect 7317 9355 7385 9411
rect 7441 9355 7451 9411
rect 7127 9287 7451 9355
rect 7127 9231 7137 9287
rect 7193 9231 7261 9287
rect 7317 9231 7385 9287
rect 7441 9231 7451 9287
rect 7127 9163 7451 9231
rect 7127 9107 7137 9163
rect 7193 9107 7261 9163
rect 7317 9107 7385 9163
rect 7441 9107 7451 9163
rect 7127 9039 7451 9107
rect 7127 8983 7137 9039
rect 7193 8983 7261 9039
rect 7317 8983 7385 9039
rect 7441 8983 7451 9039
rect 7127 8915 7451 8983
rect 7127 8859 7137 8915
rect 7193 8859 7261 8915
rect 7317 8859 7385 8915
rect 7441 8859 7451 8915
rect 7127 8791 7451 8859
rect 7127 8735 7137 8791
rect 7193 8735 7261 8791
rect 7317 8735 7385 8791
rect 7441 8735 7451 8791
rect 7127 8667 7451 8735
rect 7127 8611 7137 8667
rect 7193 8611 7261 8667
rect 7317 8611 7385 8667
rect 7441 8611 7451 8667
rect 7127 8543 7451 8611
rect 7127 8487 7137 8543
rect 7193 8487 7261 8543
rect 7317 8487 7385 8543
rect 7441 8487 7451 8543
rect 7127 8419 7451 8487
rect 7127 8363 7137 8419
rect 7193 8363 7261 8419
rect 7317 8363 7385 8419
rect 7441 8363 7451 8419
rect 7127 8295 7451 8363
rect 7127 8239 7137 8295
rect 7193 8239 7261 8295
rect 7317 8239 7385 8295
rect 7441 8239 7451 8295
rect 7127 8171 7451 8239
rect 7127 8115 7137 8171
rect 7193 8115 7261 8171
rect 7317 8115 7385 8171
rect 7441 8115 7451 8171
rect 7127 8047 7451 8115
rect 7127 7991 7137 8047
rect 7193 7991 7261 8047
rect 7317 7991 7385 8047
rect 7441 7991 7451 8047
rect 7127 7923 7451 7991
rect 7127 7867 7137 7923
rect 7193 7867 7261 7923
rect 7317 7867 7385 7923
rect 7441 7867 7451 7923
rect 7127 7799 7451 7867
rect 7127 7743 7137 7799
rect 7193 7743 7261 7799
rect 7317 7743 7385 7799
rect 7441 7743 7451 7799
rect 7127 7733 7451 7743
rect 7613 10651 7937 10661
rect 7613 10595 7623 10651
rect 7679 10595 7747 10651
rect 7803 10595 7871 10651
rect 7927 10595 7937 10651
rect 7613 10527 7937 10595
rect 7613 10471 7623 10527
rect 7679 10471 7747 10527
rect 7803 10471 7871 10527
rect 7927 10471 7937 10527
rect 7613 10403 7937 10471
rect 7613 10347 7623 10403
rect 7679 10347 7747 10403
rect 7803 10347 7871 10403
rect 7927 10347 7937 10403
rect 7613 10279 7937 10347
rect 7613 10223 7623 10279
rect 7679 10223 7747 10279
rect 7803 10223 7871 10279
rect 7927 10223 7937 10279
rect 7613 10155 7937 10223
rect 7613 10099 7623 10155
rect 7679 10099 7747 10155
rect 7803 10099 7871 10155
rect 7927 10099 7937 10155
rect 7613 10031 7937 10099
rect 7613 9975 7623 10031
rect 7679 9975 7747 10031
rect 7803 9975 7871 10031
rect 7927 9975 7937 10031
rect 7613 9907 7937 9975
rect 7613 9851 7623 9907
rect 7679 9851 7747 9907
rect 7803 9851 7871 9907
rect 7927 9851 7937 9907
rect 7613 9783 7937 9851
rect 7613 9727 7623 9783
rect 7679 9727 7747 9783
rect 7803 9727 7871 9783
rect 7927 9727 7937 9783
rect 7613 9659 7937 9727
rect 7613 9603 7623 9659
rect 7679 9603 7747 9659
rect 7803 9603 7871 9659
rect 7927 9603 7937 9659
rect 7613 9535 7937 9603
rect 7613 9479 7623 9535
rect 7679 9479 7747 9535
rect 7803 9479 7871 9535
rect 7927 9479 7937 9535
rect 7613 9411 7937 9479
rect 7613 9355 7623 9411
rect 7679 9355 7747 9411
rect 7803 9355 7871 9411
rect 7927 9355 7937 9411
rect 7613 9287 7937 9355
rect 7613 9231 7623 9287
rect 7679 9231 7747 9287
rect 7803 9231 7871 9287
rect 7927 9231 7937 9287
rect 7613 9163 7937 9231
rect 7613 9107 7623 9163
rect 7679 9107 7747 9163
rect 7803 9107 7871 9163
rect 7927 9107 7937 9163
rect 7613 9039 7937 9107
rect 7613 8983 7623 9039
rect 7679 8983 7747 9039
rect 7803 8983 7871 9039
rect 7927 8983 7937 9039
rect 7613 8915 7937 8983
rect 7613 8859 7623 8915
rect 7679 8859 7747 8915
rect 7803 8859 7871 8915
rect 7927 8859 7937 8915
rect 7613 8791 7937 8859
rect 7613 8735 7623 8791
rect 7679 8735 7747 8791
rect 7803 8735 7871 8791
rect 7927 8735 7937 8791
rect 7613 8667 7937 8735
rect 7613 8611 7623 8667
rect 7679 8611 7747 8667
rect 7803 8611 7871 8667
rect 7927 8611 7937 8667
rect 7613 8543 7937 8611
rect 7613 8487 7623 8543
rect 7679 8487 7747 8543
rect 7803 8487 7871 8543
rect 7927 8487 7937 8543
rect 7613 8419 7937 8487
rect 7613 8363 7623 8419
rect 7679 8363 7747 8419
rect 7803 8363 7871 8419
rect 7927 8363 7937 8419
rect 7613 8295 7937 8363
rect 7613 8239 7623 8295
rect 7679 8239 7747 8295
rect 7803 8239 7871 8295
rect 7927 8239 7937 8295
rect 7613 8171 7937 8239
rect 7613 8115 7623 8171
rect 7679 8115 7747 8171
rect 7803 8115 7871 8171
rect 7927 8115 7937 8171
rect 7613 8047 7937 8115
rect 7613 7991 7623 8047
rect 7679 7991 7747 8047
rect 7803 7991 7871 8047
rect 7927 7991 7937 8047
rect 7613 7923 7937 7991
rect 7613 7867 7623 7923
rect 7679 7867 7747 7923
rect 7803 7867 7871 7923
rect 7927 7867 7937 7923
rect 7613 7799 7937 7867
rect 7613 7743 7623 7799
rect 7679 7743 7747 7799
rect 7803 7743 7871 7799
rect 7927 7743 7937 7799
rect 7613 7733 7937 7743
rect 9782 10651 10230 10661
rect 9782 10595 9792 10651
rect 9848 10595 9916 10651
rect 9972 10595 10040 10651
rect 10096 10595 10164 10651
rect 10220 10595 10230 10651
rect 9782 10527 10230 10595
rect 9782 10471 9792 10527
rect 9848 10471 9916 10527
rect 9972 10471 10040 10527
rect 10096 10471 10164 10527
rect 10220 10471 10230 10527
rect 9782 10403 10230 10471
rect 9782 10347 9792 10403
rect 9848 10347 9916 10403
rect 9972 10347 10040 10403
rect 10096 10347 10164 10403
rect 10220 10347 10230 10403
rect 9782 10279 10230 10347
rect 9782 10223 9792 10279
rect 9848 10223 9916 10279
rect 9972 10223 10040 10279
rect 10096 10223 10164 10279
rect 10220 10223 10230 10279
rect 9782 10155 10230 10223
rect 9782 10099 9792 10155
rect 9848 10099 9916 10155
rect 9972 10099 10040 10155
rect 10096 10099 10164 10155
rect 10220 10099 10230 10155
rect 9782 10031 10230 10099
rect 9782 9975 9792 10031
rect 9848 9975 9916 10031
rect 9972 9975 10040 10031
rect 10096 9975 10164 10031
rect 10220 9975 10230 10031
rect 9782 9907 10230 9975
rect 9782 9851 9792 9907
rect 9848 9851 9916 9907
rect 9972 9851 10040 9907
rect 10096 9851 10164 9907
rect 10220 9851 10230 9907
rect 9782 9783 10230 9851
rect 9782 9727 9792 9783
rect 9848 9727 9916 9783
rect 9972 9727 10040 9783
rect 10096 9727 10164 9783
rect 10220 9727 10230 9783
rect 9782 9659 10230 9727
rect 9782 9603 9792 9659
rect 9848 9603 9916 9659
rect 9972 9603 10040 9659
rect 10096 9603 10164 9659
rect 10220 9603 10230 9659
rect 9782 9535 10230 9603
rect 9782 9479 9792 9535
rect 9848 9479 9916 9535
rect 9972 9479 10040 9535
rect 10096 9479 10164 9535
rect 10220 9479 10230 9535
rect 9782 9411 10230 9479
rect 9782 9355 9792 9411
rect 9848 9355 9916 9411
rect 9972 9355 10040 9411
rect 10096 9355 10164 9411
rect 10220 9355 10230 9411
rect 9782 9287 10230 9355
rect 9782 9231 9792 9287
rect 9848 9231 9916 9287
rect 9972 9231 10040 9287
rect 10096 9231 10164 9287
rect 10220 9231 10230 9287
rect 9782 9163 10230 9231
rect 9782 9107 9792 9163
rect 9848 9107 9916 9163
rect 9972 9107 10040 9163
rect 10096 9107 10164 9163
rect 10220 9107 10230 9163
rect 9782 9039 10230 9107
rect 9782 8983 9792 9039
rect 9848 8983 9916 9039
rect 9972 8983 10040 9039
rect 10096 8983 10164 9039
rect 10220 8983 10230 9039
rect 9782 8915 10230 8983
rect 9782 8859 9792 8915
rect 9848 8859 9916 8915
rect 9972 8859 10040 8915
rect 10096 8859 10164 8915
rect 10220 8859 10230 8915
rect 9782 8791 10230 8859
rect 9782 8735 9792 8791
rect 9848 8735 9916 8791
rect 9972 8735 10040 8791
rect 10096 8735 10164 8791
rect 10220 8735 10230 8791
rect 9782 8667 10230 8735
rect 9782 8611 9792 8667
rect 9848 8611 9916 8667
rect 9972 8611 10040 8667
rect 10096 8611 10164 8667
rect 10220 8611 10230 8667
rect 9782 8543 10230 8611
rect 9782 8487 9792 8543
rect 9848 8487 9916 8543
rect 9972 8487 10040 8543
rect 10096 8487 10164 8543
rect 10220 8487 10230 8543
rect 9782 8419 10230 8487
rect 9782 8363 9792 8419
rect 9848 8363 9916 8419
rect 9972 8363 10040 8419
rect 10096 8363 10164 8419
rect 10220 8363 10230 8419
rect 9782 8295 10230 8363
rect 9782 8239 9792 8295
rect 9848 8239 9916 8295
rect 9972 8239 10040 8295
rect 10096 8239 10164 8295
rect 10220 8239 10230 8295
rect 9782 8171 10230 8239
rect 9782 8115 9792 8171
rect 9848 8115 9916 8171
rect 9972 8115 10040 8171
rect 10096 8115 10164 8171
rect 10220 8115 10230 8171
rect 9782 8047 10230 8115
rect 9782 7991 9792 8047
rect 9848 7991 9916 8047
rect 9972 7991 10040 8047
rect 10096 7991 10164 8047
rect 10220 7991 10230 8047
rect 9782 7923 10230 7991
rect 9782 7867 9792 7923
rect 9848 7867 9916 7923
rect 9972 7867 10040 7923
rect 10096 7867 10164 7923
rect 10220 7867 10230 7923
rect 9782 7799 10230 7867
rect 9782 7743 9792 7799
rect 9848 7743 9916 7799
rect 9972 7743 10040 7799
rect 10096 7743 10164 7799
rect 10220 7743 10230 7799
rect 9782 7733 10230 7743
rect 12054 10651 12502 10661
rect 12054 10595 12064 10651
rect 12120 10595 12188 10651
rect 12244 10595 12312 10651
rect 12368 10595 12436 10651
rect 12492 10595 12502 10651
rect 12054 10527 12502 10595
rect 12054 10471 12064 10527
rect 12120 10471 12188 10527
rect 12244 10471 12312 10527
rect 12368 10471 12436 10527
rect 12492 10471 12502 10527
rect 12054 10403 12502 10471
rect 12054 10347 12064 10403
rect 12120 10347 12188 10403
rect 12244 10347 12312 10403
rect 12368 10347 12436 10403
rect 12492 10347 12502 10403
rect 12054 10279 12502 10347
rect 12054 10223 12064 10279
rect 12120 10223 12188 10279
rect 12244 10223 12312 10279
rect 12368 10223 12436 10279
rect 12492 10223 12502 10279
rect 12054 10155 12502 10223
rect 12054 10099 12064 10155
rect 12120 10099 12188 10155
rect 12244 10099 12312 10155
rect 12368 10099 12436 10155
rect 12492 10099 12502 10155
rect 12054 10031 12502 10099
rect 12054 9975 12064 10031
rect 12120 9975 12188 10031
rect 12244 9975 12312 10031
rect 12368 9975 12436 10031
rect 12492 9975 12502 10031
rect 12054 9907 12502 9975
rect 12054 9851 12064 9907
rect 12120 9851 12188 9907
rect 12244 9851 12312 9907
rect 12368 9851 12436 9907
rect 12492 9851 12502 9907
rect 12054 9783 12502 9851
rect 12054 9727 12064 9783
rect 12120 9727 12188 9783
rect 12244 9727 12312 9783
rect 12368 9727 12436 9783
rect 12492 9727 12502 9783
rect 12054 9659 12502 9727
rect 12054 9603 12064 9659
rect 12120 9603 12188 9659
rect 12244 9603 12312 9659
rect 12368 9603 12436 9659
rect 12492 9603 12502 9659
rect 12054 9535 12502 9603
rect 12054 9479 12064 9535
rect 12120 9479 12188 9535
rect 12244 9479 12312 9535
rect 12368 9479 12436 9535
rect 12492 9479 12502 9535
rect 12054 9411 12502 9479
rect 12054 9355 12064 9411
rect 12120 9355 12188 9411
rect 12244 9355 12312 9411
rect 12368 9355 12436 9411
rect 12492 9355 12502 9411
rect 12054 9287 12502 9355
rect 12054 9231 12064 9287
rect 12120 9231 12188 9287
rect 12244 9231 12312 9287
rect 12368 9231 12436 9287
rect 12492 9231 12502 9287
rect 12054 9163 12502 9231
rect 12054 9107 12064 9163
rect 12120 9107 12188 9163
rect 12244 9107 12312 9163
rect 12368 9107 12436 9163
rect 12492 9107 12502 9163
rect 12054 9039 12502 9107
rect 12054 8983 12064 9039
rect 12120 8983 12188 9039
rect 12244 8983 12312 9039
rect 12368 8983 12436 9039
rect 12492 8983 12502 9039
rect 12054 8915 12502 8983
rect 12054 8859 12064 8915
rect 12120 8859 12188 8915
rect 12244 8859 12312 8915
rect 12368 8859 12436 8915
rect 12492 8859 12502 8915
rect 12054 8791 12502 8859
rect 12054 8735 12064 8791
rect 12120 8735 12188 8791
rect 12244 8735 12312 8791
rect 12368 8735 12436 8791
rect 12492 8735 12502 8791
rect 12054 8667 12502 8735
rect 12054 8611 12064 8667
rect 12120 8611 12188 8667
rect 12244 8611 12312 8667
rect 12368 8611 12436 8667
rect 12492 8611 12502 8667
rect 12054 8543 12502 8611
rect 12054 8487 12064 8543
rect 12120 8487 12188 8543
rect 12244 8487 12312 8543
rect 12368 8487 12436 8543
rect 12492 8487 12502 8543
rect 12054 8419 12502 8487
rect 12054 8363 12064 8419
rect 12120 8363 12188 8419
rect 12244 8363 12312 8419
rect 12368 8363 12436 8419
rect 12492 8363 12502 8419
rect 12054 8295 12502 8363
rect 12054 8239 12064 8295
rect 12120 8239 12188 8295
rect 12244 8239 12312 8295
rect 12368 8239 12436 8295
rect 12492 8239 12502 8295
rect 12054 8171 12502 8239
rect 12054 8115 12064 8171
rect 12120 8115 12188 8171
rect 12244 8115 12312 8171
rect 12368 8115 12436 8171
rect 12492 8115 12502 8171
rect 12054 8047 12502 8115
rect 12054 7991 12064 8047
rect 12120 7991 12188 8047
rect 12244 7991 12312 8047
rect 12368 7991 12436 8047
rect 12492 7991 12502 8047
rect 12054 7923 12502 7991
rect 12054 7867 12064 7923
rect 12120 7867 12188 7923
rect 12244 7867 12312 7923
rect 12368 7867 12436 7923
rect 12492 7867 12502 7923
rect 12054 7799 12502 7867
rect 12054 7743 12064 7799
rect 12120 7743 12188 7799
rect 12244 7743 12312 7799
rect 12368 7743 12436 7799
rect 12492 7743 12502 7799
rect 12054 7733 12502 7743
rect 13190 10651 13638 10661
rect 13190 10595 13200 10651
rect 13256 10595 13324 10651
rect 13380 10595 13448 10651
rect 13504 10595 13572 10651
rect 13628 10595 13638 10651
rect 13190 10527 13638 10595
rect 13190 10471 13200 10527
rect 13256 10471 13324 10527
rect 13380 10471 13448 10527
rect 13504 10471 13572 10527
rect 13628 10471 13638 10527
rect 13190 10403 13638 10471
rect 13190 10347 13200 10403
rect 13256 10347 13324 10403
rect 13380 10347 13448 10403
rect 13504 10347 13572 10403
rect 13628 10347 13638 10403
rect 13190 10279 13638 10347
rect 13190 10223 13200 10279
rect 13256 10223 13324 10279
rect 13380 10223 13448 10279
rect 13504 10223 13572 10279
rect 13628 10223 13638 10279
rect 13190 10155 13638 10223
rect 13190 10099 13200 10155
rect 13256 10099 13324 10155
rect 13380 10099 13448 10155
rect 13504 10099 13572 10155
rect 13628 10099 13638 10155
rect 13190 10031 13638 10099
rect 13190 9975 13200 10031
rect 13256 9975 13324 10031
rect 13380 9975 13448 10031
rect 13504 9975 13572 10031
rect 13628 9975 13638 10031
rect 13190 9907 13638 9975
rect 13190 9851 13200 9907
rect 13256 9851 13324 9907
rect 13380 9851 13448 9907
rect 13504 9851 13572 9907
rect 13628 9851 13638 9907
rect 13190 9783 13638 9851
rect 13190 9727 13200 9783
rect 13256 9727 13324 9783
rect 13380 9727 13448 9783
rect 13504 9727 13572 9783
rect 13628 9727 13638 9783
rect 13190 9659 13638 9727
rect 13190 9603 13200 9659
rect 13256 9603 13324 9659
rect 13380 9603 13448 9659
rect 13504 9603 13572 9659
rect 13628 9603 13638 9659
rect 13190 9535 13638 9603
rect 13190 9479 13200 9535
rect 13256 9479 13324 9535
rect 13380 9479 13448 9535
rect 13504 9479 13572 9535
rect 13628 9479 13638 9535
rect 13190 9411 13638 9479
rect 13190 9355 13200 9411
rect 13256 9355 13324 9411
rect 13380 9355 13448 9411
rect 13504 9355 13572 9411
rect 13628 9355 13638 9411
rect 13190 9287 13638 9355
rect 13190 9231 13200 9287
rect 13256 9231 13324 9287
rect 13380 9231 13448 9287
rect 13504 9231 13572 9287
rect 13628 9231 13638 9287
rect 13190 9163 13638 9231
rect 13190 9107 13200 9163
rect 13256 9107 13324 9163
rect 13380 9107 13448 9163
rect 13504 9107 13572 9163
rect 13628 9107 13638 9163
rect 13190 9039 13638 9107
rect 13190 8983 13200 9039
rect 13256 8983 13324 9039
rect 13380 8983 13448 9039
rect 13504 8983 13572 9039
rect 13628 8983 13638 9039
rect 13190 8915 13638 8983
rect 13190 8859 13200 8915
rect 13256 8859 13324 8915
rect 13380 8859 13448 8915
rect 13504 8859 13572 8915
rect 13628 8859 13638 8915
rect 13190 8791 13638 8859
rect 13190 8735 13200 8791
rect 13256 8735 13324 8791
rect 13380 8735 13448 8791
rect 13504 8735 13572 8791
rect 13628 8735 13638 8791
rect 13190 8667 13638 8735
rect 13190 8611 13200 8667
rect 13256 8611 13324 8667
rect 13380 8611 13448 8667
rect 13504 8611 13572 8667
rect 13628 8611 13638 8667
rect 13190 8543 13638 8611
rect 13190 8487 13200 8543
rect 13256 8487 13324 8543
rect 13380 8487 13448 8543
rect 13504 8487 13572 8543
rect 13628 8487 13638 8543
rect 13190 8419 13638 8487
rect 13190 8363 13200 8419
rect 13256 8363 13324 8419
rect 13380 8363 13448 8419
rect 13504 8363 13572 8419
rect 13628 8363 13638 8419
rect 13190 8295 13638 8363
rect 13190 8239 13200 8295
rect 13256 8239 13324 8295
rect 13380 8239 13448 8295
rect 13504 8239 13572 8295
rect 13628 8239 13638 8295
rect 13190 8171 13638 8239
rect 13190 8115 13200 8171
rect 13256 8115 13324 8171
rect 13380 8115 13448 8171
rect 13504 8115 13572 8171
rect 13628 8115 13638 8171
rect 13190 8047 13638 8115
rect 13190 7991 13200 8047
rect 13256 7991 13324 8047
rect 13380 7991 13448 8047
rect 13504 7991 13572 8047
rect 13628 7991 13638 8047
rect 13190 7923 13638 7991
rect 13190 7867 13200 7923
rect 13256 7867 13324 7923
rect 13380 7867 13448 7923
rect 13504 7867 13572 7923
rect 13628 7867 13638 7923
rect 13190 7799 13638 7867
rect 13190 7743 13200 7799
rect 13256 7743 13324 7799
rect 13380 7743 13448 7799
rect 13504 7743 13572 7799
rect 13628 7743 13638 7799
rect 13190 7733 13638 7743
rect 14326 10651 14774 10661
rect 14326 10595 14336 10651
rect 14392 10595 14460 10651
rect 14516 10595 14584 10651
rect 14640 10595 14708 10651
rect 14764 10595 14774 10651
rect 14326 10527 14774 10595
rect 14326 10471 14336 10527
rect 14392 10471 14460 10527
rect 14516 10471 14584 10527
rect 14640 10471 14708 10527
rect 14764 10471 14774 10527
rect 14326 10403 14774 10471
rect 14326 10347 14336 10403
rect 14392 10347 14460 10403
rect 14516 10347 14584 10403
rect 14640 10347 14708 10403
rect 14764 10347 14774 10403
rect 14326 10279 14774 10347
rect 14326 10223 14336 10279
rect 14392 10223 14460 10279
rect 14516 10223 14584 10279
rect 14640 10223 14708 10279
rect 14764 10223 14774 10279
rect 14326 10155 14774 10223
rect 14326 10099 14336 10155
rect 14392 10099 14460 10155
rect 14516 10099 14584 10155
rect 14640 10099 14708 10155
rect 14764 10099 14774 10155
rect 14326 10031 14774 10099
rect 14326 9975 14336 10031
rect 14392 9975 14460 10031
rect 14516 9975 14584 10031
rect 14640 9975 14708 10031
rect 14764 9975 14774 10031
rect 14326 9907 14774 9975
rect 14326 9851 14336 9907
rect 14392 9851 14460 9907
rect 14516 9851 14584 9907
rect 14640 9851 14708 9907
rect 14764 9851 14774 9907
rect 14326 9783 14774 9851
rect 14326 9727 14336 9783
rect 14392 9727 14460 9783
rect 14516 9727 14584 9783
rect 14640 9727 14708 9783
rect 14764 9727 14774 9783
rect 14326 9659 14774 9727
rect 14326 9603 14336 9659
rect 14392 9603 14460 9659
rect 14516 9603 14584 9659
rect 14640 9603 14708 9659
rect 14764 9603 14774 9659
rect 14326 9535 14774 9603
rect 14326 9479 14336 9535
rect 14392 9479 14460 9535
rect 14516 9479 14584 9535
rect 14640 9479 14708 9535
rect 14764 9479 14774 9535
rect 14326 9411 14774 9479
rect 14326 9355 14336 9411
rect 14392 9355 14460 9411
rect 14516 9355 14584 9411
rect 14640 9355 14708 9411
rect 14764 9355 14774 9411
rect 14326 9287 14774 9355
rect 14326 9231 14336 9287
rect 14392 9231 14460 9287
rect 14516 9231 14584 9287
rect 14640 9231 14708 9287
rect 14764 9231 14774 9287
rect 14326 9163 14774 9231
rect 14326 9107 14336 9163
rect 14392 9107 14460 9163
rect 14516 9107 14584 9163
rect 14640 9107 14708 9163
rect 14764 9107 14774 9163
rect 14326 9039 14774 9107
rect 14326 8983 14336 9039
rect 14392 8983 14460 9039
rect 14516 8983 14584 9039
rect 14640 8983 14708 9039
rect 14764 8983 14774 9039
rect 14326 8915 14774 8983
rect 14326 8859 14336 8915
rect 14392 8859 14460 8915
rect 14516 8859 14584 8915
rect 14640 8859 14708 8915
rect 14764 8859 14774 8915
rect 14326 8791 14774 8859
rect 14326 8735 14336 8791
rect 14392 8735 14460 8791
rect 14516 8735 14584 8791
rect 14640 8735 14708 8791
rect 14764 8735 14774 8791
rect 14326 8667 14774 8735
rect 14326 8611 14336 8667
rect 14392 8611 14460 8667
rect 14516 8611 14584 8667
rect 14640 8611 14708 8667
rect 14764 8611 14774 8667
rect 14326 8543 14774 8611
rect 14326 8487 14336 8543
rect 14392 8487 14460 8543
rect 14516 8487 14584 8543
rect 14640 8487 14708 8543
rect 14764 8487 14774 8543
rect 14326 8419 14774 8487
rect 14326 8363 14336 8419
rect 14392 8363 14460 8419
rect 14516 8363 14584 8419
rect 14640 8363 14708 8419
rect 14764 8363 14774 8419
rect 14326 8295 14774 8363
rect 14326 8239 14336 8295
rect 14392 8239 14460 8295
rect 14516 8239 14584 8295
rect 14640 8239 14708 8295
rect 14764 8239 14774 8295
rect 14326 8171 14774 8239
rect 14326 8115 14336 8171
rect 14392 8115 14460 8171
rect 14516 8115 14584 8171
rect 14640 8115 14708 8171
rect 14764 8115 14774 8171
rect 14326 8047 14774 8115
rect 14326 7991 14336 8047
rect 14392 7991 14460 8047
rect 14516 7991 14584 8047
rect 14640 7991 14708 8047
rect 14764 7991 14774 8047
rect 14326 7923 14774 7991
rect 14326 7867 14336 7923
rect 14392 7867 14460 7923
rect 14516 7867 14584 7923
rect 14640 7867 14708 7923
rect 14764 7867 14774 7923
rect 14326 7799 14774 7867
rect 14326 7743 14336 7799
rect 14392 7743 14460 7799
rect 14516 7743 14584 7799
rect 14640 7743 14708 7799
rect 14764 7743 14774 7799
rect 14326 7733 14774 7743
rect 290 7451 738 7461
rect 290 7395 300 7451
rect 356 7395 424 7451
rect 480 7395 548 7451
rect 604 7395 672 7451
rect 728 7395 738 7451
rect 290 7327 738 7395
rect 290 7271 300 7327
rect 356 7271 424 7327
rect 480 7271 548 7327
rect 604 7271 672 7327
rect 728 7271 738 7327
rect 290 7203 738 7271
rect 290 7147 300 7203
rect 356 7147 424 7203
rect 480 7147 548 7203
rect 604 7147 672 7203
rect 728 7147 738 7203
rect 290 7079 738 7147
rect 290 7023 300 7079
rect 356 7023 424 7079
rect 480 7023 548 7079
rect 604 7023 672 7079
rect 728 7023 738 7079
rect 290 6955 738 7023
rect 290 6899 300 6955
rect 356 6899 424 6955
rect 480 6899 548 6955
rect 604 6899 672 6955
rect 728 6899 738 6955
rect 290 6831 738 6899
rect 290 6775 300 6831
rect 356 6775 424 6831
rect 480 6775 548 6831
rect 604 6775 672 6831
rect 728 6775 738 6831
rect 290 6707 738 6775
rect 290 6651 300 6707
rect 356 6651 424 6707
rect 480 6651 548 6707
rect 604 6651 672 6707
rect 728 6651 738 6707
rect 290 6583 738 6651
rect 290 6527 300 6583
rect 356 6527 424 6583
rect 480 6527 548 6583
rect 604 6527 672 6583
rect 728 6527 738 6583
rect 290 6459 738 6527
rect 290 6403 300 6459
rect 356 6403 424 6459
rect 480 6403 548 6459
rect 604 6403 672 6459
rect 728 6403 738 6459
rect 290 6335 738 6403
rect 290 6279 300 6335
rect 356 6279 424 6335
rect 480 6279 548 6335
rect 604 6279 672 6335
rect 728 6279 738 6335
rect 290 6211 738 6279
rect 290 6155 300 6211
rect 356 6155 424 6211
rect 480 6155 548 6211
rect 604 6155 672 6211
rect 728 6155 738 6211
rect 290 6087 738 6155
rect 290 6031 300 6087
rect 356 6031 424 6087
rect 480 6031 548 6087
rect 604 6031 672 6087
rect 728 6031 738 6087
rect 290 5963 738 6031
rect 290 5907 300 5963
rect 356 5907 424 5963
rect 480 5907 548 5963
rect 604 5907 672 5963
rect 728 5907 738 5963
rect 290 5839 738 5907
rect 290 5783 300 5839
rect 356 5783 424 5839
rect 480 5783 548 5839
rect 604 5783 672 5839
rect 728 5783 738 5839
rect 290 5715 738 5783
rect 290 5659 300 5715
rect 356 5659 424 5715
rect 480 5659 548 5715
rect 604 5659 672 5715
rect 728 5659 738 5715
rect 290 5591 738 5659
rect 290 5535 300 5591
rect 356 5535 424 5591
rect 480 5535 548 5591
rect 604 5535 672 5591
rect 728 5535 738 5591
rect 290 5467 738 5535
rect 290 5411 300 5467
rect 356 5411 424 5467
rect 480 5411 548 5467
rect 604 5411 672 5467
rect 728 5411 738 5467
rect 290 5343 738 5411
rect 290 5287 300 5343
rect 356 5287 424 5343
rect 480 5287 548 5343
rect 604 5287 672 5343
rect 728 5287 738 5343
rect 290 5219 738 5287
rect 290 5163 300 5219
rect 356 5163 424 5219
rect 480 5163 548 5219
rect 604 5163 672 5219
rect 728 5163 738 5219
rect 290 5095 738 5163
rect 290 5039 300 5095
rect 356 5039 424 5095
rect 480 5039 548 5095
rect 604 5039 672 5095
rect 728 5039 738 5095
rect 290 4971 738 5039
rect 290 4915 300 4971
rect 356 4915 424 4971
rect 480 4915 548 4971
rect 604 4915 672 4971
rect 728 4915 738 4971
rect 290 4847 738 4915
rect 290 4791 300 4847
rect 356 4791 424 4847
rect 480 4791 548 4847
rect 604 4791 672 4847
rect 728 4791 738 4847
rect 290 4723 738 4791
rect 290 4667 300 4723
rect 356 4667 424 4723
rect 480 4667 548 4723
rect 604 4667 672 4723
rect 728 4667 738 4723
rect 290 4599 738 4667
rect 290 4543 300 4599
rect 356 4543 424 4599
rect 480 4543 548 4599
rect 604 4543 672 4599
rect 728 4543 738 4599
rect 290 4533 738 4543
rect 1426 7451 1874 7461
rect 1426 7395 1436 7451
rect 1492 7395 1560 7451
rect 1616 7395 1684 7451
rect 1740 7395 1808 7451
rect 1864 7395 1874 7451
rect 1426 7327 1874 7395
rect 1426 7271 1436 7327
rect 1492 7271 1560 7327
rect 1616 7271 1684 7327
rect 1740 7271 1808 7327
rect 1864 7271 1874 7327
rect 1426 7203 1874 7271
rect 1426 7147 1436 7203
rect 1492 7147 1560 7203
rect 1616 7147 1684 7203
rect 1740 7147 1808 7203
rect 1864 7147 1874 7203
rect 1426 7079 1874 7147
rect 1426 7023 1436 7079
rect 1492 7023 1560 7079
rect 1616 7023 1684 7079
rect 1740 7023 1808 7079
rect 1864 7023 1874 7079
rect 1426 6955 1874 7023
rect 1426 6899 1436 6955
rect 1492 6899 1560 6955
rect 1616 6899 1684 6955
rect 1740 6899 1808 6955
rect 1864 6899 1874 6955
rect 1426 6831 1874 6899
rect 1426 6775 1436 6831
rect 1492 6775 1560 6831
rect 1616 6775 1684 6831
rect 1740 6775 1808 6831
rect 1864 6775 1874 6831
rect 1426 6707 1874 6775
rect 1426 6651 1436 6707
rect 1492 6651 1560 6707
rect 1616 6651 1684 6707
rect 1740 6651 1808 6707
rect 1864 6651 1874 6707
rect 1426 6583 1874 6651
rect 1426 6527 1436 6583
rect 1492 6527 1560 6583
rect 1616 6527 1684 6583
rect 1740 6527 1808 6583
rect 1864 6527 1874 6583
rect 1426 6459 1874 6527
rect 1426 6403 1436 6459
rect 1492 6403 1560 6459
rect 1616 6403 1684 6459
rect 1740 6403 1808 6459
rect 1864 6403 1874 6459
rect 1426 6335 1874 6403
rect 1426 6279 1436 6335
rect 1492 6279 1560 6335
rect 1616 6279 1684 6335
rect 1740 6279 1808 6335
rect 1864 6279 1874 6335
rect 1426 6211 1874 6279
rect 1426 6155 1436 6211
rect 1492 6155 1560 6211
rect 1616 6155 1684 6211
rect 1740 6155 1808 6211
rect 1864 6155 1874 6211
rect 1426 6087 1874 6155
rect 1426 6031 1436 6087
rect 1492 6031 1560 6087
rect 1616 6031 1684 6087
rect 1740 6031 1808 6087
rect 1864 6031 1874 6087
rect 1426 5963 1874 6031
rect 1426 5907 1436 5963
rect 1492 5907 1560 5963
rect 1616 5907 1684 5963
rect 1740 5907 1808 5963
rect 1864 5907 1874 5963
rect 1426 5839 1874 5907
rect 1426 5783 1436 5839
rect 1492 5783 1560 5839
rect 1616 5783 1684 5839
rect 1740 5783 1808 5839
rect 1864 5783 1874 5839
rect 1426 5715 1874 5783
rect 1426 5659 1436 5715
rect 1492 5659 1560 5715
rect 1616 5659 1684 5715
rect 1740 5659 1808 5715
rect 1864 5659 1874 5715
rect 1426 5591 1874 5659
rect 1426 5535 1436 5591
rect 1492 5535 1560 5591
rect 1616 5535 1684 5591
rect 1740 5535 1808 5591
rect 1864 5535 1874 5591
rect 1426 5467 1874 5535
rect 1426 5411 1436 5467
rect 1492 5411 1560 5467
rect 1616 5411 1684 5467
rect 1740 5411 1808 5467
rect 1864 5411 1874 5467
rect 1426 5343 1874 5411
rect 1426 5287 1436 5343
rect 1492 5287 1560 5343
rect 1616 5287 1684 5343
rect 1740 5287 1808 5343
rect 1864 5287 1874 5343
rect 1426 5219 1874 5287
rect 1426 5163 1436 5219
rect 1492 5163 1560 5219
rect 1616 5163 1684 5219
rect 1740 5163 1808 5219
rect 1864 5163 1874 5219
rect 1426 5095 1874 5163
rect 1426 5039 1436 5095
rect 1492 5039 1560 5095
rect 1616 5039 1684 5095
rect 1740 5039 1808 5095
rect 1864 5039 1874 5095
rect 1426 4971 1874 5039
rect 1426 4915 1436 4971
rect 1492 4915 1560 4971
rect 1616 4915 1684 4971
rect 1740 4915 1808 4971
rect 1864 4915 1874 4971
rect 1426 4847 1874 4915
rect 1426 4791 1436 4847
rect 1492 4791 1560 4847
rect 1616 4791 1684 4847
rect 1740 4791 1808 4847
rect 1864 4791 1874 4847
rect 1426 4723 1874 4791
rect 1426 4667 1436 4723
rect 1492 4667 1560 4723
rect 1616 4667 1684 4723
rect 1740 4667 1808 4723
rect 1864 4667 1874 4723
rect 1426 4599 1874 4667
rect 1426 4543 1436 4599
rect 1492 4543 1560 4599
rect 1616 4543 1684 4599
rect 1740 4543 1808 4599
rect 1864 4543 1874 4599
rect 1426 4533 1874 4543
rect 2562 7451 3010 7461
rect 2562 7395 2572 7451
rect 2628 7395 2696 7451
rect 2752 7395 2820 7451
rect 2876 7395 2944 7451
rect 3000 7395 3010 7451
rect 2562 7327 3010 7395
rect 2562 7271 2572 7327
rect 2628 7271 2696 7327
rect 2752 7271 2820 7327
rect 2876 7271 2944 7327
rect 3000 7271 3010 7327
rect 2562 7203 3010 7271
rect 2562 7147 2572 7203
rect 2628 7147 2696 7203
rect 2752 7147 2820 7203
rect 2876 7147 2944 7203
rect 3000 7147 3010 7203
rect 2562 7079 3010 7147
rect 2562 7023 2572 7079
rect 2628 7023 2696 7079
rect 2752 7023 2820 7079
rect 2876 7023 2944 7079
rect 3000 7023 3010 7079
rect 2562 6955 3010 7023
rect 2562 6899 2572 6955
rect 2628 6899 2696 6955
rect 2752 6899 2820 6955
rect 2876 6899 2944 6955
rect 3000 6899 3010 6955
rect 2562 6831 3010 6899
rect 2562 6775 2572 6831
rect 2628 6775 2696 6831
rect 2752 6775 2820 6831
rect 2876 6775 2944 6831
rect 3000 6775 3010 6831
rect 2562 6707 3010 6775
rect 2562 6651 2572 6707
rect 2628 6651 2696 6707
rect 2752 6651 2820 6707
rect 2876 6651 2944 6707
rect 3000 6651 3010 6707
rect 2562 6583 3010 6651
rect 2562 6527 2572 6583
rect 2628 6527 2696 6583
rect 2752 6527 2820 6583
rect 2876 6527 2944 6583
rect 3000 6527 3010 6583
rect 2562 6459 3010 6527
rect 2562 6403 2572 6459
rect 2628 6403 2696 6459
rect 2752 6403 2820 6459
rect 2876 6403 2944 6459
rect 3000 6403 3010 6459
rect 2562 6335 3010 6403
rect 2562 6279 2572 6335
rect 2628 6279 2696 6335
rect 2752 6279 2820 6335
rect 2876 6279 2944 6335
rect 3000 6279 3010 6335
rect 2562 6211 3010 6279
rect 2562 6155 2572 6211
rect 2628 6155 2696 6211
rect 2752 6155 2820 6211
rect 2876 6155 2944 6211
rect 3000 6155 3010 6211
rect 2562 6087 3010 6155
rect 2562 6031 2572 6087
rect 2628 6031 2696 6087
rect 2752 6031 2820 6087
rect 2876 6031 2944 6087
rect 3000 6031 3010 6087
rect 2562 5963 3010 6031
rect 2562 5907 2572 5963
rect 2628 5907 2696 5963
rect 2752 5907 2820 5963
rect 2876 5907 2944 5963
rect 3000 5907 3010 5963
rect 2562 5839 3010 5907
rect 2562 5783 2572 5839
rect 2628 5783 2696 5839
rect 2752 5783 2820 5839
rect 2876 5783 2944 5839
rect 3000 5783 3010 5839
rect 2562 5715 3010 5783
rect 2562 5659 2572 5715
rect 2628 5659 2696 5715
rect 2752 5659 2820 5715
rect 2876 5659 2944 5715
rect 3000 5659 3010 5715
rect 2562 5591 3010 5659
rect 2562 5535 2572 5591
rect 2628 5535 2696 5591
rect 2752 5535 2820 5591
rect 2876 5535 2944 5591
rect 3000 5535 3010 5591
rect 2562 5467 3010 5535
rect 2562 5411 2572 5467
rect 2628 5411 2696 5467
rect 2752 5411 2820 5467
rect 2876 5411 2944 5467
rect 3000 5411 3010 5467
rect 2562 5343 3010 5411
rect 2562 5287 2572 5343
rect 2628 5287 2696 5343
rect 2752 5287 2820 5343
rect 2876 5287 2944 5343
rect 3000 5287 3010 5343
rect 2562 5219 3010 5287
rect 2562 5163 2572 5219
rect 2628 5163 2696 5219
rect 2752 5163 2820 5219
rect 2876 5163 2944 5219
rect 3000 5163 3010 5219
rect 2562 5095 3010 5163
rect 2562 5039 2572 5095
rect 2628 5039 2696 5095
rect 2752 5039 2820 5095
rect 2876 5039 2944 5095
rect 3000 5039 3010 5095
rect 2562 4971 3010 5039
rect 2562 4915 2572 4971
rect 2628 4915 2696 4971
rect 2752 4915 2820 4971
rect 2876 4915 2944 4971
rect 3000 4915 3010 4971
rect 2562 4847 3010 4915
rect 2562 4791 2572 4847
rect 2628 4791 2696 4847
rect 2752 4791 2820 4847
rect 2876 4791 2944 4847
rect 3000 4791 3010 4847
rect 2562 4723 3010 4791
rect 2562 4667 2572 4723
rect 2628 4667 2696 4723
rect 2752 4667 2820 4723
rect 2876 4667 2944 4723
rect 3000 4667 3010 4723
rect 2562 4599 3010 4667
rect 2562 4543 2572 4599
rect 2628 4543 2696 4599
rect 2752 4543 2820 4599
rect 2876 4543 2944 4599
rect 3000 4543 3010 4599
rect 2562 4533 3010 4543
rect 4834 7451 5282 7461
rect 4834 7395 4844 7451
rect 4900 7395 4968 7451
rect 5024 7395 5092 7451
rect 5148 7395 5216 7451
rect 5272 7395 5282 7451
rect 4834 7327 5282 7395
rect 4834 7271 4844 7327
rect 4900 7271 4968 7327
rect 5024 7271 5092 7327
rect 5148 7271 5216 7327
rect 5272 7271 5282 7327
rect 4834 7203 5282 7271
rect 4834 7147 4844 7203
rect 4900 7147 4968 7203
rect 5024 7147 5092 7203
rect 5148 7147 5216 7203
rect 5272 7147 5282 7203
rect 4834 7079 5282 7147
rect 4834 7023 4844 7079
rect 4900 7023 4968 7079
rect 5024 7023 5092 7079
rect 5148 7023 5216 7079
rect 5272 7023 5282 7079
rect 4834 6955 5282 7023
rect 4834 6899 4844 6955
rect 4900 6899 4968 6955
rect 5024 6899 5092 6955
rect 5148 6899 5216 6955
rect 5272 6899 5282 6955
rect 4834 6831 5282 6899
rect 4834 6775 4844 6831
rect 4900 6775 4968 6831
rect 5024 6775 5092 6831
rect 5148 6775 5216 6831
rect 5272 6775 5282 6831
rect 4834 6707 5282 6775
rect 4834 6651 4844 6707
rect 4900 6651 4968 6707
rect 5024 6651 5092 6707
rect 5148 6651 5216 6707
rect 5272 6651 5282 6707
rect 4834 6583 5282 6651
rect 4834 6527 4844 6583
rect 4900 6527 4968 6583
rect 5024 6527 5092 6583
rect 5148 6527 5216 6583
rect 5272 6527 5282 6583
rect 4834 6459 5282 6527
rect 4834 6403 4844 6459
rect 4900 6403 4968 6459
rect 5024 6403 5092 6459
rect 5148 6403 5216 6459
rect 5272 6403 5282 6459
rect 4834 6335 5282 6403
rect 4834 6279 4844 6335
rect 4900 6279 4968 6335
rect 5024 6279 5092 6335
rect 5148 6279 5216 6335
rect 5272 6279 5282 6335
rect 4834 6211 5282 6279
rect 4834 6155 4844 6211
rect 4900 6155 4968 6211
rect 5024 6155 5092 6211
rect 5148 6155 5216 6211
rect 5272 6155 5282 6211
rect 4834 6087 5282 6155
rect 4834 6031 4844 6087
rect 4900 6031 4968 6087
rect 5024 6031 5092 6087
rect 5148 6031 5216 6087
rect 5272 6031 5282 6087
rect 4834 5963 5282 6031
rect 4834 5907 4844 5963
rect 4900 5907 4968 5963
rect 5024 5907 5092 5963
rect 5148 5907 5216 5963
rect 5272 5907 5282 5963
rect 4834 5839 5282 5907
rect 4834 5783 4844 5839
rect 4900 5783 4968 5839
rect 5024 5783 5092 5839
rect 5148 5783 5216 5839
rect 5272 5783 5282 5839
rect 4834 5715 5282 5783
rect 4834 5659 4844 5715
rect 4900 5659 4968 5715
rect 5024 5659 5092 5715
rect 5148 5659 5216 5715
rect 5272 5659 5282 5715
rect 4834 5591 5282 5659
rect 4834 5535 4844 5591
rect 4900 5535 4968 5591
rect 5024 5535 5092 5591
rect 5148 5535 5216 5591
rect 5272 5535 5282 5591
rect 4834 5467 5282 5535
rect 4834 5411 4844 5467
rect 4900 5411 4968 5467
rect 5024 5411 5092 5467
rect 5148 5411 5216 5467
rect 5272 5411 5282 5467
rect 4834 5343 5282 5411
rect 4834 5287 4844 5343
rect 4900 5287 4968 5343
rect 5024 5287 5092 5343
rect 5148 5287 5216 5343
rect 5272 5287 5282 5343
rect 4834 5219 5282 5287
rect 4834 5163 4844 5219
rect 4900 5163 4968 5219
rect 5024 5163 5092 5219
rect 5148 5163 5216 5219
rect 5272 5163 5282 5219
rect 4834 5095 5282 5163
rect 4834 5039 4844 5095
rect 4900 5039 4968 5095
rect 5024 5039 5092 5095
rect 5148 5039 5216 5095
rect 5272 5039 5282 5095
rect 4834 4971 5282 5039
rect 4834 4915 4844 4971
rect 4900 4915 4968 4971
rect 5024 4915 5092 4971
rect 5148 4915 5216 4971
rect 5272 4915 5282 4971
rect 4834 4847 5282 4915
rect 4834 4791 4844 4847
rect 4900 4791 4968 4847
rect 5024 4791 5092 4847
rect 5148 4791 5216 4847
rect 5272 4791 5282 4847
rect 4834 4723 5282 4791
rect 4834 4667 4844 4723
rect 4900 4667 4968 4723
rect 5024 4667 5092 4723
rect 5148 4667 5216 4723
rect 5272 4667 5282 4723
rect 4834 4599 5282 4667
rect 4834 4543 4844 4599
rect 4900 4543 4968 4599
rect 5024 4543 5092 4599
rect 5148 4543 5216 4599
rect 5272 4543 5282 4599
rect 4834 4533 5282 4543
rect 7127 7451 7451 7461
rect 7127 7395 7137 7451
rect 7193 7395 7261 7451
rect 7317 7395 7385 7451
rect 7441 7395 7451 7451
rect 7127 7327 7451 7395
rect 7127 7271 7137 7327
rect 7193 7271 7261 7327
rect 7317 7271 7385 7327
rect 7441 7271 7451 7327
rect 7127 7203 7451 7271
rect 7127 7147 7137 7203
rect 7193 7147 7261 7203
rect 7317 7147 7385 7203
rect 7441 7147 7451 7203
rect 7127 7079 7451 7147
rect 7127 7023 7137 7079
rect 7193 7023 7261 7079
rect 7317 7023 7385 7079
rect 7441 7023 7451 7079
rect 7127 6955 7451 7023
rect 7127 6899 7137 6955
rect 7193 6899 7261 6955
rect 7317 6899 7385 6955
rect 7441 6899 7451 6955
rect 7127 6831 7451 6899
rect 7127 6775 7137 6831
rect 7193 6775 7261 6831
rect 7317 6775 7385 6831
rect 7441 6775 7451 6831
rect 7127 6707 7451 6775
rect 7127 6651 7137 6707
rect 7193 6651 7261 6707
rect 7317 6651 7385 6707
rect 7441 6651 7451 6707
rect 7127 6583 7451 6651
rect 7127 6527 7137 6583
rect 7193 6527 7261 6583
rect 7317 6527 7385 6583
rect 7441 6527 7451 6583
rect 7127 6459 7451 6527
rect 7127 6403 7137 6459
rect 7193 6403 7261 6459
rect 7317 6403 7385 6459
rect 7441 6403 7451 6459
rect 7127 6335 7451 6403
rect 7127 6279 7137 6335
rect 7193 6279 7261 6335
rect 7317 6279 7385 6335
rect 7441 6279 7451 6335
rect 7127 6211 7451 6279
rect 7127 6155 7137 6211
rect 7193 6155 7261 6211
rect 7317 6155 7385 6211
rect 7441 6155 7451 6211
rect 7127 6087 7451 6155
rect 7127 6031 7137 6087
rect 7193 6031 7261 6087
rect 7317 6031 7385 6087
rect 7441 6031 7451 6087
rect 7127 5963 7451 6031
rect 7127 5907 7137 5963
rect 7193 5907 7261 5963
rect 7317 5907 7385 5963
rect 7441 5907 7451 5963
rect 7127 5839 7451 5907
rect 7127 5783 7137 5839
rect 7193 5783 7261 5839
rect 7317 5783 7385 5839
rect 7441 5783 7451 5839
rect 7127 5715 7451 5783
rect 7127 5659 7137 5715
rect 7193 5659 7261 5715
rect 7317 5659 7385 5715
rect 7441 5659 7451 5715
rect 7127 5591 7451 5659
rect 7127 5535 7137 5591
rect 7193 5535 7261 5591
rect 7317 5535 7385 5591
rect 7441 5535 7451 5591
rect 7127 5467 7451 5535
rect 7127 5411 7137 5467
rect 7193 5411 7261 5467
rect 7317 5411 7385 5467
rect 7441 5411 7451 5467
rect 7127 5343 7451 5411
rect 7127 5287 7137 5343
rect 7193 5287 7261 5343
rect 7317 5287 7385 5343
rect 7441 5287 7451 5343
rect 7127 5219 7451 5287
rect 7127 5163 7137 5219
rect 7193 5163 7261 5219
rect 7317 5163 7385 5219
rect 7441 5163 7451 5219
rect 7127 5095 7451 5163
rect 7127 5039 7137 5095
rect 7193 5039 7261 5095
rect 7317 5039 7385 5095
rect 7441 5039 7451 5095
rect 7127 4971 7451 5039
rect 7127 4915 7137 4971
rect 7193 4915 7261 4971
rect 7317 4915 7385 4971
rect 7441 4915 7451 4971
rect 7127 4847 7451 4915
rect 7127 4791 7137 4847
rect 7193 4791 7261 4847
rect 7317 4791 7385 4847
rect 7441 4791 7451 4847
rect 7127 4723 7451 4791
rect 7127 4667 7137 4723
rect 7193 4667 7261 4723
rect 7317 4667 7385 4723
rect 7441 4667 7451 4723
rect 7127 4599 7451 4667
rect 7127 4543 7137 4599
rect 7193 4543 7261 4599
rect 7317 4543 7385 4599
rect 7441 4543 7451 4599
rect 7127 4533 7451 4543
rect 7613 7451 7937 7461
rect 7613 7395 7623 7451
rect 7679 7395 7747 7451
rect 7803 7395 7871 7451
rect 7927 7395 7937 7451
rect 7613 7327 7937 7395
rect 7613 7271 7623 7327
rect 7679 7271 7747 7327
rect 7803 7271 7871 7327
rect 7927 7271 7937 7327
rect 7613 7203 7937 7271
rect 7613 7147 7623 7203
rect 7679 7147 7747 7203
rect 7803 7147 7871 7203
rect 7927 7147 7937 7203
rect 7613 7079 7937 7147
rect 7613 7023 7623 7079
rect 7679 7023 7747 7079
rect 7803 7023 7871 7079
rect 7927 7023 7937 7079
rect 7613 6955 7937 7023
rect 7613 6899 7623 6955
rect 7679 6899 7747 6955
rect 7803 6899 7871 6955
rect 7927 6899 7937 6955
rect 7613 6831 7937 6899
rect 7613 6775 7623 6831
rect 7679 6775 7747 6831
rect 7803 6775 7871 6831
rect 7927 6775 7937 6831
rect 7613 6707 7937 6775
rect 7613 6651 7623 6707
rect 7679 6651 7747 6707
rect 7803 6651 7871 6707
rect 7927 6651 7937 6707
rect 7613 6583 7937 6651
rect 7613 6527 7623 6583
rect 7679 6527 7747 6583
rect 7803 6527 7871 6583
rect 7927 6527 7937 6583
rect 7613 6459 7937 6527
rect 7613 6403 7623 6459
rect 7679 6403 7747 6459
rect 7803 6403 7871 6459
rect 7927 6403 7937 6459
rect 7613 6335 7937 6403
rect 7613 6279 7623 6335
rect 7679 6279 7747 6335
rect 7803 6279 7871 6335
rect 7927 6279 7937 6335
rect 7613 6211 7937 6279
rect 7613 6155 7623 6211
rect 7679 6155 7747 6211
rect 7803 6155 7871 6211
rect 7927 6155 7937 6211
rect 7613 6087 7937 6155
rect 7613 6031 7623 6087
rect 7679 6031 7747 6087
rect 7803 6031 7871 6087
rect 7927 6031 7937 6087
rect 7613 5963 7937 6031
rect 7613 5907 7623 5963
rect 7679 5907 7747 5963
rect 7803 5907 7871 5963
rect 7927 5907 7937 5963
rect 7613 5839 7937 5907
rect 7613 5783 7623 5839
rect 7679 5783 7747 5839
rect 7803 5783 7871 5839
rect 7927 5783 7937 5839
rect 7613 5715 7937 5783
rect 7613 5659 7623 5715
rect 7679 5659 7747 5715
rect 7803 5659 7871 5715
rect 7927 5659 7937 5715
rect 7613 5591 7937 5659
rect 7613 5535 7623 5591
rect 7679 5535 7747 5591
rect 7803 5535 7871 5591
rect 7927 5535 7937 5591
rect 7613 5467 7937 5535
rect 7613 5411 7623 5467
rect 7679 5411 7747 5467
rect 7803 5411 7871 5467
rect 7927 5411 7937 5467
rect 7613 5343 7937 5411
rect 7613 5287 7623 5343
rect 7679 5287 7747 5343
rect 7803 5287 7871 5343
rect 7927 5287 7937 5343
rect 7613 5219 7937 5287
rect 7613 5163 7623 5219
rect 7679 5163 7747 5219
rect 7803 5163 7871 5219
rect 7927 5163 7937 5219
rect 7613 5095 7937 5163
rect 7613 5039 7623 5095
rect 7679 5039 7747 5095
rect 7803 5039 7871 5095
rect 7927 5039 7937 5095
rect 7613 4971 7937 5039
rect 7613 4915 7623 4971
rect 7679 4915 7747 4971
rect 7803 4915 7871 4971
rect 7927 4915 7937 4971
rect 7613 4847 7937 4915
rect 7613 4791 7623 4847
rect 7679 4791 7747 4847
rect 7803 4791 7871 4847
rect 7927 4791 7937 4847
rect 7613 4723 7937 4791
rect 7613 4667 7623 4723
rect 7679 4667 7747 4723
rect 7803 4667 7871 4723
rect 7927 4667 7937 4723
rect 7613 4599 7937 4667
rect 7613 4543 7623 4599
rect 7679 4543 7747 4599
rect 7803 4543 7871 4599
rect 7927 4543 7937 4599
rect 7613 4533 7937 4543
rect 9782 7451 10230 7461
rect 9782 7395 9792 7451
rect 9848 7395 9916 7451
rect 9972 7395 10040 7451
rect 10096 7395 10164 7451
rect 10220 7395 10230 7451
rect 9782 7327 10230 7395
rect 9782 7271 9792 7327
rect 9848 7271 9916 7327
rect 9972 7271 10040 7327
rect 10096 7271 10164 7327
rect 10220 7271 10230 7327
rect 9782 7203 10230 7271
rect 9782 7147 9792 7203
rect 9848 7147 9916 7203
rect 9972 7147 10040 7203
rect 10096 7147 10164 7203
rect 10220 7147 10230 7203
rect 9782 7079 10230 7147
rect 9782 7023 9792 7079
rect 9848 7023 9916 7079
rect 9972 7023 10040 7079
rect 10096 7023 10164 7079
rect 10220 7023 10230 7079
rect 9782 6955 10230 7023
rect 9782 6899 9792 6955
rect 9848 6899 9916 6955
rect 9972 6899 10040 6955
rect 10096 6899 10164 6955
rect 10220 6899 10230 6955
rect 9782 6831 10230 6899
rect 9782 6775 9792 6831
rect 9848 6775 9916 6831
rect 9972 6775 10040 6831
rect 10096 6775 10164 6831
rect 10220 6775 10230 6831
rect 9782 6707 10230 6775
rect 9782 6651 9792 6707
rect 9848 6651 9916 6707
rect 9972 6651 10040 6707
rect 10096 6651 10164 6707
rect 10220 6651 10230 6707
rect 9782 6583 10230 6651
rect 9782 6527 9792 6583
rect 9848 6527 9916 6583
rect 9972 6527 10040 6583
rect 10096 6527 10164 6583
rect 10220 6527 10230 6583
rect 9782 6459 10230 6527
rect 9782 6403 9792 6459
rect 9848 6403 9916 6459
rect 9972 6403 10040 6459
rect 10096 6403 10164 6459
rect 10220 6403 10230 6459
rect 9782 6335 10230 6403
rect 9782 6279 9792 6335
rect 9848 6279 9916 6335
rect 9972 6279 10040 6335
rect 10096 6279 10164 6335
rect 10220 6279 10230 6335
rect 9782 6211 10230 6279
rect 9782 6155 9792 6211
rect 9848 6155 9916 6211
rect 9972 6155 10040 6211
rect 10096 6155 10164 6211
rect 10220 6155 10230 6211
rect 9782 6087 10230 6155
rect 9782 6031 9792 6087
rect 9848 6031 9916 6087
rect 9972 6031 10040 6087
rect 10096 6031 10164 6087
rect 10220 6031 10230 6087
rect 9782 5963 10230 6031
rect 9782 5907 9792 5963
rect 9848 5907 9916 5963
rect 9972 5907 10040 5963
rect 10096 5907 10164 5963
rect 10220 5907 10230 5963
rect 9782 5839 10230 5907
rect 9782 5783 9792 5839
rect 9848 5783 9916 5839
rect 9972 5783 10040 5839
rect 10096 5783 10164 5839
rect 10220 5783 10230 5839
rect 9782 5715 10230 5783
rect 9782 5659 9792 5715
rect 9848 5659 9916 5715
rect 9972 5659 10040 5715
rect 10096 5659 10164 5715
rect 10220 5659 10230 5715
rect 9782 5591 10230 5659
rect 9782 5535 9792 5591
rect 9848 5535 9916 5591
rect 9972 5535 10040 5591
rect 10096 5535 10164 5591
rect 10220 5535 10230 5591
rect 9782 5467 10230 5535
rect 9782 5411 9792 5467
rect 9848 5411 9916 5467
rect 9972 5411 10040 5467
rect 10096 5411 10164 5467
rect 10220 5411 10230 5467
rect 9782 5343 10230 5411
rect 9782 5287 9792 5343
rect 9848 5287 9916 5343
rect 9972 5287 10040 5343
rect 10096 5287 10164 5343
rect 10220 5287 10230 5343
rect 9782 5219 10230 5287
rect 9782 5163 9792 5219
rect 9848 5163 9916 5219
rect 9972 5163 10040 5219
rect 10096 5163 10164 5219
rect 10220 5163 10230 5219
rect 9782 5095 10230 5163
rect 9782 5039 9792 5095
rect 9848 5039 9916 5095
rect 9972 5039 10040 5095
rect 10096 5039 10164 5095
rect 10220 5039 10230 5095
rect 9782 4971 10230 5039
rect 9782 4915 9792 4971
rect 9848 4915 9916 4971
rect 9972 4915 10040 4971
rect 10096 4915 10164 4971
rect 10220 4915 10230 4971
rect 9782 4847 10230 4915
rect 9782 4791 9792 4847
rect 9848 4791 9916 4847
rect 9972 4791 10040 4847
rect 10096 4791 10164 4847
rect 10220 4791 10230 4847
rect 9782 4723 10230 4791
rect 9782 4667 9792 4723
rect 9848 4667 9916 4723
rect 9972 4667 10040 4723
rect 10096 4667 10164 4723
rect 10220 4667 10230 4723
rect 9782 4599 10230 4667
rect 9782 4543 9792 4599
rect 9848 4543 9916 4599
rect 9972 4543 10040 4599
rect 10096 4543 10164 4599
rect 10220 4543 10230 4599
rect 9782 4533 10230 4543
rect 12054 7451 12502 7461
rect 12054 7395 12064 7451
rect 12120 7395 12188 7451
rect 12244 7395 12312 7451
rect 12368 7395 12436 7451
rect 12492 7395 12502 7451
rect 12054 7327 12502 7395
rect 12054 7271 12064 7327
rect 12120 7271 12188 7327
rect 12244 7271 12312 7327
rect 12368 7271 12436 7327
rect 12492 7271 12502 7327
rect 12054 7203 12502 7271
rect 12054 7147 12064 7203
rect 12120 7147 12188 7203
rect 12244 7147 12312 7203
rect 12368 7147 12436 7203
rect 12492 7147 12502 7203
rect 12054 7079 12502 7147
rect 12054 7023 12064 7079
rect 12120 7023 12188 7079
rect 12244 7023 12312 7079
rect 12368 7023 12436 7079
rect 12492 7023 12502 7079
rect 12054 6955 12502 7023
rect 12054 6899 12064 6955
rect 12120 6899 12188 6955
rect 12244 6899 12312 6955
rect 12368 6899 12436 6955
rect 12492 6899 12502 6955
rect 12054 6831 12502 6899
rect 12054 6775 12064 6831
rect 12120 6775 12188 6831
rect 12244 6775 12312 6831
rect 12368 6775 12436 6831
rect 12492 6775 12502 6831
rect 12054 6707 12502 6775
rect 12054 6651 12064 6707
rect 12120 6651 12188 6707
rect 12244 6651 12312 6707
rect 12368 6651 12436 6707
rect 12492 6651 12502 6707
rect 12054 6583 12502 6651
rect 12054 6527 12064 6583
rect 12120 6527 12188 6583
rect 12244 6527 12312 6583
rect 12368 6527 12436 6583
rect 12492 6527 12502 6583
rect 12054 6459 12502 6527
rect 12054 6403 12064 6459
rect 12120 6403 12188 6459
rect 12244 6403 12312 6459
rect 12368 6403 12436 6459
rect 12492 6403 12502 6459
rect 12054 6335 12502 6403
rect 12054 6279 12064 6335
rect 12120 6279 12188 6335
rect 12244 6279 12312 6335
rect 12368 6279 12436 6335
rect 12492 6279 12502 6335
rect 12054 6211 12502 6279
rect 12054 6155 12064 6211
rect 12120 6155 12188 6211
rect 12244 6155 12312 6211
rect 12368 6155 12436 6211
rect 12492 6155 12502 6211
rect 12054 6087 12502 6155
rect 12054 6031 12064 6087
rect 12120 6031 12188 6087
rect 12244 6031 12312 6087
rect 12368 6031 12436 6087
rect 12492 6031 12502 6087
rect 12054 5963 12502 6031
rect 12054 5907 12064 5963
rect 12120 5907 12188 5963
rect 12244 5907 12312 5963
rect 12368 5907 12436 5963
rect 12492 5907 12502 5963
rect 12054 5839 12502 5907
rect 12054 5783 12064 5839
rect 12120 5783 12188 5839
rect 12244 5783 12312 5839
rect 12368 5783 12436 5839
rect 12492 5783 12502 5839
rect 12054 5715 12502 5783
rect 12054 5659 12064 5715
rect 12120 5659 12188 5715
rect 12244 5659 12312 5715
rect 12368 5659 12436 5715
rect 12492 5659 12502 5715
rect 12054 5591 12502 5659
rect 12054 5535 12064 5591
rect 12120 5535 12188 5591
rect 12244 5535 12312 5591
rect 12368 5535 12436 5591
rect 12492 5535 12502 5591
rect 12054 5467 12502 5535
rect 12054 5411 12064 5467
rect 12120 5411 12188 5467
rect 12244 5411 12312 5467
rect 12368 5411 12436 5467
rect 12492 5411 12502 5467
rect 12054 5343 12502 5411
rect 12054 5287 12064 5343
rect 12120 5287 12188 5343
rect 12244 5287 12312 5343
rect 12368 5287 12436 5343
rect 12492 5287 12502 5343
rect 12054 5219 12502 5287
rect 12054 5163 12064 5219
rect 12120 5163 12188 5219
rect 12244 5163 12312 5219
rect 12368 5163 12436 5219
rect 12492 5163 12502 5219
rect 12054 5095 12502 5163
rect 12054 5039 12064 5095
rect 12120 5039 12188 5095
rect 12244 5039 12312 5095
rect 12368 5039 12436 5095
rect 12492 5039 12502 5095
rect 12054 4971 12502 5039
rect 12054 4915 12064 4971
rect 12120 4915 12188 4971
rect 12244 4915 12312 4971
rect 12368 4915 12436 4971
rect 12492 4915 12502 4971
rect 12054 4847 12502 4915
rect 12054 4791 12064 4847
rect 12120 4791 12188 4847
rect 12244 4791 12312 4847
rect 12368 4791 12436 4847
rect 12492 4791 12502 4847
rect 12054 4723 12502 4791
rect 12054 4667 12064 4723
rect 12120 4667 12188 4723
rect 12244 4667 12312 4723
rect 12368 4667 12436 4723
rect 12492 4667 12502 4723
rect 12054 4599 12502 4667
rect 12054 4543 12064 4599
rect 12120 4543 12188 4599
rect 12244 4543 12312 4599
rect 12368 4543 12436 4599
rect 12492 4543 12502 4599
rect 12054 4533 12502 4543
rect 13190 7451 13638 7461
rect 13190 7395 13200 7451
rect 13256 7395 13324 7451
rect 13380 7395 13448 7451
rect 13504 7395 13572 7451
rect 13628 7395 13638 7451
rect 13190 7327 13638 7395
rect 13190 7271 13200 7327
rect 13256 7271 13324 7327
rect 13380 7271 13448 7327
rect 13504 7271 13572 7327
rect 13628 7271 13638 7327
rect 13190 7203 13638 7271
rect 13190 7147 13200 7203
rect 13256 7147 13324 7203
rect 13380 7147 13448 7203
rect 13504 7147 13572 7203
rect 13628 7147 13638 7203
rect 13190 7079 13638 7147
rect 13190 7023 13200 7079
rect 13256 7023 13324 7079
rect 13380 7023 13448 7079
rect 13504 7023 13572 7079
rect 13628 7023 13638 7079
rect 13190 6955 13638 7023
rect 13190 6899 13200 6955
rect 13256 6899 13324 6955
rect 13380 6899 13448 6955
rect 13504 6899 13572 6955
rect 13628 6899 13638 6955
rect 13190 6831 13638 6899
rect 13190 6775 13200 6831
rect 13256 6775 13324 6831
rect 13380 6775 13448 6831
rect 13504 6775 13572 6831
rect 13628 6775 13638 6831
rect 13190 6707 13638 6775
rect 13190 6651 13200 6707
rect 13256 6651 13324 6707
rect 13380 6651 13448 6707
rect 13504 6651 13572 6707
rect 13628 6651 13638 6707
rect 13190 6583 13638 6651
rect 13190 6527 13200 6583
rect 13256 6527 13324 6583
rect 13380 6527 13448 6583
rect 13504 6527 13572 6583
rect 13628 6527 13638 6583
rect 13190 6459 13638 6527
rect 13190 6403 13200 6459
rect 13256 6403 13324 6459
rect 13380 6403 13448 6459
rect 13504 6403 13572 6459
rect 13628 6403 13638 6459
rect 13190 6335 13638 6403
rect 13190 6279 13200 6335
rect 13256 6279 13324 6335
rect 13380 6279 13448 6335
rect 13504 6279 13572 6335
rect 13628 6279 13638 6335
rect 13190 6211 13638 6279
rect 13190 6155 13200 6211
rect 13256 6155 13324 6211
rect 13380 6155 13448 6211
rect 13504 6155 13572 6211
rect 13628 6155 13638 6211
rect 13190 6087 13638 6155
rect 13190 6031 13200 6087
rect 13256 6031 13324 6087
rect 13380 6031 13448 6087
rect 13504 6031 13572 6087
rect 13628 6031 13638 6087
rect 13190 5963 13638 6031
rect 13190 5907 13200 5963
rect 13256 5907 13324 5963
rect 13380 5907 13448 5963
rect 13504 5907 13572 5963
rect 13628 5907 13638 5963
rect 13190 5839 13638 5907
rect 13190 5783 13200 5839
rect 13256 5783 13324 5839
rect 13380 5783 13448 5839
rect 13504 5783 13572 5839
rect 13628 5783 13638 5839
rect 13190 5715 13638 5783
rect 13190 5659 13200 5715
rect 13256 5659 13324 5715
rect 13380 5659 13448 5715
rect 13504 5659 13572 5715
rect 13628 5659 13638 5715
rect 13190 5591 13638 5659
rect 13190 5535 13200 5591
rect 13256 5535 13324 5591
rect 13380 5535 13448 5591
rect 13504 5535 13572 5591
rect 13628 5535 13638 5591
rect 13190 5467 13638 5535
rect 13190 5411 13200 5467
rect 13256 5411 13324 5467
rect 13380 5411 13448 5467
rect 13504 5411 13572 5467
rect 13628 5411 13638 5467
rect 13190 5343 13638 5411
rect 13190 5287 13200 5343
rect 13256 5287 13324 5343
rect 13380 5287 13448 5343
rect 13504 5287 13572 5343
rect 13628 5287 13638 5343
rect 13190 5219 13638 5287
rect 13190 5163 13200 5219
rect 13256 5163 13324 5219
rect 13380 5163 13448 5219
rect 13504 5163 13572 5219
rect 13628 5163 13638 5219
rect 13190 5095 13638 5163
rect 13190 5039 13200 5095
rect 13256 5039 13324 5095
rect 13380 5039 13448 5095
rect 13504 5039 13572 5095
rect 13628 5039 13638 5095
rect 13190 4971 13638 5039
rect 13190 4915 13200 4971
rect 13256 4915 13324 4971
rect 13380 4915 13448 4971
rect 13504 4915 13572 4971
rect 13628 4915 13638 4971
rect 13190 4847 13638 4915
rect 13190 4791 13200 4847
rect 13256 4791 13324 4847
rect 13380 4791 13448 4847
rect 13504 4791 13572 4847
rect 13628 4791 13638 4847
rect 13190 4723 13638 4791
rect 13190 4667 13200 4723
rect 13256 4667 13324 4723
rect 13380 4667 13448 4723
rect 13504 4667 13572 4723
rect 13628 4667 13638 4723
rect 13190 4599 13638 4667
rect 13190 4543 13200 4599
rect 13256 4543 13324 4599
rect 13380 4543 13448 4599
rect 13504 4543 13572 4599
rect 13628 4543 13638 4599
rect 13190 4533 13638 4543
rect 14326 7451 14774 7461
rect 14326 7395 14336 7451
rect 14392 7395 14460 7451
rect 14516 7395 14584 7451
rect 14640 7395 14708 7451
rect 14764 7395 14774 7451
rect 14326 7327 14774 7395
rect 14326 7271 14336 7327
rect 14392 7271 14460 7327
rect 14516 7271 14584 7327
rect 14640 7271 14708 7327
rect 14764 7271 14774 7327
rect 14326 7203 14774 7271
rect 14326 7147 14336 7203
rect 14392 7147 14460 7203
rect 14516 7147 14584 7203
rect 14640 7147 14708 7203
rect 14764 7147 14774 7203
rect 14326 7079 14774 7147
rect 14326 7023 14336 7079
rect 14392 7023 14460 7079
rect 14516 7023 14584 7079
rect 14640 7023 14708 7079
rect 14764 7023 14774 7079
rect 14326 6955 14774 7023
rect 14326 6899 14336 6955
rect 14392 6899 14460 6955
rect 14516 6899 14584 6955
rect 14640 6899 14708 6955
rect 14764 6899 14774 6955
rect 14326 6831 14774 6899
rect 14326 6775 14336 6831
rect 14392 6775 14460 6831
rect 14516 6775 14584 6831
rect 14640 6775 14708 6831
rect 14764 6775 14774 6831
rect 14326 6707 14774 6775
rect 14326 6651 14336 6707
rect 14392 6651 14460 6707
rect 14516 6651 14584 6707
rect 14640 6651 14708 6707
rect 14764 6651 14774 6707
rect 14326 6583 14774 6651
rect 14326 6527 14336 6583
rect 14392 6527 14460 6583
rect 14516 6527 14584 6583
rect 14640 6527 14708 6583
rect 14764 6527 14774 6583
rect 14326 6459 14774 6527
rect 14326 6403 14336 6459
rect 14392 6403 14460 6459
rect 14516 6403 14584 6459
rect 14640 6403 14708 6459
rect 14764 6403 14774 6459
rect 14326 6335 14774 6403
rect 14326 6279 14336 6335
rect 14392 6279 14460 6335
rect 14516 6279 14584 6335
rect 14640 6279 14708 6335
rect 14764 6279 14774 6335
rect 14326 6211 14774 6279
rect 14326 6155 14336 6211
rect 14392 6155 14460 6211
rect 14516 6155 14584 6211
rect 14640 6155 14708 6211
rect 14764 6155 14774 6211
rect 14326 6087 14774 6155
rect 14326 6031 14336 6087
rect 14392 6031 14460 6087
rect 14516 6031 14584 6087
rect 14640 6031 14708 6087
rect 14764 6031 14774 6087
rect 14326 5963 14774 6031
rect 14326 5907 14336 5963
rect 14392 5907 14460 5963
rect 14516 5907 14584 5963
rect 14640 5907 14708 5963
rect 14764 5907 14774 5963
rect 14326 5839 14774 5907
rect 14326 5783 14336 5839
rect 14392 5783 14460 5839
rect 14516 5783 14584 5839
rect 14640 5783 14708 5839
rect 14764 5783 14774 5839
rect 14326 5715 14774 5783
rect 14326 5659 14336 5715
rect 14392 5659 14460 5715
rect 14516 5659 14584 5715
rect 14640 5659 14708 5715
rect 14764 5659 14774 5715
rect 14326 5591 14774 5659
rect 14326 5535 14336 5591
rect 14392 5535 14460 5591
rect 14516 5535 14584 5591
rect 14640 5535 14708 5591
rect 14764 5535 14774 5591
rect 14326 5467 14774 5535
rect 14326 5411 14336 5467
rect 14392 5411 14460 5467
rect 14516 5411 14584 5467
rect 14640 5411 14708 5467
rect 14764 5411 14774 5467
rect 14326 5343 14774 5411
rect 14326 5287 14336 5343
rect 14392 5287 14460 5343
rect 14516 5287 14584 5343
rect 14640 5287 14708 5343
rect 14764 5287 14774 5343
rect 14326 5219 14774 5287
rect 14326 5163 14336 5219
rect 14392 5163 14460 5219
rect 14516 5163 14584 5219
rect 14640 5163 14708 5219
rect 14764 5163 14774 5219
rect 14326 5095 14774 5163
rect 14326 5039 14336 5095
rect 14392 5039 14460 5095
rect 14516 5039 14584 5095
rect 14640 5039 14708 5095
rect 14764 5039 14774 5095
rect 14326 4971 14774 5039
rect 14326 4915 14336 4971
rect 14392 4915 14460 4971
rect 14516 4915 14584 4971
rect 14640 4915 14708 4971
rect 14764 4915 14774 4971
rect 14326 4847 14774 4915
rect 14326 4791 14336 4847
rect 14392 4791 14460 4847
rect 14516 4791 14584 4847
rect 14640 4791 14708 4847
rect 14764 4791 14774 4847
rect 14326 4723 14774 4791
rect 14326 4667 14336 4723
rect 14392 4667 14460 4723
rect 14516 4667 14584 4723
rect 14640 4667 14708 4723
rect 14764 4667 14774 4723
rect 14326 4599 14774 4667
rect 14326 4543 14336 4599
rect 14392 4543 14460 4599
rect 14516 4543 14584 4599
rect 14640 4543 14708 4599
rect 14764 4543 14774 4599
rect 14326 4533 14774 4543
rect 290 4251 738 4261
rect 290 4195 300 4251
rect 356 4195 424 4251
rect 480 4195 548 4251
rect 604 4195 672 4251
rect 728 4195 738 4251
rect 290 4127 738 4195
rect 290 4071 300 4127
rect 356 4071 424 4127
rect 480 4071 548 4127
rect 604 4071 672 4127
rect 728 4071 738 4127
rect 290 4003 738 4071
rect 290 3947 300 4003
rect 356 3947 424 4003
rect 480 3947 548 4003
rect 604 3947 672 4003
rect 728 3947 738 4003
rect 290 3879 738 3947
rect 290 3823 300 3879
rect 356 3823 424 3879
rect 480 3823 548 3879
rect 604 3823 672 3879
rect 728 3823 738 3879
rect 290 3755 738 3823
rect 290 3699 300 3755
rect 356 3699 424 3755
rect 480 3699 548 3755
rect 604 3699 672 3755
rect 728 3699 738 3755
rect 290 3631 738 3699
rect 290 3575 300 3631
rect 356 3575 424 3631
rect 480 3575 548 3631
rect 604 3575 672 3631
rect 728 3575 738 3631
rect 290 3507 738 3575
rect 290 3451 300 3507
rect 356 3451 424 3507
rect 480 3451 548 3507
rect 604 3451 672 3507
rect 728 3451 738 3507
rect 290 3383 738 3451
rect 290 3327 300 3383
rect 356 3327 424 3383
rect 480 3327 548 3383
rect 604 3327 672 3383
rect 728 3327 738 3383
rect 290 3259 738 3327
rect 290 3203 300 3259
rect 356 3203 424 3259
rect 480 3203 548 3259
rect 604 3203 672 3259
rect 728 3203 738 3259
rect 290 3135 738 3203
rect 290 3079 300 3135
rect 356 3079 424 3135
rect 480 3079 548 3135
rect 604 3079 672 3135
rect 728 3079 738 3135
rect 290 3011 738 3079
rect 290 2955 300 3011
rect 356 2955 424 3011
rect 480 2955 548 3011
rect 604 2955 672 3011
rect 728 2955 738 3011
rect 290 2887 738 2955
rect 290 2831 300 2887
rect 356 2831 424 2887
rect 480 2831 548 2887
rect 604 2831 672 2887
rect 728 2831 738 2887
rect 290 2763 738 2831
rect 290 2707 300 2763
rect 356 2707 424 2763
rect 480 2707 548 2763
rect 604 2707 672 2763
rect 728 2707 738 2763
rect 290 2639 738 2707
rect 290 2583 300 2639
rect 356 2583 424 2639
rect 480 2583 548 2639
rect 604 2583 672 2639
rect 728 2583 738 2639
rect 290 2515 738 2583
rect 290 2459 300 2515
rect 356 2459 424 2515
rect 480 2459 548 2515
rect 604 2459 672 2515
rect 728 2459 738 2515
rect 290 2391 738 2459
rect 290 2335 300 2391
rect 356 2335 424 2391
rect 480 2335 548 2391
rect 604 2335 672 2391
rect 728 2335 738 2391
rect 290 2267 738 2335
rect 290 2211 300 2267
rect 356 2211 424 2267
rect 480 2211 548 2267
rect 604 2211 672 2267
rect 728 2211 738 2267
rect 290 2143 738 2211
rect 290 2087 300 2143
rect 356 2087 424 2143
rect 480 2087 548 2143
rect 604 2087 672 2143
rect 728 2087 738 2143
rect 290 2019 738 2087
rect 290 1963 300 2019
rect 356 1963 424 2019
rect 480 1963 548 2019
rect 604 1963 672 2019
rect 728 1963 738 2019
rect 290 1895 738 1963
rect 290 1839 300 1895
rect 356 1839 424 1895
rect 480 1839 548 1895
rect 604 1839 672 1895
rect 728 1839 738 1895
rect 290 1771 738 1839
rect 290 1715 300 1771
rect 356 1715 424 1771
rect 480 1715 548 1771
rect 604 1715 672 1771
rect 728 1715 738 1771
rect 290 1647 738 1715
rect 290 1591 300 1647
rect 356 1591 424 1647
rect 480 1591 548 1647
rect 604 1591 672 1647
rect 728 1591 738 1647
rect 290 1523 738 1591
rect 290 1467 300 1523
rect 356 1467 424 1523
rect 480 1467 548 1523
rect 604 1467 672 1523
rect 728 1467 738 1523
rect 290 1399 738 1467
rect 290 1343 300 1399
rect 356 1343 424 1399
rect 480 1343 548 1399
rect 604 1343 672 1399
rect 728 1343 738 1399
rect 290 1333 738 1343
rect 1426 4251 1874 4261
rect 1426 4195 1436 4251
rect 1492 4195 1560 4251
rect 1616 4195 1684 4251
rect 1740 4195 1808 4251
rect 1864 4195 1874 4251
rect 1426 4127 1874 4195
rect 1426 4071 1436 4127
rect 1492 4071 1560 4127
rect 1616 4071 1684 4127
rect 1740 4071 1808 4127
rect 1864 4071 1874 4127
rect 1426 4003 1874 4071
rect 1426 3947 1436 4003
rect 1492 3947 1560 4003
rect 1616 3947 1684 4003
rect 1740 3947 1808 4003
rect 1864 3947 1874 4003
rect 1426 3879 1874 3947
rect 1426 3823 1436 3879
rect 1492 3823 1560 3879
rect 1616 3823 1684 3879
rect 1740 3823 1808 3879
rect 1864 3823 1874 3879
rect 1426 3755 1874 3823
rect 1426 3699 1436 3755
rect 1492 3699 1560 3755
rect 1616 3699 1684 3755
rect 1740 3699 1808 3755
rect 1864 3699 1874 3755
rect 1426 3631 1874 3699
rect 1426 3575 1436 3631
rect 1492 3575 1560 3631
rect 1616 3575 1684 3631
rect 1740 3575 1808 3631
rect 1864 3575 1874 3631
rect 1426 3507 1874 3575
rect 1426 3451 1436 3507
rect 1492 3451 1560 3507
rect 1616 3451 1684 3507
rect 1740 3451 1808 3507
rect 1864 3451 1874 3507
rect 1426 3383 1874 3451
rect 1426 3327 1436 3383
rect 1492 3327 1560 3383
rect 1616 3327 1684 3383
rect 1740 3327 1808 3383
rect 1864 3327 1874 3383
rect 1426 3259 1874 3327
rect 1426 3203 1436 3259
rect 1492 3203 1560 3259
rect 1616 3203 1684 3259
rect 1740 3203 1808 3259
rect 1864 3203 1874 3259
rect 1426 3135 1874 3203
rect 1426 3079 1436 3135
rect 1492 3079 1560 3135
rect 1616 3079 1684 3135
rect 1740 3079 1808 3135
rect 1864 3079 1874 3135
rect 1426 3011 1874 3079
rect 1426 2955 1436 3011
rect 1492 2955 1560 3011
rect 1616 2955 1684 3011
rect 1740 2955 1808 3011
rect 1864 2955 1874 3011
rect 1426 2887 1874 2955
rect 1426 2831 1436 2887
rect 1492 2831 1560 2887
rect 1616 2831 1684 2887
rect 1740 2831 1808 2887
rect 1864 2831 1874 2887
rect 1426 2763 1874 2831
rect 1426 2707 1436 2763
rect 1492 2707 1560 2763
rect 1616 2707 1684 2763
rect 1740 2707 1808 2763
rect 1864 2707 1874 2763
rect 1426 2639 1874 2707
rect 1426 2583 1436 2639
rect 1492 2583 1560 2639
rect 1616 2583 1684 2639
rect 1740 2583 1808 2639
rect 1864 2583 1874 2639
rect 1426 2515 1874 2583
rect 1426 2459 1436 2515
rect 1492 2459 1560 2515
rect 1616 2459 1684 2515
rect 1740 2459 1808 2515
rect 1864 2459 1874 2515
rect 1426 2391 1874 2459
rect 1426 2335 1436 2391
rect 1492 2335 1560 2391
rect 1616 2335 1684 2391
rect 1740 2335 1808 2391
rect 1864 2335 1874 2391
rect 1426 2267 1874 2335
rect 1426 2211 1436 2267
rect 1492 2211 1560 2267
rect 1616 2211 1684 2267
rect 1740 2211 1808 2267
rect 1864 2211 1874 2267
rect 1426 2143 1874 2211
rect 1426 2087 1436 2143
rect 1492 2087 1560 2143
rect 1616 2087 1684 2143
rect 1740 2087 1808 2143
rect 1864 2087 1874 2143
rect 1426 2019 1874 2087
rect 1426 1963 1436 2019
rect 1492 1963 1560 2019
rect 1616 1963 1684 2019
rect 1740 1963 1808 2019
rect 1864 1963 1874 2019
rect 1426 1895 1874 1963
rect 1426 1839 1436 1895
rect 1492 1839 1560 1895
rect 1616 1839 1684 1895
rect 1740 1839 1808 1895
rect 1864 1839 1874 1895
rect 1426 1771 1874 1839
rect 1426 1715 1436 1771
rect 1492 1715 1560 1771
rect 1616 1715 1684 1771
rect 1740 1715 1808 1771
rect 1864 1715 1874 1771
rect 1426 1647 1874 1715
rect 1426 1591 1436 1647
rect 1492 1591 1560 1647
rect 1616 1591 1684 1647
rect 1740 1591 1808 1647
rect 1864 1591 1874 1647
rect 1426 1523 1874 1591
rect 1426 1467 1436 1523
rect 1492 1467 1560 1523
rect 1616 1467 1684 1523
rect 1740 1467 1808 1523
rect 1864 1467 1874 1523
rect 1426 1399 1874 1467
rect 1426 1343 1436 1399
rect 1492 1343 1560 1399
rect 1616 1343 1684 1399
rect 1740 1343 1808 1399
rect 1864 1343 1874 1399
rect 1426 1333 1874 1343
rect 2562 4251 3010 4261
rect 2562 4195 2572 4251
rect 2628 4195 2696 4251
rect 2752 4195 2820 4251
rect 2876 4195 2944 4251
rect 3000 4195 3010 4251
rect 2562 4127 3010 4195
rect 2562 4071 2572 4127
rect 2628 4071 2696 4127
rect 2752 4071 2820 4127
rect 2876 4071 2944 4127
rect 3000 4071 3010 4127
rect 2562 4003 3010 4071
rect 2562 3947 2572 4003
rect 2628 3947 2696 4003
rect 2752 3947 2820 4003
rect 2876 3947 2944 4003
rect 3000 3947 3010 4003
rect 2562 3879 3010 3947
rect 2562 3823 2572 3879
rect 2628 3823 2696 3879
rect 2752 3823 2820 3879
rect 2876 3823 2944 3879
rect 3000 3823 3010 3879
rect 2562 3755 3010 3823
rect 2562 3699 2572 3755
rect 2628 3699 2696 3755
rect 2752 3699 2820 3755
rect 2876 3699 2944 3755
rect 3000 3699 3010 3755
rect 2562 3631 3010 3699
rect 2562 3575 2572 3631
rect 2628 3575 2696 3631
rect 2752 3575 2820 3631
rect 2876 3575 2944 3631
rect 3000 3575 3010 3631
rect 2562 3507 3010 3575
rect 2562 3451 2572 3507
rect 2628 3451 2696 3507
rect 2752 3451 2820 3507
rect 2876 3451 2944 3507
rect 3000 3451 3010 3507
rect 2562 3383 3010 3451
rect 2562 3327 2572 3383
rect 2628 3327 2696 3383
rect 2752 3327 2820 3383
rect 2876 3327 2944 3383
rect 3000 3327 3010 3383
rect 2562 3259 3010 3327
rect 2562 3203 2572 3259
rect 2628 3203 2696 3259
rect 2752 3203 2820 3259
rect 2876 3203 2944 3259
rect 3000 3203 3010 3259
rect 2562 3135 3010 3203
rect 2562 3079 2572 3135
rect 2628 3079 2696 3135
rect 2752 3079 2820 3135
rect 2876 3079 2944 3135
rect 3000 3079 3010 3135
rect 2562 3011 3010 3079
rect 2562 2955 2572 3011
rect 2628 2955 2696 3011
rect 2752 2955 2820 3011
rect 2876 2955 2944 3011
rect 3000 2955 3010 3011
rect 2562 2887 3010 2955
rect 2562 2831 2572 2887
rect 2628 2831 2696 2887
rect 2752 2831 2820 2887
rect 2876 2831 2944 2887
rect 3000 2831 3010 2887
rect 2562 2763 3010 2831
rect 2562 2707 2572 2763
rect 2628 2707 2696 2763
rect 2752 2707 2820 2763
rect 2876 2707 2944 2763
rect 3000 2707 3010 2763
rect 2562 2639 3010 2707
rect 2562 2583 2572 2639
rect 2628 2583 2696 2639
rect 2752 2583 2820 2639
rect 2876 2583 2944 2639
rect 3000 2583 3010 2639
rect 2562 2515 3010 2583
rect 2562 2459 2572 2515
rect 2628 2459 2696 2515
rect 2752 2459 2820 2515
rect 2876 2459 2944 2515
rect 3000 2459 3010 2515
rect 2562 2391 3010 2459
rect 2562 2335 2572 2391
rect 2628 2335 2696 2391
rect 2752 2335 2820 2391
rect 2876 2335 2944 2391
rect 3000 2335 3010 2391
rect 2562 2267 3010 2335
rect 2562 2211 2572 2267
rect 2628 2211 2696 2267
rect 2752 2211 2820 2267
rect 2876 2211 2944 2267
rect 3000 2211 3010 2267
rect 2562 2143 3010 2211
rect 2562 2087 2572 2143
rect 2628 2087 2696 2143
rect 2752 2087 2820 2143
rect 2876 2087 2944 2143
rect 3000 2087 3010 2143
rect 2562 2019 3010 2087
rect 2562 1963 2572 2019
rect 2628 1963 2696 2019
rect 2752 1963 2820 2019
rect 2876 1963 2944 2019
rect 3000 1963 3010 2019
rect 2562 1895 3010 1963
rect 2562 1839 2572 1895
rect 2628 1839 2696 1895
rect 2752 1839 2820 1895
rect 2876 1839 2944 1895
rect 3000 1839 3010 1895
rect 2562 1771 3010 1839
rect 2562 1715 2572 1771
rect 2628 1715 2696 1771
rect 2752 1715 2820 1771
rect 2876 1715 2944 1771
rect 3000 1715 3010 1771
rect 2562 1647 3010 1715
rect 2562 1591 2572 1647
rect 2628 1591 2696 1647
rect 2752 1591 2820 1647
rect 2876 1591 2944 1647
rect 3000 1591 3010 1647
rect 2562 1523 3010 1591
rect 2562 1467 2572 1523
rect 2628 1467 2696 1523
rect 2752 1467 2820 1523
rect 2876 1467 2944 1523
rect 3000 1467 3010 1523
rect 2562 1399 3010 1467
rect 2562 1343 2572 1399
rect 2628 1343 2696 1399
rect 2752 1343 2820 1399
rect 2876 1343 2944 1399
rect 3000 1343 3010 1399
rect 2562 1333 3010 1343
rect 4834 4251 5282 4261
rect 4834 4195 4844 4251
rect 4900 4195 4968 4251
rect 5024 4195 5092 4251
rect 5148 4195 5216 4251
rect 5272 4195 5282 4251
rect 4834 4127 5282 4195
rect 4834 4071 4844 4127
rect 4900 4071 4968 4127
rect 5024 4071 5092 4127
rect 5148 4071 5216 4127
rect 5272 4071 5282 4127
rect 4834 4003 5282 4071
rect 4834 3947 4844 4003
rect 4900 3947 4968 4003
rect 5024 3947 5092 4003
rect 5148 3947 5216 4003
rect 5272 3947 5282 4003
rect 4834 3879 5282 3947
rect 4834 3823 4844 3879
rect 4900 3823 4968 3879
rect 5024 3823 5092 3879
rect 5148 3823 5216 3879
rect 5272 3823 5282 3879
rect 4834 3755 5282 3823
rect 4834 3699 4844 3755
rect 4900 3699 4968 3755
rect 5024 3699 5092 3755
rect 5148 3699 5216 3755
rect 5272 3699 5282 3755
rect 4834 3631 5282 3699
rect 4834 3575 4844 3631
rect 4900 3575 4968 3631
rect 5024 3575 5092 3631
rect 5148 3575 5216 3631
rect 5272 3575 5282 3631
rect 4834 3507 5282 3575
rect 4834 3451 4844 3507
rect 4900 3451 4968 3507
rect 5024 3451 5092 3507
rect 5148 3451 5216 3507
rect 5272 3451 5282 3507
rect 4834 3383 5282 3451
rect 4834 3327 4844 3383
rect 4900 3327 4968 3383
rect 5024 3327 5092 3383
rect 5148 3327 5216 3383
rect 5272 3327 5282 3383
rect 4834 3259 5282 3327
rect 4834 3203 4844 3259
rect 4900 3203 4968 3259
rect 5024 3203 5092 3259
rect 5148 3203 5216 3259
rect 5272 3203 5282 3259
rect 4834 3135 5282 3203
rect 4834 3079 4844 3135
rect 4900 3079 4968 3135
rect 5024 3079 5092 3135
rect 5148 3079 5216 3135
rect 5272 3079 5282 3135
rect 4834 3011 5282 3079
rect 4834 2955 4844 3011
rect 4900 2955 4968 3011
rect 5024 2955 5092 3011
rect 5148 2955 5216 3011
rect 5272 2955 5282 3011
rect 4834 2887 5282 2955
rect 4834 2831 4844 2887
rect 4900 2831 4968 2887
rect 5024 2831 5092 2887
rect 5148 2831 5216 2887
rect 5272 2831 5282 2887
rect 4834 2763 5282 2831
rect 4834 2707 4844 2763
rect 4900 2707 4968 2763
rect 5024 2707 5092 2763
rect 5148 2707 5216 2763
rect 5272 2707 5282 2763
rect 4834 2639 5282 2707
rect 4834 2583 4844 2639
rect 4900 2583 4968 2639
rect 5024 2583 5092 2639
rect 5148 2583 5216 2639
rect 5272 2583 5282 2639
rect 4834 2515 5282 2583
rect 4834 2459 4844 2515
rect 4900 2459 4968 2515
rect 5024 2459 5092 2515
rect 5148 2459 5216 2515
rect 5272 2459 5282 2515
rect 4834 2391 5282 2459
rect 4834 2335 4844 2391
rect 4900 2335 4968 2391
rect 5024 2335 5092 2391
rect 5148 2335 5216 2391
rect 5272 2335 5282 2391
rect 4834 2267 5282 2335
rect 4834 2211 4844 2267
rect 4900 2211 4968 2267
rect 5024 2211 5092 2267
rect 5148 2211 5216 2267
rect 5272 2211 5282 2267
rect 4834 2143 5282 2211
rect 4834 2087 4844 2143
rect 4900 2087 4968 2143
rect 5024 2087 5092 2143
rect 5148 2087 5216 2143
rect 5272 2087 5282 2143
rect 4834 2019 5282 2087
rect 4834 1963 4844 2019
rect 4900 1963 4968 2019
rect 5024 1963 5092 2019
rect 5148 1963 5216 2019
rect 5272 1963 5282 2019
rect 4834 1895 5282 1963
rect 4834 1839 4844 1895
rect 4900 1839 4968 1895
rect 5024 1839 5092 1895
rect 5148 1839 5216 1895
rect 5272 1839 5282 1895
rect 4834 1771 5282 1839
rect 4834 1715 4844 1771
rect 4900 1715 4968 1771
rect 5024 1715 5092 1771
rect 5148 1715 5216 1771
rect 5272 1715 5282 1771
rect 4834 1647 5282 1715
rect 4834 1591 4844 1647
rect 4900 1591 4968 1647
rect 5024 1591 5092 1647
rect 5148 1591 5216 1647
rect 5272 1591 5282 1647
rect 4834 1523 5282 1591
rect 4834 1467 4844 1523
rect 4900 1467 4968 1523
rect 5024 1467 5092 1523
rect 5148 1467 5216 1523
rect 5272 1467 5282 1523
rect 4834 1399 5282 1467
rect 4834 1343 4844 1399
rect 4900 1343 4968 1399
rect 5024 1343 5092 1399
rect 5148 1343 5216 1399
rect 5272 1343 5282 1399
rect 4834 1333 5282 1343
rect 7127 4251 7451 4261
rect 7127 4195 7137 4251
rect 7193 4195 7261 4251
rect 7317 4195 7385 4251
rect 7441 4195 7451 4251
rect 7127 4127 7451 4195
rect 7127 4071 7137 4127
rect 7193 4071 7261 4127
rect 7317 4071 7385 4127
rect 7441 4071 7451 4127
rect 7127 4003 7451 4071
rect 7127 3947 7137 4003
rect 7193 3947 7261 4003
rect 7317 3947 7385 4003
rect 7441 3947 7451 4003
rect 7127 3879 7451 3947
rect 7127 3823 7137 3879
rect 7193 3823 7261 3879
rect 7317 3823 7385 3879
rect 7441 3823 7451 3879
rect 7127 3755 7451 3823
rect 7127 3699 7137 3755
rect 7193 3699 7261 3755
rect 7317 3699 7385 3755
rect 7441 3699 7451 3755
rect 7127 3631 7451 3699
rect 7127 3575 7137 3631
rect 7193 3575 7261 3631
rect 7317 3575 7385 3631
rect 7441 3575 7451 3631
rect 7127 3507 7451 3575
rect 7127 3451 7137 3507
rect 7193 3451 7261 3507
rect 7317 3451 7385 3507
rect 7441 3451 7451 3507
rect 7127 3383 7451 3451
rect 7127 3327 7137 3383
rect 7193 3327 7261 3383
rect 7317 3327 7385 3383
rect 7441 3327 7451 3383
rect 7127 3259 7451 3327
rect 7127 3203 7137 3259
rect 7193 3203 7261 3259
rect 7317 3203 7385 3259
rect 7441 3203 7451 3259
rect 7127 3135 7451 3203
rect 7127 3079 7137 3135
rect 7193 3079 7261 3135
rect 7317 3079 7385 3135
rect 7441 3079 7451 3135
rect 7127 3011 7451 3079
rect 7127 2955 7137 3011
rect 7193 2955 7261 3011
rect 7317 2955 7385 3011
rect 7441 2955 7451 3011
rect 7127 2887 7451 2955
rect 7127 2831 7137 2887
rect 7193 2831 7261 2887
rect 7317 2831 7385 2887
rect 7441 2831 7451 2887
rect 7127 2763 7451 2831
rect 7127 2707 7137 2763
rect 7193 2707 7261 2763
rect 7317 2707 7385 2763
rect 7441 2707 7451 2763
rect 7127 2639 7451 2707
rect 7127 2583 7137 2639
rect 7193 2583 7261 2639
rect 7317 2583 7385 2639
rect 7441 2583 7451 2639
rect 7127 2515 7451 2583
rect 7127 2459 7137 2515
rect 7193 2459 7261 2515
rect 7317 2459 7385 2515
rect 7441 2459 7451 2515
rect 7127 2391 7451 2459
rect 7127 2335 7137 2391
rect 7193 2335 7261 2391
rect 7317 2335 7385 2391
rect 7441 2335 7451 2391
rect 7127 2267 7451 2335
rect 7127 2211 7137 2267
rect 7193 2211 7261 2267
rect 7317 2211 7385 2267
rect 7441 2211 7451 2267
rect 7127 2143 7451 2211
rect 7127 2087 7137 2143
rect 7193 2087 7261 2143
rect 7317 2087 7385 2143
rect 7441 2087 7451 2143
rect 7127 2019 7451 2087
rect 7127 1963 7137 2019
rect 7193 1963 7261 2019
rect 7317 1963 7385 2019
rect 7441 1963 7451 2019
rect 7127 1895 7451 1963
rect 7127 1839 7137 1895
rect 7193 1839 7261 1895
rect 7317 1839 7385 1895
rect 7441 1839 7451 1895
rect 7127 1771 7451 1839
rect 7127 1715 7137 1771
rect 7193 1715 7261 1771
rect 7317 1715 7385 1771
rect 7441 1715 7451 1771
rect 7127 1647 7451 1715
rect 7127 1591 7137 1647
rect 7193 1591 7261 1647
rect 7317 1591 7385 1647
rect 7441 1591 7451 1647
rect 7127 1523 7451 1591
rect 7127 1467 7137 1523
rect 7193 1467 7261 1523
rect 7317 1467 7385 1523
rect 7441 1467 7451 1523
rect 7127 1399 7451 1467
rect 7127 1343 7137 1399
rect 7193 1343 7261 1399
rect 7317 1343 7385 1399
rect 7441 1343 7451 1399
rect 7127 1333 7451 1343
rect 7613 4251 7937 4261
rect 7613 4195 7623 4251
rect 7679 4195 7747 4251
rect 7803 4195 7871 4251
rect 7927 4195 7937 4251
rect 7613 4127 7937 4195
rect 7613 4071 7623 4127
rect 7679 4071 7747 4127
rect 7803 4071 7871 4127
rect 7927 4071 7937 4127
rect 7613 4003 7937 4071
rect 7613 3947 7623 4003
rect 7679 3947 7747 4003
rect 7803 3947 7871 4003
rect 7927 3947 7937 4003
rect 7613 3879 7937 3947
rect 7613 3823 7623 3879
rect 7679 3823 7747 3879
rect 7803 3823 7871 3879
rect 7927 3823 7937 3879
rect 7613 3755 7937 3823
rect 7613 3699 7623 3755
rect 7679 3699 7747 3755
rect 7803 3699 7871 3755
rect 7927 3699 7937 3755
rect 7613 3631 7937 3699
rect 7613 3575 7623 3631
rect 7679 3575 7747 3631
rect 7803 3575 7871 3631
rect 7927 3575 7937 3631
rect 7613 3507 7937 3575
rect 7613 3451 7623 3507
rect 7679 3451 7747 3507
rect 7803 3451 7871 3507
rect 7927 3451 7937 3507
rect 7613 3383 7937 3451
rect 7613 3327 7623 3383
rect 7679 3327 7747 3383
rect 7803 3327 7871 3383
rect 7927 3327 7937 3383
rect 7613 3259 7937 3327
rect 7613 3203 7623 3259
rect 7679 3203 7747 3259
rect 7803 3203 7871 3259
rect 7927 3203 7937 3259
rect 7613 3135 7937 3203
rect 7613 3079 7623 3135
rect 7679 3079 7747 3135
rect 7803 3079 7871 3135
rect 7927 3079 7937 3135
rect 7613 3011 7937 3079
rect 7613 2955 7623 3011
rect 7679 2955 7747 3011
rect 7803 2955 7871 3011
rect 7927 2955 7937 3011
rect 7613 2887 7937 2955
rect 7613 2831 7623 2887
rect 7679 2831 7747 2887
rect 7803 2831 7871 2887
rect 7927 2831 7937 2887
rect 7613 2763 7937 2831
rect 7613 2707 7623 2763
rect 7679 2707 7747 2763
rect 7803 2707 7871 2763
rect 7927 2707 7937 2763
rect 7613 2639 7937 2707
rect 7613 2583 7623 2639
rect 7679 2583 7747 2639
rect 7803 2583 7871 2639
rect 7927 2583 7937 2639
rect 7613 2515 7937 2583
rect 7613 2459 7623 2515
rect 7679 2459 7747 2515
rect 7803 2459 7871 2515
rect 7927 2459 7937 2515
rect 7613 2391 7937 2459
rect 7613 2335 7623 2391
rect 7679 2335 7747 2391
rect 7803 2335 7871 2391
rect 7927 2335 7937 2391
rect 7613 2267 7937 2335
rect 7613 2211 7623 2267
rect 7679 2211 7747 2267
rect 7803 2211 7871 2267
rect 7927 2211 7937 2267
rect 7613 2143 7937 2211
rect 7613 2087 7623 2143
rect 7679 2087 7747 2143
rect 7803 2087 7871 2143
rect 7927 2087 7937 2143
rect 7613 2019 7937 2087
rect 7613 1963 7623 2019
rect 7679 1963 7747 2019
rect 7803 1963 7871 2019
rect 7927 1963 7937 2019
rect 7613 1895 7937 1963
rect 7613 1839 7623 1895
rect 7679 1839 7747 1895
rect 7803 1839 7871 1895
rect 7927 1839 7937 1895
rect 7613 1771 7937 1839
rect 7613 1715 7623 1771
rect 7679 1715 7747 1771
rect 7803 1715 7871 1771
rect 7927 1715 7937 1771
rect 7613 1647 7937 1715
rect 7613 1591 7623 1647
rect 7679 1591 7747 1647
rect 7803 1591 7871 1647
rect 7927 1591 7937 1647
rect 7613 1523 7937 1591
rect 7613 1467 7623 1523
rect 7679 1467 7747 1523
rect 7803 1467 7871 1523
rect 7927 1467 7937 1523
rect 7613 1399 7937 1467
rect 7613 1343 7623 1399
rect 7679 1343 7747 1399
rect 7803 1343 7871 1399
rect 7927 1343 7937 1399
rect 7613 1333 7937 1343
rect 9782 4251 10230 4261
rect 9782 4195 9792 4251
rect 9848 4195 9916 4251
rect 9972 4195 10040 4251
rect 10096 4195 10164 4251
rect 10220 4195 10230 4251
rect 9782 4127 10230 4195
rect 9782 4071 9792 4127
rect 9848 4071 9916 4127
rect 9972 4071 10040 4127
rect 10096 4071 10164 4127
rect 10220 4071 10230 4127
rect 9782 4003 10230 4071
rect 9782 3947 9792 4003
rect 9848 3947 9916 4003
rect 9972 3947 10040 4003
rect 10096 3947 10164 4003
rect 10220 3947 10230 4003
rect 9782 3879 10230 3947
rect 9782 3823 9792 3879
rect 9848 3823 9916 3879
rect 9972 3823 10040 3879
rect 10096 3823 10164 3879
rect 10220 3823 10230 3879
rect 9782 3755 10230 3823
rect 9782 3699 9792 3755
rect 9848 3699 9916 3755
rect 9972 3699 10040 3755
rect 10096 3699 10164 3755
rect 10220 3699 10230 3755
rect 9782 3631 10230 3699
rect 9782 3575 9792 3631
rect 9848 3575 9916 3631
rect 9972 3575 10040 3631
rect 10096 3575 10164 3631
rect 10220 3575 10230 3631
rect 9782 3507 10230 3575
rect 9782 3451 9792 3507
rect 9848 3451 9916 3507
rect 9972 3451 10040 3507
rect 10096 3451 10164 3507
rect 10220 3451 10230 3507
rect 9782 3383 10230 3451
rect 9782 3327 9792 3383
rect 9848 3327 9916 3383
rect 9972 3327 10040 3383
rect 10096 3327 10164 3383
rect 10220 3327 10230 3383
rect 9782 3259 10230 3327
rect 9782 3203 9792 3259
rect 9848 3203 9916 3259
rect 9972 3203 10040 3259
rect 10096 3203 10164 3259
rect 10220 3203 10230 3259
rect 9782 3135 10230 3203
rect 9782 3079 9792 3135
rect 9848 3079 9916 3135
rect 9972 3079 10040 3135
rect 10096 3079 10164 3135
rect 10220 3079 10230 3135
rect 9782 3011 10230 3079
rect 9782 2955 9792 3011
rect 9848 2955 9916 3011
rect 9972 2955 10040 3011
rect 10096 2955 10164 3011
rect 10220 2955 10230 3011
rect 9782 2887 10230 2955
rect 9782 2831 9792 2887
rect 9848 2831 9916 2887
rect 9972 2831 10040 2887
rect 10096 2831 10164 2887
rect 10220 2831 10230 2887
rect 9782 2763 10230 2831
rect 9782 2707 9792 2763
rect 9848 2707 9916 2763
rect 9972 2707 10040 2763
rect 10096 2707 10164 2763
rect 10220 2707 10230 2763
rect 9782 2639 10230 2707
rect 9782 2583 9792 2639
rect 9848 2583 9916 2639
rect 9972 2583 10040 2639
rect 10096 2583 10164 2639
rect 10220 2583 10230 2639
rect 9782 2515 10230 2583
rect 9782 2459 9792 2515
rect 9848 2459 9916 2515
rect 9972 2459 10040 2515
rect 10096 2459 10164 2515
rect 10220 2459 10230 2515
rect 9782 2391 10230 2459
rect 9782 2335 9792 2391
rect 9848 2335 9916 2391
rect 9972 2335 10040 2391
rect 10096 2335 10164 2391
rect 10220 2335 10230 2391
rect 9782 2267 10230 2335
rect 9782 2211 9792 2267
rect 9848 2211 9916 2267
rect 9972 2211 10040 2267
rect 10096 2211 10164 2267
rect 10220 2211 10230 2267
rect 9782 2143 10230 2211
rect 9782 2087 9792 2143
rect 9848 2087 9916 2143
rect 9972 2087 10040 2143
rect 10096 2087 10164 2143
rect 10220 2087 10230 2143
rect 9782 2019 10230 2087
rect 9782 1963 9792 2019
rect 9848 1963 9916 2019
rect 9972 1963 10040 2019
rect 10096 1963 10164 2019
rect 10220 1963 10230 2019
rect 9782 1895 10230 1963
rect 9782 1839 9792 1895
rect 9848 1839 9916 1895
rect 9972 1839 10040 1895
rect 10096 1839 10164 1895
rect 10220 1839 10230 1895
rect 9782 1771 10230 1839
rect 9782 1715 9792 1771
rect 9848 1715 9916 1771
rect 9972 1715 10040 1771
rect 10096 1715 10164 1771
rect 10220 1715 10230 1771
rect 9782 1647 10230 1715
rect 9782 1591 9792 1647
rect 9848 1591 9916 1647
rect 9972 1591 10040 1647
rect 10096 1591 10164 1647
rect 10220 1591 10230 1647
rect 9782 1523 10230 1591
rect 9782 1467 9792 1523
rect 9848 1467 9916 1523
rect 9972 1467 10040 1523
rect 10096 1467 10164 1523
rect 10220 1467 10230 1523
rect 9782 1399 10230 1467
rect 9782 1343 9792 1399
rect 9848 1343 9916 1399
rect 9972 1343 10040 1399
rect 10096 1343 10164 1399
rect 10220 1343 10230 1399
rect 9782 1333 10230 1343
rect 12054 4251 12502 4261
rect 12054 4195 12064 4251
rect 12120 4195 12188 4251
rect 12244 4195 12312 4251
rect 12368 4195 12436 4251
rect 12492 4195 12502 4251
rect 12054 4127 12502 4195
rect 12054 4071 12064 4127
rect 12120 4071 12188 4127
rect 12244 4071 12312 4127
rect 12368 4071 12436 4127
rect 12492 4071 12502 4127
rect 12054 4003 12502 4071
rect 12054 3947 12064 4003
rect 12120 3947 12188 4003
rect 12244 3947 12312 4003
rect 12368 3947 12436 4003
rect 12492 3947 12502 4003
rect 12054 3879 12502 3947
rect 12054 3823 12064 3879
rect 12120 3823 12188 3879
rect 12244 3823 12312 3879
rect 12368 3823 12436 3879
rect 12492 3823 12502 3879
rect 12054 3755 12502 3823
rect 12054 3699 12064 3755
rect 12120 3699 12188 3755
rect 12244 3699 12312 3755
rect 12368 3699 12436 3755
rect 12492 3699 12502 3755
rect 12054 3631 12502 3699
rect 12054 3575 12064 3631
rect 12120 3575 12188 3631
rect 12244 3575 12312 3631
rect 12368 3575 12436 3631
rect 12492 3575 12502 3631
rect 12054 3507 12502 3575
rect 12054 3451 12064 3507
rect 12120 3451 12188 3507
rect 12244 3451 12312 3507
rect 12368 3451 12436 3507
rect 12492 3451 12502 3507
rect 12054 3383 12502 3451
rect 12054 3327 12064 3383
rect 12120 3327 12188 3383
rect 12244 3327 12312 3383
rect 12368 3327 12436 3383
rect 12492 3327 12502 3383
rect 12054 3259 12502 3327
rect 12054 3203 12064 3259
rect 12120 3203 12188 3259
rect 12244 3203 12312 3259
rect 12368 3203 12436 3259
rect 12492 3203 12502 3259
rect 12054 3135 12502 3203
rect 12054 3079 12064 3135
rect 12120 3079 12188 3135
rect 12244 3079 12312 3135
rect 12368 3079 12436 3135
rect 12492 3079 12502 3135
rect 12054 3011 12502 3079
rect 12054 2955 12064 3011
rect 12120 2955 12188 3011
rect 12244 2955 12312 3011
rect 12368 2955 12436 3011
rect 12492 2955 12502 3011
rect 12054 2887 12502 2955
rect 12054 2831 12064 2887
rect 12120 2831 12188 2887
rect 12244 2831 12312 2887
rect 12368 2831 12436 2887
rect 12492 2831 12502 2887
rect 12054 2763 12502 2831
rect 12054 2707 12064 2763
rect 12120 2707 12188 2763
rect 12244 2707 12312 2763
rect 12368 2707 12436 2763
rect 12492 2707 12502 2763
rect 12054 2639 12502 2707
rect 12054 2583 12064 2639
rect 12120 2583 12188 2639
rect 12244 2583 12312 2639
rect 12368 2583 12436 2639
rect 12492 2583 12502 2639
rect 12054 2515 12502 2583
rect 12054 2459 12064 2515
rect 12120 2459 12188 2515
rect 12244 2459 12312 2515
rect 12368 2459 12436 2515
rect 12492 2459 12502 2515
rect 12054 2391 12502 2459
rect 12054 2335 12064 2391
rect 12120 2335 12188 2391
rect 12244 2335 12312 2391
rect 12368 2335 12436 2391
rect 12492 2335 12502 2391
rect 12054 2267 12502 2335
rect 12054 2211 12064 2267
rect 12120 2211 12188 2267
rect 12244 2211 12312 2267
rect 12368 2211 12436 2267
rect 12492 2211 12502 2267
rect 12054 2143 12502 2211
rect 12054 2087 12064 2143
rect 12120 2087 12188 2143
rect 12244 2087 12312 2143
rect 12368 2087 12436 2143
rect 12492 2087 12502 2143
rect 12054 2019 12502 2087
rect 12054 1963 12064 2019
rect 12120 1963 12188 2019
rect 12244 1963 12312 2019
rect 12368 1963 12436 2019
rect 12492 1963 12502 2019
rect 12054 1895 12502 1963
rect 12054 1839 12064 1895
rect 12120 1839 12188 1895
rect 12244 1839 12312 1895
rect 12368 1839 12436 1895
rect 12492 1839 12502 1895
rect 12054 1771 12502 1839
rect 12054 1715 12064 1771
rect 12120 1715 12188 1771
rect 12244 1715 12312 1771
rect 12368 1715 12436 1771
rect 12492 1715 12502 1771
rect 12054 1647 12502 1715
rect 12054 1591 12064 1647
rect 12120 1591 12188 1647
rect 12244 1591 12312 1647
rect 12368 1591 12436 1647
rect 12492 1591 12502 1647
rect 12054 1523 12502 1591
rect 12054 1467 12064 1523
rect 12120 1467 12188 1523
rect 12244 1467 12312 1523
rect 12368 1467 12436 1523
rect 12492 1467 12502 1523
rect 12054 1399 12502 1467
rect 12054 1343 12064 1399
rect 12120 1343 12188 1399
rect 12244 1343 12312 1399
rect 12368 1343 12436 1399
rect 12492 1343 12502 1399
rect 12054 1333 12502 1343
rect 13190 4251 13638 4261
rect 13190 4195 13200 4251
rect 13256 4195 13324 4251
rect 13380 4195 13448 4251
rect 13504 4195 13572 4251
rect 13628 4195 13638 4251
rect 13190 4127 13638 4195
rect 13190 4071 13200 4127
rect 13256 4071 13324 4127
rect 13380 4071 13448 4127
rect 13504 4071 13572 4127
rect 13628 4071 13638 4127
rect 13190 4003 13638 4071
rect 13190 3947 13200 4003
rect 13256 3947 13324 4003
rect 13380 3947 13448 4003
rect 13504 3947 13572 4003
rect 13628 3947 13638 4003
rect 13190 3879 13638 3947
rect 13190 3823 13200 3879
rect 13256 3823 13324 3879
rect 13380 3823 13448 3879
rect 13504 3823 13572 3879
rect 13628 3823 13638 3879
rect 13190 3755 13638 3823
rect 13190 3699 13200 3755
rect 13256 3699 13324 3755
rect 13380 3699 13448 3755
rect 13504 3699 13572 3755
rect 13628 3699 13638 3755
rect 13190 3631 13638 3699
rect 13190 3575 13200 3631
rect 13256 3575 13324 3631
rect 13380 3575 13448 3631
rect 13504 3575 13572 3631
rect 13628 3575 13638 3631
rect 13190 3507 13638 3575
rect 13190 3451 13200 3507
rect 13256 3451 13324 3507
rect 13380 3451 13448 3507
rect 13504 3451 13572 3507
rect 13628 3451 13638 3507
rect 13190 3383 13638 3451
rect 13190 3327 13200 3383
rect 13256 3327 13324 3383
rect 13380 3327 13448 3383
rect 13504 3327 13572 3383
rect 13628 3327 13638 3383
rect 13190 3259 13638 3327
rect 13190 3203 13200 3259
rect 13256 3203 13324 3259
rect 13380 3203 13448 3259
rect 13504 3203 13572 3259
rect 13628 3203 13638 3259
rect 13190 3135 13638 3203
rect 13190 3079 13200 3135
rect 13256 3079 13324 3135
rect 13380 3079 13448 3135
rect 13504 3079 13572 3135
rect 13628 3079 13638 3135
rect 13190 3011 13638 3079
rect 13190 2955 13200 3011
rect 13256 2955 13324 3011
rect 13380 2955 13448 3011
rect 13504 2955 13572 3011
rect 13628 2955 13638 3011
rect 13190 2887 13638 2955
rect 13190 2831 13200 2887
rect 13256 2831 13324 2887
rect 13380 2831 13448 2887
rect 13504 2831 13572 2887
rect 13628 2831 13638 2887
rect 13190 2763 13638 2831
rect 13190 2707 13200 2763
rect 13256 2707 13324 2763
rect 13380 2707 13448 2763
rect 13504 2707 13572 2763
rect 13628 2707 13638 2763
rect 13190 2639 13638 2707
rect 13190 2583 13200 2639
rect 13256 2583 13324 2639
rect 13380 2583 13448 2639
rect 13504 2583 13572 2639
rect 13628 2583 13638 2639
rect 13190 2515 13638 2583
rect 13190 2459 13200 2515
rect 13256 2459 13324 2515
rect 13380 2459 13448 2515
rect 13504 2459 13572 2515
rect 13628 2459 13638 2515
rect 13190 2391 13638 2459
rect 13190 2335 13200 2391
rect 13256 2335 13324 2391
rect 13380 2335 13448 2391
rect 13504 2335 13572 2391
rect 13628 2335 13638 2391
rect 13190 2267 13638 2335
rect 13190 2211 13200 2267
rect 13256 2211 13324 2267
rect 13380 2211 13448 2267
rect 13504 2211 13572 2267
rect 13628 2211 13638 2267
rect 13190 2143 13638 2211
rect 13190 2087 13200 2143
rect 13256 2087 13324 2143
rect 13380 2087 13448 2143
rect 13504 2087 13572 2143
rect 13628 2087 13638 2143
rect 13190 2019 13638 2087
rect 13190 1963 13200 2019
rect 13256 1963 13324 2019
rect 13380 1963 13448 2019
rect 13504 1963 13572 2019
rect 13628 1963 13638 2019
rect 13190 1895 13638 1963
rect 13190 1839 13200 1895
rect 13256 1839 13324 1895
rect 13380 1839 13448 1895
rect 13504 1839 13572 1895
rect 13628 1839 13638 1895
rect 13190 1771 13638 1839
rect 13190 1715 13200 1771
rect 13256 1715 13324 1771
rect 13380 1715 13448 1771
rect 13504 1715 13572 1771
rect 13628 1715 13638 1771
rect 13190 1647 13638 1715
rect 13190 1591 13200 1647
rect 13256 1591 13324 1647
rect 13380 1591 13448 1647
rect 13504 1591 13572 1647
rect 13628 1591 13638 1647
rect 13190 1523 13638 1591
rect 13190 1467 13200 1523
rect 13256 1467 13324 1523
rect 13380 1467 13448 1523
rect 13504 1467 13572 1523
rect 13628 1467 13638 1523
rect 13190 1399 13638 1467
rect 13190 1343 13200 1399
rect 13256 1343 13324 1399
rect 13380 1343 13448 1399
rect 13504 1343 13572 1399
rect 13628 1343 13638 1399
rect 13190 1333 13638 1343
rect 14326 4251 14774 4261
rect 14326 4195 14336 4251
rect 14392 4195 14460 4251
rect 14516 4195 14584 4251
rect 14640 4195 14708 4251
rect 14764 4195 14774 4251
rect 14326 4127 14774 4195
rect 14326 4071 14336 4127
rect 14392 4071 14460 4127
rect 14516 4071 14584 4127
rect 14640 4071 14708 4127
rect 14764 4071 14774 4127
rect 14326 4003 14774 4071
rect 14326 3947 14336 4003
rect 14392 3947 14460 4003
rect 14516 3947 14584 4003
rect 14640 3947 14708 4003
rect 14764 3947 14774 4003
rect 14326 3879 14774 3947
rect 14326 3823 14336 3879
rect 14392 3823 14460 3879
rect 14516 3823 14584 3879
rect 14640 3823 14708 3879
rect 14764 3823 14774 3879
rect 14326 3755 14774 3823
rect 14326 3699 14336 3755
rect 14392 3699 14460 3755
rect 14516 3699 14584 3755
rect 14640 3699 14708 3755
rect 14764 3699 14774 3755
rect 14326 3631 14774 3699
rect 14326 3575 14336 3631
rect 14392 3575 14460 3631
rect 14516 3575 14584 3631
rect 14640 3575 14708 3631
rect 14764 3575 14774 3631
rect 14326 3507 14774 3575
rect 14326 3451 14336 3507
rect 14392 3451 14460 3507
rect 14516 3451 14584 3507
rect 14640 3451 14708 3507
rect 14764 3451 14774 3507
rect 14326 3383 14774 3451
rect 14326 3327 14336 3383
rect 14392 3327 14460 3383
rect 14516 3327 14584 3383
rect 14640 3327 14708 3383
rect 14764 3327 14774 3383
rect 14326 3259 14774 3327
rect 14326 3203 14336 3259
rect 14392 3203 14460 3259
rect 14516 3203 14584 3259
rect 14640 3203 14708 3259
rect 14764 3203 14774 3259
rect 14326 3135 14774 3203
rect 14326 3079 14336 3135
rect 14392 3079 14460 3135
rect 14516 3079 14584 3135
rect 14640 3079 14708 3135
rect 14764 3079 14774 3135
rect 14326 3011 14774 3079
rect 14326 2955 14336 3011
rect 14392 2955 14460 3011
rect 14516 2955 14584 3011
rect 14640 2955 14708 3011
rect 14764 2955 14774 3011
rect 14326 2887 14774 2955
rect 14326 2831 14336 2887
rect 14392 2831 14460 2887
rect 14516 2831 14584 2887
rect 14640 2831 14708 2887
rect 14764 2831 14774 2887
rect 14326 2763 14774 2831
rect 14326 2707 14336 2763
rect 14392 2707 14460 2763
rect 14516 2707 14584 2763
rect 14640 2707 14708 2763
rect 14764 2707 14774 2763
rect 14326 2639 14774 2707
rect 14326 2583 14336 2639
rect 14392 2583 14460 2639
rect 14516 2583 14584 2639
rect 14640 2583 14708 2639
rect 14764 2583 14774 2639
rect 14326 2515 14774 2583
rect 14326 2459 14336 2515
rect 14392 2459 14460 2515
rect 14516 2459 14584 2515
rect 14640 2459 14708 2515
rect 14764 2459 14774 2515
rect 14326 2391 14774 2459
rect 14326 2335 14336 2391
rect 14392 2335 14460 2391
rect 14516 2335 14584 2391
rect 14640 2335 14708 2391
rect 14764 2335 14774 2391
rect 14326 2267 14774 2335
rect 14326 2211 14336 2267
rect 14392 2211 14460 2267
rect 14516 2211 14584 2267
rect 14640 2211 14708 2267
rect 14764 2211 14774 2267
rect 14326 2143 14774 2211
rect 14326 2087 14336 2143
rect 14392 2087 14460 2143
rect 14516 2087 14584 2143
rect 14640 2087 14708 2143
rect 14764 2087 14774 2143
rect 14326 2019 14774 2087
rect 14326 1963 14336 2019
rect 14392 1963 14460 2019
rect 14516 1963 14584 2019
rect 14640 1963 14708 2019
rect 14764 1963 14774 2019
rect 14326 1895 14774 1963
rect 14326 1839 14336 1895
rect 14392 1839 14460 1895
rect 14516 1839 14584 1895
rect 14640 1839 14708 1895
rect 14764 1839 14774 1895
rect 14326 1771 14774 1839
rect 14326 1715 14336 1771
rect 14392 1715 14460 1771
rect 14516 1715 14584 1771
rect 14640 1715 14708 1771
rect 14764 1715 14774 1771
rect 14326 1647 14774 1715
rect 14326 1591 14336 1647
rect 14392 1591 14460 1647
rect 14516 1591 14584 1647
rect 14640 1591 14708 1647
rect 14764 1591 14774 1647
rect 14326 1523 14774 1591
rect 14326 1467 14336 1523
rect 14392 1467 14460 1523
rect 14516 1467 14584 1523
rect 14640 1467 14708 1523
rect 14764 1467 14774 1523
rect 14326 1399 14774 1467
rect 14326 1343 14336 1399
rect 14392 1343 14460 1399
rect 14516 1343 14584 1399
rect 14640 1343 14708 1399
rect 14764 1343 14774 1399
rect 14326 1333 14774 1343
use comp018green_esd_hbm  comp018green_esd_hbm_0
timestamp 1759194789
transform 1 0 1401 0 1 857
box -51 -857 12313 56440
use M1_NWELL_CDNS_40661953145380  M1_NWELL_CDNS_40661953145380_0
timestamp 1759194789
transform 1 0 12386 0 1 18196
box 0 0 1 1
use M1_NWELL_CDNS_40661953145380  M1_NWELL_CDNS_40661953145380_1
timestamp 1759194789
transform 1 0 2678 0 1 18196
box 0 0 1 1
use M1_NWELL_CDNS_40661953145384  M1_NWELL_CDNS_40661953145384_0
timestamp 1759194789
transform 1 0 7532 0 1 20446
box 0 0 1 1
use M1_NWELL_CDNS_40661953145384  M1_NWELL_CDNS_40661953145384_1
timestamp 1759194789
transform 1 0 7532 0 1 15946
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_0
timestamp 1759194789
transform 1 0 7532 0 1 56722
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_1
timestamp 1759194789
transform 1 0 7532 0 1 52774
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_2
timestamp 1759194789
transform 1 0 7532 0 1 21190
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_3
timestamp 1759194789
transform 1 0 7532 0 1 29086
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_4
timestamp 1759194789
transform 1 0 7532 0 1 33034
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_5
timestamp 1759194789
transform 1 0 7532 0 1 36982
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_6
timestamp 1759194789
transform 1 0 7532 0 1 40930
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_7
timestamp 1759194789
transform 1 0 7532 0 1 44878
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_8
timestamp 1759194789
transform 1 0 7532 0 1 48826
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_9
timestamp 1759194789
transform 1 0 7532 0 1 25138
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_0
timestamp 1759194789
transform 1 0 11749 0 1 18632
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_1
timestamp 1759194789
transform 1 0 11749 0 1 17760
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_2
timestamp 1759194789
transform 1 0 11749 0 1 19504
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_3
timestamp 1759194789
transform 1 0 11749 0 1 16888
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_4
timestamp 1759194789
transform 1 0 3315 0 1 18632
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_5
timestamp 1759194789
transform 1 0 3315 0 1 17760
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_6
timestamp 1759194789
transform 1 0 3315 0 1 19504
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_7
timestamp 1759194789
transform 1 0 3315 0 1 16888
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_0
timestamp 1759194789
transform 1 0 7532 0 1 18914
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_1
timestamp 1759194789
transform 1 0 7532 0 1 17170
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_2
timestamp 1759194789
transform 1 0 7532 0 1 16598
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_3
timestamp 1759194789
transform 1 0 7532 0 1 19794
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_4
timestamp 1759194789
transform 1 0 7532 0 1 18042
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_5
timestamp 1759194789
transform 1 0 7532 0 1 17478
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_6
timestamp 1759194789
transform 1 0 7532 0 1 18350
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_7
timestamp 1759194789
transform 1 0 7532 0 1 19222
box 0 0 1 1
use M1_PSUB_CDNS_40661953145379  M1_PSUB_CDNS_40661953145379_0
timestamp 1759194789
transform 1 0 14642 0 1 38956
box 0 0 1 1
use M1_PSUB_CDNS_40661953145379  M1_PSUB_CDNS_40661953145379_1
timestamp 1759194789
transform 1 0 422 0 1 38956
box 0 0 1 1
use M1_PSUB_CDNS_40661953145381  M1_PSUB_CDNS_40661953145381_0
timestamp 1759194789
transform 1 0 11903 0 1 18196
box 0 0 1 1
use M1_PSUB_CDNS_40661953145381  M1_PSUB_CDNS_40661953145381_1
timestamp 1759194789
transform 1 0 3161 0 1 18196
box 0 0 1 1
use M1_PSUB_CDNS_40661953145382  M1_PSUB_CDNS_40661953145382_0
timestamp 1759194789
transform 1 0 7532 0 1 18196
box 0 0 1 1
use M1_PSUB_CDNS_40661953145382  M1_PSUB_CDNS_40661953145382_1
timestamp 1759194789
transform 1 0 7532 0 1 19068
box 0 0 1 1
use M1_PSUB_CDNS_40661953145382  M1_PSUB_CDNS_40661953145382_2
timestamp 1759194789
transform 1 0 7532 0 1 17324
box 0 0 1 1
use M1_PSUB_CDNS_40661953145383  M1_PSUB_CDNS_40661953145383_0
timestamp 1759194789
transform 1 0 7532 0 1 19948
box 0 0 1 1
use M1_PSUB_CDNS_40661953145383  M1_PSUB_CDNS_40661953145383_1
timestamp 1759194789
transform 1 0 7532 0 1 16444
box 0 0 1 1
use M1_PSUB_CDNS_40661953145396  M1_PSUB_CDNS_40661953145396_0
timestamp 1759194789
transform -1 0 14380 0 1 10634
box 0 0 1 1
use M1_PSUB_CDNS_40661953145396  M1_PSUB_CDNS_40661953145396_1
timestamp 1759194789
transform 1 0 684 0 1 10634
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_0
timestamp 1759194789
transform 1 0 8870 0 1 15949
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_1
timestamp 1759194789
transform 1 0 8870 0 1 20443
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_2
timestamp 1759194789
transform 1 0 11142 0 1 15949
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_3
timestamp 1759194789
transform 1 0 11142 0 1 20443
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_4
timestamp 1759194789
transform 1 0 10006 0 1 17324
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_5
timestamp 1759194789
transform 1 0 10006 0 1 19068
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_6
timestamp 1759194789
transform 1 0 13414 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_7
timestamp 1759194789
transform 1 0 12278 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_8
timestamp 1759194789
transform 1 0 10006 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_9
timestamp 1759194789
transform 1 0 10006 0 1 18196
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_10
timestamp 1759194789
transform 1 0 3922 0 1 15949
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_11
timestamp 1759194789
transform 1 0 3922 0 1 20443
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_12
timestamp 1759194789
transform 1 0 6194 0 1 15949
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_13
timestamp 1759194789
transform 1 0 6194 0 1 20443
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_14
timestamp 1759194789
transform 1 0 5058 0 1 17324
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_15
timestamp 1759194789
transform 1 0 5058 0 1 18196
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_16
timestamp 1759194789
transform 1 0 5058 0 1 19068
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_17
timestamp 1759194789
transform 1 0 5058 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_18
timestamp 1759194789
transform 1 0 2786 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_19
timestamp 1759194789
transform 1 0 1650 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_20
timestamp 1759194789
transform 1 0 2786 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_21
timestamp 1759194789
transform 1 0 1650 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_22
timestamp 1759194789
transform 1 0 5058 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_23
timestamp 1759194789
transform 1 0 10006 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_24
timestamp 1759194789
transform 1 0 13414 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_25
timestamp 1759194789
transform 1 0 12278 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_0
timestamp 1759194789
transform 1 0 84 0 1 37197
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_1
timestamp 1759194789
transform 1 0 84 0 1 51597
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_2
timestamp 1759194789
transform 1 0 14980 0 1 37197
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_3
timestamp 1759194789
transform 1 0 14980 0 1 51597
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_0
timestamp 1759194789
transform 1 0 8870 0 1 16888
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_1
timestamp 1759194789
transform 1 0 8870 0 1 17760
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_2
timestamp 1759194789
transform 1 0 8870 0 1 18632
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_3
timestamp 1759194789
transform 1 0 11142 0 1 16888
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_4
timestamp 1759194789
transform 1 0 11142 0 1 19504
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_5
timestamp 1759194789
transform 1 0 11142 0 1 17760
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_6
timestamp 1759194789
transform 1 0 11142 0 1 18632
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_7
timestamp 1759194789
transform 1 0 10006 0 1 16521
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_8
timestamp 1759194789
transform 1 0 10006 0 1 19871
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_9
timestamp 1759194789
transform 1 0 8870 0 1 19504
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_10
timestamp 1759194789
transform 1 0 6194 0 1 16888
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_11
timestamp 1759194789
transform 1 0 6194 0 1 19504
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_12
timestamp 1759194789
transform 1 0 6194 0 1 17760
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_13
timestamp 1759194789
transform 1 0 6194 0 1 18632
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_14
timestamp 1759194789
transform 1 0 5058 0 1 16521
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_15
timestamp 1759194789
transform 1 0 5058 0 1 19871
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_16
timestamp 1759194789
transform 1 0 3922 0 1 16888
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_17
timestamp 1759194789
transform 1 0 3922 0 1 17760
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_18
timestamp 1759194789
transform 1 0 3922 0 1 18632
box 0 0 1 1
use M2_M1_CDNS_40661953145141  M2_M1_CDNS_40661953145141_19
timestamp 1759194789
transform 1 0 3922 0 1 19504
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_0
timestamp 1759194789
transform -1 0 7650 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_1
timestamp 1759194789
transform -1 0 7650 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_2
timestamp 1759194789
transform 1 0 7414 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_3
timestamp 1759194789
transform 1 0 7414 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_4
timestamp 1759194789
transform 1 0 7414 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_5
timestamp 1759194789
transform 1 0 7414 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_6
timestamp 1759194789
transform 1 0 7414 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_7
timestamp 1759194789
transform 1 0 7414 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_8
timestamp 1759194789
transform 1 0 7414 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_9
timestamp 1759194789
transform 1 0 7414 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_10
timestamp 1759194789
transform 1 0 7414 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_11
timestamp 1759194789
transform -1 0 7650 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_12
timestamp 1759194789
transform -1 0 7650 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_13
timestamp 1759194789
transform -1 0 7650 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_14
timestamp 1759194789
transform -1 0 7650 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_15
timestamp 1759194789
transform -1 0 7650 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_16
timestamp 1759194789
transform -1 0 7650 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145151  M2_M1_CDNS_40661953145151_17
timestamp 1759194789
transform -1 0 7650 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_0
timestamp 1759194789
transform 1 0 7775 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_1
timestamp 1759194789
transform 1 0 7289 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_2
timestamp 1759194789
transform 1 0 7289 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_3
timestamp 1759194789
transform 1 0 7289 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_4
timestamp 1759194789
transform 1 0 7289 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_5
timestamp 1759194789
transform 1 0 7289 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_6
timestamp 1759194789
transform 1 0 7289 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_7
timestamp 1759194789
transform 1 0 7289 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_8
timestamp 1759194789
transform 1 0 7289 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_9
timestamp 1759194789
transform 1 0 7775 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_10
timestamp 1759194789
transform 1 0 7775 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_11
timestamp 1759194789
transform 1 0 7775 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_12
timestamp 1759194789
transform 1 0 7775 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_13
timestamp 1759194789
transform 1 0 7775 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_14
timestamp 1759194789
transform 1 0 7775 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145359  M2_M1_CDNS_40661953145359_15
timestamp 1759194789
transform 1 0 7775 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_0
timestamp 1759194789
transform 1 0 7775 0 1 16521
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_1
timestamp 1759194789
transform 1 0 7775 0 1 19871
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_2
timestamp 1759194789
transform 1 0 7289 0 1 16521
box 0 0 1 1
use M2_M1_CDNS_40661953145385  M2_M1_CDNS_40661953145385_3
timestamp 1759194789
transform 1 0 7289 0 1 19871
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_0
timestamp 1759194789
transform 1 0 7775 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_1
timestamp 1759194789
transform 1 0 7775 0 1 18196
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_2
timestamp 1759194789
transform 1 0 7775 0 1 17324
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_3
timestamp 1759194789
transform 1 0 7775 0 1 19068
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_4
timestamp 1759194789
transform 1 0 7289 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_5
timestamp 1759194789
transform 1 0 7289 0 1 19068
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_6
timestamp 1759194789
transform 1 0 7289 0 1 18196
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_7
timestamp 1759194789
transform 1 0 7289 0 1 17324
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_8
timestamp 1759194789
transform 1 0 7289 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_40661953145386  M2_M1_CDNS_40661953145386_9
timestamp 1759194789
transform 1 0 7775 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_40661953145389  M2_M1_CDNS_40661953145389_0
timestamp 1759194789
transform 1 0 1236 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145389  M2_M1_CDNS_40661953145389_1
timestamp 1759194789
transform 1 0 1236 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145389  M2_M1_CDNS_40661953145389_2
timestamp 1759194789
transform 1 0 1236 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145389  M2_M1_CDNS_40661953145389_3
timestamp 1759194789
transform 1 0 1236 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145390  M2_M1_CDNS_40661953145390_0
timestamp 1759194789
transform -1 0 14486 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_40661953145390  M2_M1_CDNS_40661953145390_1
timestamp 1759194789
transform 1 0 578 0 1 21335
box 0 0 1 1
use M2_M1_CDNS_40661953145390  M2_M1_CDNS_40661953145390_2
timestamp 1759194789
transform 1 0 578 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_40661953145390  M2_M1_CDNS_40661953145390_3
timestamp 1759194789
transform -1 0 14486 0 1 56577
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_0
timestamp 1759194789
transform -1 0 13936 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_1
timestamp 1759194789
transform 1 0 1128 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_2
timestamp 1759194789
transform 1 0 1128 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_3
timestamp 1759194789
transform 1 0 1128 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_4
timestamp 1759194789
transform 1 0 1128 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_5
timestamp 1759194789
transform -1 0 13936 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_6
timestamp 1759194789
transform -1 0 13936 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_7
timestamp 1759194789
transform -1 0 13936 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_8
timestamp 1759194789
transform -1 0 13936 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_9
timestamp 1759194789
transform -1 0 13936 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_10
timestamp 1759194789
transform -1 0 13936 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_11
timestamp 1759194789
transform -1 0 13936 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_12
timestamp 1759194789
transform -1 0 13936 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145391  M2_M1_CDNS_40661953145391_13
timestamp 1759194789
transform 1 0 1128 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_0
timestamp 1759194789
transform -1 0 8703 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_1
timestamp 1759194789
transform -1 0 11309 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_2
timestamp 1759194789
transform 1 0 3755 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_3
timestamp 1759194789
transform 1 0 6361 0 1 23164
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_4
timestamp 1759194789
transform 1 0 6361 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_5
timestamp 1759194789
transform 1 0 6361 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_6
timestamp 1759194789
transform 1 0 6361 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_7
timestamp 1759194789
transform 1 0 6361 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_8
timestamp 1759194789
transform 1 0 6361 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_9
timestamp 1759194789
transform 1 0 6361 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_10
timestamp 1759194789
transform 1 0 3755 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_11
timestamp 1759194789
transform 1 0 3755 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_12
timestamp 1759194789
transform 1 0 3755 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_13
timestamp 1759194789
transform 1 0 6361 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_14
timestamp 1759194789
transform 1 0 3755 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_15
timestamp 1759194789
transform 1 0 3755 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_16
timestamp 1759194789
transform 1 0 3755 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_17
timestamp 1759194789
transform 1 0 3755 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_18
timestamp 1759194789
transform -1 0 8703 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_19
timestamp 1759194789
transform -1 0 8703 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_20
timestamp 1759194789
transform -1 0 8703 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_21
timestamp 1759194789
transform -1 0 8703 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_22
timestamp 1759194789
transform -1 0 8703 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_23
timestamp 1759194789
transform -1 0 8703 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_24
timestamp 1759194789
transform -1 0 11309 0 1 35008
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_25
timestamp 1759194789
transform -1 0 11309 0 1 38956
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_26
timestamp 1759194789
transform -1 0 11309 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_27
timestamp 1759194789
transform -1 0 8703 0 1 42904
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_28
timestamp 1759194789
transform -1 0 11309 0 1 46852
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_29
timestamp 1759194789
transform -1 0 11309 0 1 50800
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_30
timestamp 1759194789
transform -1 0 11309 0 1 54748
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_31
timestamp 1759194789
transform -1 0 11309 0 1 31060
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_32
timestamp 1759194789
transform -1 0 8703 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_33
timestamp 1759194789
transform -1 0 11309 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_34
timestamp 1759194789
transform 1 0 6361 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145392  M2_M1_CDNS_40661953145392_35
timestamp 1759194789
transform 1 0 3755 0 1 27112
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_0
timestamp 1759194789
transform 1 0 13414 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_1
timestamp 1759194789
transform 1 0 12278 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_2
timestamp 1759194789
transform 1 0 10006 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_3
timestamp 1759194789
transform 1 0 5058 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_4
timestamp 1759194789
transform 1 0 2786 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_5
timestamp 1759194789
transform 1 0 1650 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_6
timestamp 1759194789
transform 1 0 5058 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_7
timestamp 1759194789
transform 1 0 5058 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_8
timestamp 1759194789
transform 1 0 5058 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_9
timestamp 1759194789
transform 1 0 5058 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_10
timestamp 1759194789
transform 1 0 1650 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_11
timestamp 1759194789
transform 1 0 2786 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_12
timestamp 1759194789
transform 1 0 1650 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_13
timestamp 1759194789
transform 1 0 2786 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_14
timestamp 1759194789
transform 1 0 1650 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_15
timestamp 1759194789
transform 1 0 2786 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_16
timestamp 1759194789
transform 1 0 1650 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_17
timestamp 1759194789
transform 1 0 2786 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_18
timestamp 1759194789
transform 1 0 2786 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_19
timestamp 1759194789
transform 1 0 1650 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_20
timestamp 1759194789
transform 1 0 1650 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_21
timestamp 1759194789
transform 1 0 2786 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_22
timestamp 1759194789
transform 1 0 1650 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_23
timestamp 1759194789
transform 1 0 2786 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_24
timestamp 1759194789
transform 1 0 5058 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_25
timestamp 1759194789
transform 1 0 5058 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_26
timestamp 1759194789
transform 1 0 5058 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_27
timestamp 1759194789
transform 1 0 13414 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_28
timestamp 1759194789
transform 1 0 12278 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_29
timestamp 1759194789
transform 1 0 13414 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_30
timestamp 1759194789
transform 1 0 12278 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_31
timestamp 1759194789
transform 1 0 12278 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_32
timestamp 1759194789
transform 1 0 12278 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_33
timestamp 1759194789
transform 1 0 10006 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_34
timestamp 1759194789
transform 1 0 10006 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_35
timestamp 1759194789
transform 1 0 10006 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_36
timestamp 1759194789
transform 1 0 10006 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_37
timestamp 1759194789
transform 1 0 10006 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_38
timestamp 1759194789
transform 1 0 10006 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_39
timestamp 1759194789
transform 1 0 10006 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_40
timestamp 1759194789
transform 1 0 12278 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_41
timestamp 1759194789
transform 1 0 12278 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_42
timestamp 1759194789
transform 1 0 12278 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145393  M2_M1_CDNS_40661953145393_43
timestamp 1759194789
transform 1 0 13414 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_0
timestamp 1759194789
transform -1 0 14486 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_1
timestamp 1759194789
transform 1 0 578 0 1 25138
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_2
timestamp 1759194789
transform 1 0 578 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_3
timestamp 1759194789
transform 1 0 578 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_4
timestamp 1759194789
transform 1 0 578 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_5
timestamp 1759194789
transform 1 0 578 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_6
timestamp 1759194789
transform 1 0 578 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_7
timestamp 1759194789
transform 1 0 578 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_8
timestamp 1759194789
transform 1 0 578 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_9
timestamp 1759194789
transform -1 0 14486 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_10
timestamp 1759194789
transform -1 0 14486 0 1 33034
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_11
timestamp 1759194789
transform -1 0 14486 0 1 29086
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_12
timestamp 1759194789
transform -1 0 14486 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_13
timestamp 1759194789
transform -1 0 14486 0 1 52774
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_14
timestamp 1759194789
transform -1 0 14486 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145394  M2_M1_CDNS_40661953145394_15
timestamp 1759194789
transform -1 0 14486 0 1 44878
box 0 0 1 1
use M2_M1_CDNS_40661953145395  M2_M1_CDNS_40661953145395_0
timestamp 1759194789
transform 1 0 13568 0 1 40930
box 0 0 1 1
use M2_M1_CDNS_40661953145395  M2_M1_CDNS_40661953145395_1
timestamp 1759194789
transform 1 0 13568 0 1 36982
box 0 0 1 1
use M2_M1_CDNS_40661953145395  M2_M1_CDNS_40661953145395_2
timestamp 1759194789
transform 1 0 13568 0 1 48826
box 0 0 1 1
use M2_M1_CDNS_40661953145395  M2_M1_CDNS_40661953145395_3
timestamp 1759194789
transform 1 0 13568 0 1 44878
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_0
timestamp 1759194789
transform 1 0 84 0 1 37197
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_1
timestamp 1759194789
transform 1 0 84 0 1 51597
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_2
timestamp 1759194789
transform 1 0 14980 0 1 37197
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_3
timestamp 1759194789
transform 1 0 14980 0 1 51597
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_0
timestamp 1759194789
transform 1 0 928 0 1 38797
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_1
timestamp 1759194789
transform 1 0 1236 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_2
timestamp 1759194789
transform 1 0 1236 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_3
timestamp 1759194789
transform 1 0 1236 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_4
timestamp 1759194789
transform 1 0 928 0 1 49997
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_5
timestamp 1759194789
transform 1 0 1236 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_6
timestamp 1759194789
transform -1 0 13260 0 1 37197
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_7
timestamp 1759194789
transform -1 0 13568 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_8
timestamp 1759194789
transform -1 0 13568 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_9
timestamp 1759194789
transform -1 0 13260 0 1 51597
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_0
timestamp 1759194789
transform 1 0 514 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_1
timestamp 1759194789
transform 1 0 1650 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_2
timestamp 1759194789
transform 1 0 2786 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_3
timestamp 1759194789
transform 1 0 5058 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_4
timestamp 1759194789
transform -1 0 10006 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_5
timestamp 1759194789
transform -1 0 12278 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_6
timestamp 1759194789
transform -1 0 14550 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_7
timestamp 1759194789
transform -1 0 13414 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_0
timestamp 1759194789
transform -1 0 13414 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_1
timestamp 1759194789
transform -1 0 12278 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_2
timestamp 1759194789
transform -1 0 10006 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_3
timestamp 1759194789
transform -1 0 14550 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_4
timestamp 1759194789
transform -1 0 13414 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_5
timestamp 1759194789
transform -1 0 12278 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_6
timestamp 1759194789
transform -1 0 10006 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_7
timestamp 1759194789
transform -1 0 14550 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_8
timestamp 1759194789
transform -1 0 13982 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_9
timestamp 1759194789
transform -1 0 12846 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_10
timestamp 1759194789
transform -1 0 11142 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_11
timestamp 1759194789
transform -1 0 8870 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_12
timestamp 1759194789
transform 1 0 514 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_13
timestamp 1759194789
transform 1 0 5058 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_14
timestamp 1759194789
transform 1 0 2786 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_15
timestamp 1759194789
transform 1 0 1650 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_16
timestamp 1759194789
transform 1 0 514 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_17
timestamp 1759194789
transform 1 0 2786 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_18
timestamp 1759194789
transform 1 0 1650 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_19
timestamp 1759194789
transform 1 0 6194 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_20
timestamp 1759194789
transform 1 0 3922 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_21
timestamp 1759194789
transform 1 0 2218 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_22
timestamp 1759194789
transform 1 0 1082 0 1 11597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_23
timestamp 1759194789
transform 1 0 5058 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_24
timestamp 1759194789
transform 1 0 6194 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_25
timestamp 1759194789
transform 1 0 6194 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_26
timestamp 1759194789
transform 1 0 2218 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_27
timestamp 1759194789
transform 1 0 2218 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_28
timestamp 1759194789
transform 1 0 514 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_29
timestamp 1759194789
transform 1 0 2218 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_30
timestamp 1759194789
transform 1 0 2218 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_31
timestamp 1759194789
transform 1 0 1082 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_32
timestamp 1759194789
transform 1 0 2786 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_33
timestamp 1759194789
transform 1 0 2786 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_34
timestamp 1759194789
transform 1 0 1650 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_35
timestamp 1759194789
transform 1 0 514 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_36
timestamp 1759194789
transform 1 0 2786 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_37
timestamp 1759194789
transform 1 0 1650 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_38
timestamp 1759194789
transform 1 0 514 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_39
timestamp 1759194789
transform 1 0 1650 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_40
timestamp 1759194789
transform 1 0 5058 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_41
timestamp 1759194789
transform 1 0 5058 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_42
timestamp 1759194789
transform 1 0 5058 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_43
timestamp 1759194789
transform 1 0 6194 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_44
timestamp 1759194789
transform 1 0 6194 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_45
timestamp 1759194789
transform 1 0 3922 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_46
timestamp 1759194789
transform 1 0 3922 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_47
timestamp 1759194789
transform 1 0 3922 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_48
timestamp 1759194789
transform 1 0 2218 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_49
timestamp 1759194789
transform 1 0 3922 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_50
timestamp 1759194789
transform 1 0 6194 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_51
timestamp 1759194789
transform 1 0 3922 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_52
timestamp 1759194789
transform -1 0 13982 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_53
timestamp 1759194789
transform -1 0 12846 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_54
timestamp 1759194789
transform -1 0 13982 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_55
timestamp 1759194789
transform -1 0 12846 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_56
timestamp 1759194789
transform -1 0 8870 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_57
timestamp 1759194789
transform -1 0 8870 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_58
timestamp 1759194789
transform -1 0 10006 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_59
timestamp 1759194789
transform -1 0 10006 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_60
timestamp 1759194789
transform -1 0 8870 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_61
timestamp 1759194789
transform -1 0 8870 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_62
timestamp 1759194789
transform -1 0 10006 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_63
timestamp 1759194789
transform -1 0 12846 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_64
timestamp 1759194789
transform -1 0 13982 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_65
timestamp 1759194789
transform -1 0 13414 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_66
timestamp 1759194789
transform -1 0 14550 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_67
timestamp 1759194789
transform -1 0 13982 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_68
timestamp 1759194789
transform -1 0 12846 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_69
timestamp 1759194789
transform -1 0 12278 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_70
timestamp 1759194789
transform -1 0 14550 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_71
timestamp 1759194789
transform -1 0 12278 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_72
timestamp 1759194789
transform -1 0 14550 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_73
timestamp 1759194789
transform -1 0 12278 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_74
timestamp 1759194789
transform -1 0 11142 0 1 46797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_75
timestamp 1759194789
transform -1 0 8870 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_76
timestamp 1759194789
transform -1 0 11142 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_77
timestamp 1759194789
transform -1 0 12846 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_78
timestamp 1759194789
transform -1 0 13982 0 1 43597
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_79
timestamp 1759194789
transform -1 0 11142 0 1 41997
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_80
timestamp 1759194789
transform -1 0 11142 0 1 54797
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_81
timestamp 1759194789
transform -1 0 11142 0 1 40397
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_82
timestamp 1759194789
transform -1 0 13982 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_83
timestamp 1759194789
transform -1 0 12846 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_84
timestamp 1759194789
transform -1 0 11142 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_85
timestamp 1759194789
transform -1 0 8870 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_86
timestamp 1759194789
transform 1 0 6194 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_87
timestamp 1759194789
transform 1 0 3922 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_88
timestamp 1759194789
transform 1 0 2218 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_89
timestamp 1759194789
transform 1 0 1082 0 1 29197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_0
timestamp 1759194789
transform -1 0 8870 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_1
timestamp 1759194789
transform -1 0 13982 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_2
timestamp 1759194789
transform -1 0 12846 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_3
timestamp 1759194789
transform -1 0 11142 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_4
timestamp 1759194789
transform -1 0 8870 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_5
timestamp 1759194789
transform -1 0 13982 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_6
timestamp 1759194789
transform -1 0 12846 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_7
timestamp 1759194789
transform -1 0 11142 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_8
timestamp 1759194789
transform -1 0 8870 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_9
timestamp 1759194789
transform -1 0 13982 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_10
timestamp 1759194789
transform -1 0 12846 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_11
timestamp 1759194789
transform -1 0 11142 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_12
timestamp 1759194789
transform -1 0 8870 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_13
timestamp 1759194789
transform -1 0 13982 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_14
timestamp 1759194789
transform -1 0 12846 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_15
timestamp 1759194789
transform -1 0 11142 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_16
timestamp 1759194789
transform -1 0 13414 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_17
timestamp 1759194789
transform -1 0 10006 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_18
timestamp 1759194789
transform -1 0 12278 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_19
timestamp 1759194789
transform -1 0 13414 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_20
timestamp 1759194789
transform -1 0 14550 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_21
timestamp 1759194789
transform -1 0 10006 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_22
timestamp 1759194789
transform -1 0 12278 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_23
timestamp 1759194789
transform -1 0 14550 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_24
timestamp 1759194789
transform -1 0 10006 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_25
timestamp 1759194789
transform -1 0 12278 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_26
timestamp 1759194789
transform -1 0 13414 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_27
timestamp 1759194789
transform -1 0 14550 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_28
timestamp 1759194789
transform 1 0 5058 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_29
timestamp 1759194789
transform 1 0 514 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_30
timestamp 1759194789
transform 1 0 1650 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_31
timestamp 1759194789
transform 1 0 2786 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_32
timestamp 1759194789
transform 1 0 5058 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_33
timestamp 1759194789
transform 1 0 1650 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_34
timestamp 1759194789
transform 1 0 2786 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_35
timestamp 1759194789
transform 1 0 514 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_36
timestamp 1759194789
transform 1 0 5058 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_37
timestamp 1759194789
transform 1 0 2786 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_38
timestamp 1759194789
transform 1 0 1650 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_39
timestamp 1759194789
transform 1 0 514 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_40
timestamp 1759194789
transform 1 0 2218 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_41
timestamp 1759194789
transform 1 0 6194 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_42
timestamp 1759194789
transform 1 0 3922 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_43
timestamp 1759194789
transform 1 0 2218 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_44
timestamp 1759194789
transform 1 0 1082 0 1 15597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_45
timestamp 1759194789
transform 1 0 6194 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_46
timestamp 1759194789
transform 1 0 3922 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_47
timestamp 1759194789
transform 1 0 2218 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_48
timestamp 1759194789
transform 1 0 1082 0 1 18797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_49
timestamp 1759194789
transform 1 0 6194 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_50
timestamp 1759194789
transform 1 0 3922 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_51
timestamp 1759194789
transform 1 0 2218 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_52
timestamp 1759194789
transform 1 0 1082 0 1 21997
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_53
timestamp 1759194789
transform 1 0 6194 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_54
timestamp 1759194789
transform 1 0 3922 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_55
timestamp 1759194789
transform 1 0 1082 0 1 25197
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_56
timestamp 1759194789
transform 1 0 5058 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_57
timestamp 1759194789
transform 1 0 6194 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_58
timestamp 1759194789
transform 1 0 514 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_59
timestamp 1759194789
transform 1 0 2786 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_60
timestamp 1759194789
transform 1 0 1650 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_61
timestamp 1759194789
transform 1 0 2218 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_62
timestamp 1759194789
transform 1 0 1082 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_63
timestamp 1759194789
transform 1 0 3922 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_64
timestamp 1759194789
transform -1 0 12278 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_65
timestamp 1759194789
transform -1 0 13414 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_66
timestamp 1759194789
transform -1 0 14550 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_67
timestamp 1759194789
transform -1 0 13982 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_68
timestamp 1759194789
transform -1 0 12846 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_69
timestamp 1759194789
transform -1 0 10006 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_70
timestamp 1759194789
transform -1 0 8870 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_71
timestamp 1759194789
transform -1 0 11142 0 1 31597
box 0 0 1 1
use M3_M2_CDNS_40661953145175  M3_M2_CDNS_40661953145175_0
timestamp 1759194789
transform 1 0 7289 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_40661953145175  M3_M2_CDNS_40661953145175_1
timestamp 1759194789
transform -1 0 7775 0 1 56336
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_0
timestamp 1759194789
transform -1 0 7775 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_1
timestamp 1759194789
transform -1 0 7775 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_2
timestamp 1759194789
transform 1 0 7289 0 1 27597
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_3
timestamp 1759194789
transform 1 0 7289 0 1 13197
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_4
timestamp 1759194789
transform 1 0 7289 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_5
timestamp 1759194789
transform 1 0 7289 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_6
timestamp 1759194789
transform 1 0 7289 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_7
timestamp 1759194789
transform -1 0 7775 0 1 48397
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_8
timestamp 1759194789
transform -1 0 7775 0 1 53197
box 0 0 1 1
use M3_M2_CDNS_40661953145387  M3_M2_CDNS_40661953145387_9
timestamp 1759194789
transform -1 0 7775 0 1 45197
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_0
timestamp 1759194789
transform -1 0 7775 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_1
timestamp 1759194789
transform -1 0 7775 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_2
timestamp 1759194789
transform -1 0 7775 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_3
timestamp 1759194789
transform 1 0 7289 0 1 9197
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_4
timestamp 1759194789
transform 1 0 7289 0 1 2797
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_5
timestamp 1759194789
transform 1 0 7289 0 1 5997
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_6
timestamp 1759194789
transform 1 0 7289 0 1 34797
box 0 0 1 1
use M3_M2_CDNS_40661953145388  M3_M2_CDNS_40661953145388_7
timestamp 1759194789
transform -1 0 7775 0 1 34797
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_0
timestamp 1759194789
transform 1 0 11186 0 1 21664
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_1
timestamp 1759194789
transform 1 0 878 0 1 21664
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_2
timestamp 1759194789
transform 1 0 878 0 1 49300
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_3
timestamp 1759194789
transform 1 0 878 0 1 45352
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_4
timestamp 1759194789
transform 1 0 878 0 1 41404
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_5
timestamp 1759194789
transform 1 0 878 0 1 37456
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_6
timestamp 1759194789
transform 1 0 878 0 1 33508
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_7
timestamp 1759194789
transform 1 0 878 0 1 29560
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_8
timestamp 1759194789
transform 1 0 878 0 1 53248
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_9
timestamp 1759194789
transform 1 0 11186 0 1 33508
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_10
timestamp 1759194789
transform 1 0 11186 0 1 29560
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_11
timestamp 1759194789
transform 1 0 11186 0 1 49300
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_12
timestamp 1759194789
transform 1 0 11186 0 1 53248
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_13
timestamp 1759194789
transform 1 0 11186 0 1 45352
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_14
timestamp 1759194789
transform 1 0 11186 0 1 41404
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_15
timestamp 1759194789
transform 1 0 11186 0 1 37456
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_16
timestamp 1759194789
transform 1 0 4314 0 1 21664
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_17
timestamp 1759194789
transform 1 0 4314 0 1 53248
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_18
timestamp 1759194789
transform 1 0 4314 0 1 29560
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_19
timestamp 1759194789
transform 1 0 4314 0 1 33508
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_20
timestamp 1759194789
transform 1 0 4314 0 1 37456
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_21
timestamp 1759194789
transform 1 0 4314 0 1 41404
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_22
timestamp 1759194789
transform 1 0 4314 0 1 49300
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_23
timestamp 1759194789
transform 1 0 4314 0 1 25612
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_24
timestamp 1759194789
transform 1 0 878 0 1 25612
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_25
timestamp 1759194789
transform 1 0 4314 0 1 45352
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_26
timestamp 1759194789
transform 1 0 11186 0 1 25612
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_27
timestamp 1759194789
transform 1 0 7750 0 1 49300
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_28
timestamp 1759194789
transform 1 0 7750 0 1 45352
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_29
timestamp 1759194789
transform 1 0 7750 0 1 41404
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_30
timestamp 1759194789
transform 1 0 7750 0 1 37456
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_31
timestamp 1759194789
transform 1 0 7750 0 1 33508
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_32
timestamp 1759194789
transform 1 0 7750 0 1 53248
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_33
timestamp 1759194789
transform 1 0 7750 0 1 25612
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_34
timestamp 1759194789
transform 1 0 7750 0 1 29560
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_35
timestamp 1759194789
transform 1 0 7750 0 1 21664
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_0
timestamp 1759194789
transform 1 0 3532 0 1 19404
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_1
timestamp 1759194789
transform 1 0 3532 0 1 17660
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_2
timestamp 1759194789
transform 1 0 3532 0 1 16788
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_3
timestamp 1759194789
transform 1 0 3532 0 1 18532
box 0 0 1 1
<< properties >>
string GDS_END 1461524
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1426402
string path 339.200 906.250 339.200 1311.500 
<< end >>
