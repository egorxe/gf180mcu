VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__dvss
  CLASS PAD POWER ;
  FOREIGN gf180mcu_fd_io__dvss ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 25.000 20.000 50.000 45.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 1.360 349.000 10.860 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 13.760 349.000 24.010 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 25.610 349.000 35.860 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 39.140 349.000 49.390 350.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 50.990 349.000 61.240 350.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal2 ;
        RECT 64.140 349.000 73.640 350.000 ;
    END
  END DVSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
  END VDD
  OBS
      LAYER Nwell ;
        RECT 3.060 67.195 71.940 345.275 ;
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 348.700 1.060 349.000 ;
        RECT 11.160 348.700 13.460 349.000 ;
        RECT 24.310 348.700 25.310 349.000 ;
        RECT 36.160 348.700 38.840 349.000 ;
        RECT 49.690 348.700 50.690 349.000 ;
        RECT 61.540 348.700 63.840 349.000 ;
        RECT 73.940 348.700 75.000 349.000 ;
        RECT 0.000 0.000 75.000 348.700 ;
      LAYER Metal3 ;
        RECT 1.300 341.700 73.700 348.390 ;
        RECT 1.000 341.300 74.000 341.700 ;
        RECT 1.300 333.700 73.700 341.300 ;
        RECT 1.000 333.300 74.000 333.700 ;
        RECT 1.300 325.700 73.700 333.300 ;
        RECT 1.000 325.300 74.000 325.700 ;
        RECT 1.300 317.700 73.700 325.300 ;
        RECT 1.000 317.300 74.000 317.700 ;
        RECT 1.300 309.700 73.700 317.300 ;
        RECT 1.000 309.300 74.000 309.700 ;
        RECT 1.300 301.700 73.700 309.300 ;
        RECT 1.000 301.300 74.000 301.700 ;
        RECT 1.300 293.700 73.700 301.300 ;
        RECT 1.000 293.300 74.000 293.700 ;
        RECT 1.300 285.700 73.700 293.300 ;
        RECT 1.000 285.300 74.000 285.700 ;
        RECT 1.300 277.700 73.700 285.300 ;
        RECT 1.000 277.300 74.000 277.700 ;
        RECT 1.300 269.700 73.700 277.300 ;
        RECT 1.000 269.300 74.000 269.700 ;
        RECT 1.300 261.700 73.700 269.300 ;
        RECT 1.000 261.300 74.000 261.700 ;
        RECT 1.300 253.700 73.700 261.300 ;
        RECT 1.000 253.300 74.000 253.700 ;
        RECT 1.300 245.700 73.700 253.300 ;
        RECT 1.000 245.300 74.000 245.700 ;
        RECT 1.300 229.700 73.700 245.300 ;
        RECT 1.000 229.300 74.000 229.700 ;
        RECT 1.300 213.700 73.700 229.300 ;
        RECT 1.000 213.300 74.000 213.700 ;
        RECT 1.300 205.700 73.700 213.300 ;
        RECT 1.000 205.300 74.000 205.700 ;
        RECT 1.300 197.700 73.700 205.300 ;
        RECT 1.000 197.300 74.000 197.700 ;
        RECT 1.300 181.700 73.700 197.300 ;
        RECT 1.000 181.300 74.000 181.700 ;
        RECT 1.300 165.700 73.700 181.300 ;
        RECT 1.000 165.300 74.000 165.700 ;
        RECT 1.300 149.700 73.700 165.300 ;
        RECT 1.000 149.300 74.000 149.700 ;
        RECT 1.300 133.700 73.700 149.300 ;
        RECT 1.000 133.300 74.000 133.700 ;
        RECT 1.300 125.700 73.700 133.300 ;
        RECT 1.000 125.300 74.000 125.700 ;
        RECT 1.300 117.700 73.700 125.300 ;
        RECT 1.000 117.300 74.000 117.700 ;
        RECT 1.300 101.700 73.700 117.300 ;
        RECT 1.000 101.300 74.000 101.700 ;
        RECT 1.300 85.700 73.700 101.300 ;
        RECT 1.000 85.300 74.000 85.700 ;
        RECT 1.300 69.700 73.700 85.300 ;
        RECT 1.000 0.000 74.000 69.700 ;
      LAYER Metal4 ;
        RECT 1.300 341.700 73.700 348.390 ;
        RECT 1.000 341.300 74.000 341.700 ;
        RECT 1.300 333.700 73.700 341.300 ;
        RECT 1.000 333.300 74.000 333.700 ;
        RECT 1.300 325.700 73.700 333.300 ;
        RECT 1.000 325.300 74.000 325.700 ;
        RECT 1.300 317.700 73.700 325.300 ;
        RECT 1.000 317.300 74.000 317.700 ;
        RECT 1.300 309.700 73.700 317.300 ;
        RECT 1.000 309.300 74.000 309.700 ;
        RECT 1.300 301.700 73.700 309.300 ;
        RECT 1.000 301.300 74.000 301.700 ;
        RECT 1.300 293.700 73.700 301.300 ;
        RECT 1.000 293.300 74.000 293.700 ;
        RECT 1.300 285.700 73.700 293.300 ;
        RECT 1.000 285.300 74.000 285.700 ;
        RECT 1.300 277.700 73.700 285.300 ;
        RECT 1.000 277.300 74.000 277.700 ;
        RECT 1.300 269.700 73.700 277.300 ;
        RECT 1.000 269.300 74.000 269.700 ;
        RECT 1.300 261.700 73.700 269.300 ;
        RECT 1.000 261.300 74.000 261.700 ;
        RECT 1.300 253.700 73.700 261.300 ;
        RECT 1.000 253.300 74.000 253.700 ;
        RECT 1.300 245.700 73.700 253.300 ;
        RECT 1.000 245.300 74.000 245.700 ;
        RECT 1.300 229.700 73.700 245.300 ;
        RECT 1.000 229.300 74.000 229.700 ;
        RECT 1.300 213.700 73.700 229.300 ;
        RECT 1.000 213.300 74.000 213.700 ;
        RECT 1.300 205.700 73.700 213.300 ;
        RECT 1.000 205.300 74.000 205.700 ;
        RECT 1.300 197.700 73.700 205.300 ;
        RECT 1.000 197.300 74.000 197.700 ;
        RECT 1.300 181.700 73.700 197.300 ;
        RECT 1.000 181.300 74.000 181.700 ;
        RECT 1.300 165.700 73.700 181.300 ;
        RECT 1.000 165.300 74.000 165.700 ;
        RECT 1.300 149.700 73.700 165.300 ;
        RECT 1.000 149.300 74.000 149.700 ;
        RECT 1.300 133.700 73.700 149.300 ;
        RECT 1.000 133.300 74.000 133.700 ;
        RECT 1.300 125.700 73.700 133.300 ;
        RECT 1.000 125.300 74.000 125.700 ;
        RECT 1.300 117.700 73.700 125.300 ;
        RECT 1.000 117.300 74.000 117.700 ;
        RECT 1.300 101.700 73.700 117.300 ;
        RECT 1.000 101.300 74.000 101.700 ;
        RECT 1.300 85.700 73.700 101.300 ;
        RECT 1.000 85.300 74.000 85.700 ;
        RECT 1.300 69.700 73.700 85.300 ;
        RECT 1.000 0.000 74.000 69.700 ;
      LAYER Metal5 ;
        RECT 1.600 69.400 73.400 348.390 ;
        RECT 1.000 0.000 74.000 69.400 ;
  END
END gf180mcu_fd_io__dvss
END LIBRARY

