magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
<< polysilicon >>
rect 22811 16197 23124 16216
rect 22811 16062 23059 16197
rect 23040 16057 23059 16062
rect 23105 16057 23124 16197
rect 23040 16038 23124 16057
rect 22811 14573 23179 14674
rect 22811 14527 23060 14573
rect 23106 14527 23179 14573
rect 22811 14520 23179 14527
rect 22987 14416 23179 14520
rect 22811 14409 23179 14416
rect 22811 14363 23060 14409
rect 23106 14363 23179 14409
rect 22811 14262 23179 14363
rect 22811 12773 23179 12874
rect 22811 12727 23060 12773
rect 23106 12727 23179 12773
rect 22811 12720 23179 12727
rect 22987 12616 23179 12720
rect 22811 12609 23179 12616
rect 22811 12563 23060 12609
rect 23106 12563 23179 12609
rect 22811 12462 23179 12563
rect 22811 10973 23179 11074
rect 22811 10927 23060 10973
rect 23106 10927 23179 10973
rect 22811 10920 23179 10927
rect 22987 10816 23179 10920
rect 22811 10809 23179 10816
rect 22811 10763 23060 10809
rect 23106 10763 23179 10809
rect 22811 10662 23179 10763
rect 22811 9173 23179 9274
rect 22811 9127 23060 9173
rect 23106 9127 23179 9173
rect 22811 9120 23179 9127
rect 22987 9016 23179 9120
rect 22811 9009 23179 9016
rect 22811 8963 23060 9009
rect 23106 8963 23179 9009
rect 22811 8862 23179 8963
rect 22811 7373 23179 7474
rect 22811 7327 23060 7373
rect 23106 7327 23179 7373
rect 22811 7320 23179 7327
rect 22987 7216 23179 7320
rect 22811 7209 23179 7216
rect 22811 7163 23060 7209
rect 23106 7163 23179 7209
rect 22811 7062 23179 7163
rect 22811 5573 23179 5674
rect 22811 5527 23060 5573
rect 23106 5527 23179 5573
rect 22811 5520 23179 5527
rect 22987 5416 23179 5520
rect 22811 5409 23179 5416
rect 22811 5363 23060 5409
rect 23106 5363 23179 5409
rect 22811 5262 23179 5363
rect 22811 3773 23179 3874
rect 22811 3727 23060 3773
rect 23106 3727 23179 3773
rect 22811 3720 23179 3727
rect 22987 3616 23179 3720
rect 22811 3609 23179 3616
rect 22811 3563 23060 3609
rect 23106 3563 23179 3609
rect 22811 3462 23179 3563
rect 22811 1973 23179 2074
rect 22811 1927 23060 1973
rect 23106 1927 23179 1973
rect 22811 1920 23179 1927
rect 22987 1816 23179 1920
rect 22811 1809 23179 1816
rect 22811 1763 23060 1809
rect 23106 1763 23179 1809
rect 22811 1662 23179 1763
rect 22987 413 23179 459
rect 22987 367 23060 413
rect 23106 367 23179 413
rect 22987 274 23179 367
rect 22811 249 23179 274
rect 22811 203 23060 249
rect 23106 203 23179 249
rect 22811 120 23179 203
<< polycontact >>
rect 23059 16057 23105 16197
rect 23060 14527 23106 14573
rect 23060 14363 23106 14409
rect 23060 12727 23106 12773
rect 23060 12563 23106 12609
rect 23060 10927 23106 10973
rect 23060 10763 23106 10809
rect 23060 9127 23106 9173
rect 23060 8963 23106 9009
rect 23060 7327 23106 7373
rect 23060 7163 23106 7209
rect 23060 5527 23106 5573
rect 23060 5363 23106 5409
rect 23060 3727 23106 3773
rect 23060 3563 23106 3609
rect 23060 1927 23106 1973
rect 23060 1763 23106 1809
rect 23060 367 23106 413
rect 23060 203 23106 249
<< metal1 >>
rect 23044 16197 23120 16208
rect 23044 16196 23059 16197
rect 23105 16196 23120 16197
rect 23044 15936 23056 16196
rect 23108 15936 23120 16196
rect 23044 15924 23120 15936
rect 23019 14605 23143 14645
rect 23019 14553 23055 14605
rect 23107 14553 23143 14605
rect 23019 14527 23060 14553
rect 23106 14527 23143 14553
rect 23019 14409 23143 14527
rect 23019 14387 23060 14409
rect 23106 14387 23143 14409
rect 23019 14335 23055 14387
rect 23107 14335 23143 14387
rect 23019 14295 23143 14335
rect 23019 12801 23143 12841
rect 23019 12749 23055 12801
rect 23107 12749 23143 12801
rect 23019 12727 23060 12749
rect 23106 12727 23143 12749
rect 23019 12609 23143 12727
rect 23019 12583 23060 12609
rect 23106 12583 23143 12609
rect 23019 12531 23055 12583
rect 23107 12531 23143 12583
rect 23019 12491 23143 12531
rect 23019 11005 23143 11045
rect 23019 10953 23055 11005
rect 23107 10953 23143 11005
rect 23019 10927 23060 10953
rect 23106 10927 23143 10953
rect 23019 10809 23143 10927
rect 23019 10787 23060 10809
rect 23106 10787 23143 10809
rect 23019 10735 23055 10787
rect 23107 10735 23143 10787
rect 23019 10695 23143 10735
rect 23019 9201 23143 9241
rect 23019 9149 23055 9201
rect 23107 9149 23143 9201
rect 23019 9127 23060 9149
rect 23106 9127 23143 9149
rect 23019 9009 23143 9127
rect 23019 8983 23060 9009
rect 23106 8983 23143 9009
rect 23019 8931 23055 8983
rect 23107 8931 23143 8983
rect 23019 8891 23143 8931
rect 23019 7405 23143 7445
rect 23019 7353 23055 7405
rect 23107 7353 23143 7405
rect 23019 7327 23060 7353
rect 23106 7327 23143 7353
rect 23019 7209 23143 7327
rect 23019 7187 23060 7209
rect 23106 7187 23143 7209
rect 23019 7135 23055 7187
rect 23107 7135 23143 7187
rect 23019 7095 23143 7135
rect 23019 5601 23143 5641
rect 23019 5549 23055 5601
rect 23107 5549 23143 5601
rect 23019 5527 23060 5549
rect 23106 5527 23143 5549
rect 23019 5409 23143 5527
rect 23019 5383 23060 5409
rect 23106 5383 23143 5409
rect 23019 5331 23055 5383
rect 23107 5331 23143 5383
rect 23019 5291 23143 5331
rect 23019 3805 23143 3845
rect 23019 3753 23055 3805
rect 23107 3753 23143 3805
rect 23019 3727 23060 3753
rect 23106 3727 23143 3753
rect 23019 3609 23143 3727
rect 23019 3587 23060 3609
rect 23106 3587 23143 3609
rect 23019 3535 23055 3587
rect 23107 3535 23143 3587
rect 23019 3495 23143 3535
rect 23019 2001 23143 2041
rect 23019 1949 23055 2001
rect 23107 1949 23143 2001
rect 23019 1927 23060 1949
rect 23106 1927 23143 1949
rect 23019 1809 23143 1927
rect 23019 1783 23060 1809
rect 23106 1783 23143 1809
rect 23019 1731 23055 1783
rect 23107 1731 23143 1783
rect 23019 1691 23143 1731
rect 23027 413 23139 450
rect 23027 367 23060 413
rect 23106 367 23139 413
rect 23027 346 23139 367
rect 23027 190 23055 346
rect 23107 190 23139 346
rect 23027 167 23139 190
<< via1 >>
rect 23056 16057 23059 16196
rect 23059 16057 23105 16196
rect 23105 16057 23108 16196
rect 23056 15936 23108 16057
rect 23055 14573 23107 14605
rect 23055 14553 23060 14573
rect 23060 14553 23106 14573
rect 23106 14553 23107 14573
rect 23055 14363 23060 14387
rect 23060 14363 23106 14387
rect 23106 14363 23107 14387
rect 23055 14335 23107 14363
rect 23055 12773 23107 12801
rect 23055 12749 23060 12773
rect 23060 12749 23106 12773
rect 23106 12749 23107 12773
rect 23055 12563 23060 12583
rect 23060 12563 23106 12583
rect 23106 12563 23107 12583
rect 23055 12531 23107 12563
rect 23055 10973 23107 11005
rect 23055 10953 23060 10973
rect 23060 10953 23106 10973
rect 23106 10953 23107 10973
rect 23055 10763 23060 10787
rect 23060 10763 23106 10787
rect 23106 10763 23107 10787
rect 23055 10735 23107 10763
rect 23055 9173 23107 9201
rect 23055 9149 23060 9173
rect 23060 9149 23106 9173
rect 23106 9149 23107 9173
rect 23055 8963 23060 8983
rect 23060 8963 23106 8983
rect 23106 8963 23107 8983
rect 23055 8931 23107 8963
rect 23055 7373 23107 7405
rect 23055 7353 23060 7373
rect 23060 7353 23106 7373
rect 23106 7353 23107 7373
rect 23055 7163 23060 7187
rect 23060 7163 23106 7187
rect 23106 7163 23107 7187
rect 23055 7135 23107 7163
rect 23055 5573 23107 5601
rect 23055 5549 23060 5573
rect 23060 5549 23106 5573
rect 23106 5549 23107 5573
rect 23055 5363 23060 5383
rect 23060 5363 23106 5383
rect 23106 5363 23107 5383
rect 23055 5331 23107 5363
rect 23055 3773 23107 3805
rect 23055 3753 23060 3773
rect 23060 3753 23106 3773
rect 23106 3753 23107 3773
rect 23055 3563 23060 3587
rect 23060 3563 23106 3587
rect 23106 3563 23107 3587
rect 23055 3535 23107 3563
rect 23055 1973 23107 2001
rect 23055 1949 23060 1973
rect 23060 1949 23106 1973
rect 23106 1949 23107 1973
rect 23055 1763 23060 1783
rect 23060 1763 23106 1783
rect 23106 1763 23107 1783
rect 23055 1731 23107 1763
rect 23055 249 23107 346
rect 23055 203 23060 249
rect 23060 203 23106 249
rect 23106 203 23107 249
rect 23055 190 23107 203
<< metal2 >>
rect 23018 16347 23143 16368
rect 23018 16187 23054 16347
rect 23110 16187 23143 16347
rect 23018 15936 23056 16187
rect 23108 15936 23143 16187
rect 23018 14605 23143 15936
rect 23018 14553 23055 14605
rect 23107 14553 23143 14605
rect 23018 14387 23143 14553
rect 23018 14335 23055 14387
rect 23107 14335 23143 14387
rect 23018 12801 23143 14335
rect 23018 12749 23055 12801
rect 23107 12749 23143 12801
rect 23018 12583 23143 12749
rect 23018 12531 23055 12583
rect 23107 12531 23143 12583
rect 23018 11005 23143 12531
rect 23018 10953 23055 11005
rect 23107 10953 23143 11005
rect 23018 10787 23143 10953
rect 23018 10735 23055 10787
rect 23107 10735 23143 10787
rect 23018 9201 23143 10735
rect 23018 9149 23055 9201
rect 23107 9149 23143 9201
rect 23018 8983 23143 9149
rect 23018 8931 23055 8983
rect 23107 8931 23143 8983
rect 23018 7405 23143 8931
rect 23018 7353 23055 7405
rect 23107 7353 23143 7405
rect 23018 7187 23143 7353
rect 23018 7135 23055 7187
rect 23107 7135 23143 7187
rect 23018 5601 23143 7135
rect 23018 5549 23055 5601
rect 23107 5549 23143 5601
rect 23018 5383 23143 5549
rect 23018 5331 23055 5383
rect 23107 5331 23143 5383
rect 23018 3805 23143 5331
rect 23018 3753 23055 3805
rect 23107 3753 23143 3805
rect 23018 3587 23143 3753
rect 23018 3535 23055 3587
rect 23107 3535 23143 3587
rect 23018 2001 23143 3535
rect 23018 1949 23055 2001
rect 23107 1949 23143 2001
rect 23018 1783 23143 1949
rect 23018 1731 23055 1783
rect 23107 1731 23143 1783
rect 23018 346 23143 1731
rect 23018 190 23055 346
rect 23107 190 23143 346
rect 23018 144 23143 190
rect 23018 -16 23053 144
rect 23109 -16 23143 144
rect 23018 -33 23143 -16
<< via2 >>
rect 23054 16196 23110 16347
rect 23054 16187 23056 16196
rect 23056 16187 23108 16196
rect 23108 16187 23110 16196
rect 23053 -16 23109 144
<< metal3 >>
rect -30 16347 23144 16368
rect -30 16187 23054 16347
rect 23110 16187 23144 16347
rect -30 16168 23144 16187
rect -30 144 23143 168
rect -30 -16 23053 144
rect 23109 -16 23143 144
rect -30 -32 23143 -16
use 018SRAM_cell1_128x8m81  018SRAM_cell1_128x8m81_0
timestamp 1762296095
transform -1 0 22868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_128x8m81  018SRAM_cell1_128x8m81_1
timestamp 1762296095
transform -1 0 22868 0 -1 16268
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_0
timestamp 1762296095
transform -1 0 22868 0 1 14468
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_1
timestamp 1762296095
transform -1 0 22868 0 1 9068
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_2
timestamp 1762296095
transform -1 0 22868 0 1 10868
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_3
timestamp 1762296095
transform -1 0 22868 0 1 7268
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_4
timestamp 1762296095
transform -1 0 22868 0 1 1868
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_5
timestamp 1762296095
transform -1 0 22868 0 1 3668
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_6
timestamp 1762296095
transform -1 0 22868 0 1 5468
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_7
timestamp 1762296095
transform -1 0 22868 0 1 12668
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_8
timestamp 1762296095
transform -1 0 22868 0 -1 14468
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_9
timestamp 1762296095
transform -1 0 22868 0 -1 12668
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_10
timestamp 1762296095
transform -1 0 22868 0 -1 10868
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_11
timestamp 1762296095
transform -1 0 22868 0 -1 7268
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_12
timestamp 1762296095
transform -1 0 22868 0 -1 9068
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_13
timestamp 1762296095
transform -1 0 22868 0 -1 5468
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_14
timestamp 1762296095
transform -1 0 22868 0 -1 1868
box -68 -68 668 968
use 018SRAM_cell1_cutPC_128x8m81  018SRAM_cell1_cutPC_128x8m81_15
timestamp 1762296095
transform -1 0 22868 0 -1 3668
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_0
timestamp 1762296095
transform -1 0 17468 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_1
timestamp 1762296095
transform -1 0 18068 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_2
timestamp 1762296095
transform -1 0 19268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_3
timestamp 1762296095
transform -1 0 18668 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_4
timestamp 1762296095
transform -1 0 19868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_5
timestamp 1762296095
transform -1 0 20468 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_6
timestamp 1762296095
transform -1 0 21068 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_7
timestamp 1762296095
transform -1 0 21668 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_8
timestamp 1762296095
transform -1 0 16268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_9
timestamp 1762296095
transform -1 0 15668 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_10
timestamp 1762296095
transform -1 0 15068 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_11
timestamp 1762296095
transform -1 0 14468 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_12
timestamp 1762296095
transform -1 0 13268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_13
timestamp 1762296095
transform -1 0 13868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_14
timestamp 1762296095
transform -1 0 12668 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_15
timestamp 1762296095
transform -1 0 12068 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_16
timestamp 1762296095
transform -1 0 7268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_17
timestamp 1762296095
transform -1 0 8468 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_18
timestamp 1762296095
transform -1 0 7868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_19
timestamp 1762296095
transform -1 0 9068 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_20
timestamp 1762296095
transform -1 0 9668 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_21
timestamp 1762296095
transform -1 0 10268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_22
timestamp 1762296095
transform -1 0 10868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_23
timestamp 1762296095
transform -1 0 5468 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_24
timestamp 1762296095
transform -1 0 4868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_25
timestamp 1762296095
transform -1 0 4268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_26
timestamp 1762296095
transform -1 0 3668 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_27
timestamp 1762296095
transform -1 0 2468 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_28
timestamp 1762296095
transform -1 0 3068 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_29
timestamp 1762296095
transform -1 0 1868 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_30
timestamp 1762296095
transform -1 0 1268 0 1 68
box -68 -68 668 968
use 018SRAM_cell1_dummy_128x8m81  018SRAM_cell1_dummy_128x8m81_31
timestamp 1762296095
transform -1 0 6668 0 1 68
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_0
timestamp 1762296095
transform -1 0 16868 0 1 68
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_1
timestamp 1762296095
transform -1 0 11468 0 1 68
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_2
timestamp 1762296095
transform -1 0 6068 0 1 68
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_3
timestamp 1762296095
transform -1 0 668 0 1 68
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_4
timestamp 1762296095
transform -1 0 668 0 -1 16268
box -68 -68 668 968
use 018SRAM_strap1_128x8m81  018SRAM_strap1_128x8m81_5
timestamp 1762296095
transform 1 0 21668 0 1 68
box -68 -68 668 968
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_0
timestamp 1762296095
transform 1 0 23083 0 -1 308
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_1
timestamp 1762296095
transform 1 0 23083 0 -1 12668
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_2
timestamp 1762296095
transform 1 0 23083 0 -1 9068
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_3
timestamp 1762296095
transform 1 0 23083 0 -1 14468
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_4
timestamp 1762296095
transform 1 0 23083 0 -1 10868
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_5
timestamp 1762296095
transform 1 0 23083 0 -1 7268
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_6
timestamp 1762296095
transform 1 0 23083 0 -1 5468
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_7
timestamp 1762296095
transform 1 0 23083 0 -1 1868
box 0 0 1 1
use M1_POLY2$$44754988_128x8m81  M1_POLY2$$44754988_128x8m81_8
timestamp 1762296095
transform 1 0 23083 0 -1 3668
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1762296095
transform 1 0 23082 0 1 16127
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_0
timestamp 1762296095
transform 1 0 23081 0 -1 14470
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_1
timestamp 1762296095
transform 1 0 23081 0 -1 3670
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_2
timestamp 1762296095
transform 1 0 23081 0 -1 10870
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_3
timestamp 1762296095
transform 1 0 23081 0 -1 1866
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_4
timestamp 1762296095
transform 1 0 23081 0 -1 5466
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_5
timestamp 1762296095
transform 1 0 23081 0 -1 9066
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_6
timestamp 1762296095
transform 1 0 23081 0 -1 12666
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_7
timestamp 1762296095
transform 1 0 23081 0 -1 7270
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_0
timestamp 1762296095
transform 1 0 23081 0 1 268
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_0
timestamp 1762296095
transform 1 0 23082 0 1 16066
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_0
timestamp 1762296095
transform 1 0 23082 0 1 16267
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_1
timestamp 1762296095
transform 1 0 23081 0 1 64
box 0 0 1 1
use new_dummyrow_unit_01_128x8m81  new_dummyrow_unit_01_128x8m81_0
timestamp 1762296095
transform 1 0 606 0 -1 16445
box -6 109 10930 1145
use new_dummyrow_unit_128x8m81  new_dummyrow_unit_128x8m81_0
timestamp 1762296095
transform 1 0 11406 0 -1 16445
box -6 109 10930 1145
<< labels >>
rlabel metal3 s 22802 1886 22802 1886 4 VSS
rlabel metal3 s 22802 961 22802 961 4 VDD
<< properties >>
string GDS_END 1670832
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1664152
<< end >>
