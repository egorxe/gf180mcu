magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< metal1 >>
rect -44 7926 200 8000
rect -44 7874 0 7926
rect 156 7874 200 7926
rect -44 7802 200 7874
rect -44 7750 0 7802
rect 156 7750 200 7802
rect -44 7678 200 7750
rect -44 7626 0 7678
rect 156 7626 200 7678
rect -44 7554 200 7626
rect -44 7502 0 7554
rect 156 7502 200 7554
rect -44 7430 200 7502
rect -44 7378 0 7430
rect 156 7378 200 7430
rect -44 7306 200 7378
rect -44 7254 0 7306
rect 156 7254 200 7306
rect -44 7182 200 7254
rect -44 7130 0 7182
rect 156 7130 200 7182
rect -44 7058 200 7130
rect -44 7006 0 7058
rect 156 7006 200 7058
rect -44 6934 200 7006
rect -44 6882 0 6934
rect 156 6882 200 6934
rect -44 6810 200 6882
rect -44 6758 0 6810
rect 156 6758 200 6810
rect -44 6686 200 6758
rect -44 6634 0 6686
rect 156 6634 200 6686
rect -44 6562 200 6634
rect -44 6510 0 6562
rect 156 6510 200 6562
rect -44 6438 200 6510
rect -44 6386 0 6438
rect 156 6386 200 6438
rect -44 6314 200 6386
rect -44 6262 0 6314
rect 156 6262 200 6314
rect -44 6190 200 6262
rect -44 6138 0 6190
rect 156 6138 200 6190
rect -44 6066 200 6138
rect -44 6014 0 6066
rect 156 6014 200 6066
rect -44 5942 200 6014
rect -44 5890 0 5942
rect 156 5890 200 5942
rect -44 5818 200 5890
rect -44 5766 0 5818
rect 156 5766 200 5818
rect -44 5694 200 5766
rect -44 5642 0 5694
rect 156 5642 200 5694
rect -44 5570 200 5642
rect -44 5518 0 5570
rect 156 5518 200 5570
rect -44 5446 200 5518
rect -44 5394 0 5446
rect 156 5394 200 5446
rect -44 5322 200 5394
rect -44 5270 0 5322
rect 156 5270 200 5322
rect -44 5198 200 5270
rect -44 5146 0 5198
rect 156 5146 200 5198
rect -44 5074 200 5146
rect -44 5022 0 5074
rect 156 5022 200 5074
rect -44 4950 200 5022
rect -44 4898 0 4950
rect 156 4898 200 4950
rect -44 4826 200 4898
rect -44 4774 0 4826
rect 156 4774 200 4826
rect -44 4702 200 4774
rect -44 4650 0 4702
rect 156 4650 200 4702
rect -44 4578 200 4650
rect -44 4526 0 4578
rect 156 4526 200 4578
rect -44 4454 200 4526
rect -44 4402 0 4454
rect 156 4402 200 4454
rect -44 4330 200 4402
rect -44 4278 0 4330
rect 156 4278 200 4330
rect -44 4206 200 4278
rect -44 4154 0 4206
rect 156 4154 200 4206
rect -44 4082 200 4154
rect -44 4030 0 4082
rect 156 4030 200 4082
rect -44 3958 200 4030
rect -44 3906 0 3958
rect 156 3906 200 3958
rect -44 3834 200 3906
rect -44 3782 0 3834
rect 156 3782 200 3834
rect -44 3710 200 3782
rect -44 3658 0 3710
rect 156 3658 200 3710
rect -44 3586 200 3658
rect -44 3534 0 3586
rect 156 3534 200 3586
rect -44 3462 200 3534
rect -44 3410 0 3462
rect 156 3410 200 3462
rect -44 3338 200 3410
rect -44 3286 0 3338
rect 156 3286 200 3338
rect -44 3214 200 3286
rect -44 3162 0 3214
rect 156 3162 200 3214
rect -44 3090 200 3162
rect -44 3038 0 3090
rect 156 3038 200 3090
rect -44 2966 200 3038
rect -44 2914 0 2966
rect 156 2914 200 2966
rect -44 2842 200 2914
rect -44 2790 0 2842
rect 156 2790 200 2842
rect -44 2718 200 2790
rect -44 2666 0 2718
rect 156 2666 200 2718
rect -44 2594 200 2666
rect -44 2542 0 2594
rect 156 2542 200 2594
rect -44 2470 200 2542
rect -44 2418 0 2470
rect 156 2418 200 2470
rect -44 2346 200 2418
rect -44 2294 0 2346
rect 156 2294 200 2346
rect -44 2222 200 2294
rect -44 2170 0 2222
rect 156 2170 200 2222
rect -44 2098 200 2170
rect -44 2046 0 2098
rect 156 2046 200 2098
rect -44 1974 200 2046
rect -44 1922 0 1974
rect 156 1922 200 1974
rect -44 1850 200 1922
rect -44 1798 0 1850
rect 156 1798 200 1850
rect -44 1726 200 1798
rect -44 1674 0 1726
rect 156 1674 200 1726
rect -44 1602 200 1674
rect -44 1550 0 1602
rect 156 1550 200 1602
rect -44 1478 200 1550
rect -44 1426 0 1478
rect 156 1426 200 1478
rect -44 1354 200 1426
rect -44 1302 0 1354
rect 156 1302 200 1354
rect -44 1230 200 1302
rect -44 1178 0 1230
rect 156 1178 200 1230
rect -44 1106 200 1178
rect -44 1054 0 1106
rect 156 1054 200 1106
rect -44 982 200 1054
rect -44 930 0 982
rect 156 930 200 982
rect -44 858 200 930
rect -44 806 0 858
rect 156 806 200 858
rect -44 734 200 806
rect -44 682 0 734
rect 156 682 200 734
rect -44 610 200 682
rect -44 558 0 610
rect 156 558 200 610
rect -44 486 200 558
rect -44 434 0 486
rect 156 434 200 486
rect -44 362 200 434
rect -44 310 0 362
rect 156 310 200 362
rect -44 238 200 310
rect -44 186 0 238
rect 156 186 200 238
rect -44 114 200 186
rect -44 62 0 114
rect 156 62 200 114
rect -44 0 200 62
rect 340 7926 1584 8000
rect 340 7874 378 7926
rect 430 7874 502 7926
rect 554 7874 626 7926
rect 678 7874 750 7926
rect 802 7874 874 7926
rect 926 7874 998 7926
rect 1050 7874 1122 7926
rect 1174 7874 1246 7926
rect 1298 7874 1370 7926
rect 1422 7874 1494 7926
rect 1546 7874 1584 7926
rect 340 7802 1584 7874
rect 340 7750 378 7802
rect 430 7750 502 7802
rect 554 7750 626 7802
rect 678 7750 750 7802
rect 802 7750 874 7802
rect 926 7750 998 7802
rect 1050 7750 1122 7802
rect 1174 7750 1246 7802
rect 1298 7750 1370 7802
rect 1422 7750 1494 7802
rect 1546 7750 1584 7802
rect 340 7678 1584 7750
rect 340 7626 378 7678
rect 430 7626 502 7678
rect 554 7626 626 7678
rect 678 7626 750 7678
rect 802 7626 874 7678
rect 926 7626 998 7678
rect 1050 7626 1122 7678
rect 1174 7626 1246 7678
rect 1298 7626 1370 7678
rect 1422 7626 1494 7678
rect 1546 7626 1584 7678
rect 340 7554 1584 7626
rect 340 7502 378 7554
rect 430 7502 502 7554
rect 554 7502 626 7554
rect 678 7502 750 7554
rect 802 7502 874 7554
rect 926 7502 998 7554
rect 1050 7502 1122 7554
rect 1174 7502 1246 7554
rect 1298 7502 1370 7554
rect 1422 7502 1494 7554
rect 1546 7502 1584 7554
rect 340 7430 1584 7502
rect 340 7378 378 7430
rect 430 7378 502 7430
rect 554 7378 626 7430
rect 678 7378 750 7430
rect 802 7378 874 7430
rect 926 7378 998 7430
rect 1050 7378 1122 7430
rect 1174 7378 1246 7430
rect 1298 7378 1370 7430
rect 1422 7378 1494 7430
rect 1546 7378 1584 7430
rect 340 7306 1584 7378
rect 340 7254 378 7306
rect 430 7254 502 7306
rect 554 7254 626 7306
rect 678 7254 750 7306
rect 802 7254 874 7306
rect 926 7254 998 7306
rect 1050 7254 1122 7306
rect 1174 7254 1246 7306
rect 1298 7254 1370 7306
rect 1422 7254 1494 7306
rect 1546 7254 1584 7306
rect 340 7182 1584 7254
rect 340 7130 378 7182
rect 430 7130 502 7182
rect 554 7130 626 7182
rect 678 7130 750 7182
rect 802 7130 874 7182
rect 926 7130 998 7182
rect 1050 7130 1122 7182
rect 1174 7130 1246 7182
rect 1298 7130 1370 7182
rect 1422 7130 1494 7182
rect 1546 7130 1584 7182
rect 340 7058 1584 7130
rect 340 7006 378 7058
rect 430 7006 502 7058
rect 554 7006 626 7058
rect 678 7006 750 7058
rect 802 7006 874 7058
rect 926 7006 998 7058
rect 1050 7006 1122 7058
rect 1174 7006 1246 7058
rect 1298 7006 1370 7058
rect 1422 7006 1494 7058
rect 1546 7006 1584 7058
rect 340 6934 1584 7006
rect 340 6882 378 6934
rect 430 6882 502 6934
rect 554 6882 626 6934
rect 678 6882 750 6934
rect 802 6882 874 6934
rect 926 6882 998 6934
rect 1050 6882 1122 6934
rect 1174 6882 1246 6934
rect 1298 6882 1370 6934
rect 1422 6882 1494 6934
rect 1546 6882 1584 6934
rect 340 6810 1584 6882
rect 340 6758 378 6810
rect 430 6758 502 6810
rect 554 6758 626 6810
rect 678 6758 750 6810
rect 802 6758 874 6810
rect 926 6758 998 6810
rect 1050 6758 1122 6810
rect 1174 6758 1246 6810
rect 1298 6758 1370 6810
rect 1422 6758 1494 6810
rect 1546 6758 1584 6810
rect 340 6686 1584 6758
rect 340 6634 378 6686
rect 430 6634 502 6686
rect 554 6634 626 6686
rect 678 6634 750 6686
rect 802 6634 874 6686
rect 926 6634 998 6686
rect 1050 6634 1122 6686
rect 1174 6634 1246 6686
rect 1298 6634 1370 6686
rect 1422 6634 1494 6686
rect 1546 6634 1584 6686
rect 340 6562 1584 6634
rect 340 6510 378 6562
rect 430 6510 502 6562
rect 554 6510 626 6562
rect 678 6510 750 6562
rect 802 6510 874 6562
rect 926 6510 998 6562
rect 1050 6510 1122 6562
rect 1174 6510 1246 6562
rect 1298 6510 1370 6562
rect 1422 6510 1494 6562
rect 1546 6510 1584 6562
rect 340 6438 1584 6510
rect 340 6386 378 6438
rect 430 6386 502 6438
rect 554 6386 626 6438
rect 678 6386 750 6438
rect 802 6386 874 6438
rect 926 6386 998 6438
rect 1050 6386 1122 6438
rect 1174 6386 1246 6438
rect 1298 6386 1370 6438
rect 1422 6386 1494 6438
rect 1546 6386 1584 6438
rect 340 6314 1584 6386
rect 340 6262 378 6314
rect 430 6262 502 6314
rect 554 6262 626 6314
rect 678 6262 750 6314
rect 802 6262 874 6314
rect 926 6262 998 6314
rect 1050 6262 1122 6314
rect 1174 6262 1246 6314
rect 1298 6262 1370 6314
rect 1422 6262 1494 6314
rect 1546 6262 1584 6314
rect 340 6190 1584 6262
rect 340 6138 378 6190
rect 430 6138 502 6190
rect 554 6138 626 6190
rect 678 6138 750 6190
rect 802 6138 874 6190
rect 926 6138 998 6190
rect 1050 6138 1122 6190
rect 1174 6138 1246 6190
rect 1298 6138 1370 6190
rect 1422 6138 1494 6190
rect 1546 6138 1584 6190
rect 340 6066 1584 6138
rect 340 6014 378 6066
rect 430 6014 502 6066
rect 554 6014 626 6066
rect 678 6014 750 6066
rect 802 6014 874 6066
rect 926 6014 998 6066
rect 1050 6014 1122 6066
rect 1174 6014 1246 6066
rect 1298 6014 1370 6066
rect 1422 6014 1494 6066
rect 1546 6014 1584 6066
rect 340 5942 1584 6014
rect 340 5890 378 5942
rect 430 5890 502 5942
rect 554 5890 626 5942
rect 678 5890 750 5942
rect 802 5890 874 5942
rect 926 5890 998 5942
rect 1050 5890 1122 5942
rect 1174 5890 1246 5942
rect 1298 5890 1370 5942
rect 1422 5890 1494 5942
rect 1546 5890 1584 5942
rect 340 5818 1584 5890
rect 340 5766 378 5818
rect 430 5766 502 5818
rect 554 5766 626 5818
rect 678 5766 750 5818
rect 802 5766 874 5818
rect 926 5766 998 5818
rect 1050 5766 1122 5818
rect 1174 5766 1246 5818
rect 1298 5766 1370 5818
rect 1422 5766 1494 5818
rect 1546 5766 1584 5818
rect 340 5694 1584 5766
rect 340 5642 378 5694
rect 430 5642 502 5694
rect 554 5642 626 5694
rect 678 5642 750 5694
rect 802 5642 874 5694
rect 926 5642 998 5694
rect 1050 5642 1122 5694
rect 1174 5642 1246 5694
rect 1298 5642 1370 5694
rect 1422 5642 1494 5694
rect 1546 5642 1584 5694
rect 340 5570 1584 5642
rect 340 5518 378 5570
rect 430 5518 502 5570
rect 554 5518 626 5570
rect 678 5518 750 5570
rect 802 5518 874 5570
rect 926 5518 998 5570
rect 1050 5518 1122 5570
rect 1174 5518 1246 5570
rect 1298 5518 1370 5570
rect 1422 5518 1494 5570
rect 1546 5518 1584 5570
rect 340 5446 1584 5518
rect 340 5394 378 5446
rect 430 5394 502 5446
rect 554 5394 626 5446
rect 678 5394 750 5446
rect 802 5394 874 5446
rect 926 5394 998 5446
rect 1050 5394 1122 5446
rect 1174 5394 1246 5446
rect 1298 5394 1370 5446
rect 1422 5394 1494 5446
rect 1546 5394 1584 5446
rect 340 5322 1584 5394
rect 340 5270 378 5322
rect 430 5270 502 5322
rect 554 5270 626 5322
rect 678 5270 750 5322
rect 802 5270 874 5322
rect 926 5270 998 5322
rect 1050 5270 1122 5322
rect 1174 5270 1246 5322
rect 1298 5270 1370 5322
rect 1422 5270 1494 5322
rect 1546 5270 1584 5322
rect 340 5198 1584 5270
rect 340 5146 378 5198
rect 430 5146 502 5198
rect 554 5146 626 5198
rect 678 5146 750 5198
rect 802 5146 874 5198
rect 926 5146 998 5198
rect 1050 5146 1122 5198
rect 1174 5146 1246 5198
rect 1298 5146 1370 5198
rect 1422 5146 1494 5198
rect 1546 5146 1584 5198
rect 340 5074 1584 5146
rect 340 5022 378 5074
rect 430 5022 502 5074
rect 554 5022 626 5074
rect 678 5022 750 5074
rect 802 5022 874 5074
rect 926 5022 998 5074
rect 1050 5022 1122 5074
rect 1174 5022 1246 5074
rect 1298 5022 1370 5074
rect 1422 5022 1494 5074
rect 1546 5022 1584 5074
rect 340 4950 1584 5022
rect 340 4898 378 4950
rect 430 4898 502 4950
rect 554 4898 626 4950
rect 678 4898 750 4950
rect 802 4898 874 4950
rect 926 4898 998 4950
rect 1050 4898 1122 4950
rect 1174 4898 1246 4950
rect 1298 4898 1370 4950
rect 1422 4898 1494 4950
rect 1546 4898 1584 4950
rect 340 4826 1584 4898
rect 340 4774 378 4826
rect 430 4774 502 4826
rect 554 4774 626 4826
rect 678 4774 750 4826
rect 802 4774 874 4826
rect 926 4774 998 4826
rect 1050 4774 1122 4826
rect 1174 4774 1246 4826
rect 1298 4774 1370 4826
rect 1422 4774 1494 4826
rect 1546 4774 1584 4826
rect 340 4702 1584 4774
rect 340 4650 378 4702
rect 430 4650 502 4702
rect 554 4650 626 4702
rect 678 4650 750 4702
rect 802 4650 874 4702
rect 926 4650 998 4702
rect 1050 4650 1122 4702
rect 1174 4650 1246 4702
rect 1298 4650 1370 4702
rect 1422 4650 1494 4702
rect 1546 4650 1584 4702
rect 340 4578 1584 4650
rect 340 4526 378 4578
rect 430 4526 502 4578
rect 554 4526 626 4578
rect 678 4526 750 4578
rect 802 4526 874 4578
rect 926 4526 998 4578
rect 1050 4526 1122 4578
rect 1174 4526 1246 4578
rect 1298 4526 1370 4578
rect 1422 4526 1494 4578
rect 1546 4526 1584 4578
rect 340 4454 1584 4526
rect 340 4402 378 4454
rect 430 4402 502 4454
rect 554 4402 626 4454
rect 678 4402 750 4454
rect 802 4402 874 4454
rect 926 4402 998 4454
rect 1050 4402 1122 4454
rect 1174 4402 1246 4454
rect 1298 4402 1370 4454
rect 1422 4402 1494 4454
rect 1546 4402 1584 4454
rect 340 4330 1584 4402
rect 340 4278 378 4330
rect 430 4278 502 4330
rect 554 4278 626 4330
rect 678 4278 750 4330
rect 802 4278 874 4330
rect 926 4278 998 4330
rect 1050 4278 1122 4330
rect 1174 4278 1246 4330
rect 1298 4278 1370 4330
rect 1422 4278 1494 4330
rect 1546 4278 1584 4330
rect 340 4206 1584 4278
rect 340 4154 378 4206
rect 430 4154 502 4206
rect 554 4154 626 4206
rect 678 4154 750 4206
rect 802 4154 874 4206
rect 926 4154 998 4206
rect 1050 4154 1122 4206
rect 1174 4154 1246 4206
rect 1298 4154 1370 4206
rect 1422 4154 1494 4206
rect 1546 4154 1584 4206
rect 340 4082 1584 4154
rect 340 4030 378 4082
rect 430 4030 502 4082
rect 554 4030 626 4082
rect 678 4030 750 4082
rect 802 4030 874 4082
rect 926 4030 998 4082
rect 1050 4030 1122 4082
rect 1174 4030 1246 4082
rect 1298 4030 1370 4082
rect 1422 4030 1494 4082
rect 1546 4030 1584 4082
rect 340 3958 1584 4030
rect 340 3906 378 3958
rect 430 3906 502 3958
rect 554 3906 626 3958
rect 678 3906 750 3958
rect 802 3906 874 3958
rect 926 3906 998 3958
rect 1050 3906 1122 3958
rect 1174 3906 1246 3958
rect 1298 3906 1370 3958
rect 1422 3906 1494 3958
rect 1546 3906 1584 3958
rect 340 3834 1584 3906
rect 340 3782 378 3834
rect 430 3782 502 3834
rect 554 3782 626 3834
rect 678 3782 750 3834
rect 802 3782 874 3834
rect 926 3782 998 3834
rect 1050 3782 1122 3834
rect 1174 3782 1246 3834
rect 1298 3782 1370 3834
rect 1422 3782 1494 3834
rect 1546 3782 1584 3834
rect 340 3710 1584 3782
rect 340 3658 378 3710
rect 430 3658 502 3710
rect 554 3658 626 3710
rect 678 3658 750 3710
rect 802 3658 874 3710
rect 926 3658 998 3710
rect 1050 3658 1122 3710
rect 1174 3658 1246 3710
rect 1298 3658 1370 3710
rect 1422 3658 1494 3710
rect 1546 3658 1584 3710
rect 340 3586 1584 3658
rect 340 3534 378 3586
rect 430 3534 502 3586
rect 554 3534 626 3586
rect 678 3534 750 3586
rect 802 3534 874 3586
rect 926 3534 998 3586
rect 1050 3534 1122 3586
rect 1174 3534 1246 3586
rect 1298 3534 1370 3586
rect 1422 3534 1494 3586
rect 1546 3534 1584 3586
rect 340 3462 1584 3534
rect 340 3410 378 3462
rect 430 3410 502 3462
rect 554 3410 626 3462
rect 678 3410 750 3462
rect 802 3410 874 3462
rect 926 3410 998 3462
rect 1050 3410 1122 3462
rect 1174 3410 1246 3462
rect 1298 3410 1370 3462
rect 1422 3410 1494 3462
rect 1546 3410 1584 3462
rect 340 3338 1584 3410
rect 340 3286 378 3338
rect 430 3286 502 3338
rect 554 3286 626 3338
rect 678 3286 750 3338
rect 802 3286 874 3338
rect 926 3286 998 3338
rect 1050 3286 1122 3338
rect 1174 3286 1246 3338
rect 1298 3286 1370 3338
rect 1422 3286 1494 3338
rect 1546 3286 1584 3338
rect 340 3214 1584 3286
rect 340 3162 378 3214
rect 430 3162 502 3214
rect 554 3162 626 3214
rect 678 3162 750 3214
rect 802 3162 874 3214
rect 926 3162 998 3214
rect 1050 3162 1122 3214
rect 1174 3162 1246 3214
rect 1298 3162 1370 3214
rect 1422 3162 1494 3214
rect 1546 3162 1584 3214
rect 340 3090 1584 3162
rect 340 3038 378 3090
rect 430 3038 502 3090
rect 554 3038 626 3090
rect 678 3038 750 3090
rect 802 3038 874 3090
rect 926 3038 998 3090
rect 1050 3038 1122 3090
rect 1174 3038 1246 3090
rect 1298 3038 1370 3090
rect 1422 3038 1494 3090
rect 1546 3038 1584 3090
rect 340 2966 1584 3038
rect 340 2914 378 2966
rect 430 2914 502 2966
rect 554 2914 626 2966
rect 678 2914 750 2966
rect 802 2914 874 2966
rect 926 2914 998 2966
rect 1050 2914 1122 2966
rect 1174 2914 1246 2966
rect 1298 2914 1370 2966
rect 1422 2914 1494 2966
rect 1546 2914 1584 2966
rect 340 2842 1584 2914
rect 340 2790 378 2842
rect 430 2790 502 2842
rect 554 2790 626 2842
rect 678 2790 750 2842
rect 802 2790 874 2842
rect 926 2790 998 2842
rect 1050 2790 1122 2842
rect 1174 2790 1246 2842
rect 1298 2790 1370 2842
rect 1422 2790 1494 2842
rect 1546 2790 1584 2842
rect 340 2718 1584 2790
rect 340 2666 378 2718
rect 430 2666 502 2718
rect 554 2666 626 2718
rect 678 2666 750 2718
rect 802 2666 874 2718
rect 926 2666 998 2718
rect 1050 2666 1122 2718
rect 1174 2666 1246 2718
rect 1298 2666 1370 2718
rect 1422 2666 1494 2718
rect 1546 2666 1584 2718
rect 340 2594 1584 2666
rect 340 2542 378 2594
rect 430 2542 502 2594
rect 554 2542 626 2594
rect 678 2542 750 2594
rect 802 2542 874 2594
rect 926 2542 998 2594
rect 1050 2542 1122 2594
rect 1174 2542 1246 2594
rect 1298 2542 1370 2594
rect 1422 2542 1494 2594
rect 1546 2542 1584 2594
rect 340 2470 1584 2542
rect 340 2418 378 2470
rect 430 2418 502 2470
rect 554 2418 626 2470
rect 678 2418 750 2470
rect 802 2418 874 2470
rect 926 2418 998 2470
rect 1050 2418 1122 2470
rect 1174 2418 1246 2470
rect 1298 2418 1370 2470
rect 1422 2418 1494 2470
rect 1546 2418 1584 2470
rect 340 2346 1584 2418
rect 340 2294 378 2346
rect 430 2294 502 2346
rect 554 2294 626 2346
rect 678 2294 750 2346
rect 802 2294 874 2346
rect 926 2294 998 2346
rect 1050 2294 1122 2346
rect 1174 2294 1246 2346
rect 1298 2294 1370 2346
rect 1422 2294 1494 2346
rect 1546 2294 1584 2346
rect 340 2222 1584 2294
rect 340 2170 378 2222
rect 430 2170 502 2222
rect 554 2170 626 2222
rect 678 2170 750 2222
rect 802 2170 874 2222
rect 926 2170 998 2222
rect 1050 2170 1122 2222
rect 1174 2170 1246 2222
rect 1298 2170 1370 2222
rect 1422 2170 1494 2222
rect 1546 2170 1584 2222
rect 340 2098 1584 2170
rect 340 2046 378 2098
rect 430 2046 502 2098
rect 554 2046 626 2098
rect 678 2046 750 2098
rect 802 2046 874 2098
rect 926 2046 998 2098
rect 1050 2046 1122 2098
rect 1174 2046 1246 2098
rect 1298 2046 1370 2098
rect 1422 2046 1494 2098
rect 1546 2046 1584 2098
rect 340 1974 1584 2046
rect 340 1922 378 1974
rect 430 1922 502 1974
rect 554 1922 626 1974
rect 678 1922 750 1974
rect 802 1922 874 1974
rect 926 1922 998 1974
rect 1050 1922 1122 1974
rect 1174 1922 1246 1974
rect 1298 1922 1370 1974
rect 1422 1922 1494 1974
rect 1546 1922 1584 1974
rect 340 1850 1584 1922
rect 340 1798 378 1850
rect 430 1798 502 1850
rect 554 1798 626 1850
rect 678 1798 750 1850
rect 802 1798 874 1850
rect 926 1798 998 1850
rect 1050 1798 1122 1850
rect 1174 1798 1246 1850
rect 1298 1798 1370 1850
rect 1422 1798 1494 1850
rect 1546 1798 1584 1850
rect 340 1726 1584 1798
rect 340 1674 378 1726
rect 430 1674 502 1726
rect 554 1674 626 1726
rect 678 1674 750 1726
rect 802 1674 874 1726
rect 926 1674 998 1726
rect 1050 1674 1122 1726
rect 1174 1674 1246 1726
rect 1298 1674 1370 1726
rect 1422 1674 1494 1726
rect 1546 1674 1584 1726
rect 340 1602 1584 1674
rect 340 1550 378 1602
rect 430 1550 502 1602
rect 554 1550 626 1602
rect 678 1550 750 1602
rect 802 1550 874 1602
rect 926 1550 998 1602
rect 1050 1550 1122 1602
rect 1174 1550 1246 1602
rect 1298 1550 1370 1602
rect 1422 1550 1494 1602
rect 1546 1550 1584 1602
rect 340 1478 1584 1550
rect 340 1426 378 1478
rect 430 1426 502 1478
rect 554 1426 626 1478
rect 678 1426 750 1478
rect 802 1426 874 1478
rect 926 1426 998 1478
rect 1050 1426 1122 1478
rect 1174 1426 1246 1478
rect 1298 1426 1370 1478
rect 1422 1426 1494 1478
rect 1546 1426 1584 1478
rect 340 1354 1584 1426
rect 340 1302 378 1354
rect 430 1302 502 1354
rect 554 1302 626 1354
rect 678 1302 750 1354
rect 802 1302 874 1354
rect 926 1302 998 1354
rect 1050 1302 1122 1354
rect 1174 1302 1246 1354
rect 1298 1302 1370 1354
rect 1422 1302 1494 1354
rect 1546 1302 1584 1354
rect 340 1230 1584 1302
rect 340 1178 378 1230
rect 430 1178 502 1230
rect 554 1178 626 1230
rect 678 1178 750 1230
rect 802 1178 874 1230
rect 926 1178 998 1230
rect 1050 1178 1122 1230
rect 1174 1178 1246 1230
rect 1298 1178 1370 1230
rect 1422 1178 1494 1230
rect 1546 1178 1584 1230
rect 340 1106 1584 1178
rect 340 1054 378 1106
rect 430 1054 502 1106
rect 554 1054 626 1106
rect 678 1054 750 1106
rect 802 1054 874 1106
rect 926 1054 998 1106
rect 1050 1054 1122 1106
rect 1174 1054 1246 1106
rect 1298 1054 1370 1106
rect 1422 1054 1494 1106
rect 1546 1054 1584 1106
rect 340 982 1584 1054
rect 340 930 378 982
rect 430 930 502 982
rect 554 930 626 982
rect 678 930 750 982
rect 802 930 874 982
rect 926 930 998 982
rect 1050 930 1122 982
rect 1174 930 1246 982
rect 1298 930 1370 982
rect 1422 930 1494 982
rect 1546 930 1584 982
rect 340 858 1584 930
rect 340 806 378 858
rect 430 806 502 858
rect 554 806 626 858
rect 678 806 750 858
rect 802 806 874 858
rect 926 806 998 858
rect 1050 806 1122 858
rect 1174 806 1246 858
rect 1298 806 1370 858
rect 1422 806 1494 858
rect 1546 806 1584 858
rect 340 734 1584 806
rect 340 682 378 734
rect 430 682 502 734
rect 554 682 626 734
rect 678 682 750 734
rect 802 682 874 734
rect 926 682 998 734
rect 1050 682 1122 734
rect 1174 682 1246 734
rect 1298 682 1370 734
rect 1422 682 1494 734
rect 1546 682 1584 734
rect 340 610 1584 682
rect 340 558 378 610
rect 430 558 502 610
rect 554 558 626 610
rect 678 558 750 610
rect 802 558 874 610
rect 926 558 998 610
rect 1050 558 1122 610
rect 1174 558 1246 610
rect 1298 558 1370 610
rect 1422 558 1494 610
rect 1546 558 1584 610
rect 340 486 1584 558
rect 340 434 378 486
rect 430 434 502 486
rect 554 434 626 486
rect 678 434 750 486
rect 802 434 874 486
rect 926 434 998 486
rect 1050 434 1122 486
rect 1174 434 1246 486
rect 1298 434 1370 486
rect 1422 434 1494 486
rect 1546 434 1584 486
rect 340 362 1584 434
rect 340 310 378 362
rect 430 310 502 362
rect 554 310 626 362
rect 678 310 750 362
rect 802 310 874 362
rect 926 310 998 362
rect 1050 310 1122 362
rect 1174 310 1246 362
rect 1298 310 1370 362
rect 1422 310 1494 362
rect 1546 310 1584 362
rect 340 238 1584 310
rect 340 186 378 238
rect 430 186 502 238
rect 554 186 626 238
rect 678 186 750 238
rect 802 186 874 238
rect 926 186 998 238
rect 1050 186 1122 238
rect 1174 186 1246 238
rect 1298 186 1370 238
rect 1422 186 1494 238
rect 1546 186 1584 238
rect 340 114 1584 186
rect 340 62 378 114
rect 430 62 502 114
rect 554 62 626 114
rect 678 62 750 114
rect 802 62 874 114
rect 926 62 998 114
rect 1050 62 1122 114
rect 1174 62 1246 114
rect 1298 62 1370 114
rect 1422 62 1494 114
rect 1546 62 1584 114
rect 340 0 1584 62
<< via1 >>
rect 0 7874 156 7926
rect 0 7750 156 7802
rect 0 7626 156 7678
rect 0 7502 156 7554
rect 0 7378 156 7430
rect 0 7254 156 7306
rect 0 7130 156 7182
rect 0 7006 156 7058
rect 0 6882 156 6934
rect 0 6758 156 6810
rect 0 6634 156 6686
rect 0 6510 156 6562
rect 0 6386 156 6438
rect 0 6262 156 6314
rect 0 6138 156 6190
rect 0 6014 156 6066
rect 0 5890 156 5942
rect 0 5766 156 5818
rect 0 5642 156 5694
rect 0 5518 156 5570
rect 0 5394 156 5446
rect 0 5270 156 5322
rect 0 5146 156 5198
rect 0 5022 156 5074
rect 0 4898 156 4950
rect 0 4774 156 4826
rect 0 4650 156 4702
rect 0 4526 156 4578
rect 0 4402 156 4454
rect 0 4278 156 4330
rect 0 4154 156 4206
rect 0 4030 156 4082
rect 0 3906 156 3958
rect 0 3782 156 3834
rect 0 3658 156 3710
rect 0 3534 156 3586
rect 0 3410 156 3462
rect 0 3286 156 3338
rect 0 3162 156 3214
rect 0 3038 156 3090
rect 0 2914 156 2966
rect 0 2790 156 2842
rect 0 2666 156 2718
rect 0 2542 156 2594
rect 0 2418 156 2470
rect 0 2294 156 2346
rect 0 2170 156 2222
rect 0 2046 156 2098
rect 0 1922 156 1974
rect 0 1798 156 1850
rect 0 1674 156 1726
rect 0 1550 156 1602
rect 0 1426 156 1478
rect 0 1302 156 1354
rect 0 1178 156 1230
rect 0 1054 156 1106
rect 0 930 156 982
rect 0 806 156 858
rect 0 682 156 734
rect 0 558 156 610
rect 0 434 156 486
rect 0 310 156 362
rect 0 186 156 238
rect 0 62 156 114
rect 378 7874 430 7926
rect 502 7874 554 7926
rect 626 7874 678 7926
rect 750 7874 802 7926
rect 874 7874 926 7926
rect 998 7874 1050 7926
rect 1122 7874 1174 7926
rect 1246 7874 1298 7926
rect 1370 7874 1422 7926
rect 1494 7874 1546 7926
rect 378 7750 430 7802
rect 502 7750 554 7802
rect 626 7750 678 7802
rect 750 7750 802 7802
rect 874 7750 926 7802
rect 998 7750 1050 7802
rect 1122 7750 1174 7802
rect 1246 7750 1298 7802
rect 1370 7750 1422 7802
rect 1494 7750 1546 7802
rect 378 7626 430 7678
rect 502 7626 554 7678
rect 626 7626 678 7678
rect 750 7626 802 7678
rect 874 7626 926 7678
rect 998 7626 1050 7678
rect 1122 7626 1174 7678
rect 1246 7626 1298 7678
rect 1370 7626 1422 7678
rect 1494 7626 1546 7678
rect 378 7502 430 7554
rect 502 7502 554 7554
rect 626 7502 678 7554
rect 750 7502 802 7554
rect 874 7502 926 7554
rect 998 7502 1050 7554
rect 1122 7502 1174 7554
rect 1246 7502 1298 7554
rect 1370 7502 1422 7554
rect 1494 7502 1546 7554
rect 378 7378 430 7430
rect 502 7378 554 7430
rect 626 7378 678 7430
rect 750 7378 802 7430
rect 874 7378 926 7430
rect 998 7378 1050 7430
rect 1122 7378 1174 7430
rect 1246 7378 1298 7430
rect 1370 7378 1422 7430
rect 1494 7378 1546 7430
rect 378 7254 430 7306
rect 502 7254 554 7306
rect 626 7254 678 7306
rect 750 7254 802 7306
rect 874 7254 926 7306
rect 998 7254 1050 7306
rect 1122 7254 1174 7306
rect 1246 7254 1298 7306
rect 1370 7254 1422 7306
rect 1494 7254 1546 7306
rect 378 7130 430 7182
rect 502 7130 554 7182
rect 626 7130 678 7182
rect 750 7130 802 7182
rect 874 7130 926 7182
rect 998 7130 1050 7182
rect 1122 7130 1174 7182
rect 1246 7130 1298 7182
rect 1370 7130 1422 7182
rect 1494 7130 1546 7182
rect 378 7006 430 7058
rect 502 7006 554 7058
rect 626 7006 678 7058
rect 750 7006 802 7058
rect 874 7006 926 7058
rect 998 7006 1050 7058
rect 1122 7006 1174 7058
rect 1246 7006 1298 7058
rect 1370 7006 1422 7058
rect 1494 7006 1546 7058
rect 378 6882 430 6934
rect 502 6882 554 6934
rect 626 6882 678 6934
rect 750 6882 802 6934
rect 874 6882 926 6934
rect 998 6882 1050 6934
rect 1122 6882 1174 6934
rect 1246 6882 1298 6934
rect 1370 6882 1422 6934
rect 1494 6882 1546 6934
rect 378 6758 430 6810
rect 502 6758 554 6810
rect 626 6758 678 6810
rect 750 6758 802 6810
rect 874 6758 926 6810
rect 998 6758 1050 6810
rect 1122 6758 1174 6810
rect 1246 6758 1298 6810
rect 1370 6758 1422 6810
rect 1494 6758 1546 6810
rect 378 6634 430 6686
rect 502 6634 554 6686
rect 626 6634 678 6686
rect 750 6634 802 6686
rect 874 6634 926 6686
rect 998 6634 1050 6686
rect 1122 6634 1174 6686
rect 1246 6634 1298 6686
rect 1370 6634 1422 6686
rect 1494 6634 1546 6686
rect 378 6510 430 6562
rect 502 6510 554 6562
rect 626 6510 678 6562
rect 750 6510 802 6562
rect 874 6510 926 6562
rect 998 6510 1050 6562
rect 1122 6510 1174 6562
rect 1246 6510 1298 6562
rect 1370 6510 1422 6562
rect 1494 6510 1546 6562
rect 378 6386 430 6438
rect 502 6386 554 6438
rect 626 6386 678 6438
rect 750 6386 802 6438
rect 874 6386 926 6438
rect 998 6386 1050 6438
rect 1122 6386 1174 6438
rect 1246 6386 1298 6438
rect 1370 6386 1422 6438
rect 1494 6386 1546 6438
rect 378 6262 430 6314
rect 502 6262 554 6314
rect 626 6262 678 6314
rect 750 6262 802 6314
rect 874 6262 926 6314
rect 998 6262 1050 6314
rect 1122 6262 1174 6314
rect 1246 6262 1298 6314
rect 1370 6262 1422 6314
rect 1494 6262 1546 6314
rect 378 6138 430 6190
rect 502 6138 554 6190
rect 626 6138 678 6190
rect 750 6138 802 6190
rect 874 6138 926 6190
rect 998 6138 1050 6190
rect 1122 6138 1174 6190
rect 1246 6138 1298 6190
rect 1370 6138 1422 6190
rect 1494 6138 1546 6190
rect 378 6014 430 6066
rect 502 6014 554 6066
rect 626 6014 678 6066
rect 750 6014 802 6066
rect 874 6014 926 6066
rect 998 6014 1050 6066
rect 1122 6014 1174 6066
rect 1246 6014 1298 6066
rect 1370 6014 1422 6066
rect 1494 6014 1546 6066
rect 378 5890 430 5942
rect 502 5890 554 5942
rect 626 5890 678 5942
rect 750 5890 802 5942
rect 874 5890 926 5942
rect 998 5890 1050 5942
rect 1122 5890 1174 5942
rect 1246 5890 1298 5942
rect 1370 5890 1422 5942
rect 1494 5890 1546 5942
rect 378 5766 430 5818
rect 502 5766 554 5818
rect 626 5766 678 5818
rect 750 5766 802 5818
rect 874 5766 926 5818
rect 998 5766 1050 5818
rect 1122 5766 1174 5818
rect 1246 5766 1298 5818
rect 1370 5766 1422 5818
rect 1494 5766 1546 5818
rect 378 5642 430 5694
rect 502 5642 554 5694
rect 626 5642 678 5694
rect 750 5642 802 5694
rect 874 5642 926 5694
rect 998 5642 1050 5694
rect 1122 5642 1174 5694
rect 1246 5642 1298 5694
rect 1370 5642 1422 5694
rect 1494 5642 1546 5694
rect 378 5518 430 5570
rect 502 5518 554 5570
rect 626 5518 678 5570
rect 750 5518 802 5570
rect 874 5518 926 5570
rect 998 5518 1050 5570
rect 1122 5518 1174 5570
rect 1246 5518 1298 5570
rect 1370 5518 1422 5570
rect 1494 5518 1546 5570
rect 378 5394 430 5446
rect 502 5394 554 5446
rect 626 5394 678 5446
rect 750 5394 802 5446
rect 874 5394 926 5446
rect 998 5394 1050 5446
rect 1122 5394 1174 5446
rect 1246 5394 1298 5446
rect 1370 5394 1422 5446
rect 1494 5394 1546 5446
rect 378 5270 430 5322
rect 502 5270 554 5322
rect 626 5270 678 5322
rect 750 5270 802 5322
rect 874 5270 926 5322
rect 998 5270 1050 5322
rect 1122 5270 1174 5322
rect 1246 5270 1298 5322
rect 1370 5270 1422 5322
rect 1494 5270 1546 5322
rect 378 5146 430 5198
rect 502 5146 554 5198
rect 626 5146 678 5198
rect 750 5146 802 5198
rect 874 5146 926 5198
rect 998 5146 1050 5198
rect 1122 5146 1174 5198
rect 1246 5146 1298 5198
rect 1370 5146 1422 5198
rect 1494 5146 1546 5198
rect 378 5022 430 5074
rect 502 5022 554 5074
rect 626 5022 678 5074
rect 750 5022 802 5074
rect 874 5022 926 5074
rect 998 5022 1050 5074
rect 1122 5022 1174 5074
rect 1246 5022 1298 5074
rect 1370 5022 1422 5074
rect 1494 5022 1546 5074
rect 378 4898 430 4950
rect 502 4898 554 4950
rect 626 4898 678 4950
rect 750 4898 802 4950
rect 874 4898 926 4950
rect 998 4898 1050 4950
rect 1122 4898 1174 4950
rect 1246 4898 1298 4950
rect 1370 4898 1422 4950
rect 1494 4898 1546 4950
rect 378 4774 430 4826
rect 502 4774 554 4826
rect 626 4774 678 4826
rect 750 4774 802 4826
rect 874 4774 926 4826
rect 998 4774 1050 4826
rect 1122 4774 1174 4826
rect 1246 4774 1298 4826
rect 1370 4774 1422 4826
rect 1494 4774 1546 4826
rect 378 4650 430 4702
rect 502 4650 554 4702
rect 626 4650 678 4702
rect 750 4650 802 4702
rect 874 4650 926 4702
rect 998 4650 1050 4702
rect 1122 4650 1174 4702
rect 1246 4650 1298 4702
rect 1370 4650 1422 4702
rect 1494 4650 1546 4702
rect 378 4526 430 4578
rect 502 4526 554 4578
rect 626 4526 678 4578
rect 750 4526 802 4578
rect 874 4526 926 4578
rect 998 4526 1050 4578
rect 1122 4526 1174 4578
rect 1246 4526 1298 4578
rect 1370 4526 1422 4578
rect 1494 4526 1546 4578
rect 378 4402 430 4454
rect 502 4402 554 4454
rect 626 4402 678 4454
rect 750 4402 802 4454
rect 874 4402 926 4454
rect 998 4402 1050 4454
rect 1122 4402 1174 4454
rect 1246 4402 1298 4454
rect 1370 4402 1422 4454
rect 1494 4402 1546 4454
rect 378 4278 430 4330
rect 502 4278 554 4330
rect 626 4278 678 4330
rect 750 4278 802 4330
rect 874 4278 926 4330
rect 998 4278 1050 4330
rect 1122 4278 1174 4330
rect 1246 4278 1298 4330
rect 1370 4278 1422 4330
rect 1494 4278 1546 4330
rect 378 4154 430 4206
rect 502 4154 554 4206
rect 626 4154 678 4206
rect 750 4154 802 4206
rect 874 4154 926 4206
rect 998 4154 1050 4206
rect 1122 4154 1174 4206
rect 1246 4154 1298 4206
rect 1370 4154 1422 4206
rect 1494 4154 1546 4206
rect 378 4030 430 4082
rect 502 4030 554 4082
rect 626 4030 678 4082
rect 750 4030 802 4082
rect 874 4030 926 4082
rect 998 4030 1050 4082
rect 1122 4030 1174 4082
rect 1246 4030 1298 4082
rect 1370 4030 1422 4082
rect 1494 4030 1546 4082
rect 378 3906 430 3958
rect 502 3906 554 3958
rect 626 3906 678 3958
rect 750 3906 802 3958
rect 874 3906 926 3958
rect 998 3906 1050 3958
rect 1122 3906 1174 3958
rect 1246 3906 1298 3958
rect 1370 3906 1422 3958
rect 1494 3906 1546 3958
rect 378 3782 430 3834
rect 502 3782 554 3834
rect 626 3782 678 3834
rect 750 3782 802 3834
rect 874 3782 926 3834
rect 998 3782 1050 3834
rect 1122 3782 1174 3834
rect 1246 3782 1298 3834
rect 1370 3782 1422 3834
rect 1494 3782 1546 3834
rect 378 3658 430 3710
rect 502 3658 554 3710
rect 626 3658 678 3710
rect 750 3658 802 3710
rect 874 3658 926 3710
rect 998 3658 1050 3710
rect 1122 3658 1174 3710
rect 1246 3658 1298 3710
rect 1370 3658 1422 3710
rect 1494 3658 1546 3710
rect 378 3534 430 3586
rect 502 3534 554 3586
rect 626 3534 678 3586
rect 750 3534 802 3586
rect 874 3534 926 3586
rect 998 3534 1050 3586
rect 1122 3534 1174 3586
rect 1246 3534 1298 3586
rect 1370 3534 1422 3586
rect 1494 3534 1546 3586
rect 378 3410 430 3462
rect 502 3410 554 3462
rect 626 3410 678 3462
rect 750 3410 802 3462
rect 874 3410 926 3462
rect 998 3410 1050 3462
rect 1122 3410 1174 3462
rect 1246 3410 1298 3462
rect 1370 3410 1422 3462
rect 1494 3410 1546 3462
rect 378 3286 430 3338
rect 502 3286 554 3338
rect 626 3286 678 3338
rect 750 3286 802 3338
rect 874 3286 926 3338
rect 998 3286 1050 3338
rect 1122 3286 1174 3338
rect 1246 3286 1298 3338
rect 1370 3286 1422 3338
rect 1494 3286 1546 3338
rect 378 3162 430 3214
rect 502 3162 554 3214
rect 626 3162 678 3214
rect 750 3162 802 3214
rect 874 3162 926 3214
rect 998 3162 1050 3214
rect 1122 3162 1174 3214
rect 1246 3162 1298 3214
rect 1370 3162 1422 3214
rect 1494 3162 1546 3214
rect 378 3038 430 3090
rect 502 3038 554 3090
rect 626 3038 678 3090
rect 750 3038 802 3090
rect 874 3038 926 3090
rect 998 3038 1050 3090
rect 1122 3038 1174 3090
rect 1246 3038 1298 3090
rect 1370 3038 1422 3090
rect 1494 3038 1546 3090
rect 378 2914 430 2966
rect 502 2914 554 2966
rect 626 2914 678 2966
rect 750 2914 802 2966
rect 874 2914 926 2966
rect 998 2914 1050 2966
rect 1122 2914 1174 2966
rect 1246 2914 1298 2966
rect 1370 2914 1422 2966
rect 1494 2914 1546 2966
rect 378 2790 430 2842
rect 502 2790 554 2842
rect 626 2790 678 2842
rect 750 2790 802 2842
rect 874 2790 926 2842
rect 998 2790 1050 2842
rect 1122 2790 1174 2842
rect 1246 2790 1298 2842
rect 1370 2790 1422 2842
rect 1494 2790 1546 2842
rect 378 2666 430 2718
rect 502 2666 554 2718
rect 626 2666 678 2718
rect 750 2666 802 2718
rect 874 2666 926 2718
rect 998 2666 1050 2718
rect 1122 2666 1174 2718
rect 1246 2666 1298 2718
rect 1370 2666 1422 2718
rect 1494 2666 1546 2718
rect 378 2542 430 2594
rect 502 2542 554 2594
rect 626 2542 678 2594
rect 750 2542 802 2594
rect 874 2542 926 2594
rect 998 2542 1050 2594
rect 1122 2542 1174 2594
rect 1246 2542 1298 2594
rect 1370 2542 1422 2594
rect 1494 2542 1546 2594
rect 378 2418 430 2470
rect 502 2418 554 2470
rect 626 2418 678 2470
rect 750 2418 802 2470
rect 874 2418 926 2470
rect 998 2418 1050 2470
rect 1122 2418 1174 2470
rect 1246 2418 1298 2470
rect 1370 2418 1422 2470
rect 1494 2418 1546 2470
rect 378 2294 430 2346
rect 502 2294 554 2346
rect 626 2294 678 2346
rect 750 2294 802 2346
rect 874 2294 926 2346
rect 998 2294 1050 2346
rect 1122 2294 1174 2346
rect 1246 2294 1298 2346
rect 1370 2294 1422 2346
rect 1494 2294 1546 2346
rect 378 2170 430 2222
rect 502 2170 554 2222
rect 626 2170 678 2222
rect 750 2170 802 2222
rect 874 2170 926 2222
rect 998 2170 1050 2222
rect 1122 2170 1174 2222
rect 1246 2170 1298 2222
rect 1370 2170 1422 2222
rect 1494 2170 1546 2222
rect 378 2046 430 2098
rect 502 2046 554 2098
rect 626 2046 678 2098
rect 750 2046 802 2098
rect 874 2046 926 2098
rect 998 2046 1050 2098
rect 1122 2046 1174 2098
rect 1246 2046 1298 2098
rect 1370 2046 1422 2098
rect 1494 2046 1546 2098
rect 378 1922 430 1974
rect 502 1922 554 1974
rect 626 1922 678 1974
rect 750 1922 802 1974
rect 874 1922 926 1974
rect 998 1922 1050 1974
rect 1122 1922 1174 1974
rect 1246 1922 1298 1974
rect 1370 1922 1422 1974
rect 1494 1922 1546 1974
rect 378 1798 430 1850
rect 502 1798 554 1850
rect 626 1798 678 1850
rect 750 1798 802 1850
rect 874 1798 926 1850
rect 998 1798 1050 1850
rect 1122 1798 1174 1850
rect 1246 1798 1298 1850
rect 1370 1798 1422 1850
rect 1494 1798 1546 1850
rect 378 1674 430 1726
rect 502 1674 554 1726
rect 626 1674 678 1726
rect 750 1674 802 1726
rect 874 1674 926 1726
rect 998 1674 1050 1726
rect 1122 1674 1174 1726
rect 1246 1674 1298 1726
rect 1370 1674 1422 1726
rect 1494 1674 1546 1726
rect 378 1550 430 1602
rect 502 1550 554 1602
rect 626 1550 678 1602
rect 750 1550 802 1602
rect 874 1550 926 1602
rect 998 1550 1050 1602
rect 1122 1550 1174 1602
rect 1246 1550 1298 1602
rect 1370 1550 1422 1602
rect 1494 1550 1546 1602
rect 378 1426 430 1478
rect 502 1426 554 1478
rect 626 1426 678 1478
rect 750 1426 802 1478
rect 874 1426 926 1478
rect 998 1426 1050 1478
rect 1122 1426 1174 1478
rect 1246 1426 1298 1478
rect 1370 1426 1422 1478
rect 1494 1426 1546 1478
rect 378 1302 430 1354
rect 502 1302 554 1354
rect 626 1302 678 1354
rect 750 1302 802 1354
rect 874 1302 926 1354
rect 998 1302 1050 1354
rect 1122 1302 1174 1354
rect 1246 1302 1298 1354
rect 1370 1302 1422 1354
rect 1494 1302 1546 1354
rect 378 1178 430 1230
rect 502 1178 554 1230
rect 626 1178 678 1230
rect 750 1178 802 1230
rect 874 1178 926 1230
rect 998 1178 1050 1230
rect 1122 1178 1174 1230
rect 1246 1178 1298 1230
rect 1370 1178 1422 1230
rect 1494 1178 1546 1230
rect 378 1054 430 1106
rect 502 1054 554 1106
rect 626 1054 678 1106
rect 750 1054 802 1106
rect 874 1054 926 1106
rect 998 1054 1050 1106
rect 1122 1054 1174 1106
rect 1246 1054 1298 1106
rect 1370 1054 1422 1106
rect 1494 1054 1546 1106
rect 378 930 430 982
rect 502 930 554 982
rect 626 930 678 982
rect 750 930 802 982
rect 874 930 926 982
rect 998 930 1050 982
rect 1122 930 1174 982
rect 1246 930 1298 982
rect 1370 930 1422 982
rect 1494 930 1546 982
rect 378 806 430 858
rect 502 806 554 858
rect 626 806 678 858
rect 750 806 802 858
rect 874 806 926 858
rect 998 806 1050 858
rect 1122 806 1174 858
rect 1246 806 1298 858
rect 1370 806 1422 858
rect 1494 806 1546 858
rect 378 682 430 734
rect 502 682 554 734
rect 626 682 678 734
rect 750 682 802 734
rect 874 682 926 734
rect 998 682 1050 734
rect 1122 682 1174 734
rect 1246 682 1298 734
rect 1370 682 1422 734
rect 1494 682 1546 734
rect 378 558 430 610
rect 502 558 554 610
rect 626 558 678 610
rect 750 558 802 610
rect 874 558 926 610
rect 998 558 1050 610
rect 1122 558 1174 610
rect 1246 558 1298 610
rect 1370 558 1422 610
rect 1494 558 1546 610
rect 378 434 430 486
rect 502 434 554 486
rect 626 434 678 486
rect 750 434 802 486
rect 874 434 926 486
rect 998 434 1050 486
rect 1122 434 1174 486
rect 1246 434 1298 486
rect 1370 434 1422 486
rect 1494 434 1546 486
rect 378 310 430 362
rect 502 310 554 362
rect 626 310 678 362
rect 750 310 802 362
rect 874 310 926 362
rect 998 310 1050 362
rect 1122 310 1174 362
rect 1246 310 1298 362
rect 1370 310 1422 362
rect 1494 310 1546 362
rect 378 186 430 238
rect 502 186 554 238
rect 626 186 678 238
rect 750 186 802 238
rect 874 186 926 238
rect 998 186 1050 238
rect 1122 186 1174 238
rect 1246 186 1298 238
rect 1370 186 1422 238
rect 1494 186 1546 238
rect 378 62 430 114
rect 502 62 554 114
rect 626 62 678 114
rect 750 62 802 114
rect 874 62 926 114
rect 998 62 1050 114
rect 1122 62 1174 114
rect 1246 62 1298 114
rect 1370 62 1422 114
rect 1494 62 1546 114
<< metal2 >>
rect -44 7926 200 8000
rect -44 7915 0 7926
rect 156 7915 200 7926
rect -44 7859 -21 7915
rect 35 7859 121 7874
rect 177 7859 200 7915
rect -44 7802 200 7859
rect -44 7773 0 7802
rect 156 7773 200 7802
rect -44 7717 -21 7773
rect 35 7717 121 7750
rect 177 7717 200 7773
rect -44 7678 200 7717
rect -44 7631 0 7678
rect 156 7631 200 7678
rect -44 7575 -21 7631
rect 35 7575 121 7626
rect 177 7575 200 7631
rect -44 7554 200 7575
rect -44 7502 0 7554
rect 156 7502 200 7554
rect -44 7489 200 7502
rect -44 7433 -21 7489
rect 35 7433 121 7489
rect 177 7433 200 7489
rect -44 7430 200 7433
rect -44 7378 0 7430
rect 156 7378 200 7430
rect -44 7347 200 7378
rect -44 7291 -21 7347
rect 35 7306 121 7347
rect 177 7291 200 7347
rect -44 7254 0 7291
rect 156 7254 200 7291
rect -44 7182 200 7254
rect -44 7130 0 7182
rect 156 7130 200 7182
rect -44 7058 200 7130
rect -44 7006 0 7058
rect 156 7006 200 7058
rect -44 6950 200 7006
rect -44 6894 -21 6950
rect 35 6934 121 6950
rect 177 6894 200 6950
rect -44 6882 0 6894
rect 156 6882 200 6894
rect -44 6810 200 6882
rect -44 6808 0 6810
rect 156 6808 200 6810
rect -44 6752 -21 6808
rect 35 6752 121 6758
rect 177 6752 200 6808
rect -44 6686 200 6752
rect -44 6666 0 6686
rect 156 6666 200 6686
rect -44 6610 -21 6666
rect 35 6610 121 6634
rect 177 6610 200 6666
rect -44 6562 200 6610
rect -44 6524 0 6562
rect 156 6524 200 6562
rect -44 6468 -21 6524
rect 35 6468 121 6510
rect 177 6468 200 6524
rect -44 6438 200 6468
rect -44 6386 0 6438
rect 156 6386 200 6438
rect -44 6382 200 6386
rect -44 6326 -21 6382
rect 35 6326 121 6382
rect 177 6326 200 6382
rect -44 6314 200 6326
rect -44 6262 0 6314
rect 156 6262 200 6314
rect -44 6240 200 6262
rect -44 6184 -21 6240
rect 35 6190 121 6240
rect 177 6184 200 6240
rect -44 6138 0 6184
rect 156 6138 200 6184
rect -44 6098 200 6138
rect -44 6042 -21 6098
rect 35 6066 121 6098
rect 177 6042 200 6098
rect -44 6014 0 6042
rect 156 6014 200 6042
rect -44 5956 200 6014
rect -44 5900 -21 5956
rect 35 5942 121 5956
rect 177 5900 200 5956
rect -44 5890 0 5900
rect 156 5890 200 5900
rect -44 5818 200 5890
rect -44 5814 0 5818
rect 156 5814 200 5818
rect -44 5758 -21 5814
rect 35 5758 121 5766
rect 177 5758 200 5814
rect -44 5694 200 5758
rect -44 5672 0 5694
rect 156 5672 200 5694
rect -44 5616 -21 5672
rect 35 5616 121 5642
rect 177 5616 200 5672
rect -44 5570 200 5616
rect -44 5530 0 5570
rect 156 5530 200 5570
rect -44 5474 -21 5530
rect 35 5474 121 5518
rect 177 5474 200 5530
rect -44 5446 200 5474
rect -44 5394 0 5446
rect 156 5394 200 5446
rect -44 5388 200 5394
rect -44 5332 -21 5388
rect 35 5332 121 5388
rect 177 5332 200 5388
rect -44 5322 200 5332
rect -44 5270 0 5322
rect 156 5270 200 5322
rect -44 5246 200 5270
rect -44 5190 -21 5246
rect 35 5198 121 5246
rect 177 5190 200 5246
rect -44 5146 0 5190
rect 156 5146 200 5190
rect -44 5104 200 5146
rect -44 5048 -21 5104
rect 35 5074 121 5104
rect 177 5048 200 5104
rect -44 5022 0 5048
rect 156 5022 200 5048
rect -44 4962 200 5022
rect -44 4906 -21 4962
rect 35 4950 121 4962
rect 177 4906 200 4962
rect -44 4898 0 4906
rect 156 4898 200 4906
rect -44 4826 200 4898
rect -44 4820 0 4826
rect 156 4820 200 4826
rect -44 4764 -21 4820
rect 35 4764 121 4774
rect 177 4764 200 4820
rect -44 4702 200 4764
rect -44 4678 0 4702
rect 156 4678 200 4702
rect -44 4622 -21 4678
rect 35 4622 121 4650
rect 177 4622 200 4678
rect -44 4578 200 4622
rect -44 4536 0 4578
rect 156 4536 200 4578
rect -44 4480 -21 4536
rect 35 4480 121 4526
rect 177 4480 200 4536
rect -44 4454 200 4480
rect -44 4402 0 4454
rect 156 4402 200 4454
rect -44 4394 200 4402
rect -44 4338 -21 4394
rect 35 4338 121 4394
rect 177 4338 200 4394
rect -44 4330 200 4338
rect -44 4278 0 4330
rect 156 4278 200 4330
rect -44 4252 200 4278
rect -44 4196 -21 4252
rect 35 4206 121 4252
rect 177 4196 200 4252
rect -44 4154 0 4196
rect 156 4154 200 4196
rect -44 4110 200 4154
rect -44 4054 -21 4110
rect 35 4082 121 4110
rect 177 4054 200 4110
rect -44 4030 0 4054
rect 156 4030 200 4054
rect -44 3958 200 4030
rect -44 3906 0 3958
rect 156 3906 200 3958
rect -44 3834 200 3906
rect -44 3782 0 3834
rect 156 3782 200 3834
rect -44 3763 200 3782
rect -44 3707 -21 3763
rect 35 3710 121 3763
rect 177 3707 200 3763
rect -44 3658 0 3707
rect 156 3658 200 3707
rect -44 3621 200 3658
rect -44 3565 -21 3621
rect 35 3586 121 3621
rect 177 3565 200 3621
rect -44 3534 0 3565
rect 156 3534 200 3565
rect -44 3479 200 3534
rect -44 3423 -21 3479
rect 35 3462 121 3479
rect 177 3423 200 3479
rect -44 3410 0 3423
rect 156 3410 200 3423
rect -44 3338 200 3410
rect -44 3337 0 3338
rect 156 3337 200 3338
rect -44 3281 -21 3337
rect 35 3281 121 3286
rect 177 3281 200 3337
rect -44 3214 200 3281
rect -44 3195 0 3214
rect 156 3195 200 3214
rect -44 3139 -21 3195
rect 35 3139 121 3162
rect 177 3139 200 3195
rect -44 3090 200 3139
rect -44 3053 0 3090
rect 156 3053 200 3090
rect -44 2997 -21 3053
rect 35 2997 121 3038
rect 177 2997 200 3053
rect -44 2966 200 2997
rect -44 2914 0 2966
rect 156 2914 200 2966
rect -44 2911 200 2914
rect -44 2855 -21 2911
rect 35 2855 121 2911
rect 177 2855 200 2911
rect -44 2842 200 2855
rect -44 2790 0 2842
rect 156 2790 200 2842
rect -44 2769 200 2790
rect -44 2713 -21 2769
rect 35 2718 121 2769
rect 177 2713 200 2769
rect -44 2666 0 2713
rect 156 2666 200 2713
rect -44 2627 200 2666
rect -44 2571 -21 2627
rect 35 2594 121 2627
rect 177 2571 200 2627
rect -44 2542 0 2571
rect 156 2542 200 2571
rect -44 2485 200 2542
rect -44 2429 -21 2485
rect 35 2470 121 2485
rect 177 2429 200 2485
rect -44 2418 0 2429
rect 156 2418 200 2429
rect -44 2346 200 2418
rect -44 2343 0 2346
rect 156 2343 200 2346
rect -44 2287 -21 2343
rect 35 2287 121 2294
rect 177 2287 200 2343
rect -44 2222 200 2287
rect -44 2201 0 2222
rect 156 2201 200 2222
rect -44 2145 -21 2201
rect 35 2145 121 2170
rect 177 2145 200 2201
rect -44 2098 200 2145
rect -44 2059 0 2098
rect 156 2059 200 2098
rect -44 2003 -21 2059
rect 35 2003 121 2046
rect 177 2003 200 2059
rect -44 1974 200 2003
rect -44 1922 0 1974
rect 156 1922 200 1974
rect -44 1917 200 1922
rect -44 1861 -21 1917
rect 35 1861 121 1917
rect 177 1861 200 1917
rect -44 1850 200 1861
rect -44 1798 0 1850
rect 156 1798 200 1850
rect -44 1775 200 1798
rect -44 1719 -21 1775
rect 35 1726 121 1775
rect 177 1719 200 1775
rect -44 1674 0 1719
rect 156 1674 200 1719
rect -44 1633 200 1674
rect -44 1577 -21 1633
rect 35 1602 121 1633
rect 177 1577 200 1633
rect -44 1550 0 1577
rect 156 1550 200 1577
rect -44 1491 200 1550
rect -44 1435 -21 1491
rect 35 1478 121 1491
rect 177 1435 200 1491
rect -44 1426 0 1435
rect 156 1426 200 1435
rect -44 1354 200 1426
rect -44 1349 0 1354
rect 156 1349 200 1354
rect -44 1293 -21 1349
rect 35 1293 121 1302
rect 177 1293 200 1349
rect -44 1230 200 1293
rect -44 1207 0 1230
rect 156 1207 200 1230
rect -44 1151 -21 1207
rect 35 1151 121 1178
rect 177 1151 200 1207
rect -44 1106 200 1151
rect -44 1065 0 1106
rect 156 1065 200 1106
rect -44 1009 -21 1065
rect 35 1009 121 1054
rect 177 1009 200 1065
rect -44 982 200 1009
rect -44 930 0 982
rect 156 930 200 982
rect -44 923 200 930
rect -44 867 -21 923
rect 35 867 121 923
rect 177 867 200 923
rect -44 858 200 867
rect -44 806 0 858
rect 156 806 200 858
rect -44 734 200 806
rect -44 682 0 734
rect 156 682 200 734
rect -44 610 200 682
rect -44 558 0 610
rect 156 558 200 610
rect -44 550 200 558
rect -44 494 -21 550
rect 35 494 121 550
rect 177 494 200 550
rect -44 486 200 494
rect -44 434 0 486
rect 156 434 200 486
rect -44 408 200 434
rect -44 352 -21 408
rect 35 362 121 408
rect 177 352 200 408
rect -44 310 0 352
rect 156 310 200 352
rect -44 266 200 310
rect -44 210 -21 266
rect 35 238 121 266
rect 177 210 200 266
rect -44 186 0 210
rect 156 186 200 210
rect -44 124 200 186
rect -44 68 -21 124
rect 35 114 121 124
rect 177 68 200 124
rect -44 62 0 68
rect 156 62 200 68
rect -44 0 200 62
rect 340 7926 1584 8000
rect 340 7874 378 7926
rect 430 7874 502 7926
rect 554 7874 626 7926
rect 678 7874 750 7926
rect 802 7874 874 7926
rect 926 7874 998 7926
rect 1050 7874 1122 7926
rect 1174 7874 1246 7926
rect 1298 7874 1370 7926
rect 1422 7874 1494 7926
rect 1546 7874 1584 7926
rect 340 7802 1584 7874
rect 340 7750 378 7802
rect 430 7750 502 7802
rect 554 7750 626 7802
rect 678 7750 750 7802
rect 802 7750 874 7802
rect 926 7750 998 7802
rect 1050 7750 1122 7802
rect 1174 7750 1246 7802
rect 1298 7750 1370 7802
rect 1422 7750 1494 7802
rect 1546 7750 1584 7802
rect 340 7678 1584 7750
rect 340 7626 378 7678
rect 430 7626 502 7678
rect 554 7626 626 7678
rect 678 7626 750 7678
rect 802 7626 874 7678
rect 926 7626 998 7678
rect 1050 7626 1122 7678
rect 1174 7626 1246 7678
rect 1298 7626 1370 7678
rect 1422 7626 1494 7678
rect 1546 7626 1584 7678
rect 340 7554 1584 7626
rect 340 7502 378 7554
rect 430 7502 502 7554
rect 554 7502 626 7554
rect 678 7502 750 7554
rect 802 7502 874 7554
rect 926 7502 998 7554
rect 1050 7502 1122 7554
rect 1174 7502 1246 7554
rect 1298 7502 1370 7554
rect 1422 7502 1494 7554
rect 1546 7502 1584 7554
rect 340 7430 1584 7502
rect 340 7378 378 7430
rect 430 7378 502 7430
rect 554 7378 626 7430
rect 678 7378 750 7430
rect 802 7378 874 7430
rect 926 7378 998 7430
rect 1050 7378 1122 7430
rect 1174 7378 1246 7430
rect 1298 7378 1370 7430
rect 1422 7378 1494 7430
rect 1546 7378 1584 7430
rect 340 7306 1584 7378
rect 340 7254 378 7306
rect 430 7254 502 7306
rect 554 7254 626 7306
rect 678 7254 750 7306
rect 802 7254 874 7306
rect 926 7254 998 7306
rect 1050 7254 1122 7306
rect 1174 7254 1246 7306
rect 1298 7254 1370 7306
rect 1422 7254 1494 7306
rect 1546 7254 1584 7306
rect 340 7182 1584 7254
rect 340 7130 378 7182
rect 430 7130 502 7182
rect 554 7130 626 7182
rect 678 7130 750 7182
rect 802 7130 874 7182
rect 926 7130 998 7182
rect 1050 7130 1122 7182
rect 1174 7130 1246 7182
rect 1298 7130 1370 7182
rect 1422 7130 1494 7182
rect 1546 7130 1584 7182
rect 340 7058 1584 7130
rect 340 7006 378 7058
rect 430 7006 502 7058
rect 554 7006 626 7058
rect 678 7006 750 7058
rect 802 7006 874 7058
rect 926 7006 998 7058
rect 1050 7006 1122 7058
rect 1174 7006 1246 7058
rect 1298 7006 1370 7058
rect 1422 7006 1494 7058
rect 1546 7006 1584 7058
rect 340 6934 1584 7006
rect 340 6882 378 6934
rect 430 6882 502 6934
rect 554 6882 626 6934
rect 678 6882 750 6934
rect 802 6882 874 6934
rect 926 6882 998 6934
rect 1050 6882 1122 6934
rect 1174 6882 1246 6934
rect 1298 6882 1370 6934
rect 1422 6882 1494 6934
rect 1546 6882 1584 6934
rect 340 6810 1584 6882
rect 340 6758 378 6810
rect 430 6758 502 6810
rect 554 6758 626 6810
rect 678 6758 750 6810
rect 802 6758 874 6810
rect 926 6758 998 6810
rect 1050 6758 1122 6810
rect 1174 6758 1246 6810
rect 1298 6758 1370 6810
rect 1422 6758 1494 6810
rect 1546 6758 1584 6810
rect 340 6686 1584 6758
rect 340 6634 378 6686
rect 430 6634 502 6686
rect 554 6634 626 6686
rect 678 6634 750 6686
rect 802 6634 874 6686
rect 926 6634 998 6686
rect 1050 6634 1122 6686
rect 1174 6634 1246 6686
rect 1298 6634 1370 6686
rect 1422 6634 1494 6686
rect 1546 6634 1584 6686
rect 340 6562 1584 6634
rect 340 6510 378 6562
rect 430 6510 502 6562
rect 554 6510 626 6562
rect 678 6510 750 6562
rect 802 6510 874 6562
rect 926 6510 998 6562
rect 1050 6510 1122 6562
rect 1174 6510 1246 6562
rect 1298 6510 1370 6562
rect 1422 6510 1494 6562
rect 1546 6510 1584 6562
rect 340 6438 1584 6510
rect 340 6386 378 6438
rect 430 6386 502 6438
rect 554 6386 626 6438
rect 678 6386 750 6438
rect 802 6386 874 6438
rect 926 6386 998 6438
rect 1050 6386 1122 6438
rect 1174 6386 1246 6438
rect 1298 6386 1370 6438
rect 1422 6386 1494 6438
rect 1546 6386 1584 6438
rect 340 6314 1584 6386
rect 340 6262 378 6314
rect 430 6262 502 6314
rect 554 6262 626 6314
rect 678 6262 750 6314
rect 802 6262 874 6314
rect 926 6262 998 6314
rect 1050 6262 1122 6314
rect 1174 6262 1246 6314
rect 1298 6262 1370 6314
rect 1422 6262 1494 6314
rect 1546 6262 1584 6314
rect 340 6190 1584 6262
rect 340 6138 378 6190
rect 430 6138 502 6190
rect 554 6138 626 6190
rect 678 6138 750 6190
rect 802 6138 874 6190
rect 926 6138 998 6190
rect 1050 6138 1122 6190
rect 1174 6138 1246 6190
rect 1298 6138 1370 6190
rect 1422 6138 1494 6190
rect 1546 6138 1584 6190
rect 340 6066 1584 6138
rect 340 6014 378 6066
rect 430 6014 502 6066
rect 554 6014 626 6066
rect 678 6014 750 6066
rect 802 6014 874 6066
rect 926 6014 998 6066
rect 1050 6014 1122 6066
rect 1174 6014 1246 6066
rect 1298 6014 1370 6066
rect 1422 6014 1494 6066
rect 1546 6014 1584 6066
rect 340 5942 1584 6014
rect 340 5890 378 5942
rect 430 5890 502 5942
rect 554 5890 626 5942
rect 678 5890 750 5942
rect 802 5890 874 5942
rect 926 5890 998 5942
rect 1050 5890 1122 5942
rect 1174 5890 1246 5942
rect 1298 5890 1370 5942
rect 1422 5890 1494 5942
rect 1546 5890 1584 5942
rect 340 5818 1584 5890
rect 340 5766 378 5818
rect 430 5766 502 5818
rect 554 5766 626 5818
rect 678 5766 750 5818
rect 802 5766 874 5818
rect 926 5766 998 5818
rect 1050 5766 1122 5818
rect 1174 5766 1246 5818
rect 1298 5766 1370 5818
rect 1422 5766 1494 5818
rect 1546 5766 1584 5818
rect 340 5694 1584 5766
rect 340 5642 378 5694
rect 430 5642 502 5694
rect 554 5642 626 5694
rect 678 5642 750 5694
rect 802 5642 874 5694
rect 926 5642 998 5694
rect 1050 5642 1122 5694
rect 1174 5642 1246 5694
rect 1298 5642 1370 5694
rect 1422 5642 1494 5694
rect 1546 5642 1584 5694
rect 340 5570 1584 5642
rect 340 5518 378 5570
rect 430 5518 502 5570
rect 554 5518 626 5570
rect 678 5518 750 5570
rect 802 5518 874 5570
rect 926 5518 998 5570
rect 1050 5518 1122 5570
rect 1174 5518 1246 5570
rect 1298 5518 1370 5570
rect 1422 5518 1494 5570
rect 1546 5518 1584 5570
rect 340 5446 1584 5518
rect 340 5394 378 5446
rect 430 5394 502 5446
rect 554 5394 626 5446
rect 678 5394 750 5446
rect 802 5394 874 5446
rect 926 5394 998 5446
rect 1050 5394 1122 5446
rect 1174 5394 1246 5446
rect 1298 5394 1370 5446
rect 1422 5394 1494 5446
rect 1546 5394 1584 5446
rect 340 5322 1584 5394
rect 340 5270 378 5322
rect 430 5270 502 5322
rect 554 5270 626 5322
rect 678 5270 750 5322
rect 802 5270 874 5322
rect 926 5270 998 5322
rect 1050 5270 1122 5322
rect 1174 5270 1246 5322
rect 1298 5270 1370 5322
rect 1422 5270 1494 5322
rect 1546 5270 1584 5322
rect 340 5198 1584 5270
rect 340 5146 378 5198
rect 430 5146 502 5198
rect 554 5146 626 5198
rect 678 5146 750 5198
rect 802 5146 874 5198
rect 926 5146 998 5198
rect 1050 5146 1122 5198
rect 1174 5146 1246 5198
rect 1298 5146 1370 5198
rect 1422 5146 1494 5198
rect 1546 5146 1584 5198
rect 340 5074 1584 5146
rect 340 5022 378 5074
rect 430 5022 502 5074
rect 554 5022 626 5074
rect 678 5022 750 5074
rect 802 5022 874 5074
rect 926 5022 998 5074
rect 1050 5022 1122 5074
rect 1174 5022 1246 5074
rect 1298 5022 1370 5074
rect 1422 5022 1494 5074
rect 1546 5022 1584 5074
rect 340 4950 1584 5022
rect 340 4898 378 4950
rect 430 4898 502 4950
rect 554 4898 626 4950
rect 678 4898 750 4950
rect 802 4898 874 4950
rect 926 4898 998 4950
rect 1050 4898 1122 4950
rect 1174 4898 1246 4950
rect 1298 4898 1370 4950
rect 1422 4898 1494 4950
rect 1546 4898 1584 4950
rect 340 4826 1584 4898
rect 340 4774 378 4826
rect 430 4774 502 4826
rect 554 4774 626 4826
rect 678 4774 750 4826
rect 802 4774 874 4826
rect 926 4774 998 4826
rect 1050 4774 1122 4826
rect 1174 4774 1246 4826
rect 1298 4774 1370 4826
rect 1422 4774 1494 4826
rect 1546 4774 1584 4826
rect 340 4702 1584 4774
rect 340 4650 378 4702
rect 430 4650 502 4702
rect 554 4650 626 4702
rect 678 4650 750 4702
rect 802 4650 874 4702
rect 926 4650 998 4702
rect 1050 4650 1122 4702
rect 1174 4650 1246 4702
rect 1298 4650 1370 4702
rect 1422 4650 1494 4702
rect 1546 4650 1584 4702
rect 340 4578 1584 4650
rect 340 4526 378 4578
rect 430 4526 502 4578
rect 554 4526 626 4578
rect 678 4526 750 4578
rect 802 4526 874 4578
rect 926 4526 998 4578
rect 1050 4526 1122 4578
rect 1174 4526 1246 4578
rect 1298 4526 1370 4578
rect 1422 4526 1494 4578
rect 1546 4526 1584 4578
rect 340 4454 1584 4526
rect 340 4402 378 4454
rect 430 4402 502 4454
rect 554 4402 626 4454
rect 678 4402 750 4454
rect 802 4402 874 4454
rect 926 4402 998 4454
rect 1050 4402 1122 4454
rect 1174 4402 1246 4454
rect 1298 4402 1370 4454
rect 1422 4402 1494 4454
rect 1546 4402 1584 4454
rect 340 4330 1584 4402
rect 340 4278 378 4330
rect 430 4278 502 4330
rect 554 4278 626 4330
rect 678 4278 750 4330
rect 802 4278 874 4330
rect 926 4278 998 4330
rect 1050 4278 1122 4330
rect 1174 4278 1246 4330
rect 1298 4278 1370 4330
rect 1422 4278 1494 4330
rect 1546 4278 1584 4330
rect 340 4206 1584 4278
rect 340 4154 378 4206
rect 430 4154 502 4206
rect 554 4154 626 4206
rect 678 4154 750 4206
rect 802 4154 874 4206
rect 926 4154 998 4206
rect 1050 4154 1122 4206
rect 1174 4154 1246 4206
rect 1298 4154 1370 4206
rect 1422 4154 1494 4206
rect 1546 4154 1584 4206
rect 340 4082 1584 4154
rect 340 4030 378 4082
rect 430 4030 502 4082
rect 554 4030 626 4082
rect 678 4030 750 4082
rect 802 4030 874 4082
rect 926 4030 998 4082
rect 1050 4030 1122 4082
rect 1174 4030 1246 4082
rect 1298 4030 1370 4082
rect 1422 4030 1494 4082
rect 1546 4030 1584 4082
rect 340 3958 1584 4030
rect 340 3906 378 3958
rect 430 3906 502 3958
rect 554 3906 626 3958
rect 678 3906 750 3958
rect 802 3906 874 3958
rect 926 3906 998 3958
rect 1050 3906 1122 3958
rect 1174 3906 1246 3958
rect 1298 3906 1370 3958
rect 1422 3906 1494 3958
rect 1546 3906 1584 3958
rect 340 3834 1584 3906
rect 340 3782 378 3834
rect 430 3782 502 3834
rect 554 3782 626 3834
rect 678 3782 750 3834
rect 802 3782 874 3834
rect 926 3782 998 3834
rect 1050 3782 1122 3834
rect 1174 3782 1246 3834
rect 1298 3782 1370 3834
rect 1422 3782 1494 3834
rect 1546 3782 1584 3834
rect 340 3710 1584 3782
rect 340 3658 378 3710
rect 430 3658 502 3710
rect 554 3658 626 3710
rect 678 3658 750 3710
rect 802 3658 874 3710
rect 926 3658 998 3710
rect 1050 3658 1122 3710
rect 1174 3658 1246 3710
rect 1298 3658 1370 3710
rect 1422 3658 1494 3710
rect 1546 3658 1584 3710
rect 340 3586 1584 3658
rect 340 3534 378 3586
rect 430 3534 502 3586
rect 554 3534 626 3586
rect 678 3534 750 3586
rect 802 3534 874 3586
rect 926 3534 998 3586
rect 1050 3534 1122 3586
rect 1174 3534 1246 3586
rect 1298 3534 1370 3586
rect 1422 3534 1494 3586
rect 1546 3534 1584 3586
rect 340 3462 1584 3534
rect 340 3410 378 3462
rect 430 3410 502 3462
rect 554 3410 626 3462
rect 678 3410 750 3462
rect 802 3410 874 3462
rect 926 3410 998 3462
rect 1050 3410 1122 3462
rect 1174 3410 1246 3462
rect 1298 3410 1370 3462
rect 1422 3410 1494 3462
rect 1546 3410 1584 3462
rect 340 3338 1584 3410
rect 340 3286 378 3338
rect 430 3286 502 3338
rect 554 3286 626 3338
rect 678 3286 750 3338
rect 802 3286 874 3338
rect 926 3286 998 3338
rect 1050 3286 1122 3338
rect 1174 3286 1246 3338
rect 1298 3286 1370 3338
rect 1422 3286 1494 3338
rect 1546 3286 1584 3338
rect 340 3214 1584 3286
rect 340 3162 378 3214
rect 430 3162 502 3214
rect 554 3162 626 3214
rect 678 3162 750 3214
rect 802 3162 874 3214
rect 926 3162 998 3214
rect 1050 3162 1122 3214
rect 1174 3162 1246 3214
rect 1298 3162 1370 3214
rect 1422 3162 1494 3214
rect 1546 3162 1584 3214
rect 340 3090 1584 3162
rect 340 3038 378 3090
rect 430 3038 502 3090
rect 554 3038 626 3090
rect 678 3038 750 3090
rect 802 3038 874 3090
rect 926 3038 998 3090
rect 1050 3038 1122 3090
rect 1174 3038 1246 3090
rect 1298 3038 1370 3090
rect 1422 3038 1494 3090
rect 1546 3038 1584 3090
rect 340 2966 1584 3038
rect 340 2914 378 2966
rect 430 2914 502 2966
rect 554 2914 626 2966
rect 678 2914 750 2966
rect 802 2914 874 2966
rect 926 2914 998 2966
rect 1050 2914 1122 2966
rect 1174 2914 1246 2966
rect 1298 2914 1370 2966
rect 1422 2914 1494 2966
rect 1546 2914 1584 2966
rect 340 2842 1584 2914
rect 340 2790 378 2842
rect 430 2790 502 2842
rect 554 2790 626 2842
rect 678 2790 750 2842
rect 802 2790 874 2842
rect 926 2790 998 2842
rect 1050 2790 1122 2842
rect 1174 2790 1246 2842
rect 1298 2790 1370 2842
rect 1422 2790 1494 2842
rect 1546 2790 1584 2842
rect 340 2718 1584 2790
rect 340 2666 378 2718
rect 430 2666 502 2718
rect 554 2666 626 2718
rect 678 2666 750 2718
rect 802 2666 874 2718
rect 926 2666 998 2718
rect 1050 2666 1122 2718
rect 1174 2666 1246 2718
rect 1298 2666 1370 2718
rect 1422 2666 1494 2718
rect 1546 2666 1584 2718
rect 340 2594 1584 2666
rect 340 2542 378 2594
rect 430 2542 502 2594
rect 554 2542 626 2594
rect 678 2542 750 2594
rect 802 2542 874 2594
rect 926 2542 998 2594
rect 1050 2542 1122 2594
rect 1174 2542 1246 2594
rect 1298 2542 1370 2594
rect 1422 2542 1494 2594
rect 1546 2542 1584 2594
rect 340 2470 1584 2542
rect 340 2418 378 2470
rect 430 2418 502 2470
rect 554 2418 626 2470
rect 678 2418 750 2470
rect 802 2418 874 2470
rect 926 2418 998 2470
rect 1050 2418 1122 2470
rect 1174 2418 1246 2470
rect 1298 2418 1370 2470
rect 1422 2418 1494 2470
rect 1546 2418 1584 2470
rect 340 2346 1584 2418
rect 340 2294 378 2346
rect 430 2294 502 2346
rect 554 2294 626 2346
rect 678 2294 750 2346
rect 802 2294 874 2346
rect 926 2294 998 2346
rect 1050 2294 1122 2346
rect 1174 2294 1246 2346
rect 1298 2294 1370 2346
rect 1422 2294 1494 2346
rect 1546 2294 1584 2346
rect 340 2222 1584 2294
rect 340 2170 378 2222
rect 430 2170 502 2222
rect 554 2170 626 2222
rect 678 2170 750 2222
rect 802 2170 874 2222
rect 926 2170 998 2222
rect 1050 2170 1122 2222
rect 1174 2170 1246 2222
rect 1298 2170 1370 2222
rect 1422 2170 1494 2222
rect 1546 2170 1584 2222
rect 340 2098 1584 2170
rect 340 2046 378 2098
rect 430 2046 502 2098
rect 554 2046 626 2098
rect 678 2046 750 2098
rect 802 2046 874 2098
rect 926 2046 998 2098
rect 1050 2046 1122 2098
rect 1174 2046 1246 2098
rect 1298 2046 1370 2098
rect 1422 2046 1494 2098
rect 1546 2046 1584 2098
rect 340 1974 1584 2046
rect 340 1922 378 1974
rect 430 1922 502 1974
rect 554 1922 626 1974
rect 678 1922 750 1974
rect 802 1922 874 1974
rect 926 1922 998 1974
rect 1050 1922 1122 1974
rect 1174 1922 1246 1974
rect 1298 1922 1370 1974
rect 1422 1922 1494 1974
rect 1546 1922 1584 1974
rect 340 1850 1584 1922
rect 340 1798 378 1850
rect 430 1798 502 1850
rect 554 1798 626 1850
rect 678 1798 750 1850
rect 802 1798 874 1850
rect 926 1798 998 1850
rect 1050 1798 1122 1850
rect 1174 1798 1246 1850
rect 1298 1798 1370 1850
rect 1422 1798 1494 1850
rect 1546 1798 1584 1850
rect 340 1726 1584 1798
rect 340 1674 378 1726
rect 430 1674 502 1726
rect 554 1674 626 1726
rect 678 1674 750 1726
rect 802 1674 874 1726
rect 926 1674 998 1726
rect 1050 1674 1122 1726
rect 1174 1674 1246 1726
rect 1298 1674 1370 1726
rect 1422 1674 1494 1726
rect 1546 1674 1584 1726
rect 340 1602 1584 1674
rect 340 1550 378 1602
rect 430 1550 502 1602
rect 554 1550 626 1602
rect 678 1550 750 1602
rect 802 1550 874 1602
rect 926 1550 998 1602
rect 1050 1550 1122 1602
rect 1174 1550 1246 1602
rect 1298 1550 1370 1602
rect 1422 1550 1494 1602
rect 1546 1550 1584 1602
rect 340 1478 1584 1550
rect 340 1426 378 1478
rect 430 1426 502 1478
rect 554 1426 626 1478
rect 678 1426 750 1478
rect 802 1426 874 1478
rect 926 1426 998 1478
rect 1050 1426 1122 1478
rect 1174 1426 1246 1478
rect 1298 1426 1370 1478
rect 1422 1426 1494 1478
rect 1546 1426 1584 1478
rect 340 1354 1584 1426
rect 340 1302 378 1354
rect 430 1302 502 1354
rect 554 1302 626 1354
rect 678 1302 750 1354
rect 802 1302 874 1354
rect 926 1302 998 1354
rect 1050 1302 1122 1354
rect 1174 1302 1246 1354
rect 1298 1302 1370 1354
rect 1422 1302 1494 1354
rect 1546 1302 1584 1354
rect 340 1230 1584 1302
rect 340 1178 378 1230
rect 430 1178 502 1230
rect 554 1178 626 1230
rect 678 1178 750 1230
rect 802 1178 874 1230
rect 926 1178 998 1230
rect 1050 1178 1122 1230
rect 1174 1178 1246 1230
rect 1298 1178 1370 1230
rect 1422 1178 1494 1230
rect 1546 1178 1584 1230
rect 340 1106 1584 1178
rect 340 1054 378 1106
rect 430 1054 502 1106
rect 554 1054 626 1106
rect 678 1054 750 1106
rect 802 1054 874 1106
rect 926 1054 998 1106
rect 1050 1054 1122 1106
rect 1174 1054 1246 1106
rect 1298 1054 1370 1106
rect 1422 1054 1494 1106
rect 1546 1054 1584 1106
rect 340 982 1584 1054
rect 340 930 378 982
rect 430 930 502 982
rect 554 930 626 982
rect 678 930 750 982
rect 802 930 874 982
rect 926 930 998 982
rect 1050 930 1122 982
rect 1174 930 1246 982
rect 1298 930 1370 982
rect 1422 930 1494 982
rect 1546 930 1584 982
rect 340 858 1584 930
rect 340 806 378 858
rect 430 806 502 858
rect 554 806 626 858
rect 678 806 750 858
rect 802 806 874 858
rect 926 806 998 858
rect 1050 806 1122 858
rect 1174 806 1246 858
rect 1298 806 1370 858
rect 1422 806 1494 858
rect 1546 806 1584 858
rect 340 734 1584 806
rect 340 682 378 734
rect 430 682 502 734
rect 554 682 626 734
rect 678 682 750 734
rect 802 682 874 734
rect 926 682 998 734
rect 1050 682 1122 734
rect 1174 682 1246 734
rect 1298 682 1370 734
rect 1422 682 1494 734
rect 1546 682 1584 734
rect 340 610 1584 682
rect 340 558 378 610
rect 430 558 502 610
rect 554 558 626 610
rect 678 558 750 610
rect 802 558 874 610
rect 926 558 998 610
rect 1050 558 1122 610
rect 1174 558 1246 610
rect 1298 558 1370 610
rect 1422 558 1494 610
rect 1546 558 1584 610
rect 340 486 1584 558
rect 340 434 378 486
rect 430 434 502 486
rect 554 434 626 486
rect 678 434 750 486
rect 802 434 874 486
rect 926 434 998 486
rect 1050 434 1122 486
rect 1174 434 1246 486
rect 1298 434 1370 486
rect 1422 434 1494 486
rect 1546 434 1584 486
rect 340 362 1584 434
rect 340 310 378 362
rect 430 310 502 362
rect 554 310 626 362
rect 678 310 750 362
rect 802 310 874 362
rect 926 310 998 362
rect 1050 310 1122 362
rect 1174 310 1246 362
rect 1298 310 1370 362
rect 1422 310 1494 362
rect 1546 310 1584 362
rect 340 238 1584 310
rect 340 186 378 238
rect 430 186 502 238
rect 554 186 626 238
rect 678 186 750 238
rect 802 186 874 238
rect 926 186 998 238
rect 1050 186 1122 238
rect 1174 186 1246 238
rect 1298 186 1370 238
rect 1422 186 1494 238
rect 1546 186 1584 238
rect 340 114 1584 186
rect 340 62 378 114
rect 430 62 502 114
rect 554 62 626 114
rect 678 62 750 114
rect 802 62 874 114
rect 926 62 998 114
rect 1050 62 1122 114
rect 1174 62 1246 114
rect 1298 62 1370 114
rect 1422 62 1494 114
rect 1546 62 1584 114
rect 340 0 1584 62
<< via2 >>
rect -21 7874 0 7915
rect 0 7874 35 7915
rect 121 7874 156 7915
rect 156 7874 177 7915
rect -21 7859 35 7874
rect 121 7859 177 7874
rect -21 7750 0 7773
rect 0 7750 35 7773
rect 121 7750 156 7773
rect 156 7750 177 7773
rect -21 7717 35 7750
rect 121 7717 177 7750
rect -21 7626 0 7631
rect 0 7626 35 7631
rect 121 7626 156 7631
rect 156 7626 177 7631
rect -21 7575 35 7626
rect 121 7575 177 7626
rect -21 7433 35 7489
rect 121 7433 177 7489
rect -21 7306 35 7347
rect 121 7306 177 7347
rect -21 7291 0 7306
rect 0 7291 35 7306
rect 121 7291 156 7306
rect 156 7291 177 7306
rect -21 6934 35 6950
rect 121 6934 177 6950
rect -21 6894 0 6934
rect 0 6894 35 6934
rect 121 6894 156 6934
rect 156 6894 177 6934
rect -21 6758 0 6808
rect 0 6758 35 6808
rect 121 6758 156 6808
rect 156 6758 177 6808
rect -21 6752 35 6758
rect 121 6752 177 6758
rect -21 6634 0 6666
rect 0 6634 35 6666
rect 121 6634 156 6666
rect 156 6634 177 6666
rect -21 6610 35 6634
rect 121 6610 177 6634
rect -21 6510 0 6524
rect 0 6510 35 6524
rect 121 6510 156 6524
rect 156 6510 177 6524
rect -21 6468 35 6510
rect 121 6468 177 6510
rect -21 6326 35 6382
rect 121 6326 177 6382
rect -21 6190 35 6240
rect 121 6190 177 6240
rect -21 6184 0 6190
rect 0 6184 35 6190
rect 121 6184 156 6190
rect 156 6184 177 6190
rect -21 6066 35 6098
rect 121 6066 177 6098
rect -21 6042 0 6066
rect 0 6042 35 6066
rect 121 6042 156 6066
rect 156 6042 177 6066
rect -21 5942 35 5956
rect 121 5942 177 5956
rect -21 5900 0 5942
rect 0 5900 35 5942
rect 121 5900 156 5942
rect 156 5900 177 5942
rect -21 5766 0 5814
rect 0 5766 35 5814
rect 121 5766 156 5814
rect 156 5766 177 5814
rect -21 5758 35 5766
rect 121 5758 177 5766
rect -21 5642 0 5672
rect 0 5642 35 5672
rect 121 5642 156 5672
rect 156 5642 177 5672
rect -21 5616 35 5642
rect 121 5616 177 5642
rect -21 5518 0 5530
rect 0 5518 35 5530
rect 121 5518 156 5530
rect 156 5518 177 5530
rect -21 5474 35 5518
rect 121 5474 177 5518
rect -21 5332 35 5388
rect 121 5332 177 5388
rect -21 5198 35 5246
rect 121 5198 177 5246
rect -21 5190 0 5198
rect 0 5190 35 5198
rect 121 5190 156 5198
rect 156 5190 177 5198
rect -21 5074 35 5104
rect 121 5074 177 5104
rect -21 5048 0 5074
rect 0 5048 35 5074
rect 121 5048 156 5074
rect 156 5048 177 5074
rect -21 4950 35 4962
rect 121 4950 177 4962
rect -21 4906 0 4950
rect 0 4906 35 4950
rect 121 4906 156 4950
rect 156 4906 177 4950
rect -21 4774 0 4820
rect 0 4774 35 4820
rect 121 4774 156 4820
rect 156 4774 177 4820
rect -21 4764 35 4774
rect 121 4764 177 4774
rect -21 4650 0 4678
rect 0 4650 35 4678
rect 121 4650 156 4678
rect 156 4650 177 4678
rect -21 4622 35 4650
rect 121 4622 177 4650
rect -21 4526 0 4536
rect 0 4526 35 4536
rect 121 4526 156 4536
rect 156 4526 177 4536
rect -21 4480 35 4526
rect 121 4480 177 4526
rect -21 4338 35 4394
rect 121 4338 177 4394
rect -21 4206 35 4252
rect 121 4206 177 4252
rect -21 4196 0 4206
rect 0 4196 35 4206
rect 121 4196 156 4206
rect 156 4196 177 4206
rect -21 4082 35 4110
rect 121 4082 177 4110
rect -21 4054 0 4082
rect 0 4054 35 4082
rect 121 4054 156 4082
rect 156 4054 177 4082
rect -21 3710 35 3763
rect 121 3710 177 3763
rect -21 3707 0 3710
rect 0 3707 35 3710
rect 121 3707 156 3710
rect 156 3707 177 3710
rect -21 3586 35 3621
rect 121 3586 177 3621
rect -21 3565 0 3586
rect 0 3565 35 3586
rect 121 3565 156 3586
rect 156 3565 177 3586
rect -21 3462 35 3479
rect 121 3462 177 3479
rect -21 3423 0 3462
rect 0 3423 35 3462
rect 121 3423 156 3462
rect 156 3423 177 3462
rect -21 3286 0 3337
rect 0 3286 35 3337
rect 121 3286 156 3337
rect 156 3286 177 3337
rect -21 3281 35 3286
rect 121 3281 177 3286
rect -21 3162 0 3195
rect 0 3162 35 3195
rect 121 3162 156 3195
rect 156 3162 177 3195
rect -21 3139 35 3162
rect 121 3139 177 3162
rect -21 3038 0 3053
rect 0 3038 35 3053
rect 121 3038 156 3053
rect 156 3038 177 3053
rect -21 2997 35 3038
rect 121 2997 177 3038
rect -21 2855 35 2911
rect 121 2855 177 2911
rect -21 2718 35 2769
rect 121 2718 177 2769
rect -21 2713 0 2718
rect 0 2713 35 2718
rect 121 2713 156 2718
rect 156 2713 177 2718
rect -21 2594 35 2627
rect 121 2594 177 2627
rect -21 2571 0 2594
rect 0 2571 35 2594
rect 121 2571 156 2594
rect 156 2571 177 2594
rect -21 2470 35 2485
rect 121 2470 177 2485
rect -21 2429 0 2470
rect 0 2429 35 2470
rect 121 2429 156 2470
rect 156 2429 177 2470
rect -21 2294 0 2343
rect 0 2294 35 2343
rect 121 2294 156 2343
rect 156 2294 177 2343
rect -21 2287 35 2294
rect 121 2287 177 2294
rect -21 2170 0 2201
rect 0 2170 35 2201
rect 121 2170 156 2201
rect 156 2170 177 2201
rect -21 2145 35 2170
rect 121 2145 177 2170
rect -21 2046 0 2059
rect 0 2046 35 2059
rect 121 2046 156 2059
rect 156 2046 177 2059
rect -21 2003 35 2046
rect 121 2003 177 2046
rect -21 1861 35 1917
rect 121 1861 177 1917
rect -21 1726 35 1775
rect 121 1726 177 1775
rect -21 1719 0 1726
rect 0 1719 35 1726
rect 121 1719 156 1726
rect 156 1719 177 1726
rect -21 1602 35 1633
rect 121 1602 177 1633
rect -21 1577 0 1602
rect 0 1577 35 1602
rect 121 1577 156 1602
rect 156 1577 177 1602
rect -21 1478 35 1491
rect 121 1478 177 1491
rect -21 1435 0 1478
rect 0 1435 35 1478
rect 121 1435 156 1478
rect 156 1435 177 1478
rect -21 1302 0 1349
rect 0 1302 35 1349
rect 121 1302 156 1349
rect 156 1302 177 1349
rect -21 1293 35 1302
rect 121 1293 177 1302
rect -21 1178 0 1207
rect 0 1178 35 1207
rect 121 1178 156 1207
rect 156 1178 177 1207
rect -21 1151 35 1178
rect 121 1151 177 1178
rect -21 1054 0 1065
rect 0 1054 35 1065
rect 121 1054 156 1065
rect 156 1054 177 1065
rect -21 1009 35 1054
rect 121 1009 177 1054
rect -21 867 35 923
rect 121 867 177 923
rect -21 494 35 550
rect 121 494 177 550
rect -21 362 35 408
rect 121 362 177 408
rect -21 352 0 362
rect 0 352 35 362
rect 121 352 156 362
rect 156 352 177 362
rect -21 238 35 266
rect 121 238 177 266
rect -21 210 0 238
rect 0 210 35 238
rect 121 210 156 238
rect 156 210 177 238
rect -21 114 35 124
rect 121 114 177 124
rect -21 68 0 114
rect 0 68 35 114
rect 121 68 156 114
rect 156 68 177 114
<< metal3 >>
rect -31 7915 187 7925
rect -31 7859 -21 7915
rect 35 7859 121 7915
rect 177 7859 187 7915
rect -31 7773 187 7859
rect -31 7717 -21 7773
rect 35 7717 121 7773
rect 177 7717 187 7773
rect -31 7631 187 7717
rect -31 7575 -21 7631
rect 35 7575 121 7631
rect 177 7575 187 7631
rect -31 7489 187 7575
rect -31 7433 -21 7489
rect 35 7433 121 7489
rect 177 7433 187 7489
rect -31 7347 187 7433
rect -31 7291 -21 7347
rect 35 7291 121 7347
rect 177 7291 187 7347
rect -31 7281 187 7291
rect -31 6950 187 6960
rect -31 6894 -21 6950
rect 35 6894 121 6950
rect 177 6894 187 6950
rect -31 6808 187 6894
rect -31 6752 -21 6808
rect 35 6752 121 6808
rect 177 6752 187 6808
rect -31 6666 187 6752
rect -31 6610 -21 6666
rect 35 6610 121 6666
rect 177 6610 187 6666
rect -31 6524 187 6610
rect -31 6468 -21 6524
rect 35 6468 121 6524
rect 177 6468 187 6524
rect -31 6382 187 6468
rect -31 6326 -21 6382
rect 35 6326 121 6382
rect 177 6326 187 6382
rect -31 6240 187 6326
rect -31 6184 -21 6240
rect 35 6184 121 6240
rect 177 6184 187 6240
rect -31 6098 187 6184
rect -31 6042 -21 6098
rect 35 6042 121 6098
rect 177 6042 187 6098
rect -31 5956 187 6042
rect -31 5900 -21 5956
rect 35 5900 121 5956
rect 177 5900 187 5956
rect -31 5814 187 5900
rect -31 5758 -21 5814
rect 35 5758 121 5814
rect 177 5758 187 5814
rect -31 5672 187 5758
rect -31 5616 -21 5672
rect 35 5616 121 5672
rect 177 5616 187 5672
rect -31 5530 187 5616
rect -31 5474 -21 5530
rect 35 5474 121 5530
rect 177 5474 187 5530
rect -31 5388 187 5474
rect -31 5332 -21 5388
rect 35 5332 121 5388
rect 177 5332 187 5388
rect -31 5246 187 5332
rect -31 5190 -21 5246
rect 35 5190 121 5246
rect 177 5190 187 5246
rect -31 5104 187 5190
rect -31 5048 -21 5104
rect 35 5048 121 5104
rect 177 5048 187 5104
rect -31 4962 187 5048
rect -31 4906 -21 4962
rect 35 4906 121 4962
rect 177 4906 187 4962
rect -31 4820 187 4906
rect -31 4764 -21 4820
rect 35 4764 121 4820
rect 177 4764 187 4820
rect -31 4678 187 4764
rect -31 4622 -21 4678
rect 35 4622 121 4678
rect 177 4622 187 4678
rect -31 4536 187 4622
rect -31 4480 -21 4536
rect 35 4480 121 4536
rect 177 4480 187 4536
rect -31 4394 187 4480
rect -31 4338 -21 4394
rect 35 4338 121 4394
rect 177 4338 187 4394
rect -31 4252 187 4338
rect -31 4196 -21 4252
rect 35 4196 121 4252
rect 177 4196 187 4252
rect -31 4110 187 4196
rect -31 4054 -21 4110
rect 35 4054 121 4110
rect 177 4054 187 4110
rect -31 4044 187 4054
rect -31 3763 187 3773
rect -31 3707 -21 3763
rect 35 3707 121 3763
rect 177 3707 187 3763
rect -31 3621 187 3707
rect -31 3565 -21 3621
rect 35 3565 121 3621
rect 177 3565 187 3621
rect -31 3479 187 3565
rect -31 3423 -21 3479
rect 35 3423 121 3479
rect 177 3423 187 3479
rect -31 3337 187 3423
rect -31 3281 -21 3337
rect 35 3281 121 3337
rect 177 3281 187 3337
rect -31 3195 187 3281
rect -31 3139 -21 3195
rect 35 3139 121 3195
rect 177 3139 187 3195
rect -31 3053 187 3139
rect -31 2997 -21 3053
rect 35 2997 121 3053
rect 177 2997 187 3053
rect -31 2911 187 2997
rect -31 2855 -21 2911
rect 35 2855 121 2911
rect 177 2855 187 2911
rect -31 2769 187 2855
rect -31 2713 -21 2769
rect 35 2713 121 2769
rect 177 2713 187 2769
rect -31 2627 187 2713
rect -31 2571 -21 2627
rect 35 2571 121 2627
rect 177 2571 187 2627
rect -31 2485 187 2571
rect -31 2429 -21 2485
rect 35 2429 121 2485
rect 177 2429 187 2485
rect -31 2343 187 2429
rect -31 2287 -21 2343
rect 35 2287 121 2343
rect 177 2287 187 2343
rect -31 2201 187 2287
rect -31 2145 -21 2201
rect 35 2145 121 2201
rect 177 2145 187 2201
rect -31 2059 187 2145
rect -31 2003 -21 2059
rect 35 2003 121 2059
rect 177 2003 187 2059
rect -31 1917 187 2003
rect -31 1861 -21 1917
rect 35 1861 121 1917
rect 177 1861 187 1917
rect -31 1775 187 1861
rect -31 1719 -21 1775
rect 35 1719 121 1775
rect 177 1719 187 1775
rect -31 1633 187 1719
rect -31 1577 -21 1633
rect 35 1577 121 1633
rect 177 1577 187 1633
rect -31 1491 187 1577
rect -31 1435 -21 1491
rect 35 1435 121 1491
rect 177 1435 187 1491
rect -31 1349 187 1435
rect -31 1293 -21 1349
rect 35 1293 121 1349
rect 177 1293 187 1349
rect -31 1207 187 1293
rect -31 1151 -21 1207
rect 35 1151 121 1207
rect 177 1151 187 1207
rect -31 1065 187 1151
rect -31 1009 -21 1065
rect 35 1009 121 1065
rect 177 1009 187 1065
rect -31 923 187 1009
rect -31 867 -21 923
rect 35 867 121 923
rect 177 867 187 923
rect -31 857 187 867
rect -31 550 187 560
rect -31 494 -21 550
rect 35 494 121 550
rect 177 494 187 550
rect -31 408 187 494
rect -31 352 -21 408
rect 35 352 121 408
rect 177 352 187 408
rect -31 266 187 352
rect -31 210 -21 266
rect 35 210 121 266
rect 177 210 187 266
rect -31 124 187 210
rect -31 68 -21 124
rect 35 68 121 124
rect 177 68 187 124
rect -31 58 187 68
use M2_M1_CDNS_40661953145365  M2_M1_CDNS_40661953145365_0
timestamp 1759194789
transform 1 0 78 0 1 3994
box 0 0 1 1
use M2_M1_CDNS_40661953145366  M2_M1_CDNS_40661953145366_0
timestamp 1759194789
transform 1 0 962 0 1 3994
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_0
timestamp 1759194789
transform 1 0 78 0 1 2315
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_1
timestamp 1759194789
transform 1 0 78 0 1 5502
box 0 0 1 1
use M3_M2_CDNS_40661953145264  M3_M2_CDNS_40661953145264_0
timestamp 1759194789
transform 1 0 78 0 1 309
box 0 0 1 1
use M3_M2_CDNS_40661953145353  M3_M2_CDNS_40661953145353_0
timestamp 1759194789
transform 1 0 78 0 1 7603
box 0 0 1 1
<< properties >>
string GDS_END 2947614
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2947054
<< end >>
