magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
<< nwell >>
rect 29138 95074 56005 95590
rect 29138 93521 32850 95074
rect 35260 94009 39818 95074
rect 35260 93833 39436 94009
rect 45169 93833 49764 95074
rect 52285 93833 56005 95074
<< pwell >>
rect 1774 94682 24710 94714
rect 1774 35138 24710 35170
<< mvpsubdiff >>
rect 352 96683 86098 96702
rect 352 96637 371 96683
rect 417 96637 495 96683
rect 541 96637 619 96683
rect 665 96637 743 96683
rect 789 96637 867 96683
rect 913 96637 991 96683
rect 1037 96637 1115 96683
rect 1161 96637 1239 96683
rect 1285 96637 1363 96683
rect 1409 96637 1487 96683
rect 1533 96637 1611 96683
rect 1657 96637 1735 96683
rect 1781 96637 1859 96683
rect 1905 96637 1983 96683
rect 2029 96637 2107 96683
rect 2153 96637 2231 96683
rect 2277 96637 2355 96683
rect 2401 96637 2479 96683
rect 2525 96637 2603 96683
rect 2649 96637 2727 96683
rect 2773 96637 2851 96683
rect 2897 96637 2975 96683
rect 3021 96637 3099 96683
rect 3145 96637 3223 96683
rect 3269 96637 3347 96683
rect 3393 96637 3471 96683
rect 3517 96637 3595 96683
rect 3641 96637 3719 96683
rect 3765 96637 3843 96683
rect 3889 96637 3967 96683
rect 4013 96637 4091 96683
rect 4137 96637 4215 96683
rect 4261 96637 4339 96683
rect 4385 96637 4463 96683
rect 4509 96637 4587 96683
rect 4633 96637 4711 96683
rect 4757 96637 4835 96683
rect 4881 96637 4959 96683
rect 5005 96637 5083 96683
rect 5129 96637 5207 96683
rect 5253 96637 5331 96683
rect 5377 96637 5455 96683
rect 5501 96637 5579 96683
rect 5625 96637 5703 96683
rect 5749 96637 5827 96683
rect 5873 96637 5951 96683
rect 5997 96637 6075 96683
rect 6121 96637 6199 96683
rect 6245 96637 6323 96683
rect 6369 96637 6447 96683
rect 6493 96637 6571 96683
rect 6617 96637 6695 96683
rect 6741 96637 6819 96683
rect 6865 96637 6943 96683
rect 6989 96637 7067 96683
rect 7113 96637 7191 96683
rect 7237 96637 7315 96683
rect 7361 96637 7439 96683
rect 7485 96637 7563 96683
rect 7609 96637 7687 96683
rect 7733 96637 7811 96683
rect 7857 96637 7935 96683
rect 7981 96637 8059 96683
rect 8105 96637 8183 96683
rect 8229 96637 8307 96683
rect 8353 96637 8431 96683
rect 8477 96637 8555 96683
rect 8601 96637 8679 96683
rect 8725 96637 8803 96683
rect 8849 96637 8927 96683
rect 8973 96637 9051 96683
rect 9097 96637 9175 96683
rect 9221 96637 9299 96683
rect 9345 96637 9423 96683
rect 9469 96637 9547 96683
rect 9593 96637 9671 96683
rect 9717 96637 9795 96683
rect 9841 96637 9919 96683
rect 9965 96637 10043 96683
rect 10089 96637 10167 96683
rect 10213 96637 10291 96683
rect 10337 96637 10415 96683
rect 10461 96637 10539 96683
rect 10585 96637 10663 96683
rect 10709 96637 10787 96683
rect 10833 96637 10911 96683
rect 10957 96637 11035 96683
rect 11081 96637 11159 96683
rect 11205 96637 11283 96683
rect 11329 96637 11407 96683
rect 11453 96637 11531 96683
rect 11577 96637 11655 96683
rect 11701 96637 11779 96683
rect 11825 96637 11903 96683
rect 11949 96637 12027 96683
rect 12073 96637 12151 96683
rect 12197 96637 12275 96683
rect 12321 96637 12399 96683
rect 12445 96637 12523 96683
rect 12569 96637 12647 96683
rect 12693 96637 12771 96683
rect 12817 96637 12895 96683
rect 12941 96637 13019 96683
rect 13065 96637 13143 96683
rect 13189 96637 13267 96683
rect 13313 96637 13391 96683
rect 13437 96637 13515 96683
rect 13561 96637 13639 96683
rect 13685 96637 13763 96683
rect 13809 96637 13887 96683
rect 13933 96637 14011 96683
rect 14057 96637 14135 96683
rect 14181 96637 14259 96683
rect 14305 96637 14383 96683
rect 14429 96637 14507 96683
rect 14553 96637 14631 96683
rect 14677 96637 14755 96683
rect 14801 96637 14879 96683
rect 14925 96637 15003 96683
rect 15049 96637 15127 96683
rect 15173 96637 15251 96683
rect 15297 96637 15375 96683
rect 15421 96637 15499 96683
rect 15545 96637 15623 96683
rect 15669 96637 15747 96683
rect 15793 96637 15871 96683
rect 15917 96637 15995 96683
rect 16041 96637 16119 96683
rect 16165 96637 16243 96683
rect 16289 96637 16367 96683
rect 16413 96637 16491 96683
rect 16537 96637 16615 96683
rect 16661 96637 16739 96683
rect 16785 96637 16863 96683
rect 16909 96637 16987 96683
rect 17033 96637 17111 96683
rect 17157 96637 17235 96683
rect 17281 96637 17359 96683
rect 17405 96637 17483 96683
rect 17529 96637 17607 96683
rect 17653 96637 17731 96683
rect 17777 96637 17855 96683
rect 17901 96637 17979 96683
rect 18025 96637 18103 96683
rect 18149 96637 18227 96683
rect 18273 96637 18351 96683
rect 18397 96637 18475 96683
rect 18521 96637 18599 96683
rect 18645 96637 18723 96683
rect 18769 96637 18847 96683
rect 18893 96637 18971 96683
rect 19017 96637 19095 96683
rect 19141 96637 19219 96683
rect 19265 96637 19343 96683
rect 19389 96637 19467 96683
rect 19513 96637 19591 96683
rect 19637 96637 19715 96683
rect 19761 96637 19839 96683
rect 19885 96637 19963 96683
rect 20009 96637 20087 96683
rect 20133 96637 20211 96683
rect 20257 96637 20335 96683
rect 20381 96637 20459 96683
rect 20505 96637 20583 96683
rect 20629 96637 20707 96683
rect 20753 96637 20831 96683
rect 20877 96637 20955 96683
rect 21001 96637 21079 96683
rect 21125 96637 21203 96683
rect 21249 96637 21327 96683
rect 21373 96637 21451 96683
rect 21497 96637 21575 96683
rect 21621 96637 21699 96683
rect 21745 96637 21823 96683
rect 21869 96637 21947 96683
rect 21993 96637 22071 96683
rect 22117 96637 22195 96683
rect 22241 96637 22319 96683
rect 22365 96637 22443 96683
rect 22489 96637 22567 96683
rect 22613 96637 22691 96683
rect 22737 96637 22815 96683
rect 22861 96637 22939 96683
rect 22985 96637 23063 96683
rect 23109 96637 23187 96683
rect 23233 96637 23311 96683
rect 23357 96637 23435 96683
rect 23481 96637 23559 96683
rect 23605 96637 23683 96683
rect 23729 96637 23807 96683
rect 23853 96637 23931 96683
rect 23977 96637 24055 96683
rect 24101 96637 24179 96683
rect 24225 96637 24303 96683
rect 24349 96637 24427 96683
rect 24473 96637 24551 96683
rect 24597 96637 24675 96683
rect 24721 96637 24799 96683
rect 24845 96637 24923 96683
rect 24969 96637 25047 96683
rect 25093 96637 25171 96683
rect 25217 96637 25295 96683
rect 25341 96637 25419 96683
rect 25465 96637 25543 96683
rect 25589 96637 25667 96683
rect 25713 96637 25791 96683
rect 25837 96637 25915 96683
rect 25961 96637 26039 96683
rect 26085 96637 26163 96683
rect 26209 96637 26287 96683
rect 26333 96637 26411 96683
rect 26457 96637 26535 96683
rect 26581 96637 26659 96683
rect 26705 96637 26783 96683
rect 26829 96637 26907 96683
rect 26953 96637 27031 96683
rect 27077 96637 27155 96683
rect 27201 96637 27279 96683
rect 27325 96637 27403 96683
rect 27449 96637 27527 96683
rect 27573 96637 27651 96683
rect 27697 96637 27775 96683
rect 27821 96637 27899 96683
rect 27945 96637 28023 96683
rect 28069 96637 28147 96683
rect 28193 96637 28271 96683
rect 28317 96637 28395 96683
rect 28441 96637 28519 96683
rect 28565 96637 28643 96683
rect 28689 96637 28767 96683
rect 28813 96637 28891 96683
rect 28937 96637 29015 96683
rect 29061 96637 29139 96683
rect 29185 96637 29263 96683
rect 29309 96637 29387 96683
rect 29433 96637 29511 96683
rect 29557 96637 29635 96683
rect 29681 96637 29759 96683
rect 29805 96637 29883 96683
rect 29929 96637 30007 96683
rect 30053 96637 30131 96683
rect 30177 96637 30255 96683
rect 30301 96637 30379 96683
rect 30425 96637 30503 96683
rect 30549 96637 30627 96683
rect 30673 96637 30751 96683
rect 30797 96637 30875 96683
rect 30921 96637 30999 96683
rect 31045 96637 31123 96683
rect 31169 96637 31247 96683
rect 31293 96637 31371 96683
rect 31417 96637 31495 96683
rect 31541 96637 31619 96683
rect 31665 96637 31743 96683
rect 31789 96637 31867 96683
rect 31913 96637 31991 96683
rect 32037 96637 32115 96683
rect 32161 96637 32239 96683
rect 32285 96637 32363 96683
rect 32409 96637 32487 96683
rect 32533 96637 32611 96683
rect 32657 96637 32735 96683
rect 32781 96637 32859 96683
rect 32905 96637 32983 96683
rect 33029 96637 33107 96683
rect 33153 96637 33231 96683
rect 33277 96637 33355 96683
rect 33401 96637 33479 96683
rect 33525 96637 33603 96683
rect 33649 96637 33727 96683
rect 33773 96637 33851 96683
rect 33897 96637 33975 96683
rect 34021 96637 34099 96683
rect 34145 96637 34223 96683
rect 34269 96637 34347 96683
rect 34393 96637 34471 96683
rect 34517 96637 34595 96683
rect 34641 96637 34719 96683
rect 34765 96637 34843 96683
rect 34889 96637 34967 96683
rect 35013 96637 35091 96683
rect 35137 96637 35215 96683
rect 35261 96637 35339 96683
rect 35385 96637 35463 96683
rect 35509 96637 35587 96683
rect 35633 96637 35711 96683
rect 35757 96637 35835 96683
rect 35881 96637 35959 96683
rect 36005 96637 36083 96683
rect 36129 96637 36207 96683
rect 36253 96637 36331 96683
rect 36377 96637 36455 96683
rect 36501 96637 36579 96683
rect 36625 96637 36703 96683
rect 36749 96637 36827 96683
rect 36873 96637 36951 96683
rect 36997 96637 37075 96683
rect 37121 96637 37199 96683
rect 37245 96637 37323 96683
rect 37369 96637 37447 96683
rect 37493 96637 37571 96683
rect 37617 96637 37695 96683
rect 37741 96637 37819 96683
rect 37865 96637 37943 96683
rect 37989 96637 38067 96683
rect 38113 96637 38191 96683
rect 38237 96637 38315 96683
rect 38361 96637 38439 96683
rect 38485 96637 38563 96683
rect 38609 96637 38687 96683
rect 38733 96637 38811 96683
rect 38857 96637 38935 96683
rect 38981 96637 39059 96683
rect 39105 96637 39183 96683
rect 39229 96637 39307 96683
rect 39353 96637 39431 96683
rect 39477 96637 39555 96683
rect 39601 96637 39679 96683
rect 39725 96637 39803 96683
rect 39849 96637 39927 96683
rect 39973 96637 40051 96683
rect 40097 96637 40175 96683
rect 40221 96637 40299 96683
rect 40345 96637 40423 96683
rect 40469 96637 40547 96683
rect 40593 96637 40671 96683
rect 40717 96637 40795 96683
rect 40841 96637 40919 96683
rect 40965 96637 41043 96683
rect 41089 96637 41167 96683
rect 41213 96637 41291 96683
rect 41337 96637 41415 96683
rect 41461 96637 41539 96683
rect 41585 96637 41663 96683
rect 41709 96637 41787 96683
rect 41833 96637 41911 96683
rect 41957 96637 42035 96683
rect 42081 96637 42159 96683
rect 42205 96637 42283 96683
rect 42329 96637 42407 96683
rect 42453 96637 42531 96683
rect 42577 96637 42655 96683
rect 42701 96637 42779 96683
rect 42825 96637 42903 96683
rect 42949 96637 43027 96683
rect 43073 96637 43151 96683
rect 43197 96637 43275 96683
rect 43321 96637 43399 96683
rect 43445 96637 43523 96683
rect 43569 96637 43647 96683
rect 43693 96637 43771 96683
rect 43817 96637 43895 96683
rect 43941 96637 44019 96683
rect 44065 96637 44143 96683
rect 44189 96637 44267 96683
rect 44313 96637 44391 96683
rect 44437 96637 44515 96683
rect 44561 96637 44639 96683
rect 44685 96637 44763 96683
rect 44809 96637 44887 96683
rect 44933 96637 45011 96683
rect 45057 96637 45135 96683
rect 45181 96637 45259 96683
rect 45305 96637 45383 96683
rect 45429 96637 45507 96683
rect 45553 96637 45631 96683
rect 45677 96637 45755 96683
rect 45801 96637 45879 96683
rect 45925 96637 46003 96683
rect 46049 96637 46127 96683
rect 46173 96637 46251 96683
rect 46297 96637 46375 96683
rect 46421 96637 46499 96683
rect 46545 96637 46623 96683
rect 46669 96637 46747 96683
rect 46793 96637 46871 96683
rect 46917 96637 46995 96683
rect 47041 96637 47119 96683
rect 47165 96637 47243 96683
rect 47289 96637 47367 96683
rect 47413 96637 47491 96683
rect 47537 96637 47615 96683
rect 47661 96637 47739 96683
rect 47785 96637 47863 96683
rect 47909 96637 47987 96683
rect 48033 96637 48111 96683
rect 48157 96637 48235 96683
rect 48281 96637 48359 96683
rect 48405 96637 48483 96683
rect 48529 96637 48607 96683
rect 48653 96637 48731 96683
rect 48777 96637 48855 96683
rect 48901 96637 48979 96683
rect 49025 96637 49103 96683
rect 49149 96637 49227 96683
rect 49273 96637 49351 96683
rect 49397 96637 49475 96683
rect 49521 96637 49599 96683
rect 49645 96637 49723 96683
rect 49769 96637 49847 96683
rect 49893 96637 49971 96683
rect 50017 96637 50095 96683
rect 50141 96637 50219 96683
rect 50265 96637 50343 96683
rect 50389 96637 50467 96683
rect 50513 96637 50591 96683
rect 50637 96637 50715 96683
rect 50761 96637 50839 96683
rect 50885 96637 50963 96683
rect 51009 96637 51087 96683
rect 51133 96637 51211 96683
rect 51257 96637 51335 96683
rect 51381 96637 51459 96683
rect 51505 96637 51583 96683
rect 51629 96637 51707 96683
rect 51753 96637 51831 96683
rect 51877 96637 51955 96683
rect 52001 96637 52079 96683
rect 52125 96637 52203 96683
rect 52249 96637 52327 96683
rect 52373 96637 52451 96683
rect 52497 96637 52575 96683
rect 52621 96637 52699 96683
rect 52745 96637 52823 96683
rect 52869 96637 52947 96683
rect 52993 96637 53071 96683
rect 53117 96637 53195 96683
rect 53241 96637 53319 96683
rect 53365 96637 53443 96683
rect 53489 96637 53567 96683
rect 53613 96637 53691 96683
rect 53737 96637 53815 96683
rect 53861 96637 53939 96683
rect 53985 96637 54063 96683
rect 54109 96637 54187 96683
rect 54233 96637 54311 96683
rect 54357 96637 54435 96683
rect 54481 96637 54559 96683
rect 54605 96637 54683 96683
rect 54729 96637 54807 96683
rect 54853 96637 54931 96683
rect 54977 96637 55055 96683
rect 55101 96637 55179 96683
rect 55225 96637 55303 96683
rect 55349 96637 55427 96683
rect 55473 96637 55551 96683
rect 55597 96637 55675 96683
rect 55721 96637 55799 96683
rect 55845 96637 55923 96683
rect 55969 96637 56047 96683
rect 56093 96637 56171 96683
rect 56217 96637 56295 96683
rect 56341 96637 56419 96683
rect 56465 96637 56543 96683
rect 56589 96637 56667 96683
rect 56713 96637 56791 96683
rect 56837 96637 56915 96683
rect 56961 96637 57039 96683
rect 57085 96637 57163 96683
rect 57209 96637 57287 96683
rect 57333 96637 57411 96683
rect 57457 96637 57535 96683
rect 57581 96637 57659 96683
rect 57705 96637 57783 96683
rect 57829 96637 57907 96683
rect 57953 96637 58031 96683
rect 58077 96637 58155 96683
rect 58201 96637 58279 96683
rect 58325 96637 58403 96683
rect 58449 96637 58527 96683
rect 58573 96637 58651 96683
rect 58697 96637 58775 96683
rect 58821 96637 58899 96683
rect 58945 96637 59023 96683
rect 59069 96637 59147 96683
rect 59193 96637 59271 96683
rect 59317 96637 59395 96683
rect 59441 96637 59519 96683
rect 59565 96637 59643 96683
rect 59689 96637 59767 96683
rect 59813 96637 59891 96683
rect 59937 96637 60015 96683
rect 60061 96637 60139 96683
rect 60185 96637 60263 96683
rect 60309 96637 60387 96683
rect 60433 96637 60511 96683
rect 60557 96637 60635 96683
rect 60681 96637 60759 96683
rect 60805 96637 60883 96683
rect 60929 96637 61007 96683
rect 61053 96637 61131 96683
rect 61177 96637 61255 96683
rect 61301 96637 61379 96683
rect 61425 96637 61503 96683
rect 61549 96637 61627 96683
rect 61673 96637 61751 96683
rect 61797 96637 61875 96683
rect 61921 96637 61999 96683
rect 62045 96637 62123 96683
rect 62169 96637 62247 96683
rect 62293 96637 62371 96683
rect 62417 96637 62495 96683
rect 62541 96637 62619 96683
rect 62665 96637 62743 96683
rect 62789 96637 62867 96683
rect 62913 96637 62991 96683
rect 63037 96637 63115 96683
rect 63161 96637 63239 96683
rect 63285 96637 63363 96683
rect 63409 96637 63487 96683
rect 63533 96637 63611 96683
rect 63657 96637 63735 96683
rect 63781 96637 63859 96683
rect 63905 96637 63983 96683
rect 64029 96637 64107 96683
rect 64153 96637 64231 96683
rect 64277 96637 64355 96683
rect 64401 96637 64479 96683
rect 64525 96637 64603 96683
rect 64649 96637 64727 96683
rect 64773 96637 64851 96683
rect 64897 96637 64975 96683
rect 65021 96637 65099 96683
rect 65145 96637 65223 96683
rect 65269 96637 65347 96683
rect 65393 96637 65471 96683
rect 65517 96637 65595 96683
rect 65641 96637 65719 96683
rect 65765 96637 65843 96683
rect 65889 96637 65967 96683
rect 66013 96637 66091 96683
rect 66137 96637 66215 96683
rect 66261 96637 66339 96683
rect 66385 96637 66463 96683
rect 66509 96637 66587 96683
rect 66633 96637 66711 96683
rect 66757 96637 66835 96683
rect 66881 96637 66959 96683
rect 67005 96637 67083 96683
rect 67129 96637 67207 96683
rect 67253 96637 67331 96683
rect 67377 96637 67455 96683
rect 67501 96637 67579 96683
rect 67625 96637 67703 96683
rect 67749 96637 67827 96683
rect 67873 96637 67951 96683
rect 67997 96637 68075 96683
rect 68121 96637 68199 96683
rect 68245 96637 68323 96683
rect 68369 96637 68447 96683
rect 68493 96637 68571 96683
rect 68617 96637 68695 96683
rect 68741 96637 68819 96683
rect 68865 96637 68943 96683
rect 68989 96637 69067 96683
rect 69113 96637 69191 96683
rect 69237 96637 69315 96683
rect 69361 96637 69439 96683
rect 69485 96637 69563 96683
rect 69609 96637 69687 96683
rect 69733 96637 69811 96683
rect 69857 96637 69935 96683
rect 69981 96637 70059 96683
rect 70105 96637 70183 96683
rect 70229 96637 70307 96683
rect 70353 96637 70431 96683
rect 70477 96637 70555 96683
rect 70601 96637 70679 96683
rect 70725 96637 70803 96683
rect 70849 96637 70927 96683
rect 70973 96637 71051 96683
rect 71097 96637 71175 96683
rect 71221 96637 71299 96683
rect 71345 96637 71423 96683
rect 71469 96637 71547 96683
rect 71593 96637 71671 96683
rect 71717 96637 71795 96683
rect 71841 96637 71919 96683
rect 71965 96637 72043 96683
rect 72089 96637 72167 96683
rect 72213 96637 72291 96683
rect 72337 96637 72415 96683
rect 72461 96637 72539 96683
rect 72585 96637 72663 96683
rect 72709 96637 72787 96683
rect 72833 96637 72911 96683
rect 72957 96637 73035 96683
rect 73081 96637 73159 96683
rect 73205 96637 73283 96683
rect 73329 96637 73407 96683
rect 73453 96637 73531 96683
rect 73577 96637 73655 96683
rect 73701 96637 73779 96683
rect 73825 96637 73903 96683
rect 73949 96637 74027 96683
rect 74073 96637 74151 96683
rect 74197 96637 74275 96683
rect 74321 96637 74399 96683
rect 74445 96637 74523 96683
rect 74569 96637 74647 96683
rect 74693 96637 74771 96683
rect 74817 96637 74895 96683
rect 74941 96637 75019 96683
rect 75065 96637 75143 96683
rect 75189 96637 75267 96683
rect 75313 96637 75391 96683
rect 75437 96637 75515 96683
rect 75561 96637 75639 96683
rect 75685 96637 75763 96683
rect 75809 96637 75887 96683
rect 75933 96637 76011 96683
rect 76057 96637 76135 96683
rect 76181 96637 76259 96683
rect 76305 96637 76383 96683
rect 76429 96637 76507 96683
rect 76553 96637 76631 96683
rect 76677 96637 76755 96683
rect 76801 96637 76879 96683
rect 76925 96637 77003 96683
rect 77049 96637 77127 96683
rect 77173 96637 77251 96683
rect 77297 96637 77375 96683
rect 77421 96637 77499 96683
rect 77545 96637 77623 96683
rect 77669 96637 77747 96683
rect 77793 96637 77871 96683
rect 77917 96637 77995 96683
rect 78041 96637 78119 96683
rect 78165 96637 78243 96683
rect 78289 96637 78367 96683
rect 78413 96637 78491 96683
rect 78537 96637 78615 96683
rect 78661 96637 78739 96683
rect 78785 96637 78863 96683
rect 78909 96637 78987 96683
rect 79033 96637 79111 96683
rect 79157 96637 79235 96683
rect 79281 96637 79359 96683
rect 79405 96637 79483 96683
rect 79529 96637 79607 96683
rect 79653 96637 79731 96683
rect 79777 96637 79855 96683
rect 79901 96637 79979 96683
rect 80025 96637 80103 96683
rect 80149 96637 80227 96683
rect 80273 96637 80351 96683
rect 80397 96637 80475 96683
rect 80521 96637 80599 96683
rect 80645 96637 80723 96683
rect 80769 96637 80847 96683
rect 80893 96637 80971 96683
rect 81017 96637 81095 96683
rect 81141 96637 81219 96683
rect 81265 96637 81343 96683
rect 81389 96637 81467 96683
rect 81513 96637 81591 96683
rect 81637 96637 81715 96683
rect 81761 96637 81839 96683
rect 81885 96637 81963 96683
rect 82009 96637 82087 96683
rect 82133 96637 82211 96683
rect 82257 96637 82335 96683
rect 82381 96637 82459 96683
rect 82505 96637 82583 96683
rect 82629 96637 82707 96683
rect 82753 96637 82831 96683
rect 82877 96637 82955 96683
rect 83001 96637 83079 96683
rect 83125 96637 83203 96683
rect 83249 96637 83327 96683
rect 83373 96637 83451 96683
rect 83497 96637 83575 96683
rect 83621 96637 83699 96683
rect 83745 96637 83823 96683
rect 83869 96637 83947 96683
rect 83993 96637 84071 96683
rect 84117 96637 84195 96683
rect 84241 96637 84319 96683
rect 84365 96637 84443 96683
rect 84489 96637 84567 96683
rect 84613 96637 84691 96683
rect 84737 96637 84815 96683
rect 84861 96637 84939 96683
rect 84985 96637 85063 96683
rect 85109 96637 85187 96683
rect 85233 96637 85311 96683
rect 85357 96637 85435 96683
rect 85481 96637 85559 96683
rect 85605 96637 85683 96683
rect 85729 96637 85807 96683
rect 85853 96637 85931 96683
rect 85977 96637 86098 96683
rect 352 96559 86098 96637
rect 352 96513 371 96559
rect 417 96513 495 96559
rect 541 96513 619 96559
rect 665 96513 743 96559
rect 789 96513 867 96559
rect 913 96513 991 96559
rect 1037 96513 1115 96559
rect 1161 96513 1239 96559
rect 1285 96513 1363 96559
rect 1409 96513 1487 96559
rect 1533 96513 1611 96559
rect 1657 96513 1735 96559
rect 1781 96513 1859 96559
rect 1905 96513 1983 96559
rect 2029 96513 2107 96559
rect 2153 96513 2231 96559
rect 2277 96513 2355 96559
rect 2401 96513 2479 96559
rect 2525 96513 2603 96559
rect 2649 96513 2727 96559
rect 2773 96513 2851 96559
rect 2897 96513 2975 96559
rect 3021 96513 3099 96559
rect 3145 96513 3223 96559
rect 3269 96513 3347 96559
rect 3393 96513 3471 96559
rect 3517 96513 3595 96559
rect 3641 96513 3719 96559
rect 3765 96513 3843 96559
rect 3889 96513 3967 96559
rect 4013 96513 4091 96559
rect 4137 96513 4215 96559
rect 4261 96513 4339 96559
rect 4385 96513 4463 96559
rect 4509 96513 4587 96559
rect 4633 96513 4711 96559
rect 4757 96513 4835 96559
rect 4881 96513 4959 96559
rect 5005 96513 5083 96559
rect 5129 96513 5207 96559
rect 5253 96513 5331 96559
rect 5377 96513 5455 96559
rect 5501 96513 5579 96559
rect 5625 96513 5703 96559
rect 5749 96513 5827 96559
rect 5873 96513 5951 96559
rect 5997 96513 6075 96559
rect 6121 96513 6199 96559
rect 6245 96513 6323 96559
rect 6369 96513 6447 96559
rect 6493 96513 6571 96559
rect 6617 96513 6695 96559
rect 6741 96513 6819 96559
rect 6865 96513 6943 96559
rect 6989 96513 7067 96559
rect 7113 96513 7191 96559
rect 7237 96513 7315 96559
rect 7361 96513 7439 96559
rect 7485 96513 7563 96559
rect 7609 96513 7687 96559
rect 7733 96513 7811 96559
rect 7857 96513 7935 96559
rect 7981 96513 8059 96559
rect 8105 96513 8183 96559
rect 8229 96513 8307 96559
rect 8353 96513 8431 96559
rect 8477 96513 8555 96559
rect 8601 96513 8679 96559
rect 8725 96513 8803 96559
rect 8849 96513 8927 96559
rect 8973 96513 9051 96559
rect 9097 96513 9175 96559
rect 9221 96513 9299 96559
rect 9345 96513 9423 96559
rect 9469 96513 9547 96559
rect 9593 96513 9671 96559
rect 9717 96513 9795 96559
rect 9841 96513 9919 96559
rect 9965 96513 10043 96559
rect 10089 96513 10167 96559
rect 10213 96513 10291 96559
rect 10337 96513 10415 96559
rect 10461 96513 10539 96559
rect 10585 96513 10663 96559
rect 10709 96513 10787 96559
rect 10833 96513 10911 96559
rect 10957 96513 11035 96559
rect 11081 96513 11159 96559
rect 11205 96513 11283 96559
rect 11329 96513 11407 96559
rect 11453 96513 11531 96559
rect 11577 96513 11655 96559
rect 11701 96513 11779 96559
rect 11825 96513 11903 96559
rect 11949 96513 12027 96559
rect 12073 96513 12151 96559
rect 12197 96513 12275 96559
rect 12321 96513 12399 96559
rect 12445 96513 12523 96559
rect 12569 96513 12647 96559
rect 12693 96513 12771 96559
rect 12817 96513 12895 96559
rect 12941 96513 13019 96559
rect 13065 96513 13143 96559
rect 13189 96513 13267 96559
rect 13313 96513 13391 96559
rect 13437 96513 13515 96559
rect 13561 96513 13639 96559
rect 13685 96513 13763 96559
rect 13809 96513 13887 96559
rect 13933 96513 14011 96559
rect 14057 96513 14135 96559
rect 14181 96513 14259 96559
rect 14305 96513 14383 96559
rect 14429 96513 14507 96559
rect 14553 96513 14631 96559
rect 14677 96513 14755 96559
rect 14801 96513 14879 96559
rect 14925 96513 15003 96559
rect 15049 96513 15127 96559
rect 15173 96513 15251 96559
rect 15297 96513 15375 96559
rect 15421 96513 15499 96559
rect 15545 96513 15623 96559
rect 15669 96513 15747 96559
rect 15793 96513 15871 96559
rect 15917 96513 15995 96559
rect 16041 96513 16119 96559
rect 16165 96513 16243 96559
rect 16289 96513 16367 96559
rect 16413 96513 16491 96559
rect 16537 96513 16615 96559
rect 16661 96513 16739 96559
rect 16785 96513 16863 96559
rect 16909 96513 16987 96559
rect 17033 96513 17111 96559
rect 17157 96513 17235 96559
rect 17281 96513 17359 96559
rect 17405 96513 17483 96559
rect 17529 96513 17607 96559
rect 17653 96513 17731 96559
rect 17777 96513 17855 96559
rect 17901 96513 17979 96559
rect 18025 96513 18103 96559
rect 18149 96513 18227 96559
rect 18273 96513 18351 96559
rect 18397 96513 18475 96559
rect 18521 96513 18599 96559
rect 18645 96513 18723 96559
rect 18769 96513 18847 96559
rect 18893 96513 18971 96559
rect 19017 96513 19095 96559
rect 19141 96513 19219 96559
rect 19265 96513 19343 96559
rect 19389 96513 19467 96559
rect 19513 96513 19591 96559
rect 19637 96513 19715 96559
rect 19761 96513 19839 96559
rect 19885 96513 19963 96559
rect 20009 96513 20087 96559
rect 20133 96513 20211 96559
rect 20257 96513 20335 96559
rect 20381 96513 20459 96559
rect 20505 96513 20583 96559
rect 20629 96513 20707 96559
rect 20753 96513 20831 96559
rect 20877 96513 20955 96559
rect 21001 96513 21079 96559
rect 21125 96513 21203 96559
rect 21249 96513 21327 96559
rect 21373 96513 21451 96559
rect 21497 96513 21575 96559
rect 21621 96513 21699 96559
rect 21745 96513 21823 96559
rect 21869 96513 21947 96559
rect 21993 96513 22071 96559
rect 22117 96513 22195 96559
rect 22241 96513 22319 96559
rect 22365 96513 22443 96559
rect 22489 96513 22567 96559
rect 22613 96513 22691 96559
rect 22737 96513 22815 96559
rect 22861 96513 22939 96559
rect 22985 96513 23063 96559
rect 23109 96513 23187 96559
rect 23233 96513 23311 96559
rect 23357 96513 23435 96559
rect 23481 96513 23559 96559
rect 23605 96513 23683 96559
rect 23729 96513 23807 96559
rect 23853 96513 23931 96559
rect 23977 96513 24055 96559
rect 24101 96513 24179 96559
rect 24225 96513 24303 96559
rect 24349 96513 24427 96559
rect 24473 96513 24551 96559
rect 24597 96513 24675 96559
rect 24721 96513 24799 96559
rect 24845 96513 24923 96559
rect 24969 96513 25047 96559
rect 25093 96513 25171 96559
rect 25217 96513 25295 96559
rect 25341 96513 25419 96559
rect 25465 96513 25543 96559
rect 25589 96513 25667 96559
rect 25713 96513 25791 96559
rect 25837 96513 25915 96559
rect 25961 96513 26039 96559
rect 26085 96513 26163 96559
rect 26209 96513 26287 96559
rect 26333 96513 26411 96559
rect 26457 96513 26535 96559
rect 26581 96513 26659 96559
rect 26705 96513 26783 96559
rect 26829 96513 26907 96559
rect 26953 96513 27031 96559
rect 27077 96513 27155 96559
rect 27201 96513 27279 96559
rect 27325 96513 27403 96559
rect 27449 96513 27527 96559
rect 27573 96513 27651 96559
rect 27697 96513 27775 96559
rect 27821 96513 27899 96559
rect 27945 96513 28023 96559
rect 28069 96513 28147 96559
rect 28193 96513 28271 96559
rect 28317 96513 28395 96559
rect 28441 96513 28519 96559
rect 28565 96513 28643 96559
rect 28689 96513 28767 96559
rect 28813 96513 28891 96559
rect 28937 96513 29015 96559
rect 29061 96513 29139 96559
rect 29185 96513 29263 96559
rect 29309 96513 29387 96559
rect 29433 96513 29511 96559
rect 29557 96513 29635 96559
rect 29681 96513 29759 96559
rect 29805 96513 29883 96559
rect 29929 96513 30007 96559
rect 30053 96513 30131 96559
rect 30177 96513 30255 96559
rect 30301 96513 30379 96559
rect 30425 96513 30503 96559
rect 30549 96513 30627 96559
rect 30673 96513 30751 96559
rect 30797 96513 30875 96559
rect 30921 96513 30999 96559
rect 31045 96513 31123 96559
rect 31169 96513 31247 96559
rect 31293 96513 31371 96559
rect 31417 96513 31495 96559
rect 31541 96513 31619 96559
rect 31665 96513 31743 96559
rect 31789 96513 31867 96559
rect 31913 96513 31991 96559
rect 32037 96513 32115 96559
rect 32161 96513 32239 96559
rect 32285 96513 32363 96559
rect 32409 96513 32487 96559
rect 32533 96513 32611 96559
rect 32657 96513 32735 96559
rect 32781 96513 32859 96559
rect 32905 96513 32983 96559
rect 33029 96513 33107 96559
rect 33153 96513 33231 96559
rect 33277 96513 33355 96559
rect 33401 96513 33479 96559
rect 33525 96513 33603 96559
rect 33649 96513 33727 96559
rect 33773 96513 33851 96559
rect 33897 96513 33975 96559
rect 34021 96513 34099 96559
rect 34145 96513 34223 96559
rect 34269 96513 34347 96559
rect 34393 96513 34471 96559
rect 34517 96513 34595 96559
rect 34641 96513 34719 96559
rect 34765 96513 34843 96559
rect 34889 96513 34967 96559
rect 35013 96513 35091 96559
rect 35137 96513 35215 96559
rect 35261 96513 35339 96559
rect 35385 96513 35463 96559
rect 35509 96513 35587 96559
rect 35633 96513 35711 96559
rect 35757 96513 35835 96559
rect 35881 96513 35959 96559
rect 36005 96513 36083 96559
rect 36129 96513 36207 96559
rect 36253 96513 36331 96559
rect 36377 96513 36455 96559
rect 36501 96513 36579 96559
rect 36625 96513 36703 96559
rect 36749 96513 36827 96559
rect 36873 96513 36951 96559
rect 36997 96513 37075 96559
rect 37121 96513 37199 96559
rect 37245 96513 37323 96559
rect 37369 96513 37447 96559
rect 37493 96513 37571 96559
rect 37617 96513 37695 96559
rect 37741 96513 37819 96559
rect 37865 96513 37943 96559
rect 37989 96513 38067 96559
rect 38113 96513 38191 96559
rect 38237 96513 38315 96559
rect 38361 96513 38439 96559
rect 38485 96513 38563 96559
rect 38609 96513 38687 96559
rect 38733 96513 38811 96559
rect 38857 96513 38935 96559
rect 38981 96513 39059 96559
rect 39105 96513 39183 96559
rect 39229 96513 39307 96559
rect 39353 96513 39431 96559
rect 39477 96513 39555 96559
rect 39601 96513 39679 96559
rect 39725 96513 39803 96559
rect 39849 96513 39927 96559
rect 39973 96513 40051 96559
rect 40097 96513 40175 96559
rect 40221 96513 40299 96559
rect 40345 96513 40423 96559
rect 40469 96513 40547 96559
rect 40593 96513 40671 96559
rect 40717 96513 40795 96559
rect 40841 96513 40919 96559
rect 40965 96513 41043 96559
rect 41089 96513 41167 96559
rect 41213 96513 41291 96559
rect 41337 96513 41415 96559
rect 41461 96513 41539 96559
rect 41585 96513 41663 96559
rect 41709 96513 41787 96559
rect 41833 96513 41911 96559
rect 41957 96513 42035 96559
rect 42081 96513 42159 96559
rect 42205 96513 42283 96559
rect 42329 96513 42407 96559
rect 42453 96513 42531 96559
rect 42577 96513 42655 96559
rect 42701 96513 42779 96559
rect 42825 96513 42903 96559
rect 42949 96513 43027 96559
rect 43073 96513 43151 96559
rect 43197 96513 43275 96559
rect 43321 96513 43399 96559
rect 43445 96513 43523 96559
rect 43569 96513 43647 96559
rect 43693 96513 43771 96559
rect 43817 96513 43895 96559
rect 43941 96513 44019 96559
rect 44065 96513 44143 96559
rect 44189 96513 44267 96559
rect 44313 96513 44391 96559
rect 44437 96513 44515 96559
rect 44561 96513 44639 96559
rect 44685 96513 44763 96559
rect 44809 96513 44887 96559
rect 44933 96513 45011 96559
rect 45057 96513 45135 96559
rect 45181 96513 45259 96559
rect 45305 96513 45383 96559
rect 45429 96513 45507 96559
rect 45553 96513 45631 96559
rect 45677 96513 45755 96559
rect 45801 96513 45879 96559
rect 45925 96513 46003 96559
rect 46049 96513 46127 96559
rect 46173 96513 46251 96559
rect 46297 96513 46375 96559
rect 46421 96513 46499 96559
rect 46545 96513 46623 96559
rect 46669 96513 46747 96559
rect 46793 96513 46871 96559
rect 46917 96513 46995 96559
rect 47041 96513 47119 96559
rect 47165 96513 47243 96559
rect 47289 96513 47367 96559
rect 47413 96513 47491 96559
rect 47537 96513 47615 96559
rect 47661 96513 47739 96559
rect 47785 96513 47863 96559
rect 47909 96513 47987 96559
rect 48033 96513 48111 96559
rect 48157 96513 48235 96559
rect 48281 96513 48359 96559
rect 48405 96513 48483 96559
rect 48529 96513 48607 96559
rect 48653 96513 48731 96559
rect 48777 96513 48855 96559
rect 48901 96513 48979 96559
rect 49025 96513 49103 96559
rect 49149 96513 49227 96559
rect 49273 96513 49351 96559
rect 49397 96513 49475 96559
rect 49521 96513 49599 96559
rect 49645 96513 49723 96559
rect 49769 96513 49847 96559
rect 49893 96513 49971 96559
rect 50017 96513 50095 96559
rect 50141 96513 50219 96559
rect 50265 96513 50343 96559
rect 50389 96513 50467 96559
rect 50513 96513 50591 96559
rect 50637 96513 50715 96559
rect 50761 96513 50839 96559
rect 50885 96513 50963 96559
rect 51009 96513 51087 96559
rect 51133 96513 51211 96559
rect 51257 96513 51335 96559
rect 51381 96513 51459 96559
rect 51505 96513 51583 96559
rect 51629 96513 51707 96559
rect 51753 96513 51831 96559
rect 51877 96513 51955 96559
rect 52001 96513 52079 96559
rect 52125 96513 52203 96559
rect 52249 96513 52327 96559
rect 52373 96513 52451 96559
rect 52497 96513 52575 96559
rect 52621 96513 52699 96559
rect 52745 96513 52823 96559
rect 52869 96513 52947 96559
rect 52993 96513 53071 96559
rect 53117 96513 53195 96559
rect 53241 96513 53319 96559
rect 53365 96513 53443 96559
rect 53489 96513 53567 96559
rect 53613 96513 53691 96559
rect 53737 96513 53815 96559
rect 53861 96513 53939 96559
rect 53985 96513 54063 96559
rect 54109 96513 54187 96559
rect 54233 96513 54311 96559
rect 54357 96513 54435 96559
rect 54481 96513 54559 96559
rect 54605 96513 54683 96559
rect 54729 96513 54807 96559
rect 54853 96513 54931 96559
rect 54977 96513 55055 96559
rect 55101 96513 55179 96559
rect 55225 96513 55303 96559
rect 55349 96513 55427 96559
rect 55473 96513 55551 96559
rect 55597 96513 55675 96559
rect 55721 96513 55799 96559
rect 55845 96513 55923 96559
rect 55969 96513 56047 96559
rect 56093 96513 56171 96559
rect 56217 96513 56295 96559
rect 56341 96513 56419 96559
rect 56465 96513 56543 96559
rect 56589 96513 56667 96559
rect 56713 96513 56791 96559
rect 56837 96513 56915 96559
rect 56961 96513 57039 96559
rect 57085 96513 57163 96559
rect 57209 96513 57287 96559
rect 57333 96513 57411 96559
rect 57457 96513 57535 96559
rect 57581 96513 57659 96559
rect 57705 96513 57783 96559
rect 57829 96513 57907 96559
rect 57953 96513 58031 96559
rect 58077 96513 58155 96559
rect 58201 96513 58279 96559
rect 58325 96513 58403 96559
rect 58449 96513 58527 96559
rect 58573 96513 58651 96559
rect 58697 96513 58775 96559
rect 58821 96513 58899 96559
rect 58945 96513 59023 96559
rect 59069 96513 59147 96559
rect 59193 96513 59271 96559
rect 59317 96513 59395 96559
rect 59441 96513 59519 96559
rect 59565 96513 59643 96559
rect 59689 96513 59767 96559
rect 59813 96513 59891 96559
rect 59937 96513 60015 96559
rect 60061 96513 60139 96559
rect 60185 96513 60263 96559
rect 60309 96513 60387 96559
rect 60433 96513 60511 96559
rect 60557 96513 60635 96559
rect 60681 96513 60759 96559
rect 60805 96513 60883 96559
rect 60929 96513 61007 96559
rect 61053 96513 61131 96559
rect 61177 96513 61255 96559
rect 61301 96513 61379 96559
rect 61425 96513 61503 96559
rect 61549 96513 61627 96559
rect 61673 96513 61751 96559
rect 61797 96513 61875 96559
rect 61921 96513 61999 96559
rect 62045 96513 62123 96559
rect 62169 96513 62247 96559
rect 62293 96513 62371 96559
rect 62417 96513 62495 96559
rect 62541 96513 62619 96559
rect 62665 96513 62743 96559
rect 62789 96513 62867 96559
rect 62913 96513 62991 96559
rect 63037 96513 63115 96559
rect 63161 96513 63239 96559
rect 63285 96513 63363 96559
rect 63409 96513 63487 96559
rect 63533 96513 63611 96559
rect 63657 96513 63735 96559
rect 63781 96513 63859 96559
rect 63905 96513 63983 96559
rect 64029 96513 64107 96559
rect 64153 96513 64231 96559
rect 64277 96513 64355 96559
rect 64401 96513 64479 96559
rect 64525 96513 64603 96559
rect 64649 96513 64727 96559
rect 64773 96513 64851 96559
rect 64897 96513 64975 96559
rect 65021 96513 65099 96559
rect 65145 96513 65223 96559
rect 65269 96513 65347 96559
rect 65393 96513 65471 96559
rect 65517 96513 65595 96559
rect 65641 96513 65719 96559
rect 65765 96513 65843 96559
rect 65889 96513 65967 96559
rect 66013 96513 66091 96559
rect 66137 96513 66215 96559
rect 66261 96513 66339 96559
rect 66385 96513 66463 96559
rect 66509 96513 66587 96559
rect 66633 96513 66711 96559
rect 66757 96513 66835 96559
rect 66881 96513 66959 96559
rect 67005 96513 67083 96559
rect 67129 96513 67207 96559
rect 67253 96513 67331 96559
rect 67377 96513 67455 96559
rect 67501 96513 67579 96559
rect 67625 96513 67703 96559
rect 67749 96513 67827 96559
rect 67873 96513 67951 96559
rect 67997 96513 68075 96559
rect 68121 96513 68199 96559
rect 68245 96513 68323 96559
rect 68369 96513 68447 96559
rect 68493 96513 68571 96559
rect 68617 96513 68695 96559
rect 68741 96513 68819 96559
rect 68865 96513 68943 96559
rect 68989 96513 69067 96559
rect 69113 96513 69191 96559
rect 69237 96513 69315 96559
rect 69361 96513 69439 96559
rect 69485 96513 69563 96559
rect 69609 96513 69687 96559
rect 69733 96513 69811 96559
rect 69857 96513 69935 96559
rect 69981 96513 70059 96559
rect 70105 96513 70183 96559
rect 70229 96513 70307 96559
rect 70353 96513 70431 96559
rect 70477 96513 70555 96559
rect 70601 96513 70679 96559
rect 70725 96513 70803 96559
rect 70849 96513 70927 96559
rect 70973 96513 71051 96559
rect 71097 96513 71175 96559
rect 71221 96513 71299 96559
rect 71345 96513 71423 96559
rect 71469 96513 71547 96559
rect 71593 96513 71671 96559
rect 71717 96513 71795 96559
rect 71841 96513 71919 96559
rect 71965 96513 72043 96559
rect 72089 96513 72167 96559
rect 72213 96513 72291 96559
rect 72337 96513 72415 96559
rect 72461 96513 72539 96559
rect 72585 96513 72663 96559
rect 72709 96513 72787 96559
rect 72833 96513 72911 96559
rect 72957 96513 73035 96559
rect 73081 96513 73159 96559
rect 73205 96513 73283 96559
rect 73329 96513 73407 96559
rect 73453 96513 73531 96559
rect 73577 96513 73655 96559
rect 73701 96513 73779 96559
rect 73825 96513 73903 96559
rect 73949 96513 74027 96559
rect 74073 96513 74151 96559
rect 74197 96513 74275 96559
rect 74321 96513 74399 96559
rect 74445 96513 74523 96559
rect 74569 96513 74647 96559
rect 74693 96513 74771 96559
rect 74817 96513 74895 96559
rect 74941 96513 75019 96559
rect 75065 96513 75143 96559
rect 75189 96513 75267 96559
rect 75313 96513 75391 96559
rect 75437 96513 75515 96559
rect 75561 96513 75639 96559
rect 75685 96513 75763 96559
rect 75809 96513 75887 96559
rect 75933 96513 76011 96559
rect 76057 96513 76135 96559
rect 76181 96513 76259 96559
rect 76305 96513 76383 96559
rect 76429 96513 76507 96559
rect 76553 96513 76631 96559
rect 76677 96513 76755 96559
rect 76801 96513 76879 96559
rect 76925 96513 77003 96559
rect 77049 96513 77127 96559
rect 77173 96513 77251 96559
rect 77297 96513 77375 96559
rect 77421 96513 77499 96559
rect 77545 96513 77623 96559
rect 77669 96513 77747 96559
rect 77793 96513 77871 96559
rect 77917 96513 77995 96559
rect 78041 96513 78119 96559
rect 78165 96513 78243 96559
rect 78289 96513 78367 96559
rect 78413 96513 78491 96559
rect 78537 96513 78615 96559
rect 78661 96513 78739 96559
rect 78785 96513 78863 96559
rect 78909 96513 78987 96559
rect 79033 96513 79111 96559
rect 79157 96513 79235 96559
rect 79281 96513 79359 96559
rect 79405 96513 79483 96559
rect 79529 96513 79607 96559
rect 79653 96513 79731 96559
rect 79777 96513 79855 96559
rect 79901 96513 79979 96559
rect 80025 96513 80103 96559
rect 80149 96513 80227 96559
rect 80273 96513 80351 96559
rect 80397 96513 80475 96559
rect 80521 96513 80599 96559
rect 80645 96513 80723 96559
rect 80769 96513 80847 96559
rect 80893 96513 80971 96559
rect 81017 96513 81095 96559
rect 81141 96513 81219 96559
rect 81265 96513 81343 96559
rect 81389 96513 81467 96559
rect 81513 96513 81591 96559
rect 81637 96513 81715 96559
rect 81761 96513 81839 96559
rect 81885 96513 81963 96559
rect 82009 96513 82087 96559
rect 82133 96513 82211 96559
rect 82257 96513 82335 96559
rect 82381 96513 82459 96559
rect 82505 96513 82583 96559
rect 82629 96513 82707 96559
rect 82753 96513 82831 96559
rect 82877 96513 82955 96559
rect 83001 96513 83079 96559
rect 83125 96513 83203 96559
rect 83249 96513 83327 96559
rect 83373 96513 83451 96559
rect 83497 96513 83575 96559
rect 83621 96513 83699 96559
rect 83745 96513 83823 96559
rect 83869 96513 83947 96559
rect 83993 96513 84071 96559
rect 84117 96513 84195 96559
rect 84241 96513 84319 96559
rect 84365 96513 84443 96559
rect 84489 96513 84567 96559
rect 84613 96513 84691 96559
rect 84737 96513 84815 96559
rect 84861 96513 84939 96559
rect 84985 96513 85063 96559
rect 85109 96513 85187 96559
rect 85233 96513 85311 96559
rect 85357 96513 85435 96559
rect 85481 96513 85559 96559
rect 85605 96513 85683 96559
rect 85729 96513 85807 96559
rect 85853 96513 85931 96559
rect 85977 96513 86098 96559
rect 352 96435 86098 96513
rect 352 96389 371 96435
rect 417 96389 495 96435
rect 541 96389 619 96435
rect 665 96389 743 96435
rect 789 96389 867 96435
rect 913 96389 991 96435
rect 1037 96389 1115 96435
rect 1161 96389 1239 96435
rect 1285 96389 1363 96435
rect 1409 96389 1487 96435
rect 1533 96389 1611 96435
rect 1657 96389 1735 96435
rect 1781 96389 1859 96435
rect 1905 96389 1983 96435
rect 2029 96389 2107 96435
rect 2153 96389 2231 96435
rect 2277 96389 2355 96435
rect 2401 96389 2479 96435
rect 2525 96389 2603 96435
rect 2649 96389 2727 96435
rect 2773 96389 2851 96435
rect 2897 96389 2975 96435
rect 3021 96389 3099 96435
rect 3145 96389 3223 96435
rect 3269 96389 3347 96435
rect 3393 96389 3471 96435
rect 3517 96389 3595 96435
rect 3641 96389 3719 96435
rect 3765 96389 3843 96435
rect 3889 96389 3967 96435
rect 4013 96389 4091 96435
rect 4137 96389 4215 96435
rect 4261 96389 4339 96435
rect 4385 96389 4463 96435
rect 4509 96389 4587 96435
rect 4633 96389 4711 96435
rect 4757 96389 4835 96435
rect 4881 96389 4959 96435
rect 5005 96389 5083 96435
rect 5129 96389 5207 96435
rect 5253 96389 5331 96435
rect 5377 96389 5455 96435
rect 5501 96389 5579 96435
rect 5625 96389 5703 96435
rect 5749 96389 5827 96435
rect 5873 96389 5951 96435
rect 5997 96389 6075 96435
rect 6121 96389 6199 96435
rect 6245 96389 6323 96435
rect 6369 96389 6447 96435
rect 6493 96389 6571 96435
rect 6617 96389 6695 96435
rect 6741 96389 6819 96435
rect 6865 96389 6943 96435
rect 6989 96389 7067 96435
rect 7113 96389 7191 96435
rect 7237 96389 7315 96435
rect 7361 96389 7439 96435
rect 7485 96389 7563 96435
rect 7609 96389 7687 96435
rect 7733 96389 7811 96435
rect 7857 96389 7935 96435
rect 7981 96389 8059 96435
rect 8105 96389 8183 96435
rect 8229 96389 8307 96435
rect 8353 96389 8431 96435
rect 8477 96389 8555 96435
rect 8601 96389 8679 96435
rect 8725 96389 8803 96435
rect 8849 96389 8927 96435
rect 8973 96389 9051 96435
rect 9097 96389 9175 96435
rect 9221 96389 9299 96435
rect 9345 96389 9423 96435
rect 9469 96389 9547 96435
rect 9593 96389 9671 96435
rect 9717 96389 9795 96435
rect 9841 96389 9919 96435
rect 9965 96389 10043 96435
rect 10089 96389 10167 96435
rect 10213 96389 10291 96435
rect 10337 96389 10415 96435
rect 10461 96389 10539 96435
rect 10585 96389 10663 96435
rect 10709 96389 10787 96435
rect 10833 96389 10911 96435
rect 10957 96389 11035 96435
rect 11081 96389 11159 96435
rect 11205 96389 11283 96435
rect 11329 96389 11407 96435
rect 11453 96389 11531 96435
rect 11577 96389 11655 96435
rect 11701 96389 11779 96435
rect 11825 96389 11903 96435
rect 11949 96389 12027 96435
rect 12073 96389 12151 96435
rect 12197 96389 12275 96435
rect 12321 96389 12399 96435
rect 12445 96389 12523 96435
rect 12569 96389 12647 96435
rect 12693 96389 12771 96435
rect 12817 96389 12895 96435
rect 12941 96389 13019 96435
rect 13065 96389 13143 96435
rect 13189 96389 13267 96435
rect 13313 96389 13391 96435
rect 13437 96389 13515 96435
rect 13561 96389 13639 96435
rect 13685 96389 13763 96435
rect 13809 96389 13887 96435
rect 13933 96389 14011 96435
rect 14057 96389 14135 96435
rect 14181 96389 14259 96435
rect 14305 96389 14383 96435
rect 14429 96389 14507 96435
rect 14553 96389 14631 96435
rect 14677 96389 14755 96435
rect 14801 96389 14879 96435
rect 14925 96389 15003 96435
rect 15049 96389 15127 96435
rect 15173 96389 15251 96435
rect 15297 96389 15375 96435
rect 15421 96389 15499 96435
rect 15545 96389 15623 96435
rect 15669 96389 15747 96435
rect 15793 96389 15871 96435
rect 15917 96389 15995 96435
rect 16041 96389 16119 96435
rect 16165 96389 16243 96435
rect 16289 96389 16367 96435
rect 16413 96389 16491 96435
rect 16537 96389 16615 96435
rect 16661 96389 16739 96435
rect 16785 96389 16863 96435
rect 16909 96389 16987 96435
rect 17033 96389 17111 96435
rect 17157 96389 17235 96435
rect 17281 96389 17359 96435
rect 17405 96389 17483 96435
rect 17529 96389 17607 96435
rect 17653 96389 17731 96435
rect 17777 96389 17855 96435
rect 17901 96389 17979 96435
rect 18025 96389 18103 96435
rect 18149 96389 18227 96435
rect 18273 96389 18351 96435
rect 18397 96389 18475 96435
rect 18521 96389 18599 96435
rect 18645 96389 18723 96435
rect 18769 96389 18847 96435
rect 18893 96389 18971 96435
rect 19017 96389 19095 96435
rect 19141 96389 19219 96435
rect 19265 96389 19343 96435
rect 19389 96389 19467 96435
rect 19513 96389 19591 96435
rect 19637 96389 19715 96435
rect 19761 96389 19839 96435
rect 19885 96389 19963 96435
rect 20009 96389 20087 96435
rect 20133 96389 20211 96435
rect 20257 96389 20335 96435
rect 20381 96389 20459 96435
rect 20505 96389 20583 96435
rect 20629 96389 20707 96435
rect 20753 96389 20831 96435
rect 20877 96389 20955 96435
rect 21001 96389 21079 96435
rect 21125 96389 21203 96435
rect 21249 96389 21327 96435
rect 21373 96389 21451 96435
rect 21497 96389 21575 96435
rect 21621 96389 21699 96435
rect 21745 96389 21823 96435
rect 21869 96389 21947 96435
rect 21993 96389 22071 96435
rect 22117 96389 22195 96435
rect 22241 96389 22319 96435
rect 22365 96389 22443 96435
rect 22489 96389 22567 96435
rect 22613 96389 22691 96435
rect 22737 96389 22815 96435
rect 22861 96389 22939 96435
rect 22985 96389 23063 96435
rect 23109 96389 23187 96435
rect 23233 96389 23311 96435
rect 23357 96389 23435 96435
rect 23481 96389 23559 96435
rect 23605 96389 23683 96435
rect 23729 96389 23807 96435
rect 23853 96389 23931 96435
rect 23977 96389 24055 96435
rect 24101 96389 24179 96435
rect 24225 96389 24303 96435
rect 24349 96389 24427 96435
rect 24473 96389 24551 96435
rect 24597 96389 24675 96435
rect 24721 96389 24799 96435
rect 24845 96389 24923 96435
rect 24969 96389 25047 96435
rect 25093 96389 25171 96435
rect 25217 96389 25295 96435
rect 25341 96389 25419 96435
rect 25465 96389 25543 96435
rect 25589 96389 25667 96435
rect 25713 96389 25791 96435
rect 25837 96389 25915 96435
rect 25961 96389 26039 96435
rect 26085 96389 26163 96435
rect 26209 96389 26287 96435
rect 26333 96389 26411 96435
rect 26457 96389 26535 96435
rect 26581 96389 26659 96435
rect 26705 96389 26783 96435
rect 26829 96389 26907 96435
rect 26953 96389 27031 96435
rect 27077 96389 27155 96435
rect 27201 96389 27279 96435
rect 27325 96389 27403 96435
rect 27449 96389 27527 96435
rect 27573 96389 27651 96435
rect 27697 96389 27775 96435
rect 27821 96389 27899 96435
rect 27945 96389 28023 96435
rect 28069 96389 28147 96435
rect 28193 96389 28271 96435
rect 28317 96389 28395 96435
rect 28441 96389 28519 96435
rect 28565 96389 28643 96435
rect 28689 96389 28767 96435
rect 28813 96389 28891 96435
rect 28937 96389 29015 96435
rect 29061 96389 29139 96435
rect 29185 96389 29263 96435
rect 29309 96389 29387 96435
rect 29433 96389 29511 96435
rect 29557 96389 29635 96435
rect 29681 96389 29759 96435
rect 29805 96389 29883 96435
rect 29929 96389 30007 96435
rect 30053 96389 30131 96435
rect 30177 96389 30255 96435
rect 30301 96389 30379 96435
rect 30425 96389 30503 96435
rect 30549 96389 30627 96435
rect 30673 96389 30751 96435
rect 30797 96389 30875 96435
rect 30921 96389 30999 96435
rect 31045 96389 31123 96435
rect 31169 96389 31247 96435
rect 31293 96389 31371 96435
rect 31417 96389 31495 96435
rect 31541 96389 31619 96435
rect 31665 96389 31743 96435
rect 31789 96389 31867 96435
rect 31913 96389 31991 96435
rect 32037 96389 32115 96435
rect 32161 96389 32239 96435
rect 32285 96389 32363 96435
rect 32409 96389 32487 96435
rect 32533 96389 32611 96435
rect 32657 96389 32735 96435
rect 32781 96389 32859 96435
rect 32905 96389 32983 96435
rect 33029 96389 33107 96435
rect 33153 96389 33231 96435
rect 33277 96389 33355 96435
rect 33401 96389 33479 96435
rect 33525 96389 33603 96435
rect 33649 96389 33727 96435
rect 33773 96389 33851 96435
rect 33897 96389 33975 96435
rect 34021 96389 34099 96435
rect 34145 96389 34223 96435
rect 34269 96389 34347 96435
rect 34393 96389 34471 96435
rect 34517 96389 34595 96435
rect 34641 96389 34719 96435
rect 34765 96389 34843 96435
rect 34889 96389 34967 96435
rect 35013 96389 35091 96435
rect 35137 96389 35215 96435
rect 35261 96389 35339 96435
rect 35385 96389 35463 96435
rect 35509 96389 35587 96435
rect 35633 96389 35711 96435
rect 35757 96389 35835 96435
rect 35881 96389 35959 96435
rect 36005 96389 36083 96435
rect 36129 96389 36207 96435
rect 36253 96389 36331 96435
rect 36377 96389 36455 96435
rect 36501 96389 36579 96435
rect 36625 96389 36703 96435
rect 36749 96389 36827 96435
rect 36873 96389 36951 96435
rect 36997 96389 37075 96435
rect 37121 96389 37199 96435
rect 37245 96389 37323 96435
rect 37369 96389 37447 96435
rect 37493 96389 37571 96435
rect 37617 96389 37695 96435
rect 37741 96389 37819 96435
rect 37865 96389 37943 96435
rect 37989 96389 38067 96435
rect 38113 96389 38191 96435
rect 38237 96389 38315 96435
rect 38361 96389 38439 96435
rect 38485 96389 38563 96435
rect 38609 96389 38687 96435
rect 38733 96389 38811 96435
rect 38857 96389 38935 96435
rect 38981 96389 39059 96435
rect 39105 96389 39183 96435
rect 39229 96389 39307 96435
rect 39353 96389 39431 96435
rect 39477 96389 39555 96435
rect 39601 96389 39679 96435
rect 39725 96389 39803 96435
rect 39849 96389 39927 96435
rect 39973 96389 40051 96435
rect 40097 96389 40175 96435
rect 40221 96389 40299 96435
rect 40345 96389 40423 96435
rect 40469 96389 40547 96435
rect 40593 96389 40671 96435
rect 40717 96389 40795 96435
rect 40841 96389 40919 96435
rect 40965 96389 41043 96435
rect 41089 96389 41167 96435
rect 41213 96389 41291 96435
rect 41337 96389 41415 96435
rect 41461 96389 41539 96435
rect 41585 96389 41663 96435
rect 41709 96389 41787 96435
rect 41833 96389 41911 96435
rect 41957 96389 42035 96435
rect 42081 96389 42159 96435
rect 42205 96389 42283 96435
rect 42329 96389 42407 96435
rect 42453 96389 42531 96435
rect 42577 96389 42655 96435
rect 42701 96389 42779 96435
rect 42825 96389 42903 96435
rect 42949 96389 43027 96435
rect 43073 96389 43151 96435
rect 43197 96389 43275 96435
rect 43321 96389 43399 96435
rect 43445 96389 43523 96435
rect 43569 96389 43647 96435
rect 43693 96389 43771 96435
rect 43817 96389 43895 96435
rect 43941 96389 44019 96435
rect 44065 96389 44143 96435
rect 44189 96389 44267 96435
rect 44313 96389 44391 96435
rect 44437 96389 44515 96435
rect 44561 96389 44639 96435
rect 44685 96389 44763 96435
rect 44809 96389 44887 96435
rect 44933 96389 45011 96435
rect 45057 96389 45135 96435
rect 45181 96389 45259 96435
rect 45305 96389 45383 96435
rect 45429 96389 45507 96435
rect 45553 96389 45631 96435
rect 45677 96389 45755 96435
rect 45801 96389 45879 96435
rect 45925 96389 46003 96435
rect 46049 96389 46127 96435
rect 46173 96389 46251 96435
rect 46297 96389 46375 96435
rect 46421 96389 46499 96435
rect 46545 96389 46623 96435
rect 46669 96389 46747 96435
rect 46793 96389 46871 96435
rect 46917 96389 46995 96435
rect 47041 96389 47119 96435
rect 47165 96389 47243 96435
rect 47289 96389 47367 96435
rect 47413 96389 47491 96435
rect 47537 96389 47615 96435
rect 47661 96389 47739 96435
rect 47785 96389 47863 96435
rect 47909 96389 47987 96435
rect 48033 96389 48111 96435
rect 48157 96389 48235 96435
rect 48281 96389 48359 96435
rect 48405 96389 48483 96435
rect 48529 96389 48607 96435
rect 48653 96389 48731 96435
rect 48777 96389 48855 96435
rect 48901 96389 48979 96435
rect 49025 96389 49103 96435
rect 49149 96389 49227 96435
rect 49273 96389 49351 96435
rect 49397 96389 49475 96435
rect 49521 96389 49599 96435
rect 49645 96389 49723 96435
rect 49769 96389 49847 96435
rect 49893 96389 49971 96435
rect 50017 96389 50095 96435
rect 50141 96389 50219 96435
rect 50265 96389 50343 96435
rect 50389 96389 50467 96435
rect 50513 96389 50591 96435
rect 50637 96389 50715 96435
rect 50761 96389 50839 96435
rect 50885 96389 50963 96435
rect 51009 96389 51087 96435
rect 51133 96389 51211 96435
rect 51257 96389 51335 96435
rect 51381 96389 51459 96435
rect 51505 96389 51583 96435
rect 51629 96389 51707 96435
rect 51753 96389 51831 96435
rect 51877 96389 51955 96435
rect 52001 96389 52079 96435
rect 52125 96389 52203 96435
rect 52249 96389 52327 96435
rect 52373 96389 52451 96435
rect 52497 96389 52575 96435
rect 52621 96389 52699 96435
rect 52745 96389 52823 96435
rect 52869 96389 52947 96435
rect 52993 96389 53071 96435
rect 53117 96389 53195 96435
rect 53241 96389 53319 96435
rect 53365 96389 53443 96435
rect 53489 96389 53567 96435
rect 53613 96389 53691 96435
rect 53737 96389 53815 96435
rect 53861 96389 53939 96435
rect 53985 96389 54063 96435
rect 54109 96389 54187 96435
rect 54233 96389 54311 96435
rect 54357 96389 54435 96435
rect 54481 96389 54559 96435
rect 54605 96389 54683 96435
rect 54729 96389 54807 96435
rect 54853 96389 54931 96435
rect 54977 96389 55055 96435
rect 55101 96389 55179 96435
rect 55225 96389 55303 96435
rect 55349 96389 55427 96435
rect 55473 96389 55551 96435
rect 55597 96389 55675 96435
rect 55721 96389 55799 96435
rect 55845 96389 55923 96435
rect 55969 96389 56047 96435
rect 56093 96389 56171 96435
rect 56217 96389 56295 96435
rect 56341 96389 56419 96435
rect 56465 96389 56543 96435
rect 56589 96389 56667 96435
rect 56713 96389 56791 96435
rect 56837 96389 56915 96435
rect 56961 96389 57039 96435
rect 57085 96389 57163 96435
rect 57209 96389 57287 96435
rect 57333 96389 57411 96435
rect 57457 96389 57535 96435
rect 57581 96389 57659 96435
rect 57705 96389 57783 96435
rect 57829 96389 57907 96435
rect 57953 96389 58031 96435
rect 58077 96389 58155 96435
rect 58201 96389 58279 96435
rect 58325 96389 58403 96435
rect 58449 96389 58527 96435
rect 58573 96389 58651 96435
rect 58697 96389 58775 96435
rect 58821 96389 58899 96435
rect 58945 96389 59023 96435
rect 59069 96389 59147 96435
rect 59193 96389 59271 96435
rect 59317 96389 59395 96435
rect 59441 96389 59519 96435
rect 59565 96389 59643 96435
rect 59689 96389 59767 96435
rect 59813 96389 59891 96435
rect 59937 96389 60015 96435
rect 60061 96389 60139 96435
rect 60185 96389 60263 96435
rect 60309 96389 60387 96435
rect 60433 96389 60511 96435
rect 60557 96389 60635 96435
rect 60681 96389 60759 96435
rect 60805 96389 60883 96435
rect 60929 96389 61007 96435
rect 61053 96389 61131 96435
rect 61177 96389 61255 96435
rect 61301 96389 61379 96435
rect 61425 96389 61503 96435
rect 61549 96389 61627 96435
rect 61673 96389 61751 96435
rect 61797 96389 61875 96435
rect 61921 96389 61999 96435
rect 62045 96389 62123 96435
rect 62169 96389 62247 96435
rect 62293 96389 62371 96435
rect 62417 96389 62495 96435
rect 62541 96389 62619 96435
rect 62665 96389 62743 96435
rect 62789 96389 62867 96435
rect 62913 96389 62991 96435
rect 63037 96389 63115 96435
rect 63161 96389 63239 96435
rect 63285 96389 63363 96435
rect 63409 96389 63487 96435
rect 63533 96389 63611 96435
rect 63657 96389 63735 96435
rect 63781 96389 63859 96435
rect 63905 96389 63983 96435
rect 64029 96389 64107 96435
rect 64153 96389 64231 96435
rect 64277 96389 64355 96435
rect 64401 96389 64479 96435
rect 64525 96389 64603 96435
rect 64649 96389 64727 96435
rect 64773 96389 64851 96435
rect 64897 96389 64975 96435
rect 65021 96389 65099 96435
rect 65145 96389 65223 96435
rect 65269 96389 65347 96435
rect 65393 96389 65471 96435
rect 65517 96389 65595 96435
rect 65641 96389 65719 96435
rect 65765 96389 65843 96435
rect 65889 96389 65967 96435
rect 66013 96389 66091 96435
rect 66137 96389 66215 96435
rect 66261 96389 66339 96435
rect 66385 96389 66463 96435
rect 66509 96389 66587 96435
rect 66633 96389 66711 96435
rect 66757 96389 66835 96435
rect 66881 96389 66959 96435
rect 67005 96389 67083 96435
rect 67129 96389 67207 96435
rect 67253 96389 67331 96435
rect 67377 96389 67455 96435
rect 67501 96389 67579 96435
rect 67625 96389 67703 96435
rect 67749 96389 67827 96435
rect 67873 96389 67951 96435
rect 67997 96389 68075 96435
rect 68121 96389 68199 96435
rect 68245 96389 68323 96435
rect 68369 96389 68447 96435
rect 68493 96389 68571 96435
rect 68617 96389 68695 96435
rect 68741 96389 68819 96435
rect 68865 96389 68943 96435
rect 68989 96389 69067 96435
rect 69113 96389 69191 96435
rect 69237 96389 69315 96435
rect 69361 96389 69439 96435
rect 69485 96389 69563 96435
rect 69609 96389 69687 96435
rect 69733 96389 69811 96435
rect 69857 96389 69935 96435
rect 69981 96389 70059 96435
rect 70105 96389 70183 96435
rect 70229 96389 70307 96435
rect 70353 96389 70431 96435
rect 70477 96389 70555 96435
rect 70601 96389 70679 96435
rect 70725 96389 70803 96435
rect 70849 96389 70927 96435
rect 70973 96389 71051 96435
rect 71097 96389 71175 96435
rect 71221 96389 71299 96435
rect 71345 96389 71423 96435
rect 71469 96389 71547 96435
rect 71593 96389 71671 96435
rect 71717 96389 71795 96435
rect 71841 96389 71919 96435
rect 71965 96389 72043 96435
rect 72089 96389 72167 96435
rect 72213 96389 72291 96435
rect 72337 96389 72415 96435
rect 72461 96389 72539 96435
rect 72585 96389 72663 96435
rect 72709 96389 72787 96435
rect 72833 96389 72911 96435
rect 72957 96389 73035 96435
rect 73081 96389 73159 96435
rect 73205 96389 73283 96435
rect 73329 96389 73407 96435
rect 73453 96389 73531 96435
rect 73577 96389 73655 96435
rect 73701 96389 73779 96435
rect 73825 96389 73903 96435
rect 73949 96389 74027 96435
rect 74073 96389 74151 96435
rect 74197 96389 74275 96435
rect 74321 96389 74399 96435
rect 74445 96389 74523 96435
rect 74569 96389 74647 96435
rect 74693 96389 74771 96435
rect 74817 96389 74895 96435
rect 74941 96389 75019 96435
rect 75065 96389 75143 96435
rect 75189 96389 75267 96435
rect 75313 96389 75391 96435
rect 75437 96389 75515 96435
rect 75561 96389 75639 96435
rect 75685 96389 75763 96435
rect 75809 96389 75887 96435
rect 75933 96389 76011 96435
rect 76057 96389 76135 96435
rect 76181 96389 76259 96435
rect 76305 96389 76383 96435
rect 76429 96389 76507 96435
rect 76553 96389 76631 96435
rect 76677 96389 76755 96435
rect 76801 96389 76879 96435
rect 76925 96389 77003 96435
rect 77049 96389 77127 96435
rect 77173 96389 77251 96435
rect 77297 96389 77375 96435
rect 77421 96389 77499 96435
rect 77545 96389 77623 96435
rect 77669 96389 77747 96435
rect 77793 96389 77871 96435
rect 77917 96389 77995 96435
rect 78041 96389 78119 96435
rect 78165 96389 78243 96435
rect 78289 96389 78367 96435
rect 78413 96389 78491 96435
rect 78537 96389 78615 96435
rect 78661 96389 78739 96435
rect 78785 96389 78863 96435
rect 78909 96389 78987 96435
rect 79033 96389 79111 96435
rect 79157 96389 79235 96435
rect 79281 96389 79359 96435
rect 79405 96389 79483 96435
rect 79529 96389 79607 96435
rect 79653 96389 79731 96435
rect 79777 96389 79855 96435
rect 79901 96389 79979 96435
rect 80025 96389 80103 96435
rect 80149 96389 80227 96435
rect 80273 96389 80351 96435
rect 80397 96389 80475 96435
rect 80521 96389 80599 96435
rect 80645 96389 80723 96435
rect 80769 96389 80847 96435
rect 80893 96389 80971 96435
rect 81017 96389 81095 96435
rect 81141 96389 81219 96435
rect 81265 96389 81343 96435
rect 81389 96389 81467 96435
rect 81513 96389 81591 96435
rect 81637 96389 81715 96435
rect 81761 96389 81839 96435
rect 81885 96389 81963 96435
rect 82009 96389 82087 96435
rect 82133 96389 82211 96435
rect 82257 96389 82335 96435
rect 82381 96389 82459 96435
rect 82505 96389 82583 96435
rect 82629 96389 82707 96435
rect 82753 96389 82831 96435
rect 82877 96389 82955 96435
rect 83001 96389 83079 96435
rect 83125 96389 83203 96435
rect 83249 96389 83327 96435
rect 83373 96389 83451 96435
rect 83497 96389 83575 96435
rect 83621 96389 83699 96435
rect 83745 96389 83823 96435
rect 83869 96389 83947 96435
rect 83993 96389 84071 96435
rect 84117 96389 84195 96435
rect 84241 96389 84319 96435
rect 84365 96389 84443 96435
rect 84489 96389 84567 96435
rect 84613 96389 84691 96435
rect 84737 96389 84815 96435
rect 84861 96389 84939 96435
rect 84985 96389 85063 96435
rect 85109 96389 85187 96435
rect 85233 96389 85311 96435
rect 85357 96389 85435 96435
rect 85481 96389 85559 96435
rect 85605 96389 85683 96435
rect 85729 96389 85807 96435
rect 85853 96389 85931 96435
rect 85977 96389 86098 96435
rect 352 96311 86098 96389
rect 352 96265 371 96311
rect 417 96265 495 96311
rect 541 96265 619 96311
rect 665 96265 743 96311
rect 789 96265 867 96311
rect 913 96265 991 96311
rect 1037 96265 1115 96311
rect 1161 96265 1239 96311
rect 1285 96265 1363 96311
rect 1409 96265 1487 96311
rect 1533 96265 1611 96311
rect 1657 96265 1735 96311
rect 1781 96265 1859 96311
rect 1905 96265 1983 96311
rect 2029 96265 2107 96311
rect 2153 96265 2231 96311
rect 2277 96265 2355 96311
rect 2401 96265 2479 96311
rect 2525 96265 2603 96311
rect 2649 96265 2727 96311
rect 2773 96265 2851 96311
rect 2897 96265 2975 96311
rect 3021 96265 3099 96311
rect 3145 96265 3223 96311
rect 3269 96265 3347 96311
rect 3393 96265 3471 96311
rect 3517 96265 3595 96311
rect 3641 96265 3719 96311
rect 3765 96265 3843 96311
rect 3889 96265 3967 96311
rect 4013 96265 4091 96311
rect 4137 96265 4215 96311
rect 4261 96265 4339 96311
rect 4385 96265 4463 96311
rect 4509 96265 4587 96311
rect 4633 96265 4711 96311
rect 4757 96265 4835 96311
rect 4881 96265 4959 96311
rect 5005 96265 5083 96311
rect 5129 96265 5207 96311
rect 5253 96265 5331 96311
rect 5377 96265 5455 96311
rect 5501 96265 5579 96311
rect 5625 96265 5703 96311
rect 5749 96265 5827 96311
rect 5873 96265 5951 96311
rect 5997 96265 6075 96311
rect 6121 96265 6199 96311
rect 6245 96265 6323 96311
rect 6369 96265 6447 96311
rect 6493 96265 6571 96311
rect 6617 96265 6695 96311
rect 6741 96265 6819 96311
rect 6865 96265 6943 96311
rect 6989 96265 7067 96311
rect 7113 96265 7191 96311
rect 7237 96265 7315 96311
rect 7361 96265 7439 96311
rect 7485 96265 7563 96311
rect 7609 96265 7687 96311
rect 7733 96265 7811 96311
rect 7857 96265 7935 96311
rect 7981 96265 8059 96311
rect 8105 96265 8183 96311
rect 8229 96265 8307 96311
rect 8353 96265 8431 96311
rect 8477 96265 8555 96311
rect 8601 96265 8679 96311
rect 8725 96265 8803 96311
rect 8849 96265 8927 96311
rect 8973 96265 9051 96311
rect 9097 96265 9175 96311
rect 9221 96265 9299 96311
rect 9345 96265 9423 96311
rect 9469 96265 9547 96311
rect 9593 96265 9671 96311
rect 9717 96265 9795 96311
rect 9841 96265 9919 96311
rect 9965 96265 10043 96311
rect 10089 96265 10167 96311
rect 10213 96265 10291 96311
rect 10337 96265 10415 96311
rect 10461 96265 10539 96311
rect 10585 96265 10663 96311
rect 10709 96265 10787 96311
rect 10833 96265 10911 96311
rect 10957 96265 11035 96311
rect 11081 96265 11159 96311
rect 11205 96265 11283 96311
rect 11329 96265 11407 96311
rect 11453 96265 11531 96311
rect 11577 96265 11655 96311
rect 11701 96265 11779 96311
rect 11825 96265 11903 96311
rect 11949 96265 12027 96311
rect 12073 96265 12151 96311
rect 12197 96265 12275 96311
rect 12321 96265 12399 96311
rect 12445 96265 12523 96311
rect 12569 96265 12647 96311
rect 12693 96265 12771 96311
rect 12817 96265 12895 96311
rect 12941 96265 13019 96311
rect 13065 96265 13143 96311
rect 13189 96265 13267 96311
rect 13313 96265 13391 96311
rect 13437 96265 13515 96311
rect 13561 96265 13639 96311
rect 13685 96265 13763 96311
rect 13809 96265 13887 96311
rect 13933 96265 14011 96311
rect 14057 96265 14135 96311
rect 14181 96265 14259 96311
rect 14305 96265 14383 96311
rect 14429 96265 14507 96311
rect 14553 96265 14631 96311
rect 14677 96265 14755 96311
rect 14801 96265 14879 96311
rect 14925 96265 15003 96311
rect 15049 96265 15127 96311
rect 15173 96265 15251 96311
rect 15297 96265 15375 96311
rect 15421 96265 15499 96311
rect 15545 96265 15623 96311
rect 15669 96265 15747 96311
rect 15793 96265 15871 96311
rect 15917 96265 15995 96311
rect 16041 96265 16119 96311
rect 16165 96265 16243 96311
rect 16289 96265 16367 96311
rect 16413 96265 16491 96311
rect 16537 96265 16615 96311
rect 16661 96265 16739 96311
rect 16785 96265 16863 96311
rect 16909 96265 16987 96311
rect 17033 96265 17111 96311
rect 17157 96265 17235 96311
rect 17281 96265 17359 96311
rect 17405 96265 17483 96311
rect 17529 96265 17607 96311
rect 17653 96265 17731 96311
rect 17777 96265 17855 96311
rect 17901 96265 17979 96311
rect 18025 96265 18103 96311
rect 18149 96265 18227 96311
rect 18273 96265 18351 96311
rect 18397 96265 18475 96311
rect 18521 96265 18599 96311
rect 18645 96265 18723 96311
rect 18769 96265 18847 96311
rect 18893 96265 18971 96311
rect 19017 96265 19095 96311
rect 19141 96265 19219 96311
rect 19265 96265 19343 96311
rect 19389 96265 19467 96311
rect 19513 96265 19591 96311
rect 19637 96265 19715 96311
rect 19761 96265 19839 96311
rect 19885 96265 19963 96311
rect 20009 96265 20087 96311
rect 20133 96265 20211 96311
rect 20257 96265 20335 96311
rect 20381 96265 20459 96311
rect 20505 96265 20583 96311
rect 20629 96265 20707 96311
rect 20753 96265 20831 96311
rect 20877 96265 20955 96311
rect 21001 96265 21079 96311
rect 21125 96265 21203 96311
rect 21249 96265 21327 96311
rect 21373 96265 21451 96311
rect 21497 96265 21575 96311
rect 21621 96265 21699 96311
rect 21745 96265 21823 96311
rect 21869 96265 21947 96311
rect 21993 96265 22071 96311
rect 22117 96265 22195 96311
rect 22241 96265 22319 96311
rect 22365 96265 22443 96311
rect 22489 96265 22567 96311
rect 22613 96265 22691 96311
rect 22737 96265 22815 96311
rect 22861 96265 22939 96311
rect 22985 96265 23063 96311
rect 23109 96265 23187 96311
rect 23233 96265 23311 96311
rect 23357 96265 23435 96311
rect 23481 96265 23559 96311
rect 23605 96265 23683 96311
rect 23729 96265 23807 96311
rect 23853 96265 23931 96311
rect 23977 96265 24055 96311
rect 24101 96265 24179 96311
rect 24225 96265 24303 96311
rect 24349 96265 24427 96311
rect 24473 96265 24551 96311
rect 24597 96265 24675 96311
rect 24721 96265 24799 96311
rect 24845 96265 24923 96311
rect 24969 96265 25047 96311
rect 25093 96265 25171 96311
rect 25217 96265 25295 96311
rect 25341 96265 25419 96311
rect 25465 96265 25543 96311
rect 25589 96265 25667 96311
rect 25713 96265 25791 96311
rect 25837 96265 25915 96311
rect 25961 96265 26039 96311
rect 26085 96265 26163 96311
rect 26209 96265 26287 96311
rect 26333 96265 26411 96311
rect 26457 96265 26535 96311
rect 26581 96265 26659 96311
rect 26705 96265 26783 96311
rect 26829 96265 26907 96311
rect 26953 96265 27031 96311
rect 27077 96265 27155 96311
rect 27201 96265 27279 96311
rect 27325 96265 27403 96311
rect 27449 96265 27527 96311
rect 27573 96265 27651 96311
rect 27697 96265 27775 96311
rect 27821 96265 27899 96311
rect 27945 96265 28023 96311
rect 28069 96265 28147 96311
rect 28193 96265 28271 96311
rect 28317 96265 28395 96311
rect 28441 96265 28519 96311
rect 28565 96265 28643 96311
rect 28689 96265 28767 96311
rect 28813 96265 28891 96311
rect 28937 96265 29015 96311
rect 29061 96265 29139 96311
rect 29185 96265 29263 96311
rect 29309 96265 29387 96311
rect 29433 96265 29511 96311
rect 29557 96265 29635 96311
rect 29681 96265 29759 96311
rect 29805 96265 29883 96311
rect 29929 96265 30007 96311
rect 30053 96265 30131 96311
rect 30177 96265 30255 96311
rect 30301 96265 30379 96311
rect 30425 96265 30503 96311
rect 30549 96265 30627 96311
rect 30673 96265 30751 96311
rect 30797 96265 30875 96311
rect 30921 96265 30999 96311
rect 31045 96265 31123 96311
rect 31169 96265 31247 96311
rect 31293 96265 31371 96311
rect 31417 96265 31495 96311
rect 31541 96265 31619 96311
rect 31665 96265 31743 96311
rect 31789 96265 31867 96311
rect 31913 96265 31991 96311
rect 32037 96265 32115 96311
rect 32161 96265 32239 96311
rect 32285 96265 32363 96311
rect 32409 96265 32487 96311
rect 32533 96265 32611 96311
rect 32657 96265 32735 96311
rect 32781 96265 32859 96311
rect 32905 96265 32983 96311
rect 33029 96265 33107 96311
rect 33153 96265 33231 96311
rect 33277 96265 33355 96311
rect 33401 96265 33479 96311
rect 33525 96265 33603 96311
rect 33649 96265 33727 96311
rect 33773 96265 33851 96311
rect 33897 96265 33975 96311
rect 34021 96265 34099 96311
rect 34145 96265 34223 96311
rect 34269 96265 34347 96311
rect 34393 96265 34471 96311
rect 34517 96265 34595 96311
rect 34641 96265 34719 96311
rect 34765 96265 34843 96311
rect 34889 96265 34967 96311
rect 35013 96265 35091 96311
rect 35137 96265 35215 96311
rect 35261 96265 35339 96311
rect 35385 96265 35463 96311
rect 35509 96265 35587 96311
rect 35633 96265 35711 96311
rect 35757 96265 35835 96311
rect 35881 96265 35959 96311
rect 36005 96265 36083 96311
rect 36129 96265 36207 96311
rect 36253 96265 36331 96311
rect 36377 96265 36455 96311
rect 36501 96265 36579 96311
rect 36625 96265 36703 96311
rect 36749 96265 36827 96311
rect 36873 96265 36951 96311
rect 36997 96265 37075 96311
rect 37121 96265 37199 96311
rect 37245 96265 37323 96311
rect 37369 96265 37447 96311
rect 37493 96265 37571 96311
rect 37617 96265 37695 96311
rect 37741 96265 37819 96311
rect 37865 96265 37943 96311
rect 37989 96265 38067 96311
rect 38113 96265 38191 96311
rect 38237 96265 38315 96311
rect 38361 96265 38439 96311
rect 38485 96265 38563 96311
rect 38609 96265 38687 96311
rect 38733 96265 38811 96311
rect 38857 96265 38935 96311
rect 38981 96265 39059 96311
rect 39105 96265 39183 96311
rect 39229 96265 39307 96311
rect 39353 96265 39431 96311
rect 39477 96265 39555 96311
rect 39601 96265 39679 96311
rect 39725 96265 39803 96311
rect 39849 96265 39927 96311
rect 39973 96265 40051 96311
rect 40097 96265 40175 96311
rect 40221 96265 40299 96311
rect 40345 96265 40423 96311
rect 40469 96265 40547 96311
rect 40593 96265 40671 96311
rect 40717 96265 40795 96311
rect 40841 96265 40919 96311
rect 40965 96265 41043 96311
rect 41089 96265 41167 96311
rect 41213 96265 41291 96311
rect 41337 96265 41415 96311
rect 41461 96265 41539 96311
rect 41585 96265 41663 96311
rect 41709 96265 41787 96311
rect 41833 96265 41911 96311
rect 41957 96265 42035 96311
rect 42081 96265 42159 96311
rect 42205 96265 42283 96311
rect 42329 96265 42407 96311
rect 42453 96265 42531 96311
rect 42577 96265 42655 96311
rect 42701 96265 42779 96311
rect 42825 96265 42903 96311
rect 42949 96265 43027 96311
rect 43073 96265 43151 96311
rect 43197 96265 43275 96311
rect 43321 96265 43399 96311
rect 43445 96265 43523 96311
rect 43569 96265 43647 96311
rect 43693 96265 43771 96311
rect 43817 96265 43895 96311
rect 43941 96265 44019 96311
rect 44065 96265 44143 96311
rect 44189 96265 44267 96311
rect 44313 96265 44391 96311
rect 44437 96265 44515 96311
rect 44561 96265 44639 96311
rect 44685 96265 44763 96311
rect 44809 96265 44887 96311
rect 44933 96265 45011 96311
rect 45057 96265 45135 96311
rect 45181 96265 45259 96311
rect 45305 96265 45383 96311
rect 45429 96265 45507 96311
rect 45553 96265 45631 96311
rect 45677 96265 45755 96311
rect 45801 96265 45879 96311
rect 45925 96265 46003 96311
rect 46049 96265 46127 96311
rect 46173 96265 46251 96311
rect 46297 96265 46375 96311
rect 46421 96265 46499 96311
rect 46545 96265 46623 96311
rect 46669 96265 46747 96311
rect 46793 96265 46871 96311
rect 46917 96265 46995 96311
rect 47041 96265 47119 96311
rect 47165 96265 47243 96311
rect 47289 96265 47367 96311
rect 47413 96265 47491 96311
rect 47537 96265 47615 96311
rect 47661 96265 47739 96311
rect 47785 96265 47863 96311
rect 47909 96265 47987 96311
rect 48033 96265 48111 96311
rect 48157 96265 48235 96311
rect 48281 96265 48359 96311
rect 48405 96265 48483 96311
rect 48529 96265 48607 96311
rect 48653 96265 48731 96311
rect 48777 96265 48855 96311
rect 48901 96265 48979 96311
rect 49025 96265 49103 96311
rect 49149 96265 49227 96311
rect 49273 96265 49351 96311
rect 49397 96265 49475 96311
rect 49521 96265 49599 96311
rect 49645 96265 49723 96311
rect 49769 96265 49847 96311
rect 49893 96265 49971 96311
rect 50017 96265 50095 96311
rect 50141 96265 50219 96311
rect 50265 96265 50343 96311
rect 50389 96265 50467 96311
rect 50513 96265 50591 96311
rect 50637 96265 50715 96311
rect 50761 96265 50839 96311
rect 50885 96265 50963 96311
rect 51009 96265 51087 96311
rect 51133 96265 51211 96311
rect 51257 96265 51335 96311
rect 51381 96265 51459 96311
rect 51505 96265 51583 96311
rect 51629 96265 51707 96311
rect 51753 96265 51831 96311
rect 51877 96265 51955 96311
rect 52001 96265 52079 96311
rect 52125 96265 52203 96311
rect 52249 96265 52327 96311
rect 52373 96265 52451 96311
rect 52497 96265 52575 96311
rect 52621 96265 52699 96311
rect 52745 96265 52823 96311
rect 52869 96265 52947 96311
rect 52993 96265 53071 96311
rect 53117 96265 53195 96311
rect 53241 96265 53319 96311
rect 53365 96265 53443 96311
rect 53489 96265 53567 96311
rect 53613 96265 53691 96311
rect 53737 96265 53815 96311
rect 53861 96265 53939 96311
rect 53985 96265 54063 96311
rect 54109 96265 54187 96311
rect 54233 96265 54311 96311
rect 54357 96265 54435 96311
rect 54481 96265 54559 96311
rect 54605 96265 54683 96311
rect 54729 96265 54807 96311
rect 54853 96265 54931 96311
rect 54977 96265 55055 96311
rect 55101 96265 55179 96311
rect 55225 96265 55303 96311
rect 55349 96265 55427 96311
rect 55473 96265 55551 96311
rect 55597 96265 55675 96311
rect 55721 96265 55799 96311
rect 55845 96265 55923 96311
rect 55969 96265 56047 96311
rect 56093 96265 56171 96311
rect 56217 96265 56295 96311
rect 56341 96265 56419 96311
rect 56465 96265 56543 96311
rect 56589 96265 56667 96311
rect 56713 96265 56791 96311
rect 56837 96265 56915 96311
rect 56961 96265 57039 96311
rect 57085 96265 57163 96311
rect 57209 96265 57287 96311
rect 57333 96265 57411 96311
rect 57457 96265 57535 96311
rect 57581 96265 57659 96311
rect 57705 96265 57783 96311
rect 57829 96265 57907 96311
rect 57953 96265 58031 96311
rect 58077 96265 58155 96311
rect 58201 96265 58279 96311
rect 58325 96265 58403 96311
rect 58449 96265 58527 96311
rect 58573 96265 58651 96311
rect 58697 96265 58775 96311
rect 58821 96265 58899 96311
rect 58945 96265 59023 96311
rect 59069 96265 59147 96311
rect 59193 96265 59271 96311
rect 59317 96265 59395 96311
rect 59441 96265 59519 96311
rect 59565 96265 59643 96311
rect 59689 96265 59767 96311
rect 59813 96265 59891 96311
rect 59937 96265 60015 96311
rect 60061 96265 60139 96311
rect 60185 96265 60263 96311
rect 60309 96265 60387 96311
rect 60433 96265 60511 96311
rect 60557 96265 60635 96311
rect 60681 96265 60759 96311
rect 60805 96265 60883 96311
rect 60929 96265 61007 96311
rect 61053 96265 61131 96311
rect 61177 96265 61255 96311
rect 61301 96265 61379 96311
rect 61425 96265 61503 96311
rect 61549 96265 61627 96311
rect 61673 96265 61751 96311
rect 61797 96265 61875 96311
rect 61921 96265 61999 96311
rect 62045 96265 62123 96311
rect 62169 96265 62247 96311
rect 62293 96265 62371 96311
rect 62417 96265 62495 96311
rect 62541 96265 62619 96311
rect 62665 96265 62743 96311
rect 62789 96265 62867 96311
rect 62913 96265 62991 96311
rect 63037 96265 63115 96311
rect 63161 96265 63239 96311
rect 63285 96265 63363 96311
rect 63409 96265 63487 96311
rect 63533 96265 63611 96311
rect 63657 96265 63735 96311
rect 63781 96265 63859 96311
rect 63905 96265 63983 96311
rect 64029 96265 64107 96311
rect 64153 96265 64231 96311
rect 64277 96265 64355 96311
rect 64401 96265 64479 96311
rect 64525 96265 64603 96311
rect 64649 96265 64727 96311
rect 64773 96265 64851 96311
rect 64897 96265 64975 96311
rect 65021 96265 65099 96311
rect 65145 96265 65223 96311
rect 65269 96265 65347 96311
rect 65393 96265 65471 96311
rect 65517 96265 65595 96311
rect 65641 96265 65719 96311
rect 65765 96265 65843 96311
rect 65889 96265 65967 96311
rect 66013 96265 66091 96311
rect 66137 96265 66215 96311
rect 66261 96265 66339 96311
rect 66385 96265 66463 96311
rect 66509 96265 66587 96311
rect 66633 96265 66711 96311
rect 66757 96265 66835 96311
rect 66881 96265 66959 96311
rect 67005 96265 67083 96311
rect 67129 96265 67207 96311
rect 67253 96265 67331 96311
rect 67377 96265 67455 96311
rect 67501 96265 67579 96311
rect 67625 96265 67703 96311
rect 67749 96265 67827 96311
rect 67873 96265 67951 96311
rect 67997 96265 68075 96311
rect 68121 96265 68199 96311
rect 68245 96265 68323 96311
rect 68369 96265 68447 96311
rect 68493 96265 68571 96311
rect 68617 96265 68695 96311
rect 68741 96265 68819 96311
rect 68865 96265 68943 96311
rect 68989 96265 69067 96311
rect 69113 96265 69191 96311
rect 69237 96265 69315 96311
rect 69361 96265 69439 96311
rect 69485 96265 69563 96311
rect 69609 96265 69687 96311
rect 69733 96265 69811 96311
rect 69857 96265 69935 96311
rect 69981 96265 70059 96311
rect 70105 96265 70183 96311
rect 70229 96265 70307 96311
rect 70353 96265 70431 96311
rect 70477 96265 70555 96311
rect 70601 96265 70679 96311
rect 70725 96265 70803 96311
rect 70849 96265 70927 96311
rect 70973 96265 71051 96311
rect 71097 96265 71175 96311
rect 71221 96265 71299 96311
rect 71345 96265 71423 96311
rect 71469 96265 71547 96311
rect 71593 96265 71671 96311
rect 71717 96265 71795 96311
rect 71841 96265 71919 96311
rect 71965 96265 72043 96311
rect 72089 96265 72167 96311
rect 72213 96265 72291 96311
rect 72337 96265 72415 96311
rect 72461 96265 72539 96311
rect 72585 96265 72663 96311
rect 72709 96265 72787 96311
rect 72833 96265 72911 96311
rect 72957 96265 73035 96311
rect 73081 96265 73159 96311
rect 73205 96265 73283 96311
rect 73329 96265 73407 96311
rect 73453 96265 73531 96311
rect 73577 96265 73655 96311
rect 73701 96265 73779 96311
rect 73825 96265 73903 96311
rect 73949 96265 74027 96311
rect 74073 96265 74151 96311
rect 74197 96265 74275 96311
rect 74321 96265 74399 96311
rect 74445 96265 74523 96311
rect 74569 96265 74647 96311
rect 74693 96265 74771 96311
rect 74817 96265 74895 96311
rect 74941 96265 75019 96311
rect 75065 96265 75143 96311
rect 75189 96265 75267 96311
rect 75313 96265 75391 96311
rect 75437 96265 75515 96311
rect 75561 96265 75639 96311
rect 75685 96265 75763 96311
rect 75809 96265 75887 96311
rect 75933 96265 76011 96311
rect 76057 96265 76135 96311
rect 76181 96265 76259 96311
rect 76305 96265 76383 96311
rect 76429 96265 76507 96311
rect 76553 96265 76631 96311
rect 76677 96265 76755 96311
rect 76801 96265 76879 96311
rect 76925 96265 77003 96311
rect 77049 96265 77127 96311
rect 77173 96265 77251 96311
rect 77297 96265 77375 96311
rect 77421 96265 77499 96311
rect 77545 96265 77623 96311
rect 77669 96265 77747 96311
rect 77793 96265 77871 96311
rect 77917 96265 77995 96311
rect 78041 96265 78119 96311
rect 78165 96265 78243 96311
rect 78289 96265 78367 96311
rect 78413 96265 78491 96311
rect 78537 96265 78615 96311
rect 78661 96265 78739 96311
rect 78785 96265 78863 96311
rect 78909 96265 78987 96311
rect 79033 96265 79111 96311
rect 79157 96265 79235 96311
rect 79281 96265 79359 96311
rect 79405 96265 79483 96311
rect 79529 96265 79607 96311
rect 79653 96265 79731 96311
rect 79777 96265 79855 96311
rect 79901 96265 79979 96311
rect 80025 96265 80103 96311
rect 80149 96265 80227 96311
rect 80273 96265 80351 96311
rect 80397 96265 80475 96311
rect 80521 96265 80599 96311
rect 80645 96265 80723 96311
rect 80769 96265 80847 96311
rect 80893 96265 80971 96311
rect 81017 96265 81095 96311
rect 81141 96265 81219 96311
rect 81265 96265 81343 96311
rect 81389 96265 81467 96311
rect 81513 96265 81591 96311
rect 81637 96265 81715 96311
rect 81761 96265 81839 96311
rect 81885 96265 81963 96311
rect 82009 96265 82087 96311
rect 82133 96265 82211 96311
rect 82257 96265 82335 96311
rect 82381 96265 82459 96311
rect 82505 96265 82583 96311
rect 82629 96265 82707 96311
rect 82753 96265 82831 96311
rect 82877 96265 82955 96311
rect 83001 96265 83079 96311
rect 83125 96265 83203 96311
rect 83249 96265 83327 96311
rect 83373 96265 83451 96311
rect 83497 96265 83575 96311
rect 83621 96265 83699 96311
rect 83745 96265 83823 96311
rect 83869 96265 83947 96311
rect 83993 96265 84071 96311
rect 84117 96265 84195 96311
rect 84241 96265 84319 96311
rect 84365 96265 84443 96311
rect 84489 96265 84567 96311
rect 84613 96265 84691 96311
rect 84737 96265 84815 96311
rect 84861 96265 84939 96311
rect 84985 96265 85063 96311
rect 85109 96265 85187 96311
rect 85233 96265 85311 96311
rect 85357 96265 85435 96311
rect 85481 96265 85559 96311
rect 85605 96265 85683 96311
rect 85729 96265 85807 96311
rect 85853 96265 85931 96311
rect 85977 96265 86098 96311
rect 352 96246 86098 96265
rect 352 96163 736 96246
rect 352 1117 371 96163
rect 717 1117 736 96163
rect 352 1034 736 1117
rect 27379 96163 28911 96246
rect 27379 1117 27398 96163
rect 27744 96142 28911 96163
rect 27744 35996 27822 96142
rect 28668 35996 28911 96142
rect 27744 35977 28911 35996
rect 56212 96163 57671 96246
rect 56212 96142 57306 96163
rect 56212 35996 56382 96142
rect 57228 35996 57306 96142
rect 56212 35977 57306 35996
rect 27744 34639 27763 35977
rect 57287 34639 57306 35977
rect 27744 34620 57306 34639
rect 27744 34174 27822 34620
rect 57168 34174 57306 34620
rect 27744 34155 57306 34174
rect 27744 1117 27763 34155
rect 28620 3906 40188 3925
rect 28620 3860 28639 3906
rect 28685 3860 28755 3906
rect 28801 3860 28871 3906
rect 28917 3860 28987 3906
rect 29033 3860 29103 3906
rect 29149 3860 29219 3906
rect 29265 3860 29335 3906
rect 29381 3860 29451 3906
rect 29497 3860 29567 3906
rect 29613 3860 29683 3906
rect 29729 3860 29799 3906
rect 29845 3860 29915 3906
rect 29961 3860 30031 3906
rect 30077 3860 30147 3906
rect 30193 3860 30263 3906
rect 30309 3860 30379 3906
rect 30425 3860 30495 3906
rect 30541 3860 30611 3906
rect 30657 3860 30727 3906
rect 30773 3860 30843 3906
rect 30889 3860 30959 3906
rect 31005 3860 31075 3906
rect 31121 3860 31191 3906
rect 31237 3860 31307 3906
rect 31353 3860 31423 3906
rect 31469 3860 31539 3906
rect 31585 3860 31655 3906
rect 31701 3860 31771 3906
rect 31817 3860 31887 3906
rect 31933 3860 32003 3906
rect 32049 3860 32119 3906
rect 32165 3860 32235 3906
rect 32281 3860 32351 3906
rect 32397 3860 32467 3906
rect 32513 3860 32583 3906
rect 32629 3860 32699 3906
rect 32745 3860 32815 3906
rect 32861 3860 32931 3906
rect 32977 3860 33047 3906
rect 33093 3860 33163 3906
rect 33209 3860 33279 3906
rect 33325 3860 33395 3906
rect 33441 3860 33511 3906
rect 33557 3860 33627 3906
rect 33673 3860 33743 3906
rect 33789 3860 33859 3906
rect 33905 3860 33975 3906
rect 34021 3860 34091 3906
rect 34137 3860 34207 3906
rect 34253 3860 34323 3906
rect 34369 3860 34439 3906
rect 34485 3860 34555 3906
rect 34601 3860 34671 3906
rect 34717 3860 34787 3906
rect 34833 3860 34903 3906
rect 34949 3860 35019 3906
rect 35065 3860 35135 3906
rect 35181 3860 35251 3906
rect 35297 3860 35367 3906
rect 35413 3860 35483 3906
rect 35529 3860 35599 3906
rect 35645 3860 35715 3906
rect 35761 3860 35831 3906
rect 35877 3860 35947 3906
rect 35993 3860 36063 3906
rect 36109 3860 36179 3906
rect 36225 3860 36295 3906
rect 36341 3860 36411 3906
rect 36457 3860 36527 3906
rect 36573 3860 36643 3906
rect 36689 3860 36759 3906
rect 36805 3860 36875 3906
rect 36921 3860 36991 3906
rect 37037 3860 37107 3906
rect 37153 3860 37223 3906
rect 37269 3860 37339 3906
rect 37385 3860 37455 3906
rect 37501 3860 37571 3906
rect 37617 3860 37687 3906
rect 37733 3860 37803 3906
rect 37849 3860 37919 3906
rect 37965 3860 38035 3906
rect 38081 3860 38151 3906
rect 38197 3860 38267 3906
rect 38313 3860 38383 3906
rect 38429 3860 38499 3906
rect 38545 3860 38615 3906
rect 38661 3860 38731 3906
rect 38777 3860 38847 3906
rect 38893 3860 38963 3906
rect 39009 3860 39079 3906
rect 39125 3860 39195 3906
rect 39241 3860 39311 3906
rect 39357 3860 39427 3906
rect 39473 3860 39543 3906
rect 39589 3860 39659 3906
rect 39705 3860 39775 3906
rect 39821 3860 39891 3906
rect 39937 3860 40007 3906
rect 40053 3860 40123 3906
rect 40169 3860 40188 3906
rect 28620 3790 40188 3860
rect 28620 3744 28639 3790
rect 28685 3744 28755 3790
rect 28801 3744 28871 3790
rect 28917 3744 28987 3790
rect 29033 3744 29103 3790
rect 29149 3744 29219 3790
rect 29265 3744 29335 3790
rect 29381 3744 29451 3790
rect 29497 3744 29567 3790
rect 29613 3744 29683 3790
rect 29729 3744 29799 3790
rect 29845 3744 29915 3790
rect 29961 3744 30031 3790
rect 30077 3744 30147 3790
rect 30193 3744 30263 3790
rect 30309 3744 30379 3790
rect 30425 3744 30495 3790
rect 30541 3744 30611 3790
rect 30657 3744 30727 3790
rect 30773 3744 30843 3790
rect 30889 3744 30959 3790
rect 31005 3744 31075 3790
rect 31121 3744 31191 3790
rect 31237 3744 31307 3790
rect 31353 3744 31423 3790
rect 31469 3744 31539 3790
rect 31585 3744 31655 3790
rect 31701 3744 31771 3790
rect 31817 3744 31887 3790
rect 31933 3744 32003 3790
rect 32049 3744 32119 3790
rect 32165 3744 32235 3790
rect 32281 3744 32351 3790
rect 32397 3744 32467 3790
rect 32513 3744 32583 3790
rect 32629 3744 32699 3790
rect 32745 3744 32815 3790
rect 32861 3744 32931 3790
rect 32977 3744 33047 3790
rect 33093 3744 33163 3790
rect 33209 3744 33279 3790
rect 33325 3744 33395 3790
rect 33441 3744 33511 3790
rect 33557 3744 33627 3790
rect 33673 3744 33743 3790
rect 33789 3744 33859 3790
rect 33905 3744 33975 3790
rect 34021 3744 34091 3790
rect 34137 3744 34207 3790
rect 34253 3744 34323 3790
rect 34369 3744 34439 3790
rect 34485 3744 34555 3790
rect 34601 3744 34671 3790
rect 34717 3744 34787 3790
rect 34833 3744 34903 3790
rect 34949 3744 35019 3790
rect 35065 3744 35135 3790
rect 35181 3744 35251 3790
rect 35297 3744 35367 3790
rect 35413 3744 35483 3790
rect 35529 3744 35599 3790
rect 35645 3744 35715 3790
rect 35761 3744 35831 3790
rect 35877 3744 35947 3790
rect 35993 3744 36063 3790
rect 36109 3744 36179 3790
rect 36225 3744 36295 3790
rect 36341 3744 36411 3790
rect 36457 3744 36527 3790
rect 36573 3744 36643 3790
rect 36689 3744 36759 3790
rect 36805 3744 36875 3790
rect 36921 3744 36991 3790
rect 37037 3744 37107 3790
rect 37153 3744 37223 3790
rect 37269 3744 37339 3790
rect 37385 3744 37455 3790
rect 37501 3744 37571 3790
rect 37617 3744 37687 3790
rect 37733 3744 37803 3790
rect 37849 3744 37919 3790
rect 37965 3744 38035 3790
rect 38081 3744 38151 3790
rect 38197 3744 38267 3790
rect 38313 3744 38383 3790
rect 38429 3744 38499 3790
rect 38545 3744 38615 3790
rect 38661 3744 38731 3790
rect 38777 3744 38847 3790
rect 38893 3744 38963 3790
rect 39009 3744 39079 3790
rect 39125 3744 39195 3790
rect 39241 3744 39311 3790
rect 39357 3744 39427 3790
rect 39473 3744 39543 3790
rect 39589 3744 39659 3790
rect 39705 3744 39775 3790
rect 39821 3744 39891 3790
rect 39937 3744 40007 3790
rect 40053 3744 40123 3790
rect 40169 3744 40188 3790
rect 28620 3674 40188 3744
rect 28620 3628 28639 3674
rect 28685 3628 28755 3674
rect 28801 3628 28871 3674
rect 28917 3628 28987 3674
rect 29033 3628 29103 3674
rect 29149 3628 29219 3674
rect 29265 3628 29335 3674
rect 29381 3628 29451 3674
rect 29497 3628 29567 3674
rect 29613 3628 29683 3674
rect 29729 3628 29799 3674
rect 29845 3628 29915 3674
rect 29961 3628 30031 3674
rect 30077 3628 30147 3674
rect 30193 3628 30263 3674
rect 30309 3628 30379 3674
rect 30425 3628 30495 3674
rect 30541 3628 30611 3674
rect 30657 3628 30727 3674
rect 30773 3628 30843 3674
rect 30889 3628 30959 3674
rect 31005 3628 31075 3674
rect 31121 3628 31191 3674
rect 31237 3628 31307 3674
rect 31353 3628 31423 3674
rect 31469 3628 31539 3674
rect 31585 3628 31655 3674
rect 31701 3628 31771 3674
rect 31817 3628 31887 3674
rect 31933 3628 32003 3674
rect 32049 3628 32119 3674
rect 32165 3628 32235 3674
rect 32281 3628 32351 3674
rect 32397 3628 32467 3674
rect 32513 3628 32583 3674
rect 32629 3628 32699 3674
rect 32745 3628 32815 3674
rect 32861 3628 32931 3674
rect 32977 3628 33047 3674
rect 33093 3628 33163 3674
rect 33209 3628 33279 3674
rect 33325 3628 33395 3674
rect 33441 3628 33511 3674
rect 33557 3628 33627 3674
rect 33673 3628 33743 3674
rect 33789 3628 33859 3674
rect 33905 3628 33975 3674
rect 34021 3628 34091 3674
rect 34137 3628 34207 3674
rect 34253 3628 34323 3674
rect 34369 3628 34439 3674
rect 34485 3628 34555 3674
rect 34601 3628 34671 3674
rect 34717 3628 34787 3674
rect 34833 3628 34903 3674
rect 34949 3628 35019 3674
rect 35065 3628 35135 3674
rect 35181 3628 35251 3674
rect 35297 3628 35367 3674
rect 35413 3628 35483 3674
rect 35529 3628 35599 3674
rect 35645 3628 35715 3674
rect 35761 3628 35831 3674
rect 35877 3628 35947 3674
rect 35993 3628 36063 3674
rect 36109 3628 36179 3674
rect 36225 3628 36295 3674
rect 36341 3628 36411 3674
rect 36457 3628 36527 3674
rect 36573 3628 36643 3674
rect 36689 3628 36759 3674
rect 36805 3628 36875 3674
rect 36921 3628 36991 3674
rect 37037 3628 37107 3674
rect 37153 3628 37223 3674
rect 37269 3628 37339 3674
rect 37385 3628 37455 3674
rect 37501 3628 37571 3674
rect 37617 3628 37687 3674
rect 37733 3628 37803 3674
rect 37849 3628 37919 3674
rect 37965 3628 38035 3674
rect 38081 3628 38151 3674
rect 38197 3628 38267 3674
rect 38313 3628 38383 3674
rect 38429 3628 38499 3674
rect 38545 3628 38615 3674
rect 38661 3628 38731 3674
rect 38777 3628 38847 3674
rect 38893 3628 38963 3674
rect 39009 3628 39079 3674
rect 39125 3628 39195 3674
rect 39241 3628 39311 3674
rect 39357 3628 39427 3674
rect 39473 3628 39543 3674
rect 39589 3628 39659 3674
rect 39705 3628 39775 3674
rect 39821 3628 39891 3674
rect 39937 3628 40007 3674
rect 40053 3628 40123 3674
rect 40169 3628 40188 3674
rect 28620 3558 40188 3628
rect 28620 3512 28639 3558
rect 28685 3512 28755 3558
rect 28801 3512 28871 3558
rect 28917 3512 28987 3558
rect 29033 3512 29103 3558
rect 29149 3512 29219 3558
rect 29265 3512 29335 3558
rect 29381 3512 29451 3558
rect 29497 3512 29567 3558
rect 29613 3512 29683 3558
rect 29729 3512 29799 3558
rect 29845 3512 29915 3558
rect 29961 3512 30031 3558
rect 30077 3512 30147 3558
rect 30193 3512 30263 3558
rect 30309 3512 30379 3558
rect 30425 3512 30495 3558
rect 30541 3512 30611 3558
rect 30657 3512 30727 3558
rect 30773 3512 30843 3558
rect 30889 3512 30959 3558
rect 31005 3512 31075 3558
rect 31121 3512 31191 3558
rect 31237 3512 31307 3558
rect 31353 3512 31423 3558
rect 31469 3512 31539 3558
rect 31585 3512 31655 3558
rect 31701 3512 31771 3558
rect 31817 3512 31887 3558
rect 31933 3512 32003 3558
rect 32049 3512 32119 3558
rect 32165 3512 32235 3558
rect 32281 3512 32351 3558
rect 32397 3512 32467 3558
rect 32513 3512 32583 3558
rect 32629 3512 32699 3558
rect 32745 3512 32815 3558
rect 32861 3512 32931 3558
rect 32977 3512 33047 3558
rect 33093 3512 33163 3558
rect 33209 3512 33279 3558
rect 33325 3512 33395 3558
rect 33441 3512 33511 3558
rect 33557 3512 33627 3558
rect 33673 3512 33743 3558
rect 33789 3512 33859 3558
rect 33905 3512 33975 3558
rect 34021 3512 34091 3558
rect 34137 3512 34207 3558
rect 34253 3512 34323 3558
rect 34369 3512 34439 3558
rect 34485 3512 34555 3558
rect 34601 3512 34671 3558
rect 34717 3512 34787 3558
rect 34833 3512 34903 3558
rect 34949 3512 35019 3558
rect 35065 3512 35135 3558
rect 35181 3512 35251 3558
rect 35297 3512 35367 3558
rect 35413 3512 35483 3558
rect 35529 3512 35599 3558
rect 35645 3512 35715 3558
rect 35761 3512 35831 3558
rect 35877 3512 35947 3558
rect 35993 3512 36063 3558
rect 36109 3512 36179 3558
rect 36225 3512 36295 3558
rect 36341 3512 36411 3558
rect 36457 3512 36527 3558
rect 36573 3512 36643 3558
rect 36689 3512 36759 3558
rect 36805 3512 36875 3558
rect 36921 3512 36991 3558
rect 37037 3512 37107 3558
rect 37153 3512 37223 3558
rect 37269 3512 37339 3558
rect 37385 3512 37455 3558
rect 37501 3512 37571 3558
rect 37617 3512 37687 3558
rect 37733 3512 37803 3558
rect 37849 3512 37919 3558
rect 37965 3512 38035 3558
rect 38081 3512 38151 3558
rect 38197 3512 38267 3558
rect 38313 3512 38383 3558
rect 38429 3512 38499 3558
rect 38545 3512 38615 3558
rect 38661 3512 38731 3558
rect 38777 3512 38847 3558
rect 38893 3512 38963 3558
rect 39009 3512 39079 3558
rect 39125 3512 39195 3558
rect 39241 3512 39311 3558
rect 39357 3512 39427 3558
rect 39473 3512 39543 3558
rect 39589 3512 39659 3558
rect 39705 3512 39775 3558
rect 39821 3512 39891 3558
rect 39937 3512 40007 3558
rect 40053 3512 40123 3558
rect 40169 3512 40188 3558
rect 28620 3442 40188 3512
rect 28620 3396 28639 3442
rect 28685 3396 28755 3442
rect 28801 3396 28871 3442
rect 28917 3396 28987 3442
rect 29033 3396 29103 3442
rect 29149 3396 29219 3442
rect 29265 3396 29335 3442
rect 29381 3396 29451 3442
rect 29497 3396 29567 3442
rect 29613 3396 29683 3442
rect 29729 3396 29799 3442
rect 29845 3396 29915 3442
rect 29961 3396 30031 3442
rect 30077 3396 30147 3442
rect 30193 3396 30263 3442
rect 30309 3396 30379 3442
rect 30425 3396 30495 3442
rect 30541 3396 30611 3442
rect 30657 3396 30727 3442
rect 30773 3396 30843 3442
rect 30889 3396 30959 3442
rect 31005 3396 31075 3442
rect 31121 3396 31191 3442
rect 31237 3396 31307 3442
rect 31353 3396 31423 3442
rect 31469 3396 31539 3442
rect 31585 3396 31655 3442
rect 31701 3396 31771 3442
rect 31817 3396 31887 3442
rect 31933 3396 32003 3442
rect 32049 3396 32119 3442
rect 32165 3396 32235 3442
rect 32281 3396 32351 3442
rect 32397 3396 32467 3442
rect 32513 3396 32583 3442
rect 32629 3396 32699 3442
rect 32745 3396 32815 3442
rect 32861 3396 32931 3442
rect 32977 3396 33047 3442
rect 33093 3396 33163 3442
rect 33209 3396 33279 3442
rect 33325 3396 33395 3442
rect 33441 3396 33511 3442
rect 33557 3396 33627 3442
rect 33673 3396 33743 3442
rect 33789 3396 33859 3442
rect 33905 3396 33975 3442
rect 34021 3396 34091 3442
rect 34137 3396 34207 3442
rect 34253 3396 34323 3442
rect 34369 3396 34439 3442
rect 34485 3396 34555 3442
rect 34601 3396 34671 3442
rect 34717 3396 34787 3442
rect 34833 3396 34903 3442
rect 34949 3396 35019 3442
rect 35065 3396 35135 3442
rect 35181 3396 35251 3442
rect 35297 3396 35367 3442
rect 35413 3396 35483 3442
rect 35529 3396 35599 3442
rect 35645 3396 35715 3442
rect 35761 3396 35831 3442
rect 35877 3396 35947 3442
rect 35993 3396 36063 3442
rect 36109 3396 36179 3442
rect 36225 3396 36295 3442
rect 36341 3396 36411 3442
rect 36457 3396 36527 3442
rect 36573 3396 36643 3442
rect 36689 3396 36759 3442
rect 36805 3396 36875 3442
rect 36921 3396 36991 3442
rect 37037 3396 37107 3442
rect 37153 3396 37223 3442
rect 37269 3396 37339 3442
rect 37385 3396 37455 3442
rect 37501 3396 37571 3442
rect 37617 3396 37687 3442
rect 37733 3396 37803 3442
rect 37849 3396 37919 3442
rect 37965 3396 38035 3442
rect 38081 3396 38151 3442
rect 38197 3396 38267 3442
rect 38313 3396 38383 3442
rect 38429 3396 38499 3442
rect 38545 3396 38615 3442
rect 38661 3396 38731 3442
rect 38777 3396 38847 3442
rect 38893 3396 38963 3442
rect 39009 3396 39079 3442
rect 39125 3396 39195 3442
rect 39241 3396 39311 3442
rect 39357 3396 39427 3442
rect 39473 3396 39543 3442
rect 39589 3396 39659 3442
rect 39705 3396 39775 3442
rect 39821 3396 39891 3442
rect 39937 3396 40007 3442
rect 40053 3396 40123 3442
rect 40169 3396 40188 3442
rect 28620 3326 40188 3396
rect 28620 3280 28639 3326
rect 28685 3280 28755 3326
rect 28801 3280 28871 3326
rect 28917 3280 28987 3326
rect 29033 3280 29103 3326
rect 29149 3280 29219 3326
rect 29265 3280 29335 3326
rect 29381 3280 29451 3326
rect 29497 3280 29567 3326
rect 29613 3280 29683 3326
rect 29729 3280 29799 3326
rect 29845 3280 29915 3326
rect 29961 3280 30031 3326
rect 30077 3280 30147 3326
rect 30193 3280 30263 3326
rect 30309 3280 30379 3326
rect 30425 3280 30495 3326
rect 30541 3280 30611 3326
rect 30657 3280 30727 3326
rect 30773 3280 30843 3326
rect 30889 3280 30959 3326
rect 31005 3280 31075 3326
rect 31121 3280 31191 3326
rect 31237 3280 31307 3326
rect 31353 3280 31423 3326
rect 31469 3280 31539 3326
rect 31585 3280 31655 3326
rect 31701 3280 31771 3326
rect 31817 3280 31887 3326
rect 31933 3280 32003 3326
rect 32049 3280 32119 3326
rect 32165 3280 32235 3326
rect 32281 3280 32351 3326
rect 32397 3280 32467 3326
rect 32513 3280 32583 3326
rect 32629 3280 32699 3326
rect 32745 3280 32815 3326
rect 32861 3280 32931 3326
rect 32977 3280 33047 3326
rect 33093 3280 33163 3326
rect 33209 3280 33279 3326
rect 33325 3280 33395 3326
rect 33441 3280 33511 3326
rect 33557 3280 33627 3326
rect 33673 3280 33743 3326
rect 33789 3280 33859 3326
rect 33905 3280 33975 3326
rect 34021 3280 34091 3326
rect 34137 3280 34207 3326
rect 34253 3280 34323 3326
rect 34369 3280 34439 3326
rect 34485 3280 34555 3326
rect 34601 3280 34671 3326
rect 34717 3280 34787 3326
rect 34833 3280 34903 3326
rect 34949 3280 35019 3326
rect 35065 3280 35135 3326
rect 35181 3280 35251 3326
rect 35297 3280 35367 3326
rect 35413 3280 35483 3326
rect 35529 3280 35599 3326
rect 35645 3280 35715 3326
rect 35761 3280 35831 3326
rect 35877 3280 35947 3326
rect 35993 3280 36063 3326
rect 36109 3280 36179 3326
rect 36225 3280 36295 3326
rect 36341 3280 36411 3326
rect 36457 3280 36527 3326
rect 36573 3280 36643 3326
rect 36689 3280 36759 3326
rect 36805 3280 36875 3326
rect 36921 3280 36991 3326
rect 37037 3280 37107 3326
rect 37153 3280 37223 3326
rect 37269 3280 37339 3326
rect 37385 3280 37455 3326
rect 37501 3280 37571 3326
rect 37617 3280 37687 3326
rect 37733 3280 37803 3326
rect 37849 3280 37919 3326
rect 37965 3280 38035 3326
rect 38081 3280 38151 3326
rect 38197 3280 38267 3326
rect 38313 3280 38383 3326
rect 38429 3280 38499 3326
rect 38545 3280 38615 3326
rect 38661 3280 38731 3326
rect 38777 3280 38847 3326
rect 38893 3280 38963 3326
rect 39009 3280 39079 3326
rect 39125 3280 39195 3326
rect 39241 3280 39311 3326
rect 39357 3280 39427 3326
rect 39473 3280 39543 3326
rect 39589 3280 39659 3326
rect 39705 3280 39775 3326
rect 39821 3280 39891 3326
rect 39937 3280 40007 3326
rect 40053 3280 40123 3326
rect 40169 3280 40188 3326
rect 28620 3210 40188 3280
rect 28620 3164 28639 3210
rect 28685 3164 28755 3210
rect 28801 3164 28871 3210
rect 28917 3164 28987 3210
rect 29033 3164 29103 3210
rect 29149 3164 29219 3210
rect 29265 3164 29335 3210
rect 29381 3164 29451 3210
rect 29497 3164 29567 3210
rect 29613 3164 29683 3210
rect 29729 3164 29799 3210
rect 29845 3164 29915 3210
rect 29961 3164 30031 3210
rect 30077 3164 30147 3210
rect 30193 3164 30263 3210
rect 30309 3164 30379 3210
rect 30425 3164 30495 3210
rect 30541 3164 30611 3210
rect 30657 3164 30727 3210
rect 30773 3164 30843 3210
rect 30889 3164 30959 3210
rect 31005 3164 31075 3210
rect 31121 3164 31191 3210
rect 31237 3164 31307 3210
rect 31353 3164 31423 3210
rect 31469 3164 31539 3210
rect 31585 3164 31655 3210
rect 31701 3164 31771 3210
rect 31817 3164 31887 3210
rect 31933 3164 32003 3210
rect 32049 3164 32119 3210
rect 32165 3164 32235 3210
rect 32281 3164 32351 3210
rect 32397 3164 32467 3210
rect 32513 3164 32583 3210
rect 32629 3164 32699 3210
rect 32745 3164 32815 3210
rect 32861 3164 32931 3210
rect 32977 3164 33047 3210
rect 33093 3164 33163 3210
rect 33209 3164 33279 3210
rect 33325 3164 33395 3210
rect 33441 3164 33511 3210
rect 33557 3164 33627 3210
rect 33673 3164 33743 3210
rect 33789 3164 33859 3210
rect 33905 3164 33975 3210
rect 34021 3164 34091 3210
rect 34137 3164 34207 3210
rect 34253 3164 34323 3210
rect 34369 3164 34439 3210
rect 34485 3164 34555 3210
rect 34601 3164 34671 3210
rect 34717 3164 34787 3210
rect 34833 3164 34903 3210
rect 34949 3164 35019 3210
rect 35065 3164 35135 3210
rect 35181 3164 35251 3210
rect 35297 3164 35367 3210
rect 35413 3164 35483 3210
rect 35529 3164 35599 3210
rect 35645 3164 35715 3210
rect 35761 3164 35831 3210
rect 35877 3164 35947 3210
rect 35993 3164 36063 3210
rect 36109 3164 36179 3210
rect 36225 3164 36295 3210
rect 36341 3164 36411 3210
rect 36457 3164 36527 3210
rect 36573 3164 36643 3210
rect 36689 3164 36759 3210
rect 36805 3164 36875 3210
rect 36921 3164 36991 3210
rect 37037 3164 37107 3210
rect 37153 3164 37223 3210
rect 37269 3164 37339 3210
rect 37385 3164 37455 3210
rect 37501 3164 37571 3210
rect 37617 3164 37687 3210
rect 37733 3164 37803 3210
rect 37849 3164 37919 3210
rect 37965 3164 38035 3210
rect 38081 3164 38151 3210
rect 38197 3164 38267 3210
rect 38313 3164 38383 3210
rect 38429 3164 38499 3210
rect 38545 3164 38615 3210
rect 38661 3164 38731 3210
rect 38777 3164 38847 3210
rect 38893 3164 38963 3210
rect 39009 3164 39079 3210
rect 39125 3164 39195 3210
rect 39241 3164 39311 3210
rect 39357 3164 39427 3210
rect 39473 3164 39543 3210
rect 39589 3164 39659 3210
rect 39705 3164 39775 3210
rect 39821 3164 39891 3210
rect 39937 3164 40007 3210
rect 40053 3164 40123 3210
rect 40169 3164 40188 3210
rect 28620 3094 40188 3164
rect 28620 3048 28639 3094
rect 28685 3048 28755 3094
rect 28801 3048 28871 3094
rect 28917 3048 28987 3094
rect 29033 3048 29103 3094
rect 29149 3048 29219 3094
rect 29265 3048 29335 3094
rect 29381 3048 29451 3094
rect 29497 3048 29567 3094
rect 29613 3048 29683 3094
rect 29729 3048 29799 3094
rect 29845 3048 29915 3094
rect 29961 3048 30031 3094
rect 30077 3048 30147 3094
rect 30193 3048 30263 3094
rect 30309 3048 30379 3094
rect 30425 3048 30495 3094
rect 30541 3048 30611 3094
rect 30657 3048 30727 3094
rect 30773 3048 30843 3094
rect 30889 3048 30959 3094
rect 31005 3048 31075 3094
rect 31121 3048 31191 3094
rect 31237 3048 31307 3094
rect 31353 3048 31423 3094
rect 31469 3048 31539 3094
rect 31585 3048 31655 3094
rect 31701 3048 31771 3094
rect 31817 3048 31887 3094
rect 31933 3048 32003 3094
rect 32049 3048 32119 3094
rect 32165 3048 32235 3094
rect 32281 3048 32351 3094
rect 32397 3048 32467 3094
rect 32513 3048 32583 3094
rect 32629 3048 32699 3094
rect 32745 3048 32815 3094
rect 32861 3048 32931 3094
rect 32977 3048 33047 3094
rect 33093 3048 33163 3094
rect 33209 3048 33279 3094
rect 33325 3048 33395 3094
rect 33441 3048 33511 3094
rect 33557 3048 33627 3094
rect 33673 3048 33743 3094
rect 33789 3048 33859 3094
rect 33905 3048 33975 3094
rect 34021 3048 34091 3094
rect 34137 3048 34207 3094
rect 34253 3048 34323 3094
rect 34369 3048 34439 3094
rect 34485 3048 34555 3094
rect 34601 3048 34671 3094
rect 34717 3048 34787 3094
rect 34833 3048 34903 3094
rect 34949 3048 35019 3094
rect 35065 3048 35135 3094
rect 35181 3048 35251 3094
rect 35297 3048 35367 3094
rect 35413 3048 35483 3094
rect 35529 3048 35599 3094
rect 35645 3048 35715 3094
rect 35761 3048 35831 3094
rect 35877 3048 35947 3094
rect 35993 3048 36063 3094
rect 36109 3048 36179 3094
rect 36225 3048 36295 3094
rect 36341 3048 36411 3094
rect 36457 3048 36527 3094
rect 36573 3048 36643 3094
rect 36689 3048 36759 3094
rect 36805 3048 36875 3094
rect 36921 3048 36991 3094
rect 37037 3048 37107 3094
rect 37153 3048 37223 3094
rect 37269 3048 37339 3094
rect 37385 3048 37455 3094
rect 37501 3048 37571 3094
rect 37617 3048 37687 3094
rect 37733 3048 37803 3094
rect 37849 3048 37919 3094
rect 37965 3048 38035 3094
rect 38081 3048 38151 3094
rect 38197 3048 38267 3094
rect 38313 3048 38383 3094
rect 38429 3048 38499 3094
rect 38545 3048 38615 3094
rect 38661 3048 38731 3094
rect 38777 3048 38847 3094
rect 38893 3048 38963 3094
rect 39009 3048 39079 3094
rect 39125 3048 39195 3094
rect 39241 3048 39311 3094
rect 39357 3048 39427 3094
rect 39473 3048 39543 3094
rect 39589 3048 39659 3094
rect 39705 3048 39775 3094
rect 39821 3048 39891 3094
rect 39937 3048 40007 3094
rect 40053 3048 40123 3094
rect 40169 3048 40188 3094
rect 28620 2978 40188 3048
rect 28620 2932 28639 2978
rect 28685 2932 28755 2978
rect 28801 2932 28871 2978
rect 28917 2932 28987 2978
rect 29033 2932 29103 2978
rect 29149 2932 29219 2978
rect 29265 2932 29335 2978
rect 29381 2932 29451 2978
rect 29497 2932 29567 2978
rect 29613 2932 29683 2978
rect 29729 2932 29799 2978
rect 29845 2932 29915 2978
rect 29961 2932 30031 2978
rect 30077 2932 30147 2978
rect 30193 2932 30263 2978
rect 30309 2932 30379 2978
rect 30425 2932 30495 2978
rect 30541 2932 30611 2978
rect 30657 2932 30727 2978
rect 30773 2932 30843 2978
rect 30889 2932 30959 2978
rect 31005 2932 31075 2978
rect 31121 2932 31191 2978
rect 31237 2932 31307 2978
rect 31353 2932 31423 2978
rect 31469 2932 31539 2978
rect 31585 2932 31655 2978
rect 31701 2932 31771 2978
rect 31817 2932 31887 2978
rect 31933 2932 32003 2978
rect 32049 2932 32119 2978
rect 32165 2932 32235 2978
rect 32281 2932 32351 2978
rect 32397 2932 32467 2978
rect 32513 2932 32583 2978
rect 32629 2932 32699 2978
rect 32745 2932 32815 2978
rect 32861 2932 32931 2978
rect 32977 2932 33047 2978
rect 33093 2932 33163 2978
rect 33209 2932 33279 2978
rect 33325 2932 33395 2978
rect 33441 2932 33511 2978
rect 33557 2932 33627 2978
rect 33673 2932 33743 2978
rect 33789 2932 33859 2978
rect 33905 2932 33975 2978
rect 34021 2932 34091 2978
rect 34137 2932 34207 2978
rect 34253 2932 34323 2978
rect 34369 2932 34439 2978
rect 34485 2932 34555 2978
rect 34601 2932 34671 2978
rect 34717 2932 34787 2978
rect 34833 2932 34903 2978
rect 34949 2932 35019 2978
rect 35065 2932 35135 2978
rect 35181 2932 35251 2978
rect 35297 2932 35367 2978
rect 35413 2932 35483 2978
rect 35529 2932 35599 2978
rect 35645 2932 35715 2978
rect 35761 2932 35831 2978
rect 35877 2932 35947 2978
rect 35993 2932 36063 2978
rect 36109 2932 36179 2978
rect 36225 2932 36295 2978
rect 36341 2932 36411 2978
rect 36457 2932 36527 2978
rect 36573 2932 36643 2978
rect 36689 2932 36759 2978
rect 36805 2932 36875 2978
rect 36921 2932 36991 2978
rect 37037 2932 37107 2978
rect 37153 2932 37223 2978
rect 37269 2932 37339 2978
rect 37385 2932 37455 2978
rect 37501 2932 37571 2978
rect 37617 2932 37687 2978
rect 37733 2932 37803 2978
rect 37849 2932 37919 2978
rect 37965 2932 38035 2978
rect 38081 2932 38151 2978
rect 38197 2932 38267 2978
rect 38313 2932 38383 2978
rect 38429 2932 38499 2978
rect 38545 2932 38615 2978
rect 38661 2932 38731 2978
rect 38777 2932 38847 2978
rect 38893 2932 38963 2978
rect 39009 2932 39079 2978
rect 39125 2932 39195 2978
rect 39241 2932 39311 2978
rect 39357 2932 39427 2978
rect 39473 2932 39543 2978
rect 39589 2932 39659 2978
rect 39705 2932 39775 2978
rect 39821 2932 39891 2978
rect 39937 2932 40007 2978
rect 40053 2932 40123 2978
rect 40169 2932 40188 2978
rect 28620 2862 40188 2932
rect 28620 2816 28639 2862
rect 28685 2816 28755 2862
rect 28801 2816 28871 2862
rect 28917 2816 28987 2862
rect 29033 2816 29103 2862
rect 29149 2816 29219 2862
rect 29265 2816 29335 2862
rect 29381 2816 29451 2862
rect 29497 2816 29567 2862
rect 29613 2816 29683 2862
rect 29729 2816 29799 2862
rect 29845 2816 29915 2862
rect 29961 2816 30031 2862
rect 30077 2816 30147 2862
rect 30193 2816 30263 2862
rect 30309 2816 30379 2862
rect 30425 2816 30495 2862
rect 30541 2816 30611 2862
rect 30657 2816 30727 2862
rect 30773 2816 30843 2862
rect 30889 2816 30959 2862
rect 31005 2816 31075 2862
rect 31121 2816 31191 2862
rect 31237 2816 31307 2862
rect 31353 2816 31423 2862
rect 31469 2816 31539 2862
rect 31585 2816 31655 2862
rect 31701 2816 31771 2862
rect 31817 2816 31887 2862
rect 31933 2816 32003 2862
rect 32049 2816 32119 2862
rect 32165 2816 32235 2862
rect 32281 2816 32351 2862
rect 32397 2816 32467 2862
rect 32513 2816 32583 2862
rect 32629 2816 32699 2862
rect 32745 2816 32815 2862
rect 32861 2816 32931 2862
rect 32977 2816 33047 2862
rect 33093 2816 33163 2862
rect 33209 2816 33279 2862
rect 33325 2816 33395 2862
rect 33441 2816 33511 2862
rect 33557 2816 33627 2862
rect 33673 2816 33743 2862
rect 33789 2816 33859 2862
rect 33905 2816 33975 2862
rect 34021 2816 34091 2862
rect 34137 2816 34207 2862
rect 34253 2816 34323 2862
rect 34369 2816 34439 2862
rect 34485 2816 34555 2862
rect 34601 2816 34671 2862
rect 34717 2816 34787 2862
rect 34833 2816 34903 2862
rect 34949 2816 35019 2862
rect 35065 2816 35135 2862
rect 35181 2816 35251 2862
rect 35297 2816 35367 2862
rect 35413 2816 35483 2862
rect 35529 2816 35599 2862
rect 35645 2816 35715 2862
rect 35761 2816 35831 2862
rect 35877 2816 35947 2862
rect 35993 2816 36063 2862
rect 36109 2816 36179 2862
rect 36225 2816 36295 2862
rect 36341 2816 36411 2862
rect 36457 2816 36527 2862
rect 36573 2816 36643 2862
rect 36689 2816 36759 2862
rect 36805 2816 36875 2862
rect 36921 2816 36991 2862
rect 37037 2816 37107 2862
rect 37153 2816 37223 2862
rect 37269 2816 37339 2862
rect 37385 2816 37455 2862
rect 37501 2816 37571 2862
rect 37617 2816 37687 2862
rect 37733 2816 37803 2862
rect 37849 2816 37919 2862
rect 37965 2816 38035 2862
rect 38081 2816 38151 2862
rect 38197 2816 38267 2862
rect 38313 2816 38383 2862
rect 38429 2816 38499 2862
rect 38545 2816 38615 2862
rect 38661 2816 38731 2862
rect 38777 2816 38847 2862
rect 38893 2816 38963 2862
rect 39009 2816 39079 2862
rect 39125 2816 39195 2862
rect 39241 2816 39311 2862
rect 39357 2816 39427 2862
rect 39473 2816 39543 2862
rect 39589 2816 39659 2862
rect 39705 2816 39775 2862
rect 39821 2816 39891 2862
rect 39937 2816 40007 2862
rect 40053 2816 40123 2862
rect 40169 2816 40188 2862
rect 28620 2746 40188 2816
rect 28620 2700 28639 2746
rect 28685 2700 28755 2746
rect 28801 2700 28871 2746
rect 28917 2700 28987 2746
rect 29033 2700 29103 2746
rect 29149 2700 29219 2746
rect 29265 2700 29335 2746
rect 29381 2700 29451 2746
rect 29497 2700 29567 2746
rect 29613 2700 29683 2746
rect 29729 2700 29799 2746
rect 29845 2700 29915 2746
rect 29961 2700 30031 2746
rect 30077 2700 30147 2746
rect 30193 2700 30263 2746
rect 30309 2700 30379 2746
rect 30425 2700 30495 2746
rect 30541 2700 30611 2746
rect 30657 2700 30727 2746
rect 30773 2700 30843 2746
rect 30889 2700 30959 2746
rect 31005 2700 31075 2746
rect 31121 2700 31191 2746
rect 31237 2700 31307 2746
rect 31353 2700 31423 2746
rect 31469 2700 31539 2746
rect 31585 2700 31655 2746
rect 31701 2700 31771 2746
rect 31817 2700 31887 2746
rect 31933 2700 32003 2746
rect 32049 2700 32119 2746
rect 32165 2700 32235 2746
rect 32281 2700 32351 2746
rect 32397 2700 32467 2746
rect 32513 2700 32583 2746
rect 32629 2700 32699 2746
rect 32745 2700 32815 2746
rect 32861 2700 32931 2746
rect 32977 2700 33047 2746
rect 33093 2700 33163 2746
rect 33209 2700 33279 2746
rect 33325 2700 33395 2746
rect 33441 2700 33511 2746
rect 33557 2700 33627 2746
rect 33673 2700 33743 2746
rect 33789 2700 33859 2746
rect 33905 2700 33975 2746
rect 34021 2700 34091 2746
rect 34137 2700 34207 2746
rect 34253 2700 34323 2746
rect 34369 2700 34439 2746
rect 34485 2700 34555 2746
rect 34601 2700 34671 2746
rect 34717 2700 34787 2746
rect 34833 2700 34903 2746
rect 34949 2700 35019 2746
rect 35065 2700 35135 2746
rect 35181 2700 35251 2746
rect 35297 2700 35367 2746
rect 35413 2700 35483 2746
rect 35529 2700 35599 2746
rect 35645 2700 35715 2746
rect 35761 2700 35831 2746
rect 35877 2700 35947 2746
rect 35993 2700 36063 2746
rect 36109 2700 36179 2746
rect 36225 2700 36295 2746
rect 36341 2700 36411 2746
rect 36457 2700 36527 2746
rect 36573 2700 36643 2746
rect 36689 2700 36759 2746
rect 36805 2700 36875 2746
rect 36921 2700 36991 2746
rect 37037 2700 37107 2746
rect 37153 2700 37223 2746
rect 37269 2700 37339 2746
rect 37385 2700 37455 2746
rect 37501 2700 37571 2746
rect 37617 2700 37687 2746
rect 37733 2700 37803 2746
rect 37849 2700 37919 2746
rect 37965 2700 38035 2746
rect 38081 2700 38151 2746
rect 38197 2700 38267 2746
rect 38313 2700 38383 2746
rect 38429 2700 38499 2746
rect 38545 2700 38615 2746
rect 38661 2700 38731 2746
rect 38777 2700 38847 2746
rect 38893 2700 38963 2746
rect 39009 2700 39079 2746
rect 39125 2700 39195 2746
rect 39241 2700 39311 2746
rect 39357 2700 39427 2746
rect 39473 2700 39543 2746
rect 39589 2700 39659 2746
rect 39705 2700 39775 2746
rect 39821 2700 39891 2746
rect 39937 2700 40007 2746
rect 40053 2700 40123 2746
rect 40169 2700 40188 2746
rect 28620 2630 40188 2700
rect 28620 2584 28639 2630
rect 28685 2584 28755 2630
rect 28801 2584 28871 2630
rect 28917 2584 28987 2630
rect 29033 2584 29103 2630
rect 29149 2584 29219 2630
rect 29265 2584 29335 2630
rect 29381 2584 29451 2630
rect 29497 2584 29567 2630
rect 29613 2584 29683 2630
rect 29729 2584 29799 2630
rect 29845 2584 29915 2630
rect 29961 2584 30031 2630
rect 30077 2584 30147 2630
rect 30193 2584 30263 2630
rect 30309 2584 30379 2630
rect 30425 2584 30495 2630
rect 30541 2584 30611 2630
rect 30657 2584 30727 2630
rect 30773 2584 30843 2630
rect 30889 2584 30959 2630
rect 31005 2584 31075 2630
rect 31121 2584 31191 2630
rect 31237 2584 31307 2630
rect 31353 2584 31423 2630
rect 31469 2584 31539 2630
rect 31585 2584 31655 2630
rect 31701 2584 31771 2630
rect 31817 2584 31887 2630
rect 31933 2584 32003 2630
rect 32049 2584 32119 2630
rect 32165 2584 32235 2630
rect 32281 2584 32351 2630
rect 32397 2584 32467 2630
rect 32513 2584 32583 2630
rect 32629 2584 32699 2630
rect 32745 2584 32815 2630
rect 32861 2584 32931 2630
rect 32977 2584 33047 2630
rect 33093 2584 33163 2630
rect 33209 2584 33279 2630
rect 33325 2584 33395 2630
rect 33441 2584 33511 2630
rect 33557 2584 33627 2630
rect 33673 2584 33743 2630
rect 33789 2584 33859 2630
rect 33905 2584 33975 2630
rect 34021 2584 34091 2630
rect 34137 2584 34207 2630
rect 34253 2584 34323 2630
rect 34369 2584 34439 2630
rect 34485 2584 34555 2630
rect 34601 2584 34671 2630
rect 34717 2584 34787 2630
rect 34833 2584 34903 2630
rect 34949 2584 35019 2630
rect 35065 2584 35135 2630
rect 35181 2584 35251 2630
rect 35297 2584 35367 2630
rect 35413 2584 35483 2630
rect 35529 2584 35599 2630
rect 35645 2584 35715 2630
rect 35761 2584 35831 2630
rect 35877 2584 35947 2630
rect 35993 2584 36063 2630
rect 36109 2584 36179 2630
rect 36225 2584 36295 2630
rect 36341 2584 36411 2630
rect 36457 2584 36527 2630
rect 36573 2584 36643 2630
rect 36689 2584 36759 2630
rect 36805 2584 36875 2630
rect 36921 2584 36991 2630
rect 37037 2584 37107 2630
rect 37153 2584 37223 2630
rect 37269 2584 37339 2630
rect 37385 2584 37455 2630
rect 37501 2584 37571 2630
rect 37617 2584 37687 2630
rect 37733 2584 37803 2630
rect 37849 2584 37919 2630
rect 37965 2584 38035 2630
rect 38081 2584 38151 2630
rect 38197 2584 38267 2630
rect 38313 2584 38383 2630
rect 38429 2584 38499 2630
rect 38545 2584 38615 2630
rect 38661 2584 38731 2630
rect 38777 2584 38847 2630
rect 38893 2584 38963 2630
rect 39009 2584 39079 2630
rect 39125 2584 39195 2630
rect 39241 2584 39311 2630
rect 39357 2584 39427 2630
rect 39473 2584 39543 2630
rect 39589 2584 39659 2630
rect 39705 2584 39775 2630
rect 39821 2584 39891 2630
rect 39937 2584 40007 2630
rect 40053 2584 40123 2630
rect 40169 2584 40188 2630
rect 28620 2514 40188 2584
rect 28620 2468 28639 2514
rect 28685 2468 28755 2514
rect 28801 2468 28871 2514
rect 28917 2468 28987 2514
rect 29033 2468 29103 2514
rect 29149 2468 29219 2514
rect 29265 2468 29335 2514
rect 29381 2468 29451 2514
rect 29497 2468 29567 2514
rect 29613 2468 29683 2514
rect 29729 2468 29799 2514
rect 29845 2468 29915 2514
rect 29961 2468 30031 2514
rect 30077 2468 30147 2514
rect 30193 2468 30263 2514
rect 30309 2468 30379 2514
rect 30425 2468 30495 2514
rect 30541 2468 30611 2514
rect 30657 2468 30727 2514
rect 30773 2468 30843 2514
rect 30889 2468 30959 2514
rect 31005 2468 31075 2514
rect 31121 2468 31191 2514
rect 31237 2468 31307 2514
rect 31353 2468 31423 2514
rect 31469 2468 31539 2514
rect 31585 2468 31655 2514
rect 31701 2468 31771 2514
rect 31817 2468 31887 2514
rect 31933 2468 32003 2514
rect 32049 2468 32119 2514
rect 32165 2468 32235 2514
rect 32281 2468 32351 2514
rect 32397 2468 32467 2514
rect 32513 2468 32583 2514
rect 32629 2468 32699 2514
rect 32745 2468 32815 2514
rect 32861 2468 32931 2514
rect 32977 2468 33047 2514
rect 33093 2468 33163 2514
rect 33209 2468 33279 2514
rect 33325 2468 33395 2514
rect 33441 2468 33511 2514
rect 33557 2468 33627 2514
rect 33673 2468 33743 2514
rect 33789 2468 33859 2514
rect 33905 2468 33975 2514
rect 34021 2468 34091 2514
rect 34137 2468 34207 2514
rect 34253 2468 34323 2514
rect 34369 2468 34439 2514
rect 34485 2468 34555 2514
rect 34601 2468 34671 2514
rect 34717 2468 34787 2514
rect 34833 2468 34903 2514
rect 34949 2468 35019 2514
rect 35065 2468 35135 2514
rect 35181 2468 35251 2514
rect 35297 2468 35367 2514
rect 35413 2468 35483 2514
rect 35529 2468 35599 2514
rect 35645 2468 35715 2514
rect 35761 2468 35831 2514
rect 35877 2468 35947 2514
rect 35993 2468 36063 2514
rect 36109 2468 36179 2514
rect 36225 2468 36295 2514
rect 36341 2468 36411 2514
rect 36457 2468 36527 2514
rect 36573 2468 36643 2514
rect 36689 2468 36759 2514
rect 36805 2468 36875 2514
rect 36921 2468 36991 2514
rect 37037 2468 37107 2514
rect 37153 2468 37223 2514
rect 37269 2468 37339 2514
rect 37385 2468 37455 2514
rect 37501 2468 37571 2514
rect 37617 2468 37687 2514
rect 37733 2468 37803 2514
rect 37849 2468 37919 2514
rect 37965 2468 38035 2514
rect 38081 2468 38151 2514
rect 38197 2468 38267 2514
rect 38313 2468 38383 2514
rect 38429 2468 38499 2514
rect 38545 2468 38615 2514
rect 38661 2468 38731 2514
rect 38777 2468 38847 2514
rect 38893 2468 38963 2514
rect 39009 2468 39079 2514
rect 39125 2468 39195 2514
rect 39241 2468 39311 2514
rect 39357 2468 39427 2514
rect 39473 2468 39543 2514
rect 39589 2468 39659 2514
rect 39705 2468 39775 2514
rect 39821 2468 39891 2514
rect 39937 2468 40007 2514
rect 40053 2468 40123 2514
rect 40169 2468 40188 2514
rect 28620 2398 40188 2468
rect 28620 2352 28639 2398
rect 28685 2352 28755 2398
rect 28801 2352 28871 2398
rect 28917 2352 28987 2398
rect 29033 2352 29103 2398
rect 29149 2352 29219 2398
rect 29265 2352 29335 2398
rect 29381 2352 29451 2398
rect 29497 2352 29567 2398
rect 29613 2352 29683 2398
rect 29729 2352 29799 2398
rect 29845 2352 29915 2398
rect 29961 2352 30031 2398
rect 30077 2352 30147 2398
rect 30193 2352 30263 2398
rect 30309 2352 30379 2398
rect 30425 2352 30495 2398
rect 30541 2352 30611 2398
rect 30657 2352 30727 2398
rect 30773 2352 30843 2398
rect 30889 2352 30959 2398
rect 31005 2352 31075 2398
rect 31121 2352 31191 2398
rect 31237 2352 31307 2398
rect 31353 2352 31423 2398
rect 31469 2352 31539 2398
rect 31585 2352 31655 2398
rect 31701 2352 31771 2398
rect 31817 2352 31887 2398
rect 31933 2352 32003 2398
rect 32049 2352 32119 2398
rect 32165 2352 32235 2398
rect 32281 2352 32351 2398
rect 32397 2352 32467 2398
rect 32513 2352 32583 2398
rect 32629 2352 32699 2398
rect 32745 2352 32815 2398
rect 32861 2352 32931 2398
rect 32977 2352 33047 2398
rect 33093 2352 33163 2398
rect 33209 2352 33279 2398
rect 33325 2352 33395 2398
rect 33441 2352 33511 2398
rect 33557 2352 33627 2398
rect 33673 2352 33743 2398
rect 33789 2352 33859 2398
rect 33905 2352 33975 2398
rect 34021 2352 34091 2398
rect 34137 2352 34207 2398
rect 34253 2352 34323 2398
rect 34369 2352 34439 2398
rect 34485 2352 34555 2398
rect 34601 2352 34671 2398
rect 34717 2352 34787 2398
rect 34833 2352 34903 2398
rect 34949 2352 35019 2398
rect 35065 2352 35135 2398
rect 35181 2352 35251 2398
rect 35297 2352 35367 2398
rect 35413 2352 35483 2398
rect 35529 2352 35599 2398
rect 35645 2352 35715 2398
rect 35761 2352 35831 2398
rect 35877 2352 35947 2398
rect 35993 2352 36063 2398
rect 36109 2352 36179 2398
rect 36225 2352 36295 2398
rect 36341 2352 36411 2398
rect 36457 2352 36527 2398
rect 36573 2352 36643 2398
rect 36689 2352 36759 2398
rect 36805 2352 36875 2398
rect 36921 2352 36991 2398
rect 37037 2352 37107 2398
rect 37153 2352 37223 2398
rect 37269 2352 37339 2398
rect 37385 2352 37455 2398
rect 37501 2352 37571 2398
rect 37617 2352 37687 2398
rect 37733 2352 37803 2398
rect 37849 2352 37919 2398
rect 37965 2352 38035 2398
rect 38081 2352 38151 2398
rect 38197 2352 38267 2398
rect 38313 2352 38383 2398
rect 38429 2352 38499 2398
rect 38545 2352 38615 2398
rect 38661 2352 38731 2398
rect 38777 2352 38847 2398
rect 38893 2352 38963 2398
rect 39009 2352 39079 2398
rect 39125 2352 39195 2398
rect 39241 2352 39311 2398
rect 39357 2352 39427 2398
rect 39473 2352 39543 2398
rect 39589 2352 39659 2398
rect 39705 2352 39775 2398
rect 39821 2352 39891 2398
rect 39937 2352 40007 2398
rect 40053 2352 40123 2398
rect 40169 2352 40188 2398
rect 28620 2282 40188 2352
rect 28620 2236 28639 2282
rect 28685 2236 28755 2282
rect 28801 2236 28871 2282
rect 28917 2236 28987 2282
rect 29033 2236 29103 2282
rect 29149 2236 29219 2282
rect 29265 2236 29335 2282
rect 29381 2236 29451 2282
rect 29497 2236 29567 2282
rect 29613 2236 29683 2282
rect 29729 2236 29799 2282
rect 29845 2236 29915 2282
rect 29961 2236 30031 2282
rect 30077 2236 30147 2282
rect 30193 2236 30263 2282
rect 30309 2236 30379 2282
rect 30425 2236 30495 2282
rect 30541 2236 30611 2282
rect 30657 2236 30727 2282
rect 30773 2236 30843 2282
rect 30889 2236 30959 2282
rect 31005 2236 31075 2282
rect 31121 2236 31191 2282
rect 31237 2236 31307 2282
rect 31353 2236 31423 2282
rect 31469 2236 31539 2282
rect 31585 2236 31655 2282
rect 31701 2236 31771 2282
rect 31817 2236 31887 2282
rect 31933 2236 32003 2282
rect 32049 2236 32119 2282
rect 32165 2236 32235 2282
rect 32281 2236 32351 2282
rect 32397 2236 32467 2282
rect 32513 2236 32583 2282
rect 32629 2236 32699 2282
rect 32745 2236 32815 2282
rect 32861 2236 32931 2282
rect 32977 2236 33047 2282
rect 33093 2236 33163 2282
rect 33209 2236 33279 2282
rect 33325 2236 33395 2282
rect 33441 2236 33511 2282
rect 33557 2236 33627 2282
rect 33673 2236 33743 2282
rect 33789 2236 33859 2282
rect 33905 2236 33975 2282
rect 34021 2236 34091 2282
rect 34137 2236 34207 2282
rect 34253 2236 34323 2282
rect 34369 2236 34439 2282
rect 34485 2236 34555 2282
rect 34601 2236 34671 2282
rect 34717 2236 34787 2282
rect 34833 2236 34903 2282
rect 34949 2236 35019 2282
rect 35065 2236 35135 2282
rect 35181 2236 35251 2282
rect 35297 2236 35367 2282
rect 35413 2236 35483 2282
rect 35529 2236 35599 2282
rect 35645 2236 35715 2282
rect 35761 2236 35831 2282
rect 35877 2236 35947 2282
rect 35993 2236 36063 2282
rect 36109 2236 36179 2282
rect 36225 2236 36295 2282
rect 36341 2236 36411 2282
rect 36457 2236 36527 2282
rect 36573 2236 36643 2282
rect 36689 2236 36759 2282
rect 36805 2236 36875 2282
rect 36921 2236 36991 2282
rect 37037 2236 37107 2282
rect 37153 2236 37223 2282
rect 37269 2236 37339 2282
rect 37385 2236 37455 2282
rect 37501 2236 37571 2282
rect 37617 2236 37687 2282
rect 37733 2236 37803 2282
rect 37849 2236 37919 2282
rect 37965 2236 38035 2282
rect 38081 2236 38151 2282
rect 38197 2236 38267 2282
rect 38313 2236 38383 2282
rect 38429 2236 38499 2282
rect 38545 2236 38615 2282
rect 38661 2236 38731 2282
rect 38777 2236 38847 2282
rect 38893 2236 38963 2282
rect 39009 2236 39079 2282
rect 39125 2236 39195 2282
rect 39241 2236 39311 2282
rect 39357 2236 39427 2282
rect 39473 2236 39543 2282
rect 39589 2236 39659 2282
rect 39705 2236 39775 2282
rect 39821 2236 39891 2282
rect 39937 2236 40007 2282
rect 40053 2236 40123 2282
rect 40169 2236 40188 2282
rect 28620 2166 40188 2236
rect 28620 2120 28639 2166
rect 28685 2120 28755 2166
rect 28801 2120 28871 2166
rect 28917 2120 28987 2166
rect 29033 2120 29103 2166
rect 29149 2120 29219 2166
rect 29265 2120 29335 2166
rect 29381 2120 29451 2166
rect 29497 2120 29567 2166
rect 29613 2120 29683 2166
rect 29729 2120 29799 2166
rect 29845 2120 29915 2166
rect 29961 2120 30031 2166
rect 30077 2120 30147 2166
rect 30193 2120 30263 2166
rect 30309 2120 30379 2166
rect 30425 2120 30495 2166
rect 30541 2120 30611 2166
rect 30657 2120 30727 2166
rect 30773 2120 30843 2166
rect 30889 2120 30959 2166
rect 31005 2120 31075 2166
rect 31121 2120 31191 2166
rect 31237 2120 31307 2166
rect 31353 2120 31423 2166
rect 31469 2120 31539 2166
rect 31585 2120 31655 2166
rect 31701 2120 31771 2166
rect 31817 2120 31887 2166
rect 31933 2120 32003 2166
rect 32049 2120 32119 2166
rect 32165 2120 32235 2166
rect 32281 2120 32351 2166
rect 32397 2120 32467 2166
rect 32513 2120 32583 2166
rect 32629 2120 32699 2166
rect 32745 2120 32815 2166
rect 32861 2120 32931 2166
rect 32977 2120 33047 2166
rect 33093 2120 33163 2166
rect 33209 2120 33279 2166
rect 33325 2120 33395 2166
rect 33441 2120 33511 2166
rect 33557 2120 33627 2166
rect 33673 2120 33743 2166
rect 33789 2120 33859 2166
rect 33905 2120 33975 2166
rect 34021 2120 34091 2166
rect 34137 2120 34207 2166
rect 34253 2120 34323 2166
rect 34369 2120 34439 2166
rect 34485 2120 34555 2166
rect 34601 2120 34671 2166
rect 34717 2120 34787 2166
rect 34833 2120 34903 2166
rect 34949 2120 35019 2166
rect 35065 2120 35135 2166
rect 35181 2120 35251 2166
rect 35297 2120 35367 2166
rect 35413 2120 35483 2166
rect 35529 2120 35599 2166
rect 35645 2120 35715 2166
rect 35761 2120 35831 2166
rect 35877 2120 35947 2166
rect 35993 2120 36063 2166
rect 36109 2120 36179 2166
rect 36225 2120 36295 2166
rect 36341 2120 36411 2166
rect 36457 2120 36527 2166
rect 36573 2120 36643 2166
rect 36689 2120 36759 2166
rect 36805 2120 36875 2166
rect 36921 2120 36991 2166
rect 37037 2120 37107 2166
rect 37153 2120 37223 2166
rect 37269 2120 37339 2166
rect 37385 2120 37455 2166
rect 37501 2120 37571 2166
rect 37617 2120 37687 2166
rect 37733 2120 37803 2166
rect 37849 2120 37919 2166
rect 37965 2120 38035 2166
rect 38081 2120 38151 2166
rect 38197 2120 38267 2166
rect 38313 2120 38383 2166
rect 38429 2120 38499 2166
rect 38545 2120 38615 2166
rect 38661 2120 38731 2166
rect 38777 2120 38847 2166
rect 38893 2120 38963 2166
rect 39009 2120 39079 2166
rect 39125 2120 39195 2166
rect 39241 2120 39311 2166
rect 39357 2120 39427 2166
rect 39473 2120 39543 2166
rect 39589 2120 39659 2166
rect 39705 2120 39775 2166
rect 39821 2120 39891 2166
rect 39937 2120 40007 2166
rect 40053 2120 40123 2166
rect 40169 2120 40188 2166
rect 28620 2050 40188 2120
rect 28620 2004 28639 2050
rect 28685 2004 28755 2050
rect 28801 2004 28871 2050
rect 28917 2004 28987 2050
rect 29033 2004 29103 2050
rect 29149 2004 29219 2050
rect 29265 2004 29335 2050
rect 29381 2004 29451 2050
rect 29497 2004 29567 2050
rect 29613 2004 29683 2050
rect 29729 2004 29799 2050
rect 29845 2004 29915 2050
rect 29961 2004 30031 2050
rect 30077 2004 30147 2050
rect 30193 2004 30263 2050
rect 30309 2004 30379 2050
rect 30425 2004 30495 2050
rect 30541 2004 30611 2050
rect 30657 2004 30727 2050
rect 30773 2004 30843 2050
rect 30889 2004 30959 2050
rect 31005 2004 31075 2050
rect 31121 2004 31191 2050
rect 31237 2004 31307 2050
rect 31353 2004 31423 2050
rect 31469 2004 31539 2050
rect 31585 2004 31655 2050
rect 31701 2004 31771 2050
rect 31817 2004 31887 2050
rect 31933 2004 32003 2050
rect 32049 2004 32119 2050
rect 32165 2004 32235 2050
rect 32281 2004 32351 2050
rect 32397 2004 32467 2050
rect 32513 2004 32583 2050
rect 32629 2004 32699 2050
rect 32745 2004 32815 2050
rect 32861 2004 32931 2050
rect 32977 2004 33047 2050
rect 33093 2004 33163 2050
rect 33209 2004 33279 2050
rect 33325 2004 33395 2050
rect 33441 2004 33511 2050
rect 33557 2004 33627 2050
rect 33673 2004 33743 2050
rect 33789 2004 33859 2050
rect 33905 2004 33975 2050
rect 34021 2004 34091 2050
rect 34137 2004 34207 2050
rect 34253 2004 34323 2050
rect 34369 2004 34439 2050
rect 34485 2004 34555 2050
rect 34601 2004 34671 2050
rect 34717 2004 34787 2050
rect 34833 2004 34903 2050
rect 34949 2004 35019 2050
rect 35065 2004 35135 2050
rect 35181 2004 35251 2050
rect 35297 2004 35367 2050
rect 35413 2004 35483 2050
rect 35529 2004 35599 2050
rect 35645 2004 35715 2050
rect 35761 2004 35831 2050
rect 35877 2004 35947 2050
rect 35993 2004 36063 2050
rect 36109 2004 36179 2050
rect 36225 2004 36295 2050
rect 36341 2004 36411 2050
rect 36457 2004 36527 2050
rect 36573 2004 36643 2050
rect 36689 2004 36759 2050
rect 36805 2004 36875 2050
rect 36921 2004 36991 2050
rect 37037 2004 37107 2050
rect 37153 2004 37223 2050
rect 37269 2004 37339 2050
rect 37385 2004 37455 2050
rect 37501 2004 37571 2050
rect 37617 2004 37687 2050
rect 37733 2004 37803 2050
rect 37849 2004 37919 2050
rect 37965 2004 38035 2050
rect 38081 2004 38151 2050
rect 38197 2004 38267 2050
rect 38313 2004 38383 2050
rect 38429 2004 38499 2050
rect 38545 2004 38615 2050
rect 38661 2004 38731 2050
rect 38777 2004 38847 2050
rect 38893 2004 38963 2050
rect 39009 2004 39079 2050
rect 39125 2004 39195 2050
rect 39241 2004 39311 2050
rect 39357 2004 39427 2050
rect 39473 2004 39543 2050
rect 39589 2004 39659 2050
rect 39705 2004 39775 2050
rect 39821 2004 39891 2050
rect 39937 2004 40007 2050
rect 40053 2004 40123 2050
rect 40169 2004 40188 2050
rect 28620 1934 40188 2004
rect 28620 1888 28639 1934
rect 28685 1888 28755 1934
rect 28801 1888 28871 1934
rect 28917 1888 28987 1934
rect 29033 1888 29103 1934
rect 29149 1888 29219 1934
rect 29265 1888 29335 1934
rect 29381 1888 29451 1934
rect 29497 1888 29567 1934
rect 29613 1888 29683 1934
rect 29729 1888 29799 1934
rect 29845 1888 29915 1934
rect 29961 1888 30031 1934
rect 30077 1888 30147 1934
rect 30193 1888 30263 1934
rect 30309 1888 30379 1934
rect 30425 1888 30495 1934
rect 30541 1888 30611 1934
rect 30657 1888 30727 1934
rect 30773 1888 30843 1934
rect 30889 1888 30959 1934
rect 31005 1888 31075 1934
rect 31121 1888 31191 1934
rect 31237 1888 31307 1934
rect 31353 1888 31423 1934
rect 31469 1888 31539 1934
rect 31585 1888 31655 1934
rect 31701 1888 31771 1934
rect 31817 1888 31887 1934
rect 31933 1888 32003 1934
rect 32049 1888 32119 1934
rect 32165 1888 32235 1934
rect 32281 1888 32351 1934
rect 32397 1888 32467 1934
rect 32513 1888 32583 1934
rect 32629 1888 32699 1934
rect 32745 1888 32815 1934
rect 32861 1888 32931 1934
rect 32977 1888 33047 1934
rect 33093 1888 33163 1934
rect 33209 1888 33279 1934
rect 33325 1888 33395 1934
rect 33441 1888 33511 1934
rect 33557 1888 33627 1934
rect 33673 1888 33743 1934
rect 33789 1888 33859 1934
rect 33905 1888 33975 1934
rect 34021 1888 34091 1934
rect 34137 1888 34207 1934
rect 34253 1888 34323 1934
rect 34369 1888 34439 1934
rect 34485 1888 34555 1934
rect 34601 1888 34671 1934
rect 34717 1888 34787 1934
rect 34833 1888 34903 1934
rect 34949 1888 35019 1934
rect 35065 1888 35135 1934
rect 35181 1888 35251 1934
rect 35297 1888 35367 1934
rect 35413 1888 35483 1934
rect 35529 1888 35599 1934
rect 35645 1888 35715 1934
rect 35761 1888 35831 1934
rect 35877 1888 35947 1934
rect 35993 1888 36063 1934
rect 36109 1888 36179 1934
rect 36225 1888 36295 1934
rect 36341 1888 36411 1934
rect 36457 1888 36527 1934
rect 36573 1888 36643 1934
rect 36689 1888 36759 1934
rect 36805 1888 36875 1934
rect 36921 1888 36991 1934
rect 37037 1888 37107 1934
rect 37153 1888 37223 1934
rect 37269 1888 37339 1934
rect 37385 1888 37455 1934
rect 37501 1888 37571 1934
rect 37617 1888 37687 1934
rect 37733 1888 37803 1934
rect 37849 1888 37919 1934
rect 37965 1888 38035 1934
rect 38081 1888 38151 1934
rect 38197 1888 38267 1934
rect 38313 1888 38383 1934
rect 38429 1888 38499 1934
rect 38545 1888 38615 1934
rect 38661 1888 38731 1934
rect 38777 1888 38847 1934
rect 38893 1888 38963 1934
rect 39009 1888 39079 1934
rect 39125 1888 39195 1934
rect 39241 1888 39311 1934
rect 39357 1888 39427 1934
rect 39473 1888 39543 1934
rect 39589 1888 39659 1934
rect 39705 1888 39775 1934
rect 39821 1888 39891 1934
rect 39937 1888 40007 1934
rect 40053 1888 40123 1934
rect 40169 1888 40188 1934
rect 28620 1818 40188 1888
rect 28620 1772 28639 1818
rect 28685 1772 28755 1818
rect 28801 1772 28871 1818
rect 28917 1772 28987 1818
rect 29033 1772 29103 1818
rect 29149 1772 29219 1818
rect 29265 1772 29335 1818
rect 29381 1772 29451 1818
rect 29497 1772 29567 1818
rect 29613 1772 29683 1818
rect 29729 1772 29799 1818
rect 29845 1772 29915 1818
rect 29961 1772 30031 1818
rect 30077 1772 30147 1818
rect 30193 1772 30263 1818
rect 30309 1772 30379 1818
rect 30425 1772 30495 1818
rect 30541 1772 30611 1818
rect 30657 1772 30727 1818
rect 30773 1772 30843 1818
rect 30889 1772 30959 1818
rect 31005 1772 31075 1818
rect 31121 1772 31191 1818
rect 31237 1772 31307 1818
rect 31353 1772 31423 1818
rect 31469 1772 31539 1818
rect 31585 1772 31655 1818
rect 31701 1772 31771 1818
rect 31817 1772 31887 1818
rect 31933 1772 32003 1818
rect 32049 1772 32119 1818
rect 32165 1772 32235 1818
rect 32281 1772 32351 1818
rect 32397 1772 32467 1818
rect 32513 1772 32583 1818
rect 32629 1772 32699 1818
rect 32745 1772 32815 1818
rect 32861 1772 32931 1818
rect 32977 1772 33047 1818
rect 33093 1772 33163 1818
rect 33209 1772 33279 1818
rect 33325 1772 33395 1818
rect 33441 1772 33511 1818
rect 33557 1772 33627 1818
rect 33673 1772 33743 1818
rect 33789 1772 33859 1818
rect 33905 1772 33975 1818
rect 34021 1772 34091 1818
rect 34137 1772 34207 1818
rect 34253 1772 34323 1818
rect 34369 1772 34439 1818
rect 34485 1772 34555 1818
rect 34601 1772 34671 1818
rect 34717 1772 34787 1818
rect 34833 1772 34903 1818
rect 34949 1772 35019 1818
rect 35065 1772 35135 1818
rect 35181 1772 35251 1818
rect 35297 1772 35367 1818
rect 35413 1772 35483 1818
rect 35529 1772 35599 1818
rect 35645 1772 35715 1818
rect 35761 1772 35831 1818
rect 35877 1772 35947 1818
rect 35993 1772 36063 1818
rect 36109 1772 36179 1818
rect 36225 1772 36295 1818
rect 36341 1772 36411 1818
rect 36457 1772 36527 1818
rect 36573 1772 36643 1818
rect 36689 1772 36759 1818
rect 36805 1772 36875 1818
rect 36921 1772 36991 1818
rect 37037 1772 37107 1818
rect 37153 1772 37223 1818
rect 37269 1772 37339 1818
rect 37385 1772 37455 1818
rect 37501 1772 37571 1818
rect 37617 1772 37687 1818
rect 37733 1772 37803 1818
rect 37849 1772 37919 1818
rect 37965 1772 38035 1818
rect 38081 1772 38151 1818
rect 38197 1772 38267 1818
rect 38313 1772 38383 1818
rect 38429 1772 38499 1818
rect 38545 1772 38615 1818
rect 38661 1772 38731 1818
rect 38777 1772 38847 1818
rect 38893 1772 38963 1818
rect 39009 1772 39079 1818
rect 39125 1772 39195 1818
rect 39241 1772 39311 1818
rect 39357 1772 39427 1818
rect 39473 1772 39543 1818
rect 39589 1772 39659 1818
rect 39705 1772 39775 1818
rect 39821 1772 39891 1818
rect 39937 1772 40007 1818
rect 40053 1772 40123 1818
rect 40169 1772 40188 1818
rect 28620 1702 40188 1772
rect 28620 1656 28639 1702
rect 28685 1656 28755 1702
rect 28801 1656 28871 1702
rect 28917 1656 28987 1702
rect 29033 1656 29103 1702
rect 29149 1656 29219 1702
rect 29265 1656 29335 1702
rect 29381 1656 29451 1702
rect 29497 1656 29567 1702
rect 29613 1656 29683 1702
rect 29729 1656 29799 1702
rect 29845 1656 29915 1702
rect 29961 1656 30031 1702
rect 30077 1656 30147 1702
rect 30193 1656 30263 1702
rect 30309 1656 30379 1702
rect 30425 1656 30495 1702
rect 30541 1656 30611 1702
rect 30657 1656 30727 1702
rect 30773 1656 30843 1702
rect 30889 1656 30959 1702
rect 31005 1656 31075 1702
rect 31121 1656 31191 1702
rect 31237 1656 31307 1702
rect 31353 1656 31423 1702
rect 31469 1656 31539 1702
rect 31585 1656 31655 1702
rect 31701 1656 31771 1702
rect 31817 1656 31887 1702
rect 31933 1656 32003 1702
rect 32049 1656 32119 1702
rect 32165 1656 32235 1702
rect 32281 1656 32351 1702
rect 32397 1656 32467 1702
rect 32513 1656 32583 1702
rect 32629 1656 32699 1702
rect 32745 1656 32815 1702
rect 32861 1656 32931 1702
rect 32977 1656 33047 1702
rect 33093 1656 33163 1702
rect 33209 1656 33279 1702
rect 33325 1656 33395 1702
rect 33441 1656 33511 1702
rect 33557 1656 33627 1702
rect 33673 1656 33743 1702
rect 33789 1656 33859 1702
rect 33905 1656 33975 1702
rect 34021 1656 34091 1702
rect 34137 1656 34207 1702
rect 34253 1656 34323 1702
rect 34369 1656 34439 1702
rect 34485 1656 34555 1702
rect 34601 1656 34671 1702
rect 34717 1656 34787 1702
rect 34833 1656 34903 1702
rect 34949 1656 35019 1702
rect 35065 1656 35135 1702
rect 35181 1656 35251 1702
rect 35297 1656 35367 1702
rect 35413 1656 35483 1702
rect 35529 1656 35599 1702
rect 35645 1656 35715 1702
rect 35761 1656 35831 1702
rect 35877 1656 35947 1702
rect 35993 1656 36063 1702
rect 36109 1656 36179 1702
rect 36225 1656 36295 1702
rect 36341 1656 36411 1702
rect 36457 1656 36527 1702
rect 36573 1656 36643 1702
rect 36689 1656 36759 1702
rect 36805 1656 36875 1702
rect 36921 1656 36991 1702
rect 37037 1656 37107 1702
rect 37153 1656 37223 1702
rect 37269 1656 37339 1702
rect 37385 1656 37455 1702
rect 37501 1656 37571 1702
rect 37617 1656 37687 1702
rect 37733 1656 37803 1702
rect 37849 1656 37919 1702
rect 37965 1656 38035 1702
rect 38081 1656 38151 1702
rect 38197 1656 38267 1702
rect 38313 1656 38383 1702
rect 38429 1656 38499 1702
rect 38545 1656 38615 1702
rect 38661 1656 38731 1702
rect 38777 1656 38847 1702
rect 38893 1656 38963 1702
rect 39009 1656 39079 1702
rect 39125 1656 39195 1702
rect 39241 1656 39311 1702
rect 39357 1656 39427 1702
rect 39473 1656 39543 1702
rect 39589 1656 39659 1702
rect 39705 1656 39775 1702
rect 39821 1656 39891 1702
rect 39937 1656 40007 1702
rect 40053 1656 40123 1702
rect 40169 1656 40188 1702
rect 28620 1637 40188 1656
rect 50826 3906 56594 3925
rect 50826 3860 50845 3906
rect 50891 3860 50961 3906
rect 51007 3860 51077 3906
rect 51123 3860 51193 3906
rect 51239 3860 51309 3906
rect 51355 3860 51425 3906
rect 51471 3860 51541 3906
rect 51587 3860 51657 3906
rect 51703 3860 51773 3906
rect 51819 3860 51889 3906
rect 51935 3860 52005 3906
rect 52051 3860 52121 3906
rect 52167 3860 52237 3906
rect 52283 3860 52353 3906
rect 52399 3860 52469 3906
rect 52515 3860 52585 3906
rect 52631 3860 52701 3906
rect 52747 3860 52817 3906
rect 52863 3860 52933 3906
rect 52979 3860 53049 3906
rect 53095 3860 53165 3906
rect 53211 3860 53281 3906
rect 53327 3860 53397 3906
rect 53443 3860 53513 3906
rect 53559 3860 53629 3906
rect 53675 3860 53745 3906
rect 53791 3860 53861 3906
rect 53907 3860 53977 3906
rect 54023 3860 54093 3906
rect 54139 3860 54209 3906
rect 54255 3860 54325 3906
rect 54371 3860 54441 3906
rect 54487 3860 54557 3906
rect 54603 3860 54673 3906
rect 54719 3860 54789 3906
rect 54835 3860 54905 3906
rect 54951 3860 55021 3906
rect 55067 3860 55137 3906
rect 55183 3860 55253 3906
rect 55299 3860 55369 3906
rect 55415 3860 55485 3906
rect 55531 3860 55601 3906
rect 55647 3860 55717 3906
rect 55763 3860 55833 3906
rect 55879 3860 55949 3906
rect 55995 3860 56065 3906
rect 56111 3860 56181 3906
rect 56227 3860 56297 3906
rect 56343 3860 56413 3906
rect 56459 3860 56529 3906
rect 56575 3860 56594 3906
rect 50826 3790 56594 3860
rect 50826 3744 50845 3790
rect 50891 3744 50961 3790
rect 51007 3744 51077 3790
rect 51123 3744 51193 3790
rect 51239 3744 51309 3790
rect 51355 3744 51425 3790
rect 51471 3744 51541 3790
rect 51587 3744 51657 3790
rect 51703 3744 51773 3790
rect 51819 3744 51889 3790
rect 51935 3744 52005 3790
rect 52051 3744 52121 3790
rect 52167 3744 52237 3790
rect 52283 3744 52353 3790
rect 52399 3744 52469 3790
rect 52515 3744 52585 3790
rect 52631 3744 52701 3790
rect 52747 3744 52817 3790
rect 52863 3744 52933 3790
rect 52979 3744 53049 3790
rect 53095 3744 53165 3790
rect 53211 3744 53281 3790
rect 53327 3744 53397 3790
rect 53443 3744 53513 3790
rect 53559 3744 53629 3790
rect 53675 3744 53745 3790
rect 53791 3744 53861 3790
rect 53907 3744 53977 3790
rect 54023 3744 54093 3790
rect 54139 3744 54209 3790
rect 54255 3744 54325 3790
rect 54371 3744 54441 3790
rect 54487 3744 54557 3790
rect 54603 3744 54673 3790
rect 54719 3744 54789 3790
rect 54835 3744 54905 3790
rect 54951 3744 55021 3790
rect 55067 3744 55137 3790
rect 55183 3744 55253 3790
rect 55299 3744 55369 3790
rect 55415 3744 55485 3790
rect 55531 3744 55601 3790
rect 55647 3744 55717 3790
rect 55763 3744 55833 3790
rect 55879 3744 55949 3790
rect 55995 3744 56065 3790
rect 56111 3744 56181 3790
rect 56227 3744 56297 3790
rect 56343 3744 56413 3790
rect 56459 3744 56529 3790
rect 56575 3744 56594 3790
rect 50826 3674 56594 3744
rect 50826 3628 50845 3674
rect 50891 3628 50961 3674
rect 51007 3628 51077 3674
rect 51123 3628 51193 3674
rect 51239 3628 51309 3674
rect 51355 3628 51425 3674
rect 51471 3628 51541 3674
rect 51587 3628 51657 3674
rect 51703 3628 51773 3674
rect 51819 3628 51889 3674
rect 51935 3628 52005 3674
rect 52051 3628 52121 3674
rect 52167 3628 52237 3674
rect 52283 3628 52353 3674
rect 52399 3628 52469 3674
rect 52515 3628 52585 3674
rect 52631 3628 52701 3674
rect 52747 3628 52817 3674
rect 52863 3628 52933 3674
rect 52979 3628 53049 3674
rect 53095 3628 53165 3674
rect 53211 3628 53281 3674
rect 53327 3628 53397 3674
rect 53443 3628 53513 3674
rect 53559 3628 53629 3674
rect 53675 3628 53745 3674
rect 53791 3628 53861 3674
rect 53907 3628 53977 3674
rect 54023 3628 54093 3674
rect 54139 3628 54209 3674
rect 54255 3628 54325 3674
rect 54371 3628 54441 3674
rect 54487 3628 54557 3674
rect 54603 3628 54673 3674
rect 54719 3628 54789 3674
rect 54835 3628 54905 3674
rect 54951 3628 55021 3674
rect 55067 3628 55137 3674
rect 55183 3628 55253 3674
rect 55299 3628 55369 3674
rect 55415 3628 55485 3674
rect 55531 3628 55601 3674
rect 55647 3628 55717 3674
rect 55763 3628 55833 3674
rect 55879 3628 55949 3674
rect 55995 3628 56065 3674
rect 56111 3628 56181 3674
rect 56227 3628 56297 3674
rect 56343 3628 56413 3674
rect 56459 3628 56529 3674
rect 56575 3628 56594 3674
rect 50826 3558 56594 3628
rect 50826 3512 50845 3558
rect 50891 3512 50961 3558
rect 51007 3512 51077 3558
rect 51123 3512 51193 3558
rect 51239 3512 51309 3558
rect 51355 3512 51425 3558
rect 51471 3512 51541 3558
rect 51587 3512 51657 3558
rect 51703 3512 51773 3558
rect 51819 3512 51889 3558
rect 51935 3512 52005 3558
rect 52051 3512 52121 3558
rect 52167 3512 52237 3558
rect 52283 3512 52353 3558
rect 52399 3512 52469 3558
rect 52515 3512 52585 3558
rect 52631 3512 52701 3558
rect 52747 3512 52817 3558
rect 52863 3512 52933 3558
rect 52979 3512 53049 3558
rect 53095 3512 53165 3558
rect 53211 3512 53281 3558
rect 53327 3512 53397 3558
rect 53443 3512 53513 3558
rect 53559 3512 53629 3558
rect 53675 3512 53745 3558
rect 53791 3512 53861 3558
rect 53907 3512 53977 3558
rect 54023 3512 54093 3558
rect 54139 3512 54209 3558
rect 54255 3512 54325 3558
rect 54371 3512 54441 3558
rect 54487 3512 54557 3558
rect 54603 3512 54673 3558
rect 54719 3512 54789 3558
rect 54835 3512 54905 3558
rect 54951 3512 55021 3558
rect 55067 3512 55137 3558
rect 55183 3512 55253 3558
rect 55299 3512 55369 3558
rect 55415 3512 55485 3558
rect 55531 3512 55601 3558
rect 55647 3512 55717 3558
rect 55763 3512 55833 3558
rect 55879 3512 55949 3558
rect 55995 3512 56065 3558
rect 56111 3512 56181 3558
rect 56227 3512 56297 3558
rect 56343 3512 56413 3558
rect 56459 3512 56529 3558
rect 56575 3512 56594 3558
rect 50826 3442 56594 3512
rect 50826 3396 50845 3442
rect 50891 3396 50961 3442
rect 51007 3396 51077 3442
rect 51123 3396 51193 3442
rect 51239 3396 51309 3442
rect 51355 3396 51425 3442
rect 51471 3396 51541 3442
rect 51587 3396 51657 3442
rect 51703 3396 51773 3442
rect 51819 3396 51889 3442
rect 51935 3396 52005 3442
rect 52051 3396 52121 3442
rect 52167 3396 52237 3442
rect 52283 3396 52353 3442
rect 52399 3396 52469 3442
rect 52515 3396 52585 3442
rect 52631 3396 52701 3442
rect 52747 3396 52817 3442
rect 52863 3396 52933 3442
rect 52979 3396 53049 3442
rect 53095 3396 53165 3442
rect 53211 3396 53281 3442
rect 53327 3396 53397 3442
rect 53443 3396 53513 3442
rect 53559 3396 53629 3442
rect 53675 3396 53745 3442
rect 53791 3396 53861 3442
rect 53907 3396 53977 3442
rect 54023 3396 54093 3442
rect 54139 3396 54209 3442
rect 54255 3396 54325 3442
rect 54371 3396 54441 3442
rect 54487 3396 54557 3442
rect 54603 3396 54673 3442
rect 54719 3396 54789 3442
rect 54835 3396 54905 3442
rect 54951 3396 55021 3442
rect 55067 3396 55137 3442
rect 55183 3396 55253 3442
rect 55299 3396 55369 3442
rect 55415 3396 55485 3442
rect 55531 3396 55601 3442
rect 55647 3396 55717 3442
rect 55763 3396 55833 3442
rect 55879 3396 55949 3442
rect 55995 3396 56065 3442
rect 56111 3396 56181 3442
rect 56227 3396 56297 3442
rect 56343 3396 56413 3442
rect 56459 3396 56529 3442
rect 56575 3396 56594 3442
rect 50826 3326 56594 3396
rect 50826 3280 50845 3326
rect 50891 3280 50961 3326
rect 51007 3280 51077 3326
rect 51123 3280 51193 3326
rect 51239 3280 51309 3326
rect 51355 3280 51425 3326
rect 51471 3280 51541 3326
rect 51587 3280 51657 3326
rect 51703 3280 51773 3326
rect 51819 3280 51889 3326
rect 51935 3280 52005 3326
rect 52051 3280 52121 3326
rect 52167 3280 52237 3326
rect 52283 3280 52353 3326
rect 52399 3280 52469 3326
rect 52515 3280 52585 3326
rect 52631 3280 52701 3326
rect 52747 3280 52817 3326
rect 52863 3280 52933 3326
rect 52979 3280 53049 3326
rect 53095 3280 53165 3326
rect 53211 3280 53281 3326
rect 53327 3280 53397 3326
rect 53443 3280 53513 3326
rect 53559 3280 53629 3326
rect 53675 3280 53745 3326
rect 53791 3280 53861 3326
rect 53907 3280 53977 3326
rect 54023 3280 54093 3326
rect 54139 3280 54209 3326
rect 54255 3280 54325 3326
rect 54371 3280 54441 3326
rect 54487 3280 54557 3326
rect 54603 3280 54673 3326
rect 54719 3280 54789 3326
rect 54835 3280 54905 3326
rect 54951 3280 55021 3326
rect 55067 3280 55137 3326
rect 55183 3280 55253 3326
rect 55299 3280 55369 3326
rect 55415 3280 55485 3326
rect 55531 3280 55601 3326
rect 55647 3280 55717 3326
rect 55763 3280 55833 3326
rect 55879 3280 55949 3326
rect 55995 3280 56065 3326
rect 56111 3280 56181 3326
rect 56227 3280 56297 3326
rect 56343 3280 56413 3326
rect 56459 3280 56529 3326
rect 56575 3280 56594 3326
rect 50826 3210 56594 3280
rect 50826 3164 50845 3210
rect 50891 3164 50961 3210
rect 51007 3164 51077 3210
rect 51123 3164 51193 3210
rect 51239 3164 51309 3210
rect 51355 3164 51425 3210
rect 51471 3164 51541 3210
rect 51587 3164 51657 3210
rect 51703 3164 51773 3210
rect 51819 3164 51889 3210
rect 51935 3164 52005 3210
rect 52051 3164 52121 3210
rect 52167 3164 52237 3210
rect 52283 3164 52353 3210
rect 52399 3164 52469 3210
rect 52515 3164 52585 3210
rect 52631 3164 52701 3210
rect 52747 3164 52817 3210
rect 52863 3164 52933 3210
rect 52979 3164 53049 3210
rect 53095 3164 53165 3210
rect 53211 3164 53281 3210
rect 53327 3164 53397 3210
rect 53443 3164 53513 3210
rect 53559 3164 53629 3210
rect 53675 3164 53745 3210
rect 53791 3164 53861 3210
rect 53907 3164 53977 3210
rect 54023 3164 54093 3210
rect 54139 3164 54209 3210
rect 54255 3164 54325 3210
rect 54371 3164 54441 3210
rect 54487 3164 54557 3210
rect 54603 3164 54673 3210
rect 54719 3164 54789 3210
rect 54835 3164 54905 3210
rect 54951 3164 55021 3210
rect 55067 3164 55137 3210
rect 55183 3164 55253 3210
rect 55299 3164 55369 3210
rect 55415 3164 55485 3210
rect 55531 3164 55601 3210
rect 55647 3164 55717 3210
rect 55763 3164 55833 3210
rect 55879 3164 55949 3210
rect 55995 3164 56065 3210
rect 56111 3164 56181 3210
rect 56227 3164 56297 3210
rect 56343 3164 56413 3210
rect 56459 3164 56529 3210
rect 56575 3164 56594 3210
rect 50826 3094 56594 3164
rect 50826 3048 50845 3094
rect 50891 3048 50961 3094
rect 51007 3048 51077 3094
rect 51123 3048 51193 3094
rect 51239 3048 51309 3094
rect 51355 3048 51425 3094
rect 51471 3048 51541 3094
rect 51587 3048 51657 3094
rect 51703 3048 51773 3094
rect 51819 3048 51889 3094
rect 51935 3048 52005 3094
rect 52051 3048 52121 3094
rect 52167 3048 52237 3094
rect 52283 3048 52353 3094
rect 52399 3048 52469 3094
rect 52515 3048 52585 3094
rect 52631 3048 52701 3094
rect 52747 3048 52817 3094
rect 52863 3048 52933 3094
rect 52979 3048 53049 3094
rect 53095 3048 53165 3094
rect 53211 3048 53281 3094
rect 53327 3048 53397 3094
rect 53443 3048 53513 3094
rect 53559 3048 53629 3094
rect 53675 3048 53745 3094
rect 53791 3048 53861 3094
rect 53907 3048 53977 3094
rect 54023 3048 54093 3094
rect 54139 3048 54209 3094
rect 54255 3048 54325 3094
rect 54371 3048 54441 3094
rect 54487 3048 54557 3094
rect 54603 3048 54673 3094
rect 54719 3048 54789 3094
rect 54835 3048 54905 3094
rect 54951 3048 55021 3094
rect 55067 3048 55137 3094
rect 55183 3048 55253 3094
rect 55299 3048 55369 3094
rect 55415 3048 55485 3094
rect 55531 3048 55601 3094
rect 55647 3048 55717 3094
rect 55763 3048 55833 3094
rect 55879 3048 55949 3094
rect 55995 3048 56065 3094
rect 56111 3048 56181 3094
rect 56227 3048 56297 3094
rect 56343 3048 56413 3094
rect 56459 3048 56529 3094
rect 56575 3048 56594 3094
rect 50826 2978 56594 3048
rect 50826 2932 50845 2978
rect 50891 2932 50961 2978
rect 51007 2932 51077 2978
rect 51123 2932 51193 2978
rect 51239 2932 51309 2978
rect 51355 2932 51425 2978
rect 51471 2932 51541 2978
rect 51587 2932 51657 2978
rect 51703 2932 51773 2978
rect 51819 2932 51889 2978
rect 51935 2932 52005 2978
rect 52051 2932 52121 2978
rect 52167 2932 52237 2978
rect 52283 2932 52353 2978
rect 52399 2932 52469 2978
rect 52515 2932 52585 2978
rect 52631 2932 52701 2978
rect 52747 2932 52817 2978
rect 52863 2932 52933 2978
rect 52979 2932 53049 2978
rect 53095 2932 53165 2978
rect 53211 2932 53281 2978
rect 53327 2932 53397 2978
rect 53443 2932 53513 2978
rect 53559 2932 53629 2978
rect 53675 2932 53745 2978
rect 53791 2932 53861 2978
rect 53907 2932 53977 2978
rect 54023 2932 54093 2978
rect 54139 2932 54209 2978
rect 54255 2932 54325 2978
rect 54371 2932 54441 2978
rect 54487 2932 54557 2978
rect 54603 2932 54673 2978
rect 54719 2932 54789 2978
rect 54835 2932 54905 2978
rect 54951 2932 55021 2978
rect 55067 2932 55137 2978
rect 55183 2932 55253 2978
rect 55299 2932 55369 2978
rect 55415 2932 55485 2978
rect 55531 2932 55601 2978
rect 55647 2932 55717 2978
rect 55763 2932 55833 2978
rect 55879 2932 55949 2978
rect 55995 2932 56065 2978
rect 56111 2932 56181 2978
rect 56227 2932 56297 2978
rect 56343 2932 56413 2978
rect 56459 2932 56529 2978
rect 56575 2932 56594 2978
rect 50826 2862 56594 2932
rect 50826 2816 50845 2862
rect 50891 2816 50961 2862
rect 51007 2816 51077 2862
rect 51123 2816 51193 2862
rect 51239 2816 51309 2862
rect 51355 2816 51425 2862
rect 51471 2816 51541 2862
rect 51587 2816 51657 2862
rect 51703 2816 51773 2862
rect 51819 2816 51889 2862
rect 51935 2816 52005 2862
rect 52051 2816 52121 2862
rect 52167 2816 52237 2862
rect 52283 2816 52353 2862
rect 52399 2816 52469 2862
rect 52515 2816 52585 2862
rect 52631 2816 52701 2862
rect 52747 2816 52817 2862
rect 52863 2816 52933 2862
rect 52979 2816 53049 2862
rect 53095 2816 53165 2862
rect 53211 2816 53281 2862
rect 53327 2816 53397 2862
rect 53443 2816 53513 2862
rect 53559 2816 53629 2862
rect 53675 2816 53745 2862
rect 53791 2816 53861 2862
rect 53907 2816 53977 2862
rect 54023 2816 54093 2862
rect 54139 2816 54209 2862
rect 54255 2816 54325 2862
rect 54371 2816 54441 2862
rect 54487 2816 54557 2862
rect 54603 2816 54673 2862
rect 54719 2816 54789 2862
rect 54835 2816 54905 2862
rect 54951 2816 55021 2862
rect 55067 2816 55137 2862
rect 55183 2816 55253 2862
rect 55299 2816 55369 2862
rect 55415 2816 55485 2862
rect 55531 2816 55601 2862
rect 55647 2816 55717 2862
rect 55763 2816 55833 2862
rect 55879 2816 55949 2862
rect 55995 2816 56065 2862
rect 56111 2816 56181 2862
rect 56227 2816 56297 2862
rect 56343 2816 56413 2862
rect 56459 2816 56529 2862
rect 56575 2816 56594 2862
rect 50826 2746 56594 2816
rect 50826 2700 50845 2746
rect 50891 2700 50961 2746
rect 51007 2700 51077 2746
rect 51123 2700 51193 2746
rect 51239 2700 51309 2746
rect 51355 2700 51425 2746
rect 51471 2700 51541 2746
rect 51587 2700 51657 2746
rect 51703 2700 51773 2746
rect 51819 2700 51889 2746
rect 51935 2700 52005 2746
rect 52051 2700 52121 2746
rect 52167 2700 52237 2746
rect 52283 2700 52353 2746
rect 52399 2700 52469 2746
rect 52515 2700 52585 2746
rect 52631 2700 52701 2746
rect 52747 2700 52817 2746
rect 52863 2700 52933 2746
rect 52979 2700 53049 2746
rect 53095 2700 53165 2746
rect 53211 2700 53281 2746
rect 53327 2700 53397 2746
rect 53443 2700 53513 2746
rect 53559 2700 53629 2746
rect 53675 2700 53745 2746
rect 53791 2700 53861 2746
rect 53907 2700 53977 2746
rect 54023 2700 54093 2746
rect 54139 2700 54209 2746
rect 54255 2700 54325 2746
rect 54371 2700 54441 2746
rect 54487 2700 54557 2746
rect 54603 2700 54673 2746
rect 54719 2700 54789 2746
rect 54835 2700 54905 2746
rect 54951 2700 55021 2746
rect 55067 2700 55137 2746
rect 55183 2700 55253 2746
rect 55299 2700 55369 2746
rect 55415 2700 55485 2746
rect 55531 2700 55601 2746
rect 55647 2700 55717 2746
rect 55763 2700 55833 2746
rect 55879 2700 55949 2746
rect 55995 2700 56065 2746
rect 56111 2700 56181 2746
rect 56227 2700 56297 2746
rect 56343 2700 56413 2746
rect 56459 2700 56529 2746
rect 56575 2700 56594 2746
rect 50826 2630 56594 2700
rect 50826 2584 50845 2630
rect 50891 2584 50961 2630
rect 51007 2584 51077 2630
rect 51123 2584 51193 2630
rect 51239 2584 51309 2630
rect 51355 2584 51425 2630
rect 51471 2584 51541 2630
rect 51587 2584 51657 2630
rect 51703 2584 51773 2630
rect 51819 2584 51889 2630
rect 51935 2584 52005 2630
rect 52051 2584 52121 2630
rect 52167 2584 52237 2630
rect 52283 2584 52353 2630
rect 52399 2584 52469 2630
rect 52515 2584 52585 2630
rect 52631 2584 52701 2630
rect 52747 2584 52817 2630
rect 52863 2584 52933 2630
rect 52979 2584 53049 2630
rect 53095 2584 53165 2630
rect 53211 2584 53281 2630
rect 53327 2584 53397 2630
rect 53443 2584 53513 2630
rect 53559 2584 53629 2630
rect 53675 2584 53745 2630
rect 53791 2584 53861 2630
rect 53907 2584 53977 2630
rect 54023 2584 54093 2630
rect 54139 2584 54209 2630
rect 54255 2584 54325 2630
rect 54371 2584 54441 2630
rect 54487 2584 54557 2630
rect 54603 2584 54673 2630
rect 54719 2584 54789 2630
rect 54835 2584 54905 2630
rect 54951 2584 55021 2630
rect 55067 2584 55137 2630
rect 55183 2584 55253 2630
rect 55299 2584 55369 2630
rect 55415 2584 55485 2630
rect 55531 2584 55601 2630
rect 55647 2584 55717 2630
rect 55763 2584 55833 2630
rect 55879 2584 55949 2630
rect 55995 2584 56065 2630
rect 56111 2584 56181 2630
rect 56227 2584 56297 2630
rect 56343 2584 56413 2630
rect 56459 2584 56529 2630
rect 56575 2584 56594 2630
rect 50826 2514 56594 2584
rect 50826 2468 50845 2514
rect 50891 2468 50961 2514
rect 51007 2468 51077 2514
rect 51123 2468 51193 2514
rect 51239 2468 51309 2514
rect 51355 2468 51425 2514
rect 51471 2468 51541 2514
rect 51587 2468 51657 2514
rect 51703 2468 51773 2514
rect 51819 2468 51889 2514
rect 51935 2468 52005 2514
rect 52051 2468 52121 2514
rect 52167 2468 52237 2514
rect 52283 2468 52353 2514
rect 52399 2468 52469 2514
rect 52515 2468 52585 2514
rect 52631 2468 52701 2514
rect 52747 2468 52817 2514
rect 52863 2468 52933 2514
rect 52979 2468 53049 2514
rect 53095 2468 53165 2514
rect 53211 2468 53281 2514
rect 53327 2468 53397 2514
rect 53443 2468 53513 2514
rect 53559 2468 53629 2514
rect 53675 2468 53745 2514
rect 53791 2468 53861 2514
rect 53907 2468 53977 2514
rect 54023 2468 54093 2514
rect 54139 2468 54209 2514
rect 54255 2468 54325 2514
rect 54371 2468 54441 2514
rect 54487 2468 54557 2514
rect 54603 2468 54673 2514
rect 54719 2468 54789 2514
rect 54835 2468 54905 2514
rect 54951 2468 55021 2514
rect 55067 2468 55137 2514
rect 55183 2468 55253 2514
rect 55299 2468 55369 2514
rect 55415 2468 55485 2514
rect 55531 2468 55601 2514
rect 55647 2468 55717 2514
rect 55763 2468 55833 2514
rect 55879 2468 55949 2514
rect 55995 2468 56065 2514
rect 56111 2468 56181 2514
rect 56227 2468 56297 2514
rect 56343 2468 56413 2514
rect 56459 2468 56529 2514
rect 56575 2468 56594 2514
rect 50826 2398 56594 2468
rect 50826 2352 50845 2398
rect 50891 2352 50961 2398
rect 51007 2352 51077 2398
rect 51123 2352 51193 2398
rect 51239 2352 51309 2398
rect 51355 2352 51425 2398
rect 51471 2352 51541 2398
rect 51587 2352 51657 2398
rect 51703 2352 51773 2398
rect 51819 2352 51889 2398
rect 51935 2352 52005 2398
rect 52051 2352 52121 2398
rect 52167 2352 52237 2398
rect 52283 2352 52353 2398
rect 52399 2352 52469 2398
rect 52515 2352 52585 2398
rect 52631 2352 52701 2398
rect 52747 2352 52817 2398
rect 52863 2352 52933 2398
rect 52979 2352 53049 2398
rect 53095 2352 53165 2398
rect 53211 2352 53281 2398
rect 53327 2352 53397 2398
rect 53443 2352 53513 2398
rect 53559 2352 53629 2398
rect 53675 2352 53745 2398
rect 53791 2352 53861 2398
rect 53907 2352 53977 2398
rect 54023 2352 54093 2398
rect 54139 2352 54209 2398
rect 54255 2352 54325 2398
rect 54371 2352 54441 2398
rect 54487 2352 54557 2398
rect 54603 2352 54673 2398
rect 54719 2352 54789 2398
rect 54835 2352 54905 2398
rect 54951 2352 55021 2398
rect 55067 2352 55137 2398
rect 55183 2352 55253 2398
rect 55299 2352 55369 2398
rect 55415 2352 55485 2398
rect 55531 2352 55601 2398
rect 55647 2352 55717 2398
rect 55763 2352 55833 2398
rect 55879 2352 55949 2398
rect 55995 2352 56065 2398
rect 56111 2352 56181 2398
rect 56227 2352 56297 2398
rect 56343 2352 56413 2398
rect 56459 2352 56529 2398
rect 56575 2352 56594 2398
rect 50826 2282 56594 2352
rect 50826 2236 50845 2282
rect 50891 2236 50961 2282
rect 51007 2236 51077 2282
rect 51123 2236 51193 2282
rect 51239 2236 51309 2282
rect 51355 2236 51425 2282
rect 51471 2236 51541 2282
rect 51587 2236 51657 2282
rect 51703 2236 51773 2282
rect 51819 2236 51889 2282
rect 51935 2236 52005 2282
rect 52051 2236 52121 2282
rect 52167 2236 52237 2282
rect 52283 2236 52353 2282
rect 52399 2236 52469 2282
rect 52515 2236 52585 2282
rect 52631 2236 52701 2282
rect 52747 2236 52817 2282
rect 52863 2236 52933 2282
rect 52979 2236 53049 2282
rect 53095 2236 53165 2282
rect 53211 2236 53281 2282
rect 53327 2236 53397 2282
rect 53443 2236 53513 2282
rect 53559 2236 53629 2282
rect 53675 2236 53745 2282
rect 53791 2236 53861 2282
rect 53907 2236 53977 2282
rect 54023 2236 54093 2282
rect 54139 2236 54209 2282
rect 54255 2236 54325 2282
rect 54371 2236 54441 2282
rect 54487 2236 54557 2282
rect 54603 2236 54673 2282
rect 54719 2236 54789 2282
rect 54835 2236 54905 2282
rect 54951 2236 55021 2282
rect 55067 2236 55137 2282
rect 55183 2236 55253 2282
rect 55299 2236 55369 2282
rect 55415 2236 55485 2282
rect 55531 2236 55601 2282
rect 55647 2236 55717 2282
rect 55763 2236 55833 2282
rect 55879 2236 55949 2282
rect 55995 2236 56065 2282
rect 56111 2236 56181 2282
rect 56227 2236 56297 2282
rect 56343 2236 56413 2282
rect 56459 2236 56529 2282
rect 56575 2236 56594 2282
rect 50826 2166 56594 2236
rect 50826 2120 50845 2166
rect 50891 2120 50961 2166
rect 51007 2120 51077 2166
rect 51123 2120 51193 2166
rect 51239 2120 51309 2166
rect 51355 2120 51425 2166
rect 51471 2120 51541 2166
rect 51587 2120 51657 2166
rect 51703 2120 51773 2166
rect 51819 2120 51889 2166
rect 51935 2120 52005 2166
rect 52051 2120 52121 2166
rect 52167 2120 52237 2166
rect 52283 2120 52353 2166
rect 52399 2120 52469 2166
rect 52515 2120 52585 2166
rect 52631 2120 52701 2166
rect 52747 2120 52817 2166
rect 52863 2120 52933 2166
rect 52979 2120 53049 2166
rect 53095 2120 53165 2166
rect 53211 2120 53281 2166
rect 53327 2120 53397 2166
rect 53443 2120 53513 2166
rect 53559 2120 53629 2166
rect 53675 2120 53745 2166
rect 53791 2120 53861 2166
rect 53907 2120 53977 2166
rect 54023 2120 54093 2166
rect 54139 2120 54209 2166
rect 54255 2120 54325 2166
rect 54371 2120 54441 2166
rect 54487 2120 54557 2166
rect 54603 2120 54673 2166
rect 54719 2120 54789 2166
rect 54835 2120 54905 2166
rect 54951 2120 55021 2166
rect 55067 2120 55137 2166
rect 55183 2120 55253 2166
rect 55299 2120 55369 2166
rect 55415 2120 55485 2166
rect 55531 2120 55601 2166
rect 55647 2120 55717 2166
rect 55763 2120 55833 2166
rect 55879 2120 55949 2166
rect 55995 2120 56065 2166
rect 56111 2120 56181 2166
rect 56227 2120 56297 2166
rect 56343 2120 56413 2166
rect 56459 2120 56529 2166
rect 56575 2120 56594 2166
rect 50826 2050 56594 2120
rect 50826 2004 50845 2050
rect 50891 2004 50961 2050
rect 51007 2004 51077 2050
rect 51123 2004 51193 2050
rect 51239 2004 51309 2050
rect 51355 2004 51425 2050
rect 51471 2004 51541 2050
rect 51587 2004 51657 2050
rect 51703 2004 51773 2050
rect 51819 2004 51889 2050
rect 51935 2004 52005 2050
rect 52051 2004 52121 2050
rect 52167 2004 52237 2050
rect 52283 2004 52353 2050
rect 52399 2004 52469 2050
rect 52515 2004 52585 2050
rect 52631 2004 52701 2050
rect 52747 2004 52817 2050
rect 52863 2004 52933 2050
rect 52979 2004 53049 2050
rect 53095 2004 53165 2050
rect 53211 2004 53281 2050
rect 53327 2004 53397 2050
rect 53443 2004 53513 2050
rect 53559 2004 53629 2050
rect 53675 2004 53745 2050
rect 53791 2004 53861 2050
rect 53907 2004 53977 2050
rect 54023 2004 54093 2050
rect 54139 2004 54209 2050
rect 54255 2004 54325 2050
rect 54371 2004 54441 2050
rect 54487 2004 54557 2050
rect 54603 2004 54673 2050
rect 54719 2004 54789 2050
rect 54835 2004 54905 2050
rect 54951 2004 55021 2050
rect 55067 2004 55137 2050
rect 55183 2004 55253 2050
rect 55299 2004 55369 2050
rect 55415 2004 55485 2050
rect 55531 2004 55601 2050
rect 55647 2004 55717 2050
rect 55763 2004 55833 2050
rect 55879 2004 55949 2050
rect 55995 2004 56065 2050
rect 56111 2004 56181 2050
rect 56227 2004 56297 2050
rect 56343 2004 56413 2050
rect 56459 2004 56529 2050
rect 56575 2004 56594 2050
rect 50826 1934 56594 2004
rect 50826 1888 50845 1934
rect 50891 1888 50961 1934
rect 51007 1888 51077 1934
rect 51123 1888 51193 1934
rect 51239 1888 51309 1934
rect 51355 1888 51425 1934
rect 51471 1888 51541 1934
rect 51587 1888 51657 1934
rect 51703 1888 51773 1934
rect 51819 1888 51889 1934
rect 51935 1888 52005 1934
rect 52051 1888 52121 1934
rect 52167 1888 52237 1934
rect 52283 1888 52353 1934
rect 52399 1888 52469 1934
rect 52515 1888 52585 1934
rect 52631 1888 52701 1934
rect 52747 1888 52817 1934
rect 52863 1888 52933 1934
rect 52979 1888 53049 1934
rect 53095 1888 53165 1934
rect 53211 1888 53281 1934
rect 53327 1888 53397 1934
rect 53443 1888 53513 1934
rect 53559 1888 53629 1934
rect 53675 1888 53745 1934
rect 53791 1888 53861 1934
rect 53907 1888 53977 1934
rect 54023 1888 54093 1934
rect 54139 1888 54209 1934
rect 54255 1888 54325 1934
rect 54371 1888 54441 1934
rect 54487 1888 54557 1934
rect 54603 1888 54673 1934
rect 54719 1888 54789 1934
rect 54835 1888 54905 1934
rect 54951 1888 55021 1934
rect 55067 1888 55137 1934
rect 55183 1888 55253 1934
rect 55299 1888 55369 1934
rect 55415 1888 55485 1934
rect 55531 1888 55601 1934
rect 55647 1888 55717 1934
rect 55763 1888 55833 1934
rect 55879 1888 55949 1934
rect 55995 1888 56065 1934
rect 56111 1888 56181 1934
rect 56227 1888 56297 1934
rect 56343 1888 56413 1934
rect 56459 1888 56529 1934
rect 56575 1888 56594 1934
rect 50826 1818 56594 1888
rect 50826 1772 50845 1818
rect 50891 1772 50961 1818
rect 51007 1772 51077 1818
rect 51123 1772 51193 1818
rect 51239 1772 51309 1818
rect 51355 1772 51425 1818
rect 51471 1772 51541 1818
rect 51587 1772 51657 1818
rect 51703 1772 51773 1818
rect 51819 1772 51889 1818
rect 51935 1772 52005 1818
rect 52051 1772 52121 1818
rect 52167 1772 52237 1818
rect 52283 1772 52353 1818
rect 52399 1772 52469 1818
rect 52515 1772 52585 1818
rect 52631 1772 52701 1818
rect 52747 1772 52817 1818
rect 52863 1772 52933 1818
rect 52979 1772 53049 1818
rect 53095 1772 53165 1818
rect 53211 1772 53281 1818
rect 53327 1772 53397 1818
rect 53443 1772 53513 1818
rect 53559 1772 53629 1818
rect 53675 1772 53745 1818
rect 53791 1772 53861 1818
rect 53907 1772 53977 1818
rect 54023 1772 54093 1818
rect 54139 1772 54209 1818
rect 54255 1772 54325 1818
rect 54371 1772 54441 1818
rect 54487 1772 54557 1818
rect 54603 1772 54673 1818
rect 54719 1772 54789 1818
rect 54835 1772 54905 1818
rect 54951 1772 55021 1818
rect 55067 1772 55137 1818
rect 55183 1772 55253 1818
rect 55299 1772 55369 1818
rect 55415 1772 55485 1818
rect 55531 1772 55601 1818
rect 55647 1772 55717 1818
rect 55763 1772 55833 1818
rect 55879 1772 55949 1818
rect 55995 1772 56065 1818
rect 56111 1772 56181 1818
rect 56227 1772 56297 1818
rect 56343 1772 56413 1818
rect 56459 1772 56529 1818
rect 56575 1772 56594 1818
rect 50826 1702 56594 1772
rect 50826 1656 50845 1702
rect 50891 1656 50961 1702
rect 51007 1656 51077 1702
rect 51123 1656 51193 1702
rect 51239 1656 51309 1702
rect 51355 1656 51425 1702
rect 51471 1656 51541 1702
rect 51587 1656 51657 1702
rect 51703 1656 51773 1702
rect 51819 1656 51889 1702
rect 51935 1656 52005 1702
rect 52051 1656 52121 1702
rect 52167 1656 52237 1702
rect 52283 1656 52353 1702
rect 52399 1656 52469 1702
rect 52515 1656 52585 1702
rect 52631 1656 52701 1702
rect 52747 1656 52817 1702
rect 52863 1656 52933 1702
rect 52979 1656 53049 1702
rect 53095 1656 53165 1702
rect 53211 1656 53281 1702
rect 53327 1656 53397 1702
rect 53443 1656 53513 1702
rect 53559 1656 53629 1702
rect 53675 1656 53745 1702
rect 53791 1656 53861 1702
rect 53907 1656 53977 1702
rect 54023 1656 54093 1702
rect 54139 1656 54209 1702
rect 54255 1656 54325 1702
rect 54371 1656 54441 1702
rect 54487 1656 54557 1702
rect 54603 1656 54673 1702
rect 54719 1656 54789 1702
rect 54835 1656 54905 1702
rect 54951 1656 55021 1702
rect 55067 1656 55137 1702
rect 55183 1656 55253 1702
rect 55299 1656 55369 1702
rect 55415 1656 55485 1702
rect 55531 1656 55601 1702
rect 55647 1656 55717 1702
rect 55763 1656 55833 1702
rect 55879 1656 55949 1702
rect 55995 1656 56065 1702
rect 56111 1656 56181 1702
rect 56227 1656 56297 1702
rect 56343 1656 56413 1702
rect 56459 1656 56529 1702
rect 56575 1656 56594 1702
rect 50826 1637 56594 1656
rect 27379 1034 27763 1117
rect 57287 1117 57306 34155
rect 57652 1117 57671 96163
rect 57287 1034 57671 1117
rect 85714 96163 86098 96246
rect 85714 1117 85733 96163
rect 86079 1117 86098 96163
rect 85714 1034 86098 1117
rect 352 1015 86098 1034
rect 352 969 371 1015
rect 417 969 495 1015
rect 541 969 619 1015
rect 665 969 743 1015
rect 789 969 867 1015
rect 913 969 991 1015
rect 1037 969 1115 1015
rect 1161 969 1239 1015
rect 1285 969 1363 1015
rect 1409 969 1487 1015
rect 1533 969 1611 1015
rect 1657 969 1735 1015
rect 1781 969 1859 1015
rect 1905 969 1983 1015
rect 2029 969 2107 1015
rect 2153 969 2231 1015
rect 2277 969 2355 1015
rect 2401 969 2479 1015
rect 2525 969 2603 1015
rect 2649 969 2727 1015
rect 2773 969 2851 1015
rect 2897 969 2975 1015
rect 3021 969 3099 1015
rect 3145 969 3223 1015
rect 3269 969 3347 1015
rect 3393 969 3471 1015
rect 3517 969 3595 1015
rect 3641 969 3719 1015
rect 3765 969 3843 1015
rect 3889 969 3967 1015
rect 4013 969 4091 1015
rect 4137 969 4215 1015
rect 4261 969 4339 1015
rect 4385 969 4463 1015
rect 4509 969 4587 1015
rect 4633 969 4711 1015
rect 4757 969 4835 1015
rect 4881 969 4959 1015
rect 5005 969 5083 1015
rect 5129 969 5207 1015
rect 5253 969 5331 1015
rect 5377 969 5455 1015
rect 5501 969 5579 1015
rect 5625 969 5703 1015
rect 5749 969 5827 1015
rect 5873 969 5951 1015
rect 5997 969 6075 1015
rect 6121 969 6199 1015
rect 6245 969 6323 1015
rect 6369 969 6447 1015
rect 6493 969 6571 1015
rect 6617 969 6695 1015
rect 6741 969 6819 1015
rect 6865 969 6943 1015
rect 6989 969 7067 1015
rect 7113 969 7191 1015
rect 7237 969 7315 1015
rect 7361 969 7439 1015
rect 7485 969 7563 1015
rect 7609 969 7687 1015
rect 7733 969 7811 1015
rect 7857 969 7935 1015
rect 7981 969 8059 1015
rect 8105 969 8183 1015
rect 8229 969 8307 1015
rect 8353 969 8431 1015
rect 8477 969 8555 1015
rect 8601 969 8679 1015
rect 8725 969 8803 1015
rect 8849 969 8927 1015
rect 8973 969 9051 1015
rect 9097 969 9175 1015
rect 9221 969 9299 1015
rect 9345 969 9423 1015
rect 9469 969 9547 1015
rect 9593 969 9671 1015
rect 9717 969 9795 1015
rect 9841 969 9919 1015
rect 9965 969 10043 1015
rect 10089 969 10167 1015
rect 10213 969 10291 1015
rect 10337 969 10415 1015
rect 10461 969 10539 1015
rect 10585 969 10663 1015
rect 10709 969 10787 1015
rect 10833 969 10911 1015
rect 10957 969 11035 1015
rect 11081 969 11159 1015
rect 11205 969 11283 1015
rect 11329 969 11407 1015
rect 11453 969 11531 1015
rect 11577 969 11655 1015
rect 11701 969 11779 1015
rect 11825 969 11903 1015
rect 11949 969 12027 1015
rect 12073 969 12151 1015
rect 12197 969 12275 1015
rect 12321 969 12399 1015
rect 12445 969 12523 1015
rect 12569 969 12647 1015
rect 12693 969 12771 1015
rect 12817 969 12895 1015
rect 12941 969 13019 1015
rect 13065 969 13143 1015
rect 13189 969 13267 1015
rect 13313 969 13391 1015
rect 13437 969 13515 1015
rect 13561 969 13639 1015
rect 13685 969 13763 1015
rect 13809 969 13887 1015
rect 13933 969 14011 1015
rect 14057 969 14135 1015
rect 14181 969 14259 1015
rect 14305 969 14383 1015
rect 14429 969 14507 1015
rect 14553 969 14631 1015
rect 14677 969 14755 1015
rect 14801 969 14879 1015
rect 14925 969 15003 1015
rect 15049 969 15127 1015
rect 15173 969 15251 1015
rect 15297 969 15375 1015
rect 15421 969 15499 1015
rect 15545 969 15623 1015
rect 15669 969 15747 1015
rect 15793 969 15871 1015
rect 15917 969 15995 1015
rect 16041 969 16119 1015
rect 16165 969 16243 1015
rect 16289 969 16367 1015
rect 16413 969 16491 1015
rect 16537 969 16615 1015
rect 16661 969 16739 1015
rect 16785 969 16863 1015
rect 16909 969 16987 1015
rect 17033 969 17111 1015
rect 17157 969 17235 1015
rect 17281 969 17359 1015
rect 17405 969 17483 1015
rect 17529 969 17607 1015
rect 17653 969 17731 1015
rect 17777 969 17855 1015
rect 17901 969 17979 1015
rect 18025 969 18103 1015
rect 18149 969 18227 1015
rect 18273 969 18351 1015
rect 18397 969 18475 1015
rect 18521 969 18599 1015
rect 18645 969 18723 1015
rect 18769 969 18847 1015
rect 18893 969 18971 1015
rect 19017 969 19095 1015
rect 19141 969 19219 1015
rect 19265 969 19343 1015
rect 19389 969 19467 1015
rect 19513 969 19591 1015
rect 19637 969 19715 1015
rect 19761 969 19839 1015
rect 19885 969 19963 1015
rect 20009 969 20087 1015
rect 20133 969 20211 1015
rect 20257 969 20335 1015
rect 20381 969 20459 1015
rect 20505 969 20583 1015
rect 20629 969 20707 1015
rect 20753 969 20831 1015
rect 20877 969 20955 1015
rect 21001 969 21079 1015
rect 21125 969 21203 1015
rect 21249 969 21327 1015
rect 21373 969 21451 1015
rect 21497 969 21575 1015
rect 21621 969 21699 1015
rect 21745 969 21823 1015
rect 21869 969 21947 1015
rect 21993 969 22071 1015
rect 22117 969 22195 1015
rect 22241 969 22319 1015
rect 22365 969 22443 1015
rect 22489 969 22567 1015
rect 22613 969 22691 1015
rect 22737 969 22815 1015
rect 22861 969 22939 1015
rect 22985 969 23063 1015
rect 23109 969 23187 1015
rect 23233 969 23311 1015
rect 23357 969 23435 1015
rect 23481 969 23559 1015
rect 23605 969 23683 1015
rect 23729 969 23807 1015
rect 23853 969 23931 1015
rect 23977 969 24055 1015
rect 24101 969 24179 1015
rect 24225 969 24303 1015
rect 24349 969 24427 1015
rect 24473 969 24551 1015
rect 24597 969 24675 1015
rect 24721 969 24799 1015
rect 24845 969 24923 1015
rect 24969 969 25047 1015
rect 25093 969 25171 1015
rect 25217 969 25295 1015
rect 25341 969 25419 1015
rect 25465 969 25543 1015
rect 25589 969 25667 1015
rect 25713 969 25791 1015
rect 25837 969 25915 1015
rect 25961 969 26039 1015
rect 26085 969 26163 1015
rect 26209 969 26287 1015
rect 26333 969 26411 1015
rect 26457 969 26535 1015
rect 26581 969 26659 1015
rect 26705 969 26783 1015
rect 26829 969 26907 1015
rect 26953 969 27031 1015
rect 27077 969 27155 1015
rect 27201 969 27279 1015
rect 27325 969 27403 1015
rect 27449 969 27527 1015
rect 27573 969 27651 1015
rect 27697 969 27775 1015
rect 27821 969 27899 1015
rect 27945 969 28023 1015
rect 28069 969 28147 1015
rect 28193 969 28271 1015
rect 28317 969 28395 1015
rect 28441 969 28519 1015
rect 28565 969 28643 1015
rect 28689 969 28767 1015
rect 28813 969 28891 1015
rect 28937 969 29015 1015
rect 29061 969 29139 1015
rect 29185 969 29263 1015
rect 29309 969 29387 1015
rect 29433 969 29511 1015
rect 29557 969 29635 1015
rect 29681 969 29759 1015
rect 29805 969 29883 1015
rect 29929 969 30007 1015
rect 30053 969 30131 1015
rect 30177 969 30255 1015
rect 30301 969 30379 1015
rect 30425 969 30503 1015
rect 30549 969 30627 1015
rect 30673 969 30751 1015
rect 30797 969 30875 1015
rect 30921 969 30999 1015
rect 31045 969 31123 1015
rect 31169 969 31247 1015
rect 31293 969 31371 1015
rect 31417 969 31495 1015
rect 31541 969 31619 1015
rect 31665 969 31743 1015
rect 31789 969 31867 1015
rect 31913 969 31991 1015
rect 32037 969 32115 1015
rect 32161 969 32239 1015
rect 32285 969 32363 1015
rect 32409 969 32487 1015
rect 32533 969 32611 1015
rect 32657 969 32735 1015
rect 32781 969 32859 1015
rect 32905 969 32983 1015
rect 33029 969 33107 1015
rect 33153 969 33231 1015
rect 33277 969 33355 1015
rect 33401 969 33479 1015
rect 33525 969 33603 1015
rect 33649 969 33727 1015
rect 33773 969 33851 1015
rect 33897 969 33975 1015
rect 34021 969 34099 1015
rect 34145 969 34223 1015
rect 34269 969 34347 1015
rect 34393 969 34471 1015
rect 34517 969 34595 1015
rect 34641 969 34719 1015
rect 34765 969 34843 1015
rect 34889 969 34967 1015
rect 35013 969 35091 1015
rect 35137 969 35215 1015
rect 35261 969 35339 1015
rect 35385 969 35463 1015
rect 35509 969 35587 1015
rect 35633 969 35711 1015
rect 35757 969 35835 1015
rect 35881 969 35959 1015
rect 36005 969 36083 1015
rect 36129 969 36207 1015
rect 36253 969 36331 1015
rect 36377 969 36455 1015
rect 36501 969 36579 1015
rect 36625 969 36703 1015
rect 36749 969 36827 1015
rect 36873 969 36951 1015
rect 36997 969 37075 1015
rect 37121 969 37199 1015
rect 37245 969 37323 1015
rect 37369 969 37447 1015
rect 37493 969 37571 1015
rect 37617 969 37695 1015
rect 37741 969 37819 1015
rect 37865 969 37943 1015
rect 37989 969 38067 1015
rect 38113 969 38191 1015
rect 38237 969 38315 1015
rect 38361 969 38439 1015
rect 38485 969 38563 1015
rect 38609 969 38687 1015
rect 38733 969 38811 1015
rect 38857 969 38935 1015
rect 38981 969 39059 1015
rect 39105 969 39183 1015
rect 39229 969 39307 1015
rect 39353 969 39431 1015
rect 39477 969 39555 1015
rect 39601 969 39679 1015
rect 39725 969 39803 1015
rect 39849 969 39927 1015
rect 39973 969 40051 1015
rect 40097 969 40175 1015
rect 40221 969 40299 1015
rect 40345 969 40423 1015
rect 40469 969 40547 1015
rect 40593 969 40671 1015
rect 40717 969 40795 1015
rect 40841 969 40919 1015
rect 40965 969 41043 1015
rect 41089 969 41167 1015
rect 41213 969 41291 1015
rect 41337 969 41415 1015
rect 41461 969 41539 1015
rect 41585 969 41663 1015
rect 41709 969 41787 1015
rect 41833 969 41911 1015
rect 41957 969 42035 1015
rect 42081 969 42159 1015
rect 42205 969 42283 1015
rect 42329 969 42407 1015
rect 42453 969 42531 1015
rect 42577 969 42655 1015
rect 42701 969 42779 1015
rect 42825 969 42903 1015
rect 42949 969 43027 1015
rect 43073 969 43151 1015
rect 43197 969 43275 1015
rect 43321 969 43399 1015
rect 43445 969 43523 1015
rect 43569 969 43647 1015
rect 43693 969 43771 1015
rect 43817 969 43895 1015
rect 43941 969 44019 1015
rect 44065 969 44143 1015
rect 44189 969 44267 1015
rect 44313 969 44391 1015
rect 44437 969 44515 1015
rect 44561 969 44639 1015
rect 44685 969 44763 1015
rect 44809 969 44887 1015
rect 44933 969 45011 1015
rect 45057 969 45135 1015
rect 45181 969 45259 1015
rect 45305 969 45383 1015
rect 45429 969 45507 1015
rect 45553 969 45631 1015
rect 45677 969 45755 1015
rect 45801 969 45879 1015
rect 45925 969 46003 1015
rect 46049 969 46127 1015
rect 46173 969 46251 1015
rect 46297 969 46375 1015
rect 46421 969 46499 1015
rect 46545 969 46623 1015
rect 46669 969 46747 1015
rect 46793 969 46871 1015
rect 46917 969 46995 1015
rect 47041 969 47119 1015
rect 47165 969 47243 1015
rect 47289 969 47367 1015
rect 47413 969 47491 1015
rect 47537 969 47615 1015
rect 47661 969 47739 1015
rect 47785 969 47863 1015
rect 47909 969 47987 1015
rect 48033 969 48111 1015
rect 48157 969 48235 1015
rect 48281 969 48359 1015
rect 48405 969 48483 1015
rect 48529 969 48607 1015
rect 48653 969 48731 1015
rect 48777 969 48855 1015
rect 48901 969 48979 1015
rect 49025 969 49103 1015
rect 49149 969 49227 1015
rect 49273 969 49351 1015
rect 49397 969 49475 1015
rect 49521 969 49599 1015
rect 49645 969 49723 1015
rect 49769 969 49847 1015
rect 49893 969 49971 1015
rect 50017 969 50095 1015
rect 50141 969 50219 1015
rect 50265 969 50343 1015
rect 50389 969 50467 1015
rect 50513 969 50591 1015
rect 50637 969 50715 1015
rect 50761 969 50839 1015
rect 50885 969 50963 1015
rect 51009 969 51087 1015
rect 51133 969 51211 1015
rect 51257 969 51335 1015
rect 51381 969 51459 1015
rect 51505 969 51583 1015
rect 51629 969 51707 1015
rect 51753 969 51831 1015
rect 51877 969 51955 1015
rect 52001 969 52079 1015
rect 52125 969 52203 1015
rect 52249 969 52327 1015
rect 52373 969 52451 1015
rect 52497 969 52575 1015
rect 52621 969 52699 1015
rect 52745 969 52823 1015
rect 52869 969 52947 1015
rect 52993 969 53071 1015
rect 53117 969 53195 1015
rect 53241 969 53319 1015
rect 53365 969 53443 1015
rect 53489 969 53567 1015
rect 53613 969 53691 1015
rect 53737 969 53815 1015
rect 53861 969 53939 1015
rect 53985 969 54063 1015
rect 54109 969 54187 1015
rect 54233 969 54311 1015
rect 54357 969 54435 1015
rect 54481 969 54559 1015
rect 54605 969 54683 1015
rect 54729 969 54807 1015
rect 54853 969 54931 1015
rect 54977 969 55055 1015
rect 55101 969 55179 1015
rect 55225 969 55303 1015
rect 55349 969 55427 1015
rect 55473 969 55551 1015
rect 55597 969 55675 1015
rect 55721 969 55799 1015
rect 55845 969 55923 1015
rect 55969 969 56047 1015
rect 56093 969 56171 1015
rect 56217 969 56295 1015
rect 56341 969 56419 1015
rect 56465 969 56543 1015
rect 56589 969 56667 1015
rect 56713 969 56791 1015
rect 56837 969 56915 1015
rect 56961 969 57039 1015
rect 57085 969 57163 1015
rect 57209 969 57287 1015
rect 57333 969 57411 1015
rect 57457 969 57535 1015
rect 57581 969 57659 1015
rect 57705 969 57783 1015
rect 57829 969 57907 1015
rect 57953 969 58031 1015
rect 58077 969 58155 1015
rect 58201 969 58279 1015
rect 58325 969 58403 1015
rect 58449 969 58527 1015
rect 58573 969 58651 1015
rect 58697 969 58775 1015
rect 58821 969 58899 1015
rect 58945 969 59023 1015
rect 59069 969 59147 1015
rect 59193 969 59271 1015
rect 59317 969 59395 1015
rect 59441 969 59519 1015
rect 59565 969 59643 1015
rect 59689 969 59767 1015
rect 59813 969 59891 1015
rect 59937 969 60015 1015
rect 60061 969 60139 1015
rect 60185 969 60263 1015
rect 60309 969 60387 1015
rect 60433 969 60511 1015
rect 60557 969 60635 1015
rect 60681 969 60759 1015
rect 60805 969 60883 1015
rect 60929 969 61007 1015
rect 61053 969 61131 1015
rect 61177 969 61255 1015
rect 61301 969 61379 1015
rect 61425 969 61503 1015
rect 61549 969 61627 1015
rect 61673 969 61751 1015
rect 61797 969 61875 1015
rect 61921 969 61999 1015
rect 62045 969 62123 1015
rect 62169 969 62247 1015
rect 62293 969 62371 1015
rect 62417 969 62495 1015
rect 62541 969 62619 1015
rect 62665 969 62743 1015
rect 62789 969 62867 1015
rect 62913 969 62991 1015
rect 63037 969 63115 1015
rect 63161 969 63239 1015
rect 63285 969 63363 1015
rect 63409 969 63487 1015
rect 63533 969 63611 1015
rect 63657 969 63735 1015
rect 63781 969 63859 1015
rect 63905 969 63983 1015
rect 64029 969 64107 1015
rect 64153 969 64231 1015
rect 64277 969 64355 1015
rect 64401 969 64479 1015
rect 64525 969 64603 1015
rect 64649 969 64727 1015
rect 64773 969 64851 1015
rect 64897 969 64975 1015
rect 65021 969 65099 1015
rect 65145 969 65223 1015
rect 65269 969 65347 1015
rect 65393 969 65471 1015
rect 65517 969 65595 1015
rect 65641 969 65719 1015
rect 65765 969 65843 1015
rect 65889 969 65967 1015
rect 66013 969 66091 1015
rect 66137 969 66215 1015
rect 66261 969 66339 1015
rect 66385 969 66463 1015
rect 66509 969 66587 1015
rect 66633 969 66711 1015
rect 66757 969 66835 1015
rect 66881 969 66959 1015
rect 67005 969 67083 1015
rect 67129 969 67207 1015
rect 67253 969 67331 1015
rect 67377 969 67455 1015
rect 67501 969 67579 1015
rect 67625 969 67703 1015
rect 67749 969 67827 1015
rect 67873 969 67951 1015
rect 67997 969 68075 1015
rect 68121 969 68199 1015
rect 68245 969 68323 1015
rect 68369 969 68447 1015
rect 68493 969 68571 1015
rect 68617 969 68695 1015
rect 68741 969 68819 1015
rect 68865 969 68943 1015
rect 68989 969 69067 1015
rect 69113 969 69191 1015
rect 69237 969 69315 1015
rect 69361 969 69439 1015
rect 69485 969 69563 1015
rect 69609 969 69687 1015
rect 69733 969 69811 1015
rect 69857 969 69935 1015
rect 69981 969 70059 1015
rect 70105 969 70183 1015
rect 70229 969 70307 1015
rect 70353 969 70431 1015
rect 70477 969 70555 1015
rect 70601 969 70679 1015
rect 70725 969 70803 1015
rect 70849 969 70927 1015
rect 70973 969 71051 1015
rect 71097 969 71175 1015
rect 71221 969 71299 1015
rect 71345 969 71423 1015
rect 71469 969 71547 1015
rect 71593 969 71671 1015
rect 71717 969 71795 1015
rect 71841 969 71919 1015
rect 71965 969 72043 1015
rect 72089 969 72167 1015
rect 72213 969 72291 1015
rect 72337 969 72415 1015
rect 72461 969 72539 1015
rect 72585 969 72663 1015
rect 72709 969 72787 1015
rect 72833 969 72911 1015
rect 72957 969 73035 1015
rect 73081 969 73159 1015
rect 73205 969 73283 1015
rect 73329 969 73407 1015
rect 73453 969 73531 1015
rect 73577 969 73655 1015
rect 73701 969 73779 1015
rect 73825 969 73903 1015
rect 73949 969 74027 1015
rect 74073 969 74151 1015
rect 74197 969 74275 1015
rect 74321 969 74399 1015
rect 74445 969 74523 1015
rect 74569 969 74647 1015
rect 74693 969 74771 1015
rect 74817 969 74895 1015
rect 74941 969 75019 1015
rect 75065 969 75143 1015
rect 75189 969 75267 1015
rect 75313 969 75391 1015
rect 75437 969 75515 1015
rect 75561 969 75639 1015
rect 75685 969 75763 1015
rect 75809 969 75887 1015
rect 75933 969 76011 1015
rect 76057 969 76135 1015
rect 76181 969 76259 1015
rect 76305 969 76383 1015
rect 76429 969 76507 1015
rect 76553 969 76631 1015
rect 76677 969 76755 1015
rect 76801 969 76879 1015
rect 76925 969 77003 1015
rect 77049 969 77127 1015
rect 77173 969 77251 1015
rect 77297 969 77375 1015
rect 77421 969 77499 1015
rect 77545 969 77623 1015
rect 77669 969 77747 1015
rect 77793 969 77871 1015
rect 77917 969 77995 1015
rect 78041 969 78119 1015
rect 78165 969 78243 1015
rect 78289 969 78367 1015
rect 78413 969 78491 1015
rect 78537 969 78615 1015
rect 78661 969 78739 1015
rect 78785 969 78863 1015
rect 78909 969 78987 1015
rect 79033 969 79111 1015
rect 79157 969 79235 1015
rect 79281 969 79359 1015
rect 79405 969 79483 1015
rect 79529 969 79607 1015
rect 79653 969 79731 1015
rect 79777 969 79855 1015
rect 79901 969 79979 1015
rect 80025 969 80103 1015
rect 80149 969 80227 1015
rect 80273 969 80351 1015
rect 80397 969 80475 1015
rect 80521 969 80599 1015
rect 80645 969 80723 1015
rect 80769 969 80847 1015
rect 80893 969 80971 1015
rect 81017 969 81095 1015
rect 81141 969 81219 1015
rect 81265 969 81343 1015
rect 81389 969 81467 1015
rect 81513 969 81591 1015
rect 81637 969 81715 1015
rect 81761 969 81839 1015
rect 81885 969 81963 1015
rect 82009 969 82087 1015
rect 82133 969 82211 1015
rect 82257 969 82335 1015
rect 82381 969 82459 1015
rect 82505 969 82583 1015
rect 82629 969 82707 1015
rect 82753 969 82831 1015
rect 82877 969 82955 1015
rect 83001 969 83079 1015
rect 83125 969 83203 1015
rect 83249 969 83327 1015
rect 83373 969 83451 1015
rect 83497 969 83575 1015
rect 83621 969 83699 1015
rect 83745 969 83823 1015
rect 83869 969 83947 1015
rect 83993 969 84071 1015
rect 84117 969 84195 1015
rect 84241 969 84319 1015
rect 84365 969 84443 1015
rect 84489 969 84567 1015
rect 84613 969 84691 1015
rect 84737 969 84815 1015
rect 84861 969 84939 1015
rect 84985 969 85063 1015
rect 85109 969 85187 1015
rect 85233 969 85311 1015
rect 85357 969 85435 1015
rect 85481 969 85559 1015
rect 85605 969 85683 1015
rect 85729 969 85807 1015
rect 85853 969 85931 1015
rect 85977 969 86098 1015
rect 352 891 86098 969
rect 352 845 371 891
rect 417 845 495 891
rect 541 845 619 891
rect 665 845 743 891
rect 789 845 867 891
rect 913 845 991 891
rect 1037 845 1115 891
rect 1161 845 1239 891
rect 1285 845 1363 891
rect 1409 845 1487 891
rect 1533 845 1611 891
rect 1657 845 1735 891
rect 1781 845 1859 891
rect 1905 845 1983 891
rect 2029 845 2107 891
rect 2153 845 2231 891
rect 2277 845 2355 891
rect 2401 845 2479 891
rect 2525 845 2603 891
rect 2649 845 2727 891
rect 2773 845 2851 891
rect 2897 845 2975 891
rect 3021 845 3099 891
rect 3145 845 3223 891
rect 3269 845 3347 891
rect 3393 845 3471 891
rect 3517 845 3595 891
rect 3641 845 3719 891
rect 3765 845 3843 891
rect 3889 845 3967 891
rect 4013 845 4091 891
rect 4137 845 4215 891
rect 4261 845 4339 891
rect 4385 845 4463 891
rect 4509 845 4587 891
rect 4633 845 4711 891
rect 4757 845 4835 891
rect 4881 845 4959 891
rect 5005 845 5083 891
rect 5129 845 5207 891
rect 5253 845 5331 891
rect 5377 845 5455 891
rect 5501 845 5579 891
rect 5625 845 5703 891
rect 5749 845 5827 891
rect 5873 845 5951 891
rect 5997 845 6075 891
rect 6121 845 6199 891
rect 6245 845 6323 891
rect 6369 845 6447 891
rect 6493 845 6571 891
rect 6617 845 6695 891
rect 6741 845 6819 891
rect 6865 845 6943 891
rect 6989 845 7067 891
rect 7113 845 7191 891
rect 7237 845 7315 891
rect 7361 845 7439 891
rect 7485 845 7563 891
rect 7609 845 7687 891
rect 7733 845 7811 891
rect 7857 845 7935 891
rect 7981 845 8059 891
rect 8105 845 8183 891
rect 8229 845 8307 891
rect 8353 845 8431 891
rect 8477 845 8555 891
rect 8601 845 8679 891
rect 8725 845 8803 891
rect 8849 845 8927 891
rect 8973 845 9051 891
rect 9097 845 9175 891
rect 9221 845 9299 891
rect 9345 845 9423 891
rect 9469 845 9547 891
rect 9593 845 9671 891
rect 9717 845 9795 891
rect 9841 845 9919 891
rect 9965 845 10043 891
rect 10089 845 10167 891
rect 10213 845 10291 891
rect 10337 845 10415 891
rect 10461 845 10539 891
rect 10585 845 10663 891
rect 10709 845 10787 891
rect 10833 845 10911 891
rect 10957 845 11035 891
rect 11081 845 11159 891
rect 11205 845 11283 891
rect 11329 845 11407 891
rect 11453 845 11531 891
rect 11577 845 11655 891
rect 11701 845 11779 891
rect 11825 845 11903 891
rect 11949 845 12027 891
rect 12073 845 12151 891
rect 12197 845 12275 891
rect 12321 845 12399 891
rect 12445 845 12523 891
rect 12569 845 12647 891
rect 12693 845 12771 891
rect 12817 845 12895 891
rect 12941 845 13019 891
rect 13065 845 13143 891
rect 13189 845 13267 891
rect 13313 845 13391 891
rect 13437 845 13515 891
rect 13561 845 13639 891
rect 13685 845 13763 891
rect 13809 845 13887 891
rect 13933 845 14011 891
rect 14057 845 14135 891
rect 14181 845 14259 891
rect 14305 845 14383 891
rect 14429 845 14507 891
rect 14553 845 14631 891
rect 14677 845 14755 891
rect 14801 845 14879 891
rect 14925 845 15003 891
rect 15049 845 15127 891
rect 15173 845 15251 891
rect 15297 845 15375 891
rect 15421 845 15499 891
rect 15545 845 15623 891
rect 15669 845 15747 891
rect 15793 845 15871 891
rect 15917 845 15995 891
rect 16041 845 16119 891
rect 16165 845 16243 891
rect 16289 845 16367 891
rect 16413 845 16491 891
rect 16537 845 16615 891
rect 16661 845 16739 891
rect 16785 845 16863 891
rect 16909 845 16987 891
rect 17033 845 17111 891
rect 17157 845 17235 891
rect 17281 845 17359 891
rect 17405 845 17483 891
rect 17529 845 17607 891
rect 17653 845 17731 891
rect 17777 845 17855 891
rect 17901 845 17979 891
rect 18025 845 18103 891
rect 18149 845 18227 891
rect 18273 845 18351 891
rect 18397 845 18475 891
rect 18521 845 18599 891
rect 18645 845 18723 891
rect 18769 845 18847 891
rect 18893 845 18971 891
rect 19017 845 19095 891
rect 19141 845 19219 891
rect 19265 845 19343 891
rect 19389 845 19467 891
rect 19513 845 19591 891
rect 19637 845 19715 891
rect 19761 845 19839 891
rect 19885 845 19963 891
rect 20009 845 20087 891
rect 20133 845 20211 891
rect 20257 845 20335 891
rect 20381 845 20459 891
rect 20505 845 20583 891
rect 20629 845 20707 891
rect 20753 845 20831 891
rect 20877 845 20955 891
rect 21001 845 21079 891
rect 21125 845 21203 891
rect 21249 845 21327 891
rect 21373 845 21451 891
rect 21497 845 21575 891
rect 21621 845 21699 891
rect 21745 845 21823 891
rect 21869 845 21947 891
rect 21993 845 22071 891
rect 22117 845 22195 891
rect 22241 845 22319 891
rect 22365 845 22443 891
rect 22489 845 22567 891
rect 22613 845 22691 891
rect 22737 845 22815 891
rect 22861 845 22939 891
rect 22985 845 23063 891
rect 23109 845 23187 891
rect 23233 845 23311 891
rect 23357 845 23435 891
rect 23481 845 23559 891
rect 23605 845 23683 891
rect 23729 845 23807 891
rect 23853 845 23931 891
rect 23977 845 24055 891
rect 24101 845 24179 891
rect 24225 845 24303 891
rect 24349 845 24427 891
rect 24473 845 24551 891
rect 24597 845 24675 891
rect 24721 845 24799 891
rect 24845 845 24923 891
rect 24969 845 25047 891
rect 25093 845 25171 891
rect 25217 845 25295 891
rect 25341 845 25419 891
rect 25465 845 25543 891
rect 25589 845 25667 891
rect 25713 845 25791 891
rect 25837 845 25915 891
rect 25961 845 26039 891
rect 26085 845 26163 891
rect 26209 845 26287 891
rect 26333 845 26411 891
rect 26457 845 26535 891
rect 26581 845 26659 891
rect 26705 845 26783 891
rect 26829 845 26907 891
rect 26953 845 27031 891
rect 27077 845 27155 891
rect 27201 845 27279 891
rect 27325 845 27403 891
rect 27449 845 27527 891
rect 27573 845 27651 891
rect 27697 845 27775 891
rect 27821 845 27899 891
rect 27945 845 28023 891
rect 28069 845 28147 891
rect 28193 845 28271 891
rect 28317 845 28395 891
rect 28441 845 28519 891
rect 28565 845 28643 891
rect 28689 845 28767 891
rect 28813 845 28891 891
rect 28937 845 29015 891
rect 29061 845 29139 891
rect 29185 845 29263 891
rect 29309 845 29387 891
rect 29433 845 29511 891
rect 29557 845 29635 891
rect 29681 845 29759 891
rect 29805 845 29883 891
rect 29929 845 30007 891
rect 30053 845 30131 891
rect 30177 845 30255 891
rect 30301 845 30379 891
rect 30425 845 30503 891
rect 30549 845 30627 891
rect 30673 845 30751 891
rect 30797 845 30875 891
rect 30921 845 30999 891
rect 31045 845 31123 891
rect 31169 845 31247 891
rect 31293 845 31371 891
rect 31417 845 31495 891
rect 31541 845 31619 891
rect 31665 845 31743 891
rect 31789 845 31867 891
rect 31913 845 31991 891
rect 32037 845 32115 891
rect 32161 845 32239 891
rect 32285 845 32363 891
rect 32409 845 32487 891
rect 32533 845 32611 891
rect 32657 845 32735 891
rect 32781 845 32859 891
rect 32905 845 32983 891
rect 33029 845 33107 891
rect 33153 845 33231 891
rect 33277 845 33355 891
rect 33401 845 33479 891
rect 33525 845 33603 891
rect 33649 845 33727 891
rect 33773 845 33851 891
rect 33897 845 33975 891
rect 34021 845 34099 891
rect 34145 845 34223 891
rect 34269 845 34347 891
rect 34393 845 34471 891
rect 34517 845 34595 891
rect 34641 845 34719 891
rect 34765 845 34843 891
rect 34889 845 34967 891
rect 35013 845 35091 891
rect 35137 845 35215 891
rect 35261 845 35339 891
rect 35385 845 35463 891
rect 35509 845 35587 891
rect 35633 845 35711 891
rect 35757 845 35835 891
rect 35881 845 35959 891
rect 36005 845 36083 891
rect 36129 845 36207 891
rect 36253 845 36331 891
rect 36377 845 36455 891
rect 36501 845 36579 891
rect 36625 845 36703 891
rect 36749 845 36827 891
rect 36873 845 36951 891
rect 36997 845 37075 891
rect 37121 845 37199 891
rect 37245 845 37323 891
rect 37369 845 37447 891
rect 37493 845 37571 891
rect 37617 845 37695 891
rect 37741 845 37819 891
rect 37865 845 37943 891
rect 37989 845 38067 891
rect 38113 845 38191 891
rect 38237 845 38315 891
rect 38361 845 38439 891
rect 38485 845 38563 891
rect 38609 845 38687 891
rect 38733 845 38811 891
rect 38857 845 38935 891
rect 38981 845 39059 891
rect 39105 845 39183 891
rect 39229 845 39307 891
rect 39353 845 39431 891
rect 39477 845 39555 891
rect 39601 845 39679 891
rect 39725 845 39803 891
rect 39849 845 39927 891
rect 39973 845 40051 891
rect 40097 845 40175 891
rect 40221 845 40299 891
rect 40345 845 40423 891
rect 40469 845 40547 891
rect 40593 845 40671 891
rect 40717 845 40795 891
rect 40841 845 40919 891
rect 40965 845 41043 891
rect 41089 845 41167 891
rect 41213 845 41291 891
rect 41337 845 41415 891
rect 41461 845 41539 891
rect 41585 845 41663 891
rect 41709 845 41787 891
rect 41833 845 41911 891
rect 41957 845 42035 891
rect 42081 845 42159 891
rect 42205 845 42283 891
rect 42329 845 42407 891
rect 42453 845 42531 891
rect 42577 845 42655 891
rect 42701 845 42779 891
rect 42825 845 42903 891
rect 42949 845 43027 891
rect 43073 845 43151 891
rect 43197 845 43275 891
rect 43321 845 43399 891
rect 43445 845 43523 891
rect 43569 845 43647 891
rect 43693 845 43771 891
rect 43817 845 43895 891
rect 43941 845 44019 891
rect 44065 845 44143 891
rect 44189 845 44267 891
rect 44313 845 44391 891
rect 44437 845 44515 891
rect 44561 845 44639 891
rect 44685 845 44763 891
rect 44809 845 44887 891
rect 44933 845 45011 891
rect 45057 845 45135 891
rect 45181 845 45259 891
rect 45305 845 45383 891
rect 45429 845 45507 891
rect 45553 845 45631 891
rect 45677 845 45755 891
rect 45801 845 45879 891
rect 45925 845 46003 891
rect 46049 845 46127 891
rect 46173 845 46251 891
rect 46297 845 46375 891
rect 46421 845 46499 891
rect 46545 845 46623 891
rect 46669 845 46747 891
rect 46793 845 46871 891
rect 46917 845 46995 891
rect 47041 845 47119 891
rect 47165 845 47243 891
rect 47289 845 47367 891
rect 47413 845 47491 891
rect 47537 845 47615 891
rect 47661 845 47739 891
rect 47785 845 47863 891
rect 47909 845 47987 891
rect 48033 845 48111 891
rect 48157 845 48235 891
rect 48281 845 48359 891
rect 48405 845 48483 891
rect 48529 845 48607 891
rect 48653 845 48731 891
rect 48777 845 48855 891
rect 48901 845 48979 891
rect 49025 845 49103 891
rect 49149 845 49227 891
rect 49273 845 49351 891
rect 49397 845 49475 891
rect 49521 845 49599 891
rect 49645 845 49723 891
rect 49769 845 49847 891
rect 49893 845 49971 891
rect 50017 845 50095 891
rect 50141 845 50219 891
rect 50265 845 50343 891
rect 50389 845 50467 891
rect 50513 845 50591 891
rect 50637 845 50715 891
rect 50761 845 50839 891
rect 50885 845 50963 891
rect 51009 845 51087 891
rect 51133 845 51211 891
rect 51257 845 51335 891
rect 51381 845 51459 891
rect 51505 845 51583 891
rect 51629 845 51707 891
rect 51753 845 51831 891
rect 51877 845 51955 891
rect 52001 845 52079 891
rect 52125 845 52203 891
rect 52249 845 52327 891
rect 52373 845 52451 891
rect 52497 845 52575 891
rect 52621 845 52699 891
rect 52745 845 52823 891
rect 52869 845 52947 891
rect 52993 845 53071 891
rect 53117 845 53195 891
rect 53241 845 53319 891
rect 53365 845 53443 891
rect 53489 845 53567 891
rect 53613 845 53691 891
rect 53737 845 53815 891
rect 53861 845 53939 891
rect 53985 845 54063 891
rect 54109 845 54187 891
rect 54233 845 54311 891
rect 54357 845 54435 891
rect 54481 845 54559 891
rect 54605 845 54683 891
rect 54729 845 54807 891
rect 54853 845 54931 891
rect 54977 845 55055 891
rect 55101 845 55179 891
rect 55225 845 55303 891
rect 55349 845 55427 891
rect 55473 845 55551 891
rect 55597 845 55675 891
rect 55721 845 55799 891
rect 55845 845 55923 891
rect 55969 845 56047 891
rect 56093 845 56171 891
rect 56217 845 56295 891
rect 56341 845 56419 891
rect 56465 845 56543 891
rect 56589 845 56667 891
rect 56713 845 56791 891
rect 56837 845 56915 891
rect 56961 845 57039 891
rect 57085 845 57163 891
rect 57209 845 57287 891
rect 57333 845 57411 891
rect 57457 845 57535 891
rect 57581 845 57659 891
rect 57705 845 57783 891
rect 57829 845 57907 891
rect 57953 845 58031 891
rect 58077 845 58155 891
rect 58201 845 58279 891
rect 58325 845 58403 891
rect 58449 845 58527 891
rect 58573 845 58651 891
rect 58697 845 58775 891
rect 58821 845 58899 891
rect 58945 845 59023 891
rect 59069 845 59147 891
rect 59193 845 59271 891
rect 59317 845 59395 891
rect 59441 845 59519 891
rect 59565 845 59643 891
rect 59689 845 59767 891
rect 59813 845 59891 891
rect 59937 845 60015 891
rect 60061 845 60139 891
rect 60185 845 60263 891
rect 60309 845 60387 891
rect 60433 845 60511 891
rect 60557 845 60635 891
rect 60681 845 60759 891
rect 60805 845 60883 891
rect 60929 845 61007 891
rect 61053 845 61131 891
rect 61177 845 61255 891
rect 61301 845 61379 891
rect 61425 845 61503 891
rect 61549 845 61627 891
rect 61673 845 61751 891
rect 61797 845 61875 891
rect 61921 845 61999 891
rect 62045 845 62123 891
rect 62169 845 62247 891
rect 62293 845 62371 891
rect 62417 845 62495 891
rect 62541 845 62619 891
rect 62665 845 62743 891
rect 62789 845 62867 891
rect 62913 845 62991 891
rect 63037 845 63115 891
rect 63161 845 63239 891
rect 63285 845 63363 891
rect 63409 845 63487 891
rect 63533 845 63611 891
rect 63657 845 63735 891
rect 63781 845 63859 891
rect 63905 845 63983 891
rect 64029 845 64107 891
rect 64153 845 64231 891
rect 64277 845 64355 891
rect 64401 845 64479 891
rect 64525 845 64603 891
rect 64649 845 64727 891
rect 64773 845 64851 891
rect 64897 845 64975 891
rect 65021 845 65099 891
rect 65145 845 65223 891
rect 65269 845 65347 891
rect 65393 845 65471 891
rect 65517 845 65595 891
rect 65641 845 65719 891
rect 65765 845 65843 891
rect 65889 845 65967 891
rect 66013 845 66091 891
rect 66137 845 66215 891
rect 66261 845 66339 891
rect 66385 845 66463 891
rect 66509 845 66587 891
rect 66633 845 66711 891
rect 66757 845 66835 891
rect 66881 845 66959 891
rect 67005 845 67083 891
rect 67129 845 67207 891
rect 67253 845 67331 891
rect 67377 845 67455 891
rect 67501 845 67579 891
rect 67625 845 67703 891
rect 67749 845 67827 891
rect 67873 845 67951 891
rect 67997 845 68075 891
rect 68121 845 68199 891
rect 68245 845 68323 891
rect 68369 845 68447 891
rect 68493 845 68571 891
rect 68617 845 68695 891
rect 68741 845 68819 891
rect 68865 845 68943 891
rect 68989 845 69067 891
rect 69113 845 69191 891
rect 69237 845 69315 891
rect 69361 845 69439 891
rect 69485 845 69563 891
rect 69609 845 69687 891
rect 69733 845 69811 891
rect 69857 845 69935 891
rect 69981 845 70059 891
rect 70105 845 70183 891
rect 70229 845 70307 891
rect 70353 845 70431 891
rect 70477 845 70555 891
rect 70601 845 70679 891
rect 70725 845 70803 891
rect 70849 845 70927 891
rect 70973 845 71051 891
rect 71097 845 71175 891
rect 71221 845 71299 891
rect 71345 845 71423 891
rect 71469 845 71547 891
rect 71593 845 71671 891
rect 71717 845 71795 891
rect 71841 845 71919 891
rect 71965 845 72043 891
rect 72089 845 72167 891
rect 72213 845 72291 891
rect 72337 845 72415 891
rect 72461 845 72539 891
rect 72585 845 72663 891
rect 72709 845 72787 891
rect 72833 845 72911 891
rect 72957 845 73035 891
rect 73081 845 73159 891
rect 73205 845 73283 891
rect 73329 845 73407 891
rect 73453 845 73531 891
rect 73577 845 73655 891
rect 73701 845 73779 891
rect 73825 845 73903 891
rect 73949 845 74027 891
rect 74073 845 74151 891
rect 74197 845 74275 891
rect 74321 845 74399 891
rect 74445 845 74523 891
rect 74569 845 74647 891
rect 74693 845 74771 891
rect 74817 845 74895 891
rect 74941 845 75019 891
rect 75065 845 75143 891
rect 75189 845 75267 891
rect 75313 845 75391 891
rect 75437 845 75515 891
rect 75561 845 75639 891
rect 75685 845 75763 891
rect 75809 845 75887 891
rect 75933 845 76011 891
rect 76057 845 76135 891
rect 76181 845 76259 891
rect 76305 845 76383 891
rect 76429 845 76507 891
rect 76553 845 76631 891
rect 76677 845 76755 891
rect 76801 845 76879 891
rect 76925 845 77003 891
rect 77049 845 77127 891
rect 77173 845 77251 891
rect 77297 845 77375 891
rect 77421 845 77499 891
rect 77545 845 77623 891
rect 77669 845 77747 891
rect 77793 845 77871 891
rect 77917 845 77995 891
rect 78041 845 78119 891
rect 78165 845 78243 891
rect 78289 845 78367 891
rect 78413 845 78491 891
rect 78537 845 78615 891
rect 78661 845 78739 891
rect 78785 845 78863 891
rect 78909 845 78987 891
rect 79033 845 79111 891
rect 79157 845 79235 891
rect 79281 845 79359 891
rect 79405 845 79483 891
rect 79529 845 79607 891
rect 79653 845 79731 891
rect 79777 845 79855 891
rect 79901 845 79979 891
rect 80025 845 80103 891
rect 80149 845 80227 891
rect 80273 845 80351 891
rect 80397 845 80475 891
rect 80521 845 80599 891
rect 80645 845 80723 891
rect 80769 845 80847 891
rect 80893 845 80971 891
rect 81017 845 81095 891
rect 81141 845 81219 891
rect 81265 845 81343 891
rect 81389 845 81467 891
rect 81513 845 81591 891
rect 81637 845 81715 891
rect 81761 845 81839 891
rect 81885 845 81963 891
rect 82009 845 82087 891
rect 82133 845 82211 891
rect 82257 845 82335 891
rect 82381 845 82459 891
rect 82505 845 82583 891
rect 82629 845 82707 891
rect 82753 845 82831 891
rect 82877 845 82955 891
rect 83001 845 83079 891
rect 83125 845 83203 891
rect 83249 845 83327 891
rect 83373 845 83451 891
rect 83497 845 83575 891
rect 83621 845 83699 891
rect 83745 845 83823 891
rect 83869 845 83947 891
rect 83993 845 84071 891
rect 84117 845 84195 891
rect 84241 845 84319 891
rect 84365 845 84443 891
rect 84489 845 84567 891
rect 84613 845 84691 891
rect 84737 845 84815 891
rect 84861 845 84939 891
rect 84985 845 85063 891
rect 85109 845 85187 891
rect 85233 845 85311 891
rect 85357 845 85435 891
rect 85481 845 85559 891
rect 85605 845 85683 891
rect 85729 845 85807 891
rect 85853 845 85931 891
rect 85977 845 86098 891
rect 352 767 86098 845
rect 352 721 371 767
rect 417 721 495 767
rect 541 721 619 767
rect 665 721 743 767
rect 789 721 867 767
rect 913 721 991 767
rect 1037 721 1115 767
rect 1161 721 1239 767
rect 1285 721 1363 767
rect 1409 721 1487 767
rect 1533 721 1611 767
rect 1657 721 1735 767
rect 1781 721 1859 767
rect 1905 721 1983 767
rect 2029 721 2107 767
rect 2153 721 2231 767
rect 2277 721 2355 767
rect 2401 721 2479 767
rect 2525 721 2603 767
rect 2649 721 2727 767
rect 2773 721 2851 767
rect 2897 721 2975 767
rect 3021 721 3099 767
rect 3145 721 3223 767
rect 3269 721 3347 767
rect 3393 721 3471 767
rect 3517 721 3595 767
rect 3641 721 3719 767
rect 3765 721 3843 767
rect 3889 721 3967 767
rect 4013 721 4091 767
rect 4137 721 4215 767
rect 4261 721 4339 767
rect 4385 721 4463 767
rect 4509 721 4587 767
rect 4633 721 4711 767
rect 4757 721 4835 767
rect 4881 721 4959 767
rect 5005 721 5083 767
rect 5129 721 5207 767
rect 5253 721 5331 767
rect 5377 721 5455 767
rect 5501 721 5579 767
rect 5625 721 5703 767
rect 5749 721 5827 767
rect 5873 721 5951 767
rect 5997 721 6075 767
rect 6121 721 6199 767
rect 6245 721 6323 767
rect 6369 721 6447 767
rect 6493 721 6571 767
rect 6617 721 6695 767
rect 6741 721 6819 767
rect 6865 721 6943 767
rect 6989 721 7067 767
rect 7113 721 7191 767
rect 7237 721 7315 767
rect 7361 721 7439 767
rect 7485 721 7563 767
rect 7609 721 7687 767
rect 7733 721 7811 767
rect 7857 721 7935 767
rect 7981 721 8059 767
rect 8105 721 8183 767
rect 8229 721 8307 767
rect 8353 721 8431 767
rect 8477 721 8555 767
rect 8601 721 8679 767
rect 8725 721 8803 767
rect 8849 721 8927 767
rect 8973 721 9051 767
rect 9097 721 9175 767
rect 9221 721 9299 767
rect 9345 721 9423 767
rect 9469 721 9547 767
rect 9593 721 9671 767
rect 9717 721 9795 767
rect 9841 721 9919 767
rect 9965 721 10043 767
rect 10089 721 10167 767
rect 10213 721 10291 767
rect 10337 721 10415 767
rect 10461 721 10539 767
rect 10585 721 10663 767
rect 10709 721 10787 767
rect 10833 721 10911 767
rect 10957 721 11035 767
rect 11081 721 11159 767
rect 11205 721 11283 767
rect 11329 721 11407 767
rect 11453 721 11531 767
rect 11577 721 11655 767
rect 11701 721 11779 767
rect 11825 721 11903 767
rect 11949 721 12027 767
rect 12073 721 12151 767
rect 12197 721 12275 767
rect 12321 721 12399 767
rect 12445 721 12523 767
rect 12569 721 12647 767
rect 12693 721 12771 767
rect 12817 721 12895 767
rect 12941 721 13019 767
rect 13065 721 13143 767
rect 13189 721 13267 767
rect 13313 721 13391 767
rect 13437 721 13515 767
rect 13561 721 13639 767
rect 13685 721 13763 767
rect 13809 721 13887 767
rect 13933 721 14011 767
rect 14057 721 14135 767
rect 14181 721 14259 767
rect 14305 721 14383 767
rect 14429 721 14507 767
rect 14553 721 14631 767
rect 14677 721 14755 767
rect 14801 721 14879 767
rect 14925 721 15003 767
rect 15049 721 15127 767
rect 15173 721 15251 767
rect 15297 721 15375 767
rect 15421 721 15499 767
rect 15545 721 15623 767
rect 15669 721 15747 767
rect 15793 721 15871 767
rect 15917 721 15995 767
rect 16041 721 16119 767
rect 16165 721 16243 767
rect 16289 721 16367 767
rect 16413 721 16491 767
rect 16537 721 16615 767
rect 16661 721 16739 767
rect 16785 721 16863 767
rect 16909 721 16987 767
rect 17033 721 17111 767
rect 17157 721 17235 767
rect 17281 721 17359 767
rect 17405 721 17483 767
rect 17529 721 17607 767
rect 17653 721 17731 767
rect 17777 721 17855 767
rect 17901 721 17979 767
rect 18025 721 18103 767
rect 18149 721 18227 767
rect 18273 721 18351 767
rect 18397 721 18475 767
rect 18521 721 18599 767
rect 18645 721 18723 767
rect 18769 721 18847 767
rect 18893 721 18971 767
rect 19017 721 19095 767
rect 19141 721 19219 767
rect 19265 721 19343 767
rect 19389 721 19467 767
rect 19513 721 19591 767
rect 19637 721 19715 767
rect 19761 721 19839 767
rect 19885 721 19963 767
rect 20009 721 20087 767
rect 20133 721 20211 767
rect 20257 721 20335 767
rect 20381 721 20459 767
rect 20505 721 20583 767
rect 20629 721 20707 767
rect 20753 721 20831 767
rect 20877 721 20955 767
rect 21001 721 21079 767
rect 21125 721 21203 767
rect 21249 721 21327 767
rect 21373 721 21451 767
rect 21497 721 21575 767
rect 21621 721 21699 767
rect 21745 721 21823 767
rect 21869 721 21947 767
rect 21993 721 22071 767
rect 22117 721 22195 767
rect 22241 721 22319 767
rect 22365 721 22443 767
rect 22489 721 22567 767
rect 22613 721 22691 767
rect 22737 721 22815 767
rect 22861 721 22939 767
rect 22985 721 23063 767
rect 23109 721 23187 767
rect 23233 721 23311 767
rect 23357 721 23435 767
rect 23481 721 23559 767
rect 23605 721 23683 767
rect 23729 721 23807 767
rect 23853 721 23931 767
rect 23977 721 24055 767
rect 24101 721 24179 767
rect 24225 721 24303 767
rect 24349 721 24427 767
rect 24473 721 24551 767
rect 24597 721 24675 767
rect 24721 721 24799 767
rect 24845 721 24923 767
rect 24969 721 25047 767
rect 25093 721 25171 767
rect 25217 721 25295 767
rect 25341 721 25419 767
rect 25465 721 25543 767
rect 25589 721 25667 767
rect 25713 721 25791 767
rect 25837 721 25915 767
rect 25961 721 26039 767
rect 26085 721 26163 767
rect 26209 721 26287 767
rect 26333 721 26411 767
rect 26457 721 26535 767
rect 26581 721 26659 767
rect 26705 721 26783 767
rect 26829 721 26907 767
rect 26953 721 27031 767
rect 27077 721 27155 767
rect 27201 721 27279 767
rect 27325 721 27403 767
rect 27449 721 27527 767
rect 27573 721 27651 767
rect 27697 721 27775 767
rect 27821 721 27899 767
rect 27945 721 28023 767
rect 28069 721 28147 767
rect 28193 721 28271 767
rect 28317 721 28395 767
rect 28441 721 28519 767
rect 28565 721 28643 767
rect 28689 721 28767 767
rect 28813 721 28891 767
rect 28937 721 29015 767
rect 29061 721 29139 767
rect 29185 721 29263 767
rect 29309 721 29387 767
rect 29433 721 29511 767
rect 29557 721 29635 767
rect 29681 721 29759 767
rect 29805 721 29883 767
rect 29929 721 30007 767
rect 30053 721 30131 767
rect 30177 721 30255 767
rect 30301 721 30379 767
rect 30425 721 30503 767
rect 30549 721 30627 767
rect 30673 721 30751 767
rect 30797 721 30875 767
rect 30921 721 30999 767
rect 31045 721 31123 767
rect 31169 721 31247 767
rect 31293 721 31371 767
rect 31417 721 31495 767
rect 31541 721 31619 767
rect 31665 721 31743 767
rect 31789 721 31867 767
rect 31913 721 31991 767
rect 32037 721 32115 767
rect 32161 721 32239 767
rect 32285 721 32363 767
rect 32409 721 32487 767
rect 32533 721 32611 767
rect 32657 721 32735 767
rect 32781 721 32859 767
rect 32905 721 32983 767
rect 33029 721 33107 767
rect 33153 721 33231 767
rect 33277 721 33355 767
rect 33401 721 33479 767
rect 33525 721 33603 767
rect 33649 721 33727 767
rect 33773 721 33851 767
rect 33897 721 33975 767
rect 34021 721 34099 767
rect 34145 721 34223 767
rect 34269 721 34347 767
rect 34393 721 34471 767
rect 34517 721 34595 767
rect 34641 721 34719 767
rect 34765 721 34843 767
rect 34889 721 34967 767
rect 35013 721 35091 767
rect 35137 721 35215 767
rect 35261 721 35339 767
rect 35385 721 35463 767
rect 35509 721 35587 767
rect 35633 721 35711 767
rect 35757 721 35835 767
rect 35881 721 35959 767
rect 36005 721 36083 767
rect 36129 721 36207 767
rect 36253 721 36331 767
rect 36377 721 36455 767
rect 36501 721 36579 767
rect 36625 721 36703 767
rect 36749 721 36827 767
rect 36873 721 36951 767
rect 36997 721 37075 767
rect 37121 721 37199 767
rect 37245 721 37323 767
rect 37369 721 37447 767
rect 37493 721 37571 767
rect 37617 721 37695 767
rect 37741 721 37819 767
rect 37865 721 37943 767
rect 37989 721 38067 767
rect 38113 721 38191 767
rect 38237 721 38315 767
rect 38361 721 38439 767
rect 38485 721 38563 767
rect 38609 721 38687 767
rect 38733 721 38811 767
rect 38857 721 38935 767
rect 38981 721 39059 767
rect 39105 721 39183 767
rect 39229 721 39307 767
rect 39353 721 39431 767
rect 39477 721 39555 767
rect 39601 721 39679 767
rect 39725 721 39803 767
rect 39849 721 39927 767
rect 39973 721 40051 767
rect 40097 721 40175 767
rect 40221 721 40299 767
rect 40345 721 40423 767
rect 40469 721 40547 767
rect 40593 721 40671 767
rect 40717 721 40795 767
rect 40841 721 40919 767
rect 40965 721 41043 767
rect 41089 721 41167 767
rect 41213 721 41291 767
rect 41337 721 41415 767
rect 41461 721 41539 767
rect 41585 721 41663 767
rect 41709 721 41787 767
rect 41833 721 41911 767
rect 41957 721 42035 767
rect 42081 721 42159 767
rect 42205 721 42283 767
rect 42329 721 42407 767
rect 42453 721 42531 767
rect 42577 721 42655 767
rect 42701 721 42779 767
rect 42825 721 42903 767
rect 42949 721 43027 767
rect 43073 721 43151 767
rect 43197 721 43275 767
rect 43321 721 43399 767
rect 43445 721 43523 767
rect 43569 721 43647 767
rect 43693 721 43771 767
rect 43817 721 43895 767
rect 43941 721 44019 767
rect 44065 721 44143 767
rect 44189 721 44267 767
rect 44313 721 44391 767
rect 44437 721 44515 767
rect 44561 721 44639 767
rect 44685 721 44763 767
rect 44809 721 44887 767
rect 44933 721 45011 767
rect 45057 721 45135 767
rect 45181 721 45259 767
rect 45305 721 45383 767
rect 45429 721 45507 767
rect 45553 721 45631 767
rect 45677 721 45755 767
rect 45801 721 45879 767
rect 45925 721 46003 767
rect 46049 721 46127 767
rect 46173 721 46251 767
rect 46297 721 46375 767
rect 46421 721 46499 767
rect 46545 721 46623 767
rect 46669 721 46747 767
rect 46793 721 46871 767
rect 46917 721 46995 767
rect 47041 721 47119 767
rect 47165 721 47243 767
rect 47289 721 47367 767
rect 47413 721 47491 767
rect 47537 721 47615 767
rect 47661 721 47739 767
rect 47785 721 47863 767
rect 47909 721 47987 767
rect 48033 721 48111 767
rect 48157 721 48235 767
rect 48281 721 48359 767
rect 48405 721 48483 767
rect 48529 721 48607 767
rect 48653 721 48731 767
rect 48777 721 48855 767
rect 48901 721 48979 767
rect 49025 721 49103 767
rect 49149 721 49227 767
rect 49273 721 49351 767
rect 49397 721 49475 767
rect 49521 721 49599 767
rect 49645 721 49723 767
rect 49769 721 49847 767
rect 49893 721 49971 767
rect 50017 721 50095 767
rect 50141 721 50219 767
rect 50265 721 50343 767
rect 50389 721 50467 767
rect 50513 721 50591 767
rect 50637 721 50715 767
rect 50761 721 50839 767
rect 50885 721 50963 767
rect 51009 721 51087 767
rect 51133 721 51211 767
rect 51257 721 51335 767
rect 51381 721 51459 767
rect 51505 721 51583 767
rect 51629 721 51707 767
rect 51753 721 51831 767
rect 51877 721 51955 767
rect 52001 721 52079 767
rect 52125 721 52203 767
rect 52249 721 52327 767
rect 52373 721 52451 767
rect 52497 721 52575 767
rect 52621 721 52699 767
rect 52745 721 52823 767
rect 52869 721 52947 767
rect 52993 721 53071 767
rect 53117 721 53195 767
rect 53241 721 53319 767
rect 53365 721 53443 767
rect 53489 721 53567 767
rect 53613 721 53691 767
rect 53737 721 53815 767
rect 53861 721 53939 767
rect 53985 721 54063 767
rect 54109 721 54187 767
rect 54233 721 54311 767
rect 54357 721 54435 767
rect 54481 721 54559 767
rect 54605 721 54683 767
rect 54729 721 54807 767
rect 54853 721 54931 767
rect 54977 721 55055 767
rect 55101 721 55179 767
rect 55225 721 55303 767
rect 55349 721 55427 767
rect 55473 721 55551 767
rect 55597 721 55675 767
rect 55721 721 55799 767
rect 55845 721 55923 767
rect 55969 721 56047 767
rect 56093 721 56171 767
rect 56217 721 56295 767
rect 56341 721 56419 767
rect 56465 721 56543 767
rect 56589 721 56667 767
rect 56713 721 56791 767
rect 56837 721 56915 767
rect 56961 721 57039 767
rect 57085 721 57163 767
rect 57209 721 57287 767
rect 57333 721 57411 767
rect 57457 721 57535 767
rect 57581 721 57659 767
rect 57705 721 57783 767
rect 57829 721 57907 767
rect 57953 721 58031 767
rect 58077 721 58155 767
rect 58201 721 58279 767
rect 58325 721 58403 767
rect 58449 721 58527 767
rect 58573 721 58651 767
rect 58697 721 58775 767
rect 58821 721 58899 767
rect 58945 721 59023 767
rect 59069 721 59147 767
rect 59193 721 59271 767
rect 59317 721 59395 767
rect 59441 721 59519 767
rect 59565 721 59643 767
rect 59689 721 59767 767
rect 59813 721 59891 767
rect 59937 721 60015 767
rect 60061 721 60139 767
rect 60185 721 60263 767
rect 60309 721 60387 767
rect 60433 721 60511 767
rect 60557 721 60635 767
rect 60681 721 60759 767
rect 60805 721 60883 767
rect 60929 721 61007 767
rect 61053 721 61131 767
rect 61177 721 61255 767
rect 61301 721 61379 767
rect 61425 721 61503 767
rect 61549 721 61627 767
rect 61673 721 61751 767
rect 61797 721 61875 767
rect 61921 721 61999 767
rect 62045 721 62123 767
rect 62169 721 62247 767
rect 62293 721 62371 767
rect 62417 721 62495 767
rect 62541 721 62619 767
rect 62665 721 62743 767
rect 62789 721 62867 767
rect 62913 721 62991 767
rect 63037 721 63115 767
rect 63161 721 63239 767
rect 63285 721 63363 767
rect 63409 721 63487 767
rect 63533 721 63611 767
rect 63657 721 63735 767
rect 63781 721 63859 767
rect 63905 721 63983 767
rect 64029 721 64107 767
rect 64153 721 64231 767
rect 64277 721 64355 767
rect 64401 721 64479 767
rect 64525 721 64603 767
rect 64649 721 64727 767
rect 64773 721 64851 767
rect 64897 721 64975 767
rect 65021 721 65099 767
rect 65145 721 65223 767
rect 65269 721 65347 767
rect 65393 721 65471 767
rect 65517 721 65595 767
rect 65641 721 65719 767
rect 65765 721 65843 767
rect 65889 721 65967 767
rect 66013 721 66091 767
rect 66137 721 66215 767
rect 66261 721 66339 767
rect 66385 721 66463 767
rect 66509 721 66587 767
rect 66633 721 66711 767
rect 66757 721 66835 767
rect 66881 721 66959 767
rect 67005 721 67083 767
rect 67129 721 67207 767
rect 67253 721 67331 767
rect 67377 721 67455 767
rect 67501 721 67579 767
rect 67625 721 67703 767
rect 67749 721 67827 767
rect 67873 721 67951 767
rect 67997 721 68075 767
rect 68121 721 68199 767
rect 68245 721 68323 767
rect 68369 721 68447 767
rect 68493 721 68571 767
rect 68617 721 68695 767
rect 68741 721 68819 767
rect 68865 721 68943 767
rect 68989 721 69067 767
rect 69113 721 69191 767
rect 69237 721 69315 767
rect 69361 721 69439 767
rect 69485 721 69563 767
rect 69609 721 69687 767
rect 69733 721 69811 767
rect 69857 721 69935 767
rect 69981 721 70059 767
rect 70105 721 70183 767
rect 70229 721 70307 767
rect 70353 721 70431 767
rect 70477 721 70555 767
rect 70601 721 70679 767
rect 70725 721 70803 767
rect 70849 721 70927 767
rect 70973 721 71051 767
rect 71097 721 71175 767
rect 71221 721 71299 767
rect 71345 721 71423 767
rect 71469 721 71547 767
rect 71593 721 71671 767
rect 71717 721 71795 767
rect 71841 721 71919 767
rect 71965 721 72043 767
rect 72089 721 72167 767
rect 72213 721 72291 767
rect 72337 721 72415 767
rect 72461 721 72539 767
rect 72585 721 72663 767
rect 72709 721 72787 767
rect 72833 721 72911 767
rect 72957 721 73035 767
rect 73081 721 73159 767
rect 73205 721 73283 767
rect 73329 721 73407 767
rect 73453 721 73531 767
rect 73577 721 73655 767
rect 73701 721 73779 767
rect 73825 721 73903 767
rect 73949 721 74027 767
rect 74073 721 74151 767
rect 74197 721 74275 767
rect 74321 721 74399 767
rect 74445 721 74523 767
rect 74569 721 74647 767
rect 74693 721 74771 767
rect 74817 721 74895 767
rect 74941 721 75019 767
rect 75065 721 75143 767
rect 75189 721 75267 767
rect 75313 721 75391 767
rect 75437 721 75515 767
rect 75561 721 75639 767
rect 75685 721 75763 767
rect 75809 721 75887 767
rect 75933 721 76011 767
rect 76057 721 76135 767
rect 76181 721 76259 767
rect 76305 721 76383 767
rect 76429 721 76507 767
rect 76553 721 76631 767
rect 76677 721 76755 767
rect 76801 721 76879 767
rect 76925 721 77003 767
rect 77049 721 77127 767
rect 77173 721 77251 767
rect 77297 721 77375 767
rect 77421 721 77499 767
rect 77545 721 77623 767
rect 77669 721 77747 767
rect 77793 721 77871 767
rect 77917 721 77995 767
rect 78041 721 78119 767
rect 78165 721 78243 767
rect 78289 721 78367 767
rect 78413 721 78491 767
rect 78537 721 78615 767
rect 78661 721 78739 767
rect 78785 721 78863 767
rect 78909 721 78987 767
rect 79033 721 79111 767
rect 79157 721 79235 767
rect 79281 721 79359 767
rect 79405 721 79483 767
rect 79529 721 79607 767
rect 79653 721 79731 767
rect 79777 721 79855 767
rect 79901 721 79979 767
rect 80025 721 80103 767
rect 80149 721 80227 767
rect 80273 721 80351 767
rect 80397 721 80475 767
rect 80521 721 80599 767
rect 80645 721 80723 767
rect 80769 721 80847 767
rect 80893 721 80971 767
rect 81017 721 81095 767
rect 81141 721 81219 767
rect 81265 721 81343 767
rect 81389 721 81467 767
rect 81513 721 81591 767
rect 81637 721 81715 767
rect 81761 721 81839 767
rect 81885 721 81963 767
rect 82009 721 82087 767
rect 82133 721 82211 767
rect 82257 721 82335 767
rect 82381 721 82459 767
rect 82505 721 82583 767
rect 82629 721 82707 767
rect 82753 721 82831 767
rect 82877 721 82955 767
rect 83001 721 83079 767
rect 83125 721 83203 767
rect 83249 721 83327 767
rect 83373 721 83451 767
rect 83497 721 83575 767
rect 83621 721 83699 767
rect 83745 721 83823 767
rect 83869 721 83947 767
rect 83993 721 84071 767
rect 84117 721 84195 767
rect 84241 721 84319 767
rect 84365 721 84443 767
rect 84489 721 84567 767
rect 84613 721 84691 767
rect 84737 721 84815 767
rect 84861 721 84939 767
rect 84985 721 85063 767
rect 85109 721 85187 767
rect 85233 721 85311 767
rect 85357 721 85435 767
rect 85481 721 85559 767
rect 85605 721 85683 767
rect 85729 721 85807 767
rect 85853 721 85931 767
rect 85977 721 86098 767
rect 352 643 86098 721
rect 352 597 371 643
rect 417 597 495 643
rect 541 597 619 643
rect 665 597 743 643
rect 789 597 867 643
rect 913 597 991 643
rect 1037 597 1115 643
rect 1161 597 1239 643
rect 1285 597 1363 643
rect 1409 597 1487 643
rect 1533 597 1611 643
rect 1657 597 1735 643
rect 1781 597 1859 643
rect 1905 597 1983 643
rect 2029 597 2107 643
rect 2153 597 2231 643
rect 2277 597 2355 643
rect 2401 597 2479 643
rect 2525 597 2603 643
rect 2649 597 2727 643
rect 2773 597 2851 643
rect 2897 597 2975 643
rect 3021 597 3099 643
rect 3145 597 3223 643
rect 3269 597 3347 643
rect 3393 597 3471 643
rect 3517 597 3595 643
rect 3641 597 3719 643
rect 3765 597 3843 643
rect 3889 597 3967 643
rect 4013 597 4091 643
rect 4137 597 4215 643
rect 4261 597 4339 643
rect 4385 597 4463 643
rect 4509 597 4587 643
rect 4633 597 4711 643
rect 4757 597 4835 643
rect 4881 597 4959 643
rect 5005 597 5083 643
rect 5129 597 5207 643
rect 5253 597 5331 643
rect 5377 597 5455 643
rect 5501 597 5579 643
rect 5625 597 5703 643
rect 5749 597 5827 643
rect 5873 597 5951 643
rect 5997 597 6075 643
rect 6121 597 6199 643
rect 6245 597 6323 643
rect 6369 597 6447 643
rect 6493 597 6571 643
rect 6617 597 6695 643
rect 6741 597 6819 643
rect 6865 597 6943 643
rect 6989 597 7067 643
rect 7113 597 7191 643
rect 7237 597 7315 643
rect 7361 597 7439 643
rect 7485 597 7563 643
rect 7609 597 7687 643
rect 7733 597 7811 643
rect 7857 597 7935 643
rect 7981 597 8059 643
rect 8105 597 8183 643
rect 8229 597 8307 643
rect 8353 597 8431 643
rect 8477 597 8555 643
rect 8601 597 8679 643
rect 8725 597 8803 643
rect 8849 597 8927 643
rect 8973 597 9051 643
rect 9097 597 9175 643
rect 9221 597 9299 643
rect 9345 597 9423 643
rect 9469 597 9547 643
rect 9593 597 9671 643
rect 9717 597 9795 643
rect 9841 597 9919 643
rect 9965 597 10043 643
rect 10089 597 10167 643
rect 10213 597 10291 643
rect 10337 597 10415 643
rect 10461 597 10539 643
rect 10585 597 10663 643
rect 10709 597 10787 643
rect 10833 597 10911 643
rect 10957 597 11035 643
rect 11081 597 11159 643
rect 11205 597 11283 643
rect 11329 597 11407 643
rect 11453 597 11531 643
rect 11577 597 11655 643
rect 11701 597 11779 643
rect 11825 597 11903 643
rect 11949 597 12027 643
rect 12073 597 12151 643
rect 12197 597 12275 643
rect 12321 597 12399 643
rect 12445 597 12523 643
rect 12569 597 12647 643
rect 12693 597 12771 643
rect 12817 597 12895 643
rect 12941 597 13019 643
rect 13065 597 13143 643
rect 13189 597 13267 643
rect 13313 597 13391 643
rect 13437 597 13515 643
rect 13561 597 13639 643
rect 13685 597 13763 643
rect 13809 597 13887 643
rect 13933 597 14011 643
rect 14057 597 14135 643
rect 14181 597 14259 643
rect 14305 597 14383 643
rect 14429 597 14507 643
rect 14553 597 14631 643
rect 14677 597 14755 643
rect 14801 597 14879 643
rect 14925 597 15003 643
rect 15049 597 15127 643
rect 15173 597 15251 643
rect 15297 597 15375 643
rect 15421 597 15499 643
rect 15545 597 15623 643
rect 15669 597 15747 643
rect 15793 597 15871 643
rect 15917 597 15995 643
rect 16041 597 16119 643
rect 16165 597 16243 643
rect 16289 597 16367 643
rect 16413 597 16491 643
rect 16537 597 16615 643
rect 16661 597 16739 643
rect 16785 597 16863 643
rect 16909 597 16987 643
rect 17033 597 17111 643
rect 17157 597 17235 643
rect 17281 597 17359 643
rect 17405 597 17483 643
rect 17529 597 17607 643
rect 17653 597 17731 643
rect 17777 597 17855 643
rect 17901 597 17979 643
rect 18025 597 18103 643
rect 18149 597 18227 643
rect 18273 597 18351 643
rect 18397 597 18475 643
rect 18521 597 18599 643
rect 18645 597 18723 643
rect 18769 597 18847 643
rect 18893 597 18971 643
rect 19017 597 19095 643
rect 19141 597 19219 643
rect 19265 597 19343 643
rect 19389 597 19467 643
rect 19513 597 19591 643
rect 19637 597 19715 643
rect 19761 597 19839 643
rect 19885 597 19963 643
rect 20009 597 20087 643
rect 20133 597 20211 643
rect 20257 597 20335 643
rect 20381 597 20459 643
rect 20505 597 20583 643
rect 20629 597 20707 643
rect 20753 597 20831 643
rect 20877 597 20955 643
rect 21001 597 21079 643
rect 21125 597 21203 643
rect 21249 597 21327 643
rect 21373 597 21451 643
rect 21497 597 21575 643
rect 21621 597 21699 643
rect 21745 597 21823 643
rect 21869 597 21947 643
rect 21993 597 22071 643
rect 22117 597 22195 643
rect 22241 597 22319 643
rect 22365 597 22443 643
rect 22489 597 22567 643
rect 22613 597 22691 643
rect 22737 597 22815 643
rect 22861 597 22939 643
rect 22985 597 23063 643
rect 23109 597 23187 643
rect 23233 597 23311 643
rect 23357 597 23435 643
rect 23481 597 23559 643
rect 23605 597 23683 643
rect 23729 597 23807 643
rect 23853 597 23931 643
rect 23977 597 24055 643
rect 24101 597 24179 643
rect 24225 597 24303 643
rect 24349 597 24427 643
rect 24473 597 24551 643
rect 24597 597 24675 643
rect 24721 597 24799 643
rect 24845 597 24923 643
rect 24969 597 25047 643
rect 25093 597 25171 643
rect 25217 597 25295 643
rect 25341 597 25419 643
rect 25465 597 25543 643
rect 25589 597 25667 643
rect 25713 597 25791 643
rect 25837 597 25915 643
rect 25961 597 26039 643
rect 26085 597 26163 643
rect 26209 597 26287 643
rect 26333 597 26411 643
rect 26457 597 26535 643
rect 26581 597 26659 643
rect 26705 597 26783 643
rect 26829 597 26907 643
rect 26953 597 27031 643
rect 27077 597 27155 643
rect 27201 597 27279 643
rect 27325 597 27403 643
rect 27449 597 27527 643
rect 27573 597 27651 643
rect 27697 597 27775 643
rect 27821 597 27899 643
rect 27945 597 28023 643
rect 28069 597 28147 643
rect 28193 597 28271 643
rect 28317 597 28395 643
rect 28441 597 28519 643
rect 28565 597 28643 643
rect 28689 597 28767 643
rect 28813 597 28891 643
rect 28937 597 29015 643
rect 29061 597 29139 643
rect 29185 597 29263 643
rect 29309 597 29387 643
rect 29433 597 29511 643
rect 29557 597 29635 643
rect 29681 597 29759 643
rect 29805 597 29883 643
rect 29929 597 30007 643
rect 30053 597 30131 643
rect 30177 597 30255 643
rect 30301 597 30379 643
rect 30425 597 30503 643
rect 30549 597 30627 643
rect 30673 597 30751 643
rect 30797 597 30875 643
rect 30921 597 30999 643
rect 31045 597 31123 643
rect 31169 597 31247 643
rect 31293 597 31371 643
rect 31417 597 31495 643
rect 31541 597 31619 643
rect 31665 597 31743 643
rect 31789 597 31867 643
rect 31913 597 31991 643
rect 32037 597 32115 643
rect 32161 597 32239 643
rect 32285 597 32363 643
rect 32409 597 32487 643
rect 32533 597 32611 643
rect 32657 597 32735 643
rect 32781 597 32859 643
rect 32905 597 32983 643
rect 33029 597 33107 643
rect 33153 597 33231 643
rect 33277 597 33355 643
rect 33401 597 33479 643
rect 33525 597 33603 643
rect 33649 597 33727 643
rect 33773 597 33851 643
rect 33897 597 33975 643
rect 34021 597 34099 643
rect 34145 597 34223 643
rect 34269 597 34347 643
rect 34393 597 34471 643
rect 34517 597 34595 643
rect 34641 597 34719 643
rect 34765 597 34843 643
rect 34889 597 34967 643
rect 35013 597 35091 643
rect 35137 597 35215 643
rect 35261 597 35339 643
rect 35385 597 35463 643
rect 35509 597 35587 643
rect 35633 597 35711 643
rect 35757 597 35835 643
rect 35881 597 35959 643
rect 36005 597 36083 643
rect 36129 597 36207 643
rect 36253 597 36331 643
rect 36377 597 36455 643
rect 36501 597 36579 643
rect 36625 597 36703 643
rect 36749 597 36827 643
rect 36873 597 36951 643
rect 36997 597 37075 643
rect 37121 597 37199 643
rect 37245 597 37323 643
rect 37369 597 37447 643
rect 37493 597 37571 643
rect 37617 597 37695 643
rect 37741 597 37819 643
rect 37865 597 37943 643
rect 37989 597 38067 643
rect 38113 597 38191 643
rect 38237 597 38315 643
rect 38361 597 38439 643
rect 38485 597 38563 643
rect 38609 597 38687 643
rect 38733 597 38811 643
rect 38857 597 38935 643
rect 38981 597 39059 643
rect 39105 597 39183 643
rect 39229 597 39307 643
rect 39353 597 39431 643
rect 39477 597 39555 643
rect 39601 597 39679 643
rect 39725 597 39803 643
rect 39849 597 39927 643
rect 39973 597 40051 643
rect 40097 597 40175 643
rect 40221 597 40299 643
rect 40345 597 40423 643
rect 40469 597 40547 643
rect 40593 597 40671 643
rect 40717 597 40795 643
rect 40841 597 40919 643
rect 40965 597 41043 643
rect 41089 597 41167 643
rect 41213 597 41291 643
rect 41337 597 41415 643
rect 41461 597 41539 643
rect 41585 597 41663 643
rect 41709 597 41787 643
rect 41833 597 41911 643
rect 41957 597 42035 643
rect 42081 597 42159 643
rect 42205 597 42283 643
rect 42329 597 42407 643
rect 42453 597 42531 643
rect 42577 597 42655 643
rect 42701 597 42779 643
rect 42825 597 42903 643
rect 42949 597 43027 643
rect 43073 597 43151 643
rect 43197 597 43275 643
rect 43321 597 43399 643
rect 43445 597 43523 643
rect 43569 597 43647 643
rect 43693 597 43771 643
rect 43817 597 43895 643
rect 43941 597 44019 643
rect 44065 597 44143 643
rect 44189 597 44267 643
rect 44313 597 44391 643
rect 44437 597 44515 643
rect 44561 597 44639 643
rect 44685 597 44763 643
rect 44809 597 44887 643
rect 44933 597 45011 643
rect 45057 597 45135 643
rect 45181 597 45259 643
rect 45305 597 45383 643
rect 45429 597 45507 643
rect 45553 597 45631 643
rect 45677 597 45755 643
rect 45801 597 45879 643
rect 45925 597 46003 643
rect 46049 597 46127 643
rect 46173 597 46251 643
rect 46297 597 46375 643
rect 46421 597 46499 643
rect 46545 597 46623 643
rect 46669 597 46747 643
rect 46793 597 46871 643
rect 46917 597 46995 643
rect 47041 597 47119 643
rect 47165 597 47243 643
rect 47289 597 47367 643
rect 47413 597 47491 643
rect 47537 597 47615 643
rect 47661 597 47739 643
rect 47785 597 47863 643
rect 47909 597 47987 643
rect 48033 597 48111 643
rect 48157 597 48235 643
rect 48281 597 48359 643
rect 48405 597 48483 643
rect 48529 597 48607 643
rect 48653 597 48731 643
rect 48777 597 48855 643
rect 48901 597 48979 643
rect 49025 597 49103 643
rect 49149 597 49227 643
rect 49273 597 49351 643
rect 49397 597 49475 643
rect 49521 597 49599 643
rect 49645 597 49723 643
rect 49769 597 49847 643
rect 49893 597 49971 643
rect 50017 597 50095 643
rect 50141 597 50219 643
rect 50265 597 50343 643
rect 50389 597 50467 643
rect 50513 597 50591 643
rect 50637 597 50715 643
rect 50761 597 50839 643
rect 50885 597 50963 643
rect 51009 597 51087 643
rect 51133 597 51211 643
rect 51257 597 51335 643
rect 51381 597 51459 643
rect 51505 597 51583 643
rect 51629 597 51707 643
rect 51753 597 51831 643
rect 51877 597 51955 643
rect 52001 597 52079 643
rect 52125 597 52203 643
rect 52249 597 52327 643
rect 52373 597 52451 643
rect 52497 597 52575 643
rect 52621 597 52699 643
rect 52745 597 52823 643
rect 52869 597 52947 643
rect 52993 597 53071 643
rect 53117 597 53195 643
rect 53241 597 53319 643
rect 53365 597 53443 643
rect 53489 597 53567 643
rect 53613 597 53691 643
rect 53737 597 53815 643
rect 53861 597 53939 643
rect 53985 597 54063 643
rect 54109 597 54187 643
rect 54233 597 54311 643
rect 54357 597 54435 643
rect 54481 597 54559 643
rect 54605 597 54683 643
rect 54729 597 54807 643
rect 54853 597 54931 643
rect 54977 597 55055 643
rect 55101 597 55179 643
rect 55225 597 55303 643
rect 55349 597 55427 643
rect 55473 597 55551 643
rect 55597 597 55675 643
rect 55721 597 55799 643
rect 55845 597 55923 643
rect 55969 597 56047 643
rect 56093 597 56171 643
rect 56217 597 56295 643
rect 56341 597 56419 643
rect 56465 597 56543 643
rect 56589 597 56667 643
rect 56713 597 56791 643
rect 56837 597 56915 643
rect 56961 597 57039 643
rect 57085 597 57163 643
rect 57209 597 57287 643
rect 57333 597 57411 643
rect 57457 597 57535 643
rect 57581 597 57659 643
rect 57705 597 57783 643
rect 57829 597 57907 643
rect 57953 597 58031 643
rect 58077 597 58155 643
rect 58201 597 58279 643
rect 58325 597 58403 643
rect 58449 597 58527 643
rect 58573 597 58651 643
rect 58697 597 58775 643
rect 58821 597 58899 643
rect 58945 597 59023 643
rect 59069 597 59147 643
rect 59193 597 59271 643
rect 59317 597 59395 643
rect 59441 597 59519 643
rect 59565 597 59643 643
rect 59689 597 59767 643
rect 59813 597 59891 643
rect 59937 597 60015 643
rect 60061 597 60139 643
rect 60185 597 60263 643
rect 60309 597 60387 643
rect 60433 597 60511 643
rect 60557 597 60635 643
rect 60681 597 60759 643
rect 60805 597 60883 643
rect 60929 597 61007 643
rect 61053 597 61131 643
rect 61177 597 61255 643
rect 61301 597 61379 643
rect 61425 597 61503 643
rect 61549 597 61627 643
rect 61673 597 61751 643
rect 61797 597 61875 643
rect 61921 597 61999 643
rect 62045 597 62123 643
rect 62169 597 62247 643
rect 62293 597 62371 643
rect 62417 597 62495 643
rect 62541 597 62619 643
rect 62665 597 62743 643
rect 62789 597 62867 643
rect 62913 597 62991 643
rect 63037 597 63115 643
rect 63161 597 63239 643
rect 63285 597 63363 643
rect 63409 597 63487 643
rect 63533 597 63611 643
rect 63657 597 63735 643
rect 63781 597 63859 643
rect 63905 597 63983 643
rect 64029 597 64107 643
rect 64153 597 64231 643
rect 64277 597 64355 643
rect 64401 597 64479 643
rect 64525 597 64603 643
rect 64649 597 64727 643
rect 64773 597 64851 643
rect 64897 597 64975 643
rect 65021 597 65099 643
rect 65145 597 65223 643
rect 65269 597 65347 643
rect 65393 597 65471 643
rect 65517 597 65595 643
rect 65641 597 65719 643
rect 65765 597 65843 643
rect 65889 597 65967 643
rect 66013 597 66091 643
rect 66137 597 66215 643
rect 66261 597 66339 643
rect 66385 597 66463 643
rect 66509 597 66587 643
rect 66633 597 66711 643
rect 66757 597 66835 643
rect 66881 597 66959 643
rect 67005 597 67083 643
rect 67129 597 67207 643
rect 67253 597 67331 643
rect 67377 597 67455 643
rect 67501 597 67579 643
rect 67625 597 67703 643
rect 67749 597 67827 643
rect 67873 597 67951 643
rect 67997 597 68075 643
rect 68121 597 68199 643
rect 68245 597 68323 643
rect 68369 597 68447 643
rect 68493 597 68571 643
rect 68617 597 68695 643
rect 68741 597 68819 643
rect 68865 597 68943 643
rect 68989 597 69067 643
rect 69113 597 69191 643
rect 69237 597 69315 643
rect 69361 597 69439 643
rect 69485 597 69563 643
rect 69609 597 69687 643
rect 69733 597 69811 643
rect 69857 597 69935 643
rect 69981 597 70059 643
rect 70105 597 70183 643
rect 70229 597 70307 643
rect 70353 597 70431 643
rect 70477 597 70555 643
rect 70601 597 70679 643
rect 70725 597 70803 643
rect 70849 597 70927 643
rect 70973 597 71051 643
rect 71097 597 71175 643
rect 71221 597 71299 643
rect 71345 597 71423 643
rect 71469 597 71547 643
rect 71593 597 71671 643
rect 71717 597 71795 643
rect 71841 597 71919 643
rect 71965 597 72043 643
rect 72089 597 72167 643
rect 72213 597 72291 643
rect 72337 597 72415 643
rect 72461 597 72539 643
rect 72585 597 72663 643
rect 72709 597 72787 643
rect 72833 597 72911 643
rect 72957 597 73035 643
rect 73081 597 73159 643
rect 73205 597 73283 643
rect 73329 597 73407 643
rect 73453 597 73531 643
rect 73577 597 73655 643
rect 73701 597 73779 643
rect 73825 597 73903 643
rect 73949 597 74027 643
rect 74073 597 74151 643
rect 74197 597 74275 643
rect 74321 597 74399 643
rect 74445 597 74523 643
rect 74569 597 74647 643
rect 74693 597 74771 643
rect 74817 597 74895 643
rect 74941 597 75019 643
rect 75065 597 75143 643
rect 75189 597 75267 643
rect 75313 597 75391 643
rect 75437 597 75515 643
rect 75561 597 75639 643
rect 75685 597 75763 643
rect 75809 597 75887 643
rect 75933 597 76011 643
rect 76057 597 76135 643
rect 76181 597 76259 643
rect 76305 597 76383 643
rect 76429 597 76507 643
rect 76553 597 76631 643
rect 76677 597 76755 643
rect 76801 597 76879 643
rect 76925 597 77003 643
rect 77049 597 77127 643
rect 77173 597 77251 643
rect 77297 597 77375 643
rect 77421 597 77499 643
rect 77545 597 77623 643
rect 77669 597 77747 643
rect 77793 597 77871 643
rect 77917 597 77995 643
rect 78041 597 78119 643
rect 78165 597 78243 643
rect 78289 597 78367 643
rect 78413 597 78491 643
rect 78537 597 78615 643
rect 78661 597 78739 643
rect 78785 597 78863 643
rect 78909 597 78987 643
rect 79033 597 79111 643
rect 79157 597 79235 643
rect 79281 597 79359 643
rect 79405 597 79483 643
rect 79529 597 79607 643
rect 79653 597 79731 643
rect 79777 597 79855 643
rect 79901 597 79979 643
rect 80025 597 80103 643
rect 80149 597 80227 643
rect 80273 597 80351 643
rect 80397 597 80475 643
rect 80521 597 80599 643
rect 80645 597 80723 643
rect 80769 597 80847 643
rect 80893 597 80971 643
rect 81017 597 81095 643
rect 81141 597 81219 643
rect 81265 597 81343 643
rect 81389 597 81467 643
rect 81513 597 81591 643
rect 81637 597 81715 643
rect 81761 597 81839 643
rect 81885 597 81963 643
rect 82009 597 82087 643
rect 82133 597 82211 643
rect 82257 597 82335 643
rect 82381 597 82459 643
rect 82505 597 82583 643
rect 82629 597 82707 643
rect 82753 597 82831 643
rect 82877 597 82955 643
rect 83001 597 83079 643
rect 83125 597 83203 643
rect 83249 597 83327 643
rect 83373 597 83451 643
rect 83497 597 83575 643
rect 83621 597 83699 643
rect 83745 597 83823 643
rect 83869 597 83947 643
rect 83993 597 84071 643
rect 84117 597 84195 643
rect 84241 597 84319 643
rect 84365 597 84443 643
rect 84489 597 84567 643
rect 84613 597 84691 643
rect 84737 597 84815 643
rect 84861 597 84939 643
rect 84985 597 85063 643
rect 85109 597 85187 643
rect 85233 597 85311 643
rect 85357 597 85435 643
rect 85481 597 85559 643
rect 85605 597 85683 643
rect 85729 597 85807 643
rect 85853 597 85931 643
rect 85977 597 86098 643
rect 352 578 86098 597
<< mvpsubdiffcont >>
rect 371 96637 417 96683
rect 495 96637 541 96683
rect 619 96637 665 96683
rect 743 96637 789 96683
rect 867 96637 913 96683
rect 991 96637 1037 96683
rect 1115 96637 1161 96683
rect 1239 96637 1285 96683
rect 1363 96637 1409 96683
rect 1487 96637 1533 96683
rect 1611 96637 1657 96683
rect 1735 96637 1781 96683
rect 1859 96637 1905 96683
rect 1983 96637 2029 96683
rect 2107 96637 2153 96683
rect 2231 96637 2277 96683
rect 2355 96637 2401 96683
rect 2479 96637 2525 96683
rect 2603 96637 2649 96683
rect 2727 96637 2773 96683
rect 2851 96637 2897 96683
rect 2975 96637 3021 96683
rect 3099 96637 3145 96683
rect 3223 96637 3269 96683
rect 3347 96637 3393 96683
rect 3471 96637 3517 96683
rect 3595 96637 3641 96683
rect 3719 96637 3765 96683
rect 3843 96637 3889 96683
rect 3967 96637 4013 96683
rect 4091 96637 4137 96683
rect 4215 96637 4261 96683
rect 4339 96637 4385 96683
rect 4463 96637 4509 96683
rect 4587 96637 4633 96683
rect 4711 96637 4757 96683
rect 4835 96637 4881 96683
rect 4959 96637 5005 96683
rect 5083 96637 5129 96683
rect 5207 96637 5253 96683
rect 5331 96637 5377 96683
rect 5455 96637 5501 96683
rect 5579 96637 5625 96683
rect 5703 96637 5749 96683
rect 5827 96637 5873 96683
rect 5951 96637 5997 96683
rect 6075 96637 6121 96683
rect 6199 96637 6245 96683
rect 6323 96637 6369 96683
rect 6447 96637 6493 96683
rect 6571 96637 6617 96683
rect 6695 96637 6741 96683
rect 6819 96637 6865 96683
rect 6943 96637 6989 96683
rect 7067 96637 7113 96683
rect 7191 96637 7237 96683
rect 7315 96637 7361 96683
rect 7439 96637 7485 96683
rect 7563 96637 7609 96683
rect 7687 96637 7733 96683
rect 7811 96637 7857 96683
rect 7935 96637 7981 96683
rect 8059 96637 8105 96683
rect 8183 96637 8229 96683
rect 8307 96637 8353 96683
rect 8431 96637 8477 96683
rect 8555 96637 8601 96683
rect 8679 96637 8725 96683
rect 8803 96637 8849 96683
rect 8927 96637 8973 96683
rect 9051 96637 9097 96683
rect 9175 96637 9221 96683
rect 9299 96637 9345 96683
rect 9423 96637 9469 96683
rect 9547 96637 9593 96683
rect 9671 96637 9717 96683
rect 9795 96637 9841 96683
rect 9919 96637 9965 96683
rect 10043 96637 10089 96683
rect 10167 96637 10213 96683
rect 10291 96637 10337 96683
rect 10415 96637 10461 96683
rect 10539 96637 10585 96683
rect 10663 96637 10709 96683
rect 10787 96637 10833 96683
rect 10911 96637 10957 96683
rect 11035 96637 11081 96683
rect 11159 96637 11205 96683
rect 11283 96637 11329 96683
rect 11407 96637 11453 96683
rect 11531 96637 11577 96683
rect 11655 96637 11701 96683
rect 11779 96637 11825 96683
rect 11903 96637 11949 96683
rect 12027 96637 12073 96683
rect 12151 96637 12197 96683
rect 12275 96637 12321 96683
rect 12399 96637 12445 96683
rect 12523 96637 12569 96683
rect 12647 96637 12693 96683
rect 12771 96637 12817 96683
rect 12895 96637 12941 96683
rect 13019 96637 13065 96683
rect 13143 96637 13189 96683
rect 13267 96637 13313 96683
rect 13391 96637 13437 96683
rect 13515 96637 13561 96683
rect 13639 96637 13685 96683
rect 13763 96637 13809 96683
rect 13887 96637 13933 96683
rect 14011 96637 14057 96683
rect 14135 96637 14181 96683
rect 14259 96637 14305 96683
rect 14383 96637 14429 96683
rect 14507 96637 14553 96683
rect 14631 96637 14677 96683
rect 14755 96637 14801 96683
rect 14879 96637 14925 96683
rect 15003 96637 15049 96683
rect 15127 96637 15173 96683
rect 15251 96637 15297 96683
rect 15375 96637 15421 96683
rect 15499 96637 15545 96683
rect 15623 96637 15669 96683
rect 15747 96637 15793 96683
rect 15871 96637 15917 96683
rect 15995 96637 16041 96683
rect 16119 96637 16165 96683
rect 16243 96637 16289 96683
rect 16367 96637 16413 96683
rect 16491 96637 16537 96683
rect 16615 96637 16661 96683
rect 16739 96637 16785 96683
rect 16863 96637 16909 96683
rect 16987 96637 17033 96683
rect 17111 96637 17157 96683
rect 17235 96637 17281 96683
rect 17359 96637 17405 96683
rect 17483 96637 17529 96683
rect 17607 96637 17653 96683
rect 17731 96637 17777 96683
rect 17855 96637 17901 96683
rect 17979 96637 18025 96683
rect 18103 96637 18149 96683
rect 18227 96637 18273 96683
rect 18351 96637 18397 96683
rect 18475 96637 18521 96683
rect 18599 96637 18645 96683
rect 18723 96637 18769 96683
rect 18847 96637 18893 96683
rect 18971 96637 19017 96683
rect 19095 96637 19141 96683
rect 19219 96637 19265 96683
rect 19343 96637 19389 96683
rect 19467 96637 19513 96683
rect 19591 96637 19637 96683
rect 19715 96637 19761 96683
rect 19839 96637 19885 96683
rect 19963 96637 20009 96683
rect 20087 96637 20133 96683
rect 20211 96637 20257 96683
rect 20335 96637 20381 96683
rect 20459 96637 20505 96683
rect 20583 96637 20629 96683
rect 20707 96637 20753 96683
rect 20831 96637 20877 96683
rect 20955 96637 21001 96683
rect 21079 96637 21125 96683
rect 21203 96637 21249 96683
rect 21327 96637 21373 96683
rect 21451 96637 21497 96683
rect 21575 96637 21621 96683
rect 21699 96637 21745 96683
rect 21823 96637 21869 96683
rect 21947 96637 21993 96683
rect 22071 96637 22117 96683
rect 22195 96637 22241 96683
rect 22319 96637 22365 96683
rect 22443 96637 22489 96683
rect 22567 96637 22613 96683
rect 22691 96637 22737 96683
rect 22815 96637 22861 96683
rect 22939 96637 22985 96683
rect 23063 96637 23109 96683
rect 23187 96637 23233 96683
rect 23311 96637 23357 96683
rect 23435 96637 23481 96683
rect 23559 96637 23605 96683
rect 23683 96637 23729 96683
rect 23807 96637 23853 96683
rect 23931 96637 23977 96683
rect 24055 96637 24101 96683
rect 24179 96637 24225 96683
rect 24303 96637 24349 96683
rect 24427 96637 24473 96683
rect 24551 96637 24597 96683
rect 24675 96637 24721 96683
rect 24799 96637 24845 96683
rect 24923 96637 24969 96683
rect 25047 96637 25093 96683
rect 25171 96637 25217 96683
rect 25295 96637 25341 96683
rect 25419 96637 25465 96683
rect 25543 96637 25589 96683
rect 25667 96637 25713 96683
rect 25791 96637 25837 96683
rect 25915 96637 25961 96683
rect 26039 96637 26085 96683
rect 26163 96637 26209 96683
rect 26287 96637 26333 96683
rect 26411 96637 26457 96683
rect 26535 96637 26581 96683
rect 26659 96637 26705 96683
rect 26783 96637 26829 96683
rect 26907 96637 26953 96683
rect 27031 96637 27077 96683
rect 27155 96637 27201 96683
rect 27279 96637 27325 96683
rect 27403 96637 27449 96683
rect 27527 96637 27573 96683
rect 27651 96637 27697 96683
rect 27775 96637 27821 96683
rect 27899 96637 27945 96683
rect 28023 96637 28069 96683
rect 28147 96637 28193 96683
rect 28271 96637 28317 96683
rect 28395 96637 28441 96683
rect 28519 96637 28565 96683
rect 28643 96637 28689 96683
rect 28767 96637 28813 96683
rect 28891 96637 28937 96683
rect 29015 96637 29061 96683
rect 29139 96637 29185 96683
rect 29263 96637 29309 96683
rect 29387 96637 29433 96683
rect 29511 96637 29557 96683
rect 29635 96637 29681 96683
rect 29759 96637 29805 96683
rect 29883 96637 29929 96683
rect 30007 96637 30053 96683
rect 30131 96637 30177 96683
rect 30255 96637 30301 96683
rect 30379 96637 30425 96683
rect 30503 96637 30549 96683
rect 30627 96637 30673 96683
rect 30751 96637 30797 96683
rect 30875 96637 30921 96683
rect 30999 96637 31045 96683
rect 31123 96637 31169 96683
rect 31247 96637 31293 96683
rect 31371 96637 31417 96683
rect 31495 96637 31541 96683
rect 31619 96637 31665 96683
rect 31743 96637 31789 96683
rect 31867 96637 31913 96683
rect 31991 96637 32037 96683
rect 32115 96637 32161 96683
rect 32239 96637 32285 96683
rect 32363 96637 32409 96683
rect 32487 96637 32533 96683
rect 32611 96637 32657 96683
rect 32735 96637 32781 96683
rect 32859 96637 32905 96683
rect 32983 96637 33029 96683
rect 33107 96637 33153 96683
rect 33231 96637 33277 96683
rect 33355 96637 33401 96683
rect 33479 96637 33525 96683
rect 33603 96637 33649 96683
rect 33727 96637 33773 96683
rect 33851 96637 33897 96683
rect 33975 96637 34021 96683
rect 34099 96637 34145 96683
rect 34223 96637 34269 96683
rect 34347 96637 34393 96683
rect 34471 96637 34517 96683
rect 34595 96637 34641 96683
rect 34719 96637 34765 96683
rect 34843 96637 34889 96683
rect 34967 96637 35013 96683
rect 35091 96637 35137 96683
rect 35215 96637 35261 96683
rect 35339 96637 35385 96683
rect 35463 96637 35509 96683
rect 35587 96637 35633 96683
rect 35711 96637 35757 96683
rect 35835 96637 35881 96683
rect 35959 96637 36005 96683
rect 36083 96637 36129 96683
rect 36207 96637 36253 96683
rect 36331 96637 36377 96683
rect 36455 96637 36501 96683
rect 36579 96637 36625 96683
rect 36703 96637 36749 96683
rect 36827 96637 36873 96683
rect 36951 96637 36997 96683
rect 37075 96637 37121 96683
rect 37199 96637 37245 96683
rect 37323 96637 37369 96683
rect 37447 96637 37493 96683
rect 37571 96637 37617 96683
rect 37695 96637 37741 96683
rect 37819 96637 37865 96683
rect 37943 96637 37989 96683
rect 38067 96637 38113 96683
rect 38191 96637 38237 96683
rect 38315 96637 38361 96683
rect 38439 96637 38485 96683
rect 38563 96637 38609 96683
rect 38687 96637 38733 96683
rect 38811 96637 38857 96683
rect 38935 96637 38981 96683
rect 39059 96637 39105 96683
rect 39183 96637 39229 96683
rect 39307 96637 39353 96683
rect 39431 96637 39477 96683
rect 39555 96637 39601 96683
rect 39679 96637 39725 96683
rect 39803 96637 39849 96683
rect 39927 96637 39973 96683
rect 40051 96637 40097 96683
rect 40175 96637 40221 96683
rect 40299 96637 40345 96683
rect 40423 96637 40469 96683
rect 40547 96637 40593 96683
rect 40671 96637 40717 96683
rect 40795 96637 40841 96683
rect 40919 96637 40965 96683
rect 41043 96637 41089 96683
rect 41167 96637 41213 96683
rect 41291 96637 41337 96683
rect 41415 96637 41461 96683
rect 41539 96637 41585 96683
rect 41663 96637 41709 96683
rect 41787 96637 41833 96683
rect 41911 96637 41957 96683
rect 42035 96637 42081 96683
rect 42159 96637 42205 96683
rect 42283 96637 42329 96683
rect 42407 96637 42453 96683
rect 42531 96637 42577 96683
rect 42655 96637 42701 96683
rect 42779 96637 42825 96683
rect 42903 96637 42949 96683
rect 43027 96637 43073 96683
rect 43151 96637 43197 96683
rect 43275 96637 43321 96683
rect 43399 96637 43445 96683
rect 43523 96637 43569 96683
rect 43647 96637 43693 96683
rect 43771 96637 43817 96683
rect 43895 96637 43941 96683
rect 44019 96637 44065 96683
rect 44143 96637 44189 96683
rect 44267 96637 44313 96683
rect 44391 96637 44437 96683
rect 44515 96637 44561 96683
rect 44639 96637 44685 96683
rect 44763 96637 44809 96683
rect 44887 96637 44933 96683
rect 45011 96637 45057 96683
rect 45135 96637 45181 96683
rect 45259 96637 45305 96683
rect 45383 96637 45429 96683
rect 45507 96637 45553 96683
rect 45631 96637 45677 96683
rect 45755 96637 45801 96683
rect 45879 96637 45925 96683
rect 46003 96637 46049 96683
rect 46127 96637 46173 96683
rect 46251 96637 46297 96683
rect 46375 96637 46421 96683
rect 46499 96637 46545 96683
rect 46623 96637 46669 96683
rect 46747 96637 46793 96683
rect 46871 96637 46917 96683
rect 46995 96637 47041 96683
rect 47119 96637 47165 96683
rect 47243 96637 47289 96683
rect 47367 96637 47413 96683
rect 47491 96637 47537 96683
rect 47615 96637 47661 96683
rect 47739 96637 47785 96683
rect 47863 96637 47909 96683
rect 47987 96637 48033 96683
rect 48111 96637 48157 96683
rect 48235 96637 48281 96683
rect 48359 96637 48405 96683
rect 48483 96637 48529 96683
rect 48607 96637 48653 96683
rect 48731 96637 48777 96683
rect 48855 96637 48901 96683
rect 48979 96637 49025 96683
rect 49103 96637 49149 96683
rect 49227 96637 49273 96683
rect 49351 96637 49397 96683
rect 49475 96637 49521 96683
rect 49599 96637 49645 96683
rect 49723 96637 49769 96683
rect 49847 96637 49893 96683
rect 49971 96637 50017 96683
rect 50095 96637 50141 96683
rect 50219 96637 50265 96683
rect 50343 96637 50389 96683
rect 50467 96637 50513 96683
rect 50591 96637 50637 96683
rect 50715 96637 50761 96683
rect 50839 96637 50885 96683
rect 50963 96637 51009 96683
rect 51087 96637 51133 96683
rect 51211 96637 51257 96683
rect 51335 96637 51381 96683
rect 51459 96637 51505 96683
rect 51583 96637 51629 96683
rect 51707 96637 51753 96683
rect 51831 96637 51877 96683
rect 51955 96637 52001 96683
rect 52079 96637 52125 96683
rect 52203 96637 52249 96683
rect 52327 96637 52373 96683
rect 52451 96637 52497 96683
rect 52575 96637 52621 96683
rect 52699 96637 52745 96683
rect 52823 96637 52869 96683
rect 52947 96637 52993 96683
rect 53071 96637 53117 96683
rect 53195 96637 53241 96683
rect 53319 96637 53365 96683
rect 53443 96637 53489 96683
rect 53567 96637 53613 96683
rect 53691 96637 53737 96683
rect 53815 96637 53861 96683
rect 53939 96637 53985 96683
rect 54063 96637 54109 96683
rect 54187 96637 54233 96683
rect 54311 96637 54357 96683
rect 54435 96637 54481 96683
rect 54559 96637 54605 96683
rect 54683 96637 54729 96683
rect 54807 96637 54853 96683
rect 54931 96637 54977 96683
rect 55055 96637 55101 96683
rect 55179 96637 55225 96683
rect 55303 96637 55349 96683
rect 55427 96637 55473 96683
rect 55551 96637 55597 96683
rect 55675 96637 55721 96683
rect 55799 96637 55845 96683
rect 55923 96637 55969 96683
rect 56047 96637 56093 96683
rect 56171 96637 56217 96683
rect 56295 96637 56341 96683
rect 56419 96637 56465 96683
rect 56543 96637 56589 96683
rect 56667 96637 56713 96683
rect 56791 96637 56837 96683
rect 56915 96637 56961 96683
rect 57039 96637 57085 96683
rect 57163 96637 57209 96683
rect 57287 96637 57333 96683
rect 57411 96637 57457 96683
rect 57535 96637 57581 96683
rect 57659 96637 57705 96683
rect 57783 96637 57829 96683
rect 57907 96637 57953 96683
rect 58031 96637 58077 96683
rect 58155 96637 58201 96683
rect 58279 96637 58325 96683
rect 58403 96637 58449 96683
rect 58527 96637 58573 96683
rect 58651 96637 58697 96683
rect 58775 96637 58821 96683
rect 58899 96637 58945 96683
rect 59023 96637 59069 96683
rect 59147 96637 59193 96683
rect 59271 96637 59317 96683
rect 59395 96637 59441 96683
rect 59519 96637 59565 96683
rect 59643 96637 59689 96683
rect 59767 96637 59813 96683
rect 59891 96637 59937 96683
rect 60015 96637 60061 96683
rect 60139 96637 60185 96683
rect 60263 96637 60309 96683
rect 60387 96637 60433 96683
rect 60511 96637 60557 96683
rect 60635 96637 60681 96683
rect 60759 96637 60805 96683
rect 60883 96637 60929 96683
rect 61007 96637 61053 96683
rect 61131 96637 61177 96683
rect 61255 96637 61301 96683
rect 61379 96637 61425 96683
rect 61503 96637 61549 96683
rect 61627 96637 61673 96683
rect 61751 96637 61797 96683
rect 61875 96637 61921 96683
rect 61999 96637 62045 96683
rect 62123 96637 62169 96683
rect 62247 96637 62293 96683
rect 62371 96637 62417 96683
rect 62495 96637 62541 96683
rect 62619 96637 62665 96683
rect 62743 96637 62789 96683
rect 62867 96637 62913 96683
rect 62991 96637 63037 96683
rect 63115 96637 63161 96683
rect 63239 96637 63285 96683
rect 63363 96637 63409 96683
rect 63487 96637 63533 96683
rect 63611 96637 63657 96683
rect 63735 96637 63781 96683
rect 63859 96637 63905 96683
rect 63983 96637 64029 96683
rect 64107 96637 64153 96683
rect 64231 96637 64277 96683
rect 64355 96637 64401 96683
rect 64479 96637 64525 96683
rect 64603 96637 64649 96683
rect 64727 96637 64773 96683
rect 64851 96637 64897 96683
rect 64975 96637 65021 96683
rect 65099 96637 65145 96683
rect 65223 96637 65269 96683
rect 65347 96637 65393 96683
rect 65471 96637 65517 96683
rect 65595 96637 65641 96683
rect 65719 96637 65765 96683
rect 65843 96637 65889 96683
rect 65967 96637 66013 96683
rect 66091 96637 66137 96683
rect 66215 96637 66261 96683
rect 66339 96637 66385 96683
rect 66463 96637 66509 96683
rect 66587 96637 66633 96683
rect 66711 96637 66757 96683
rect 66835 96637 66881 96683
rect 66959 96637 67005 96683
rect 67083 96637 67129 96683
rect 67207 96637 67253 96683
rect 67331 96637 67377 96683
rect 67455 96637 67501 96683
rect 67579 96637 67625 96683
rect 67703 96637 67749 96683
rect 67827 96637 67873 96683
rect 67951 96637 67997 96683
rect 68075 96637 68121 96683
rect 68199 96637 68245 96683
rect 68323 96637 68369 96683
rect 68447 96637 68493 96683
rect 68571 96637 68617 96683
rect 68695 96637 68741 96683
rect 68819 96637 68865 96683
rect 68943 96637 68989 96683
rect 69067 96637 69113 96683
rect 69191 96637 69237 96683
rect 69315 96637 69361 96683
rect 69439 96637 69485 96683
rect 69563 96637 69609 96683
rect 69687 96637 69733 96683
rect 69811 96637 69857 96683
rect 69935 96637 69981 96683
rect 70059 96637 70105 96683
rect 70183 96637 70229 96683
rect 70307 96637 70353 96683
rect 70431 96637 70477 96683
rect 70555 96637 70601 96683
rect 70679 96637 70725 96683
rect 70803 96637 70849 96683
rect 70927 96637 70973 96683
rect 71051 96637 71097 96683
rect 71175 96637 71221 96683
rect 71299 96637 71345 96683
rect 71423 96637 71469 96683
rect 71547 96637 71593 96683
rect 71671 96637 71717 96683
rect 71795 96637 71841 96683
rect 71919 96637 71965 96683
rect 72043 96637 72089 96683
rect 72167 96637 72213 96683
rect 72291 96637 72337 96683
rect 72415 96637 72461 96683
rect 72539 96637 72585 96683
rect 72663 96637 72709 96683
rect 72787 96637 72833 96683
rect 72911 96637 72957 96683
rect 73035 96637 73081 96683
rect 73159 96637 73205 96683
rect 73283 96637 73329 96683
rect 73407 96637 73453 96683
rect 73531 96637 73577 96683
rect 73655 96637 73701 96683
rect 73779 96637 73825 96683
rect 73903 96637 73949 96683
rect 74027 96637 74073 96683
rect 74151 96637 74197 96683
rect 74275 96637 74321 96683
rect 74399 96637 74445 96683
rect 74523 96637 74569 96683
rect 74647 96637 74693 96683
rect 74771 96637 74817 96683
rect 74895 96637 74941 96683
rect 75019 96637 75065 96683
rect 75143 96637 75189 96683
rect 75267 96637 75313 96683
rect 75391 96637 75437 96683
rect 75515 96637 75561 96683
rect 75639 96637 75685 96683
rect 75763 96637 75809 96683
rect 75887 96637 75933 96683
rect 76011 96637 76057 96683
rect 76135 96637 76181 96683
rect 76259 96637 76305 96683
rect 76383 96637 76429 96683
rect 76507 96637 76553 96683
rect 76631 96637 76677 96683
rect 76755 96637 76801 96683
rect 76879 96637 76925 96683
rect 77003 96637 77049 96683
rect 77127 96637 77173 96683
rect 77251 96637 77297 96683
rect 77375 96637 77421 96683
rect 77499 96637 77545 96683
rect 77623 96637 77669 96683
rect 77747 96637 77793 96683
rect 77871 96637 77917 96683
rect 77995 96637 78041 96683
rect 78119 96637 78165 96683
rect 78243 96637 78289 96683
rect 78367 96637 78413 96683
rect 78491 96637 78537 96683
rect 78615 96637 78661 96683
rect 78739 96637 78785 96683
rect 78863 96637 78909 96683
rect 78987 96637 79033 96683
rect 79111 96637 79157 96683
rect 79235 96637 79281 96683
rect 79359 96637 79405 96683
rect 79483 96637 79529 96683
rect 79607 96637 79653 96683
rect 79731 96637 79777 96683
rect 79855 96637 79901 96683
rect 79979 96637 80025 96683
rect 80103 96637 80149 96683
rect 80227 96637 80273 96683
rect 80351 96637 80397 96683
rect 80475 96637 80521 96683
rect 80599 96637 80645 96683
rect 80723 96637 80769 96683
rect 80847 96637 80893 96683
rect 80971 96637 81017 96683
rect 81095 96637 81141 96683
rect 81219 96637 81265 96683
rect 81343 96637 81389 96683
rect 81467 96637 81513 96683
rect 81591 96637 81637 96683
rect 81715 96637 81761 96683
rect 81839 96637 81885 96683
rect 81963 96637 82009 96683
rect 82087 96637 82133 96683
rect 82211 96637 82257 96683
rect 82335 96637 82381 96683
rect 82459 96637 82505 96683
rect 82583 96637 82629 96683
rect 82707 96637 82753 96683
rect 82831 96637 82877 96683
rect 82955 96637 83001 96683
rect 83079 96637 83125 96683
rect 83203 96637 83249 96683
rect 83327 96637 83373 96683
rect 83451 96637 83497 96683
rect 83575 96637 83621 96683
rect 83699 96637 83745 96683
rect 83823 96637 83869 96683
rect 83947 96637 83993 96683
rect 84071 96637 84117 96683
rect 84195 96637 84241 96683
rect 84319 96637 84365 96683
rect 84443 96637 84489 96683
rect 84567 96637 84613 96683
rect 84691 96637 84737 96683
rect 84815 96637 84861 96683
rect 84939 96637 84985 96683
rect 85063 96637 85109 96683
rect 85187 96637 85233 96683
rect 85311 96637 85357 96683
rect 85435 96637 85481 96683
rect 85559 96637 85605 96683
rect 85683 96637 85729 96683
rect 85807 96637 85853 96683
rect 85931 96637 85977 96683
rect 371 96513 417 96559
rect 495 96513 541 96559
rect 619 96513 665 96559
rect 743 96513 789 96559
rect 867 96513 913 96559
rect 991 96513 1037 96559
rect 1115 96513 1161 96559
rect 1239 96513 1285 96559
rect 1363 96513 1409 96559
rect 1487 96513 1533 96559
rect 1611 96513 1657 96559
rect 1735 96513 1781 96559
rect 1859 96513 1905 96559
rect 1983 96513 2029 96559
rect 2107 96513 2153 96559
rect 2231 96513 2277 96559
rect 2355 96513 2401 96559
rect 2479 96513 2525 96559
rect 2603 96513 2649 96559
rect 2727 96513 2773 96559
rect 2851 96513 2897 96559
rect 2975 96513 3021 96559
rect 3099 96513 3145 96559
rect 3223 96513 3269 96559
rect 3347 96513 3393 96559
rect 3471 96513 3517 96559
rect 3595 96513 3641 96559
rect 3719 96513 3765 96559
rect 3843 96513 3889 96559
rect 3967 96513 4013 96559
rect 4091 96513 4137 96559
rect 4215 96513 4261 96559
rect 4339 96513 4385 96559
rect 4463 96513 4509 96559
rect 4587 96513 4633 96559
rect 4711 96513 4757 96559
rect 4835 96513 4881 96559
rect 4959 96513 5005 96559
rect 5083 96513 5129 96559
rect 5207 96513 5253 96559
rect 5331 96513 5377 96559
rect 5455 96513 5501 96559
rect 5579 96513 5625 96559
rect 5703 96513 5749 96559
rect 5827 96513 5873 96559
rect 5951 96513 5997 96559
rect 6075 96513 6121 96559
rect 6199 96513 6245 96559
rect 6323 96513 6369 96559
rect 6447 96513 6493 96559
rect 6571 96513 6617 96559
rect 6695 96513 6741 96559
rect 6819 96513 6865 96559
rect 6943 96513 6989 96559
rect 7067 96513 7113 96559
rect 7191 96513 7237 96559
rect 7315 96513 7361 96559
rect 7439 96513 7485 96559
rect 7563 96513 7609 96559
rect 7687 96513 7733 96559
rect 7811 96513 7857 96559
rect 7935 96513 7981 96559
rect 8059 96513 8105 96559
rect 8183 96513 8229 96559
rect 8307 96513 8353 96559
rect 8431 96513 8477 96559
rect 8555 96513 8601 96559
rect 8679 96513 8725 96559
rect 8803 96513 8849 96559
rect 8927 96513 8973 96559
rect 9051 96513 9097 96559
rect 9175 96513 9221 96559
rect 9299 96513 9345 96559
rect 9423 96513 9469 96559
rect 9547 96513 9593 96559
rect 9671 96513 9717 96559
rect 9795 96513 9841 96559
rect 9919 96513 9965 96559
rect 10043 96513 10089 96559
rect 10167 96513 10213 96559
rect 10291 96513 10337 96559
rect 10415 96513 10461 96559
rect 10539 96513 10585 96559
rect 10663 96513 10709 96559
rect 10787 96513 10833 96559
rect 10911 96513 10957 96559
rect 11035 96513 11081 96559
rect 11159 96513 11205 96559
rect 11283 96513 11329 96559
rect 11407 96513 11453 96559
rect 11531 96513 11577 96559
rect 11655 96513 11701 96559
rect 11779 96513 11825 96559
rect 11903 96513 11949 96559
rect 12027 96513 12073 96559
rect 12151 96513 12197 96559
rect 12275 96513 12321 96559
rect 12399 96513 12445 96559
rect 12523 96513 12569 96559
rect 12647 96513 12693 96559
rect 12771 96513 12817 96559
rect 12895 96513 12941 96559
rect 13019 96513 13065 96559
rect 13143 96513 13189 96559
rect 13267 96513 13313 96559
rect 13391 96513 13437 96559
rect 13515 96513 13561 96559
rect 13639 96513 13685 96559
rect 13763 96513 13809 96559
rect 13887 96513 13933 96559
rect 14011 96513 14057 96559
rect 14135 96513 14181 96559
rect 14259 96513 14305 96559
rect 14383 96513 14429 96559
rect 14507 96513 14553 96559
rect 14631 96513 14677 96559
rect 14755 96513 14801 96559
rect 14879 96513 14925 96559
rect 15003 96513 15049 96559
rect 15127 96513 15173 96559
rect 15251 96513 15297 96559
rect 15375 96513 15421 96559
rect 15499 96513 15545 96559
rect 15623 96513 15669 96559
rect 15747 96513 15793 96559
rect 15871 96513 15917 96559
rect 15995 96513 16041 96559
rect 16119 96513 16165 96559
rect 16243 96513 16289 96559
rect 16367 96513 16413 96559
rect 16491 96513 16537 96559
rect 16615 96513 16661 96559
rect 16739 96513 16785 96559
rect 16863 96513 16909 96559
rect 16987 96513 17033 96559
rect 17111 96513 17157 96559
rect 17235 96513 17281 96559
rect 17359 96513 17405 96559
rect 17483 96513 17529 96559
rect 17607 96513 17653 96559
rect 17731 96513 17777 96559
rect 17855 96513 17901 96559
rect 17979 96513 18025 96559
rect 18103 96513 18149 96559
rect 18227 96513 18273 96559
rect 18351 96513 18397 96559
rect 18475 96513 18521 96559
rect 18599 96513 18645 96559
rect 18723 96513 18769 96559
rect 18847 96513 18893 96559
rect 18971 96513 19017 96559
rect 19095 96513 19141 96559
rect 19219 96513 19265 96559
rect 19343 96513 19389 96559
rect 19467 96513 19513 96559
rect 19591 96513 19637 96559
rect 19715 96513 19761 96559
rect 19839 96513 19885 96559
rect 19963 96513 20009 96559
rect 20087 96513 20133 96559
rect 20211 96513 20257 96559
rect 20335 96513 20381 96559
rect 20459 96513 20505 96559
rect 20583 96513 20629 96559
rect 20707 96513 20753 96559
rect 20831 96513 20877 96559
rect 20955 96513 21001 96559
rect 21079 96513 21125 96559
rect 21203 96513 21249 96559
rect 21327 96513 21373 96559
rect 21451 96513 21497 96559
rect 21575 96513 21621 96559
rect 21699 96513 21745 96559
rect 21823 96513 21869 96559
rect 21947 96513 21993 96559
rect 22071 96513 22117 96559
rect 22195 96513 22241 96559
rect 22319 96513 22365 96559
rect 22443 96513 22489 96559
rect 22567 96513 22613 96559
rect 22691 96513 22737 96559
rect 22815 96513 22861 96559
rect 22939 96513 22985 96559
rect 23063 96513 23109 96559
rect 23187 96513 23233 96559
rect 23311 96513 23357 96559
rect 23435 96513 23481 96559
rect 23559 96513 23605 96559
rect 23683 96513 23729 96559
rect 23807 96513 23853 96559
rect 23931 96513 23977 96559
rect 24055 96513 24101 96559
rect 24179 96513 24225 96559
rect 24303 96513 24349 96559
rect 24427 96513 24473 96559
rect 24551 96513 24597 96559
rect 24675 96513 24721 96559
rect 24799 96513 24845 96559
rect 24923 96513 24969 96559
rect 25047 96513 25093 96559
rect 25171 96513 25217 96559
rect 25295 96513 25341 96559
rect 25419 96513 25465 96559
rect 25543 96513 25589 96559
rect 25667 96513 25713 96559
rect 25791 96513 25837 96559
rect 25915 96513 25961 96559
rect 26039 96513 26085 96559
rect 26163 96513 26209 96559
rect 26287 96513 26333 96559
rect 26411 96513 26457 96559
rect 26535 96513 26581 96559
rect 26659 96513 26705 96559
rect 26783 96513 26829 96559
rect 26907 96513 26953 96559
rect 27031 96513 27077 96559
rect 27155 96513 27201 96559
rect 27279 96513 27325 96559
rect 27403 96513 27449 96559
rect 27527 96513 27573 96559
rect 27651 96513 27697 96559
rect 27775 96513 27821 96559
rect 27899 96513 27945 96559
rect 28023 96513 28069 96559
rect 28147 96513 28193 96559
rect 28271 96513 28317 96559
rect 28395 96513 28441 96559
rect 28519 96513 28565 96559
rect 28643 96513 28689 96559
rect 28767 96513 28813 96559
rect 28891 96513 28937 96559
rect 29015 96513 29061 96559
rect 29139 96513 29185 96559
rect 29263 96513 29309 96559
rect 29387 96513 29433 96559
rect 29511 96513 29557 96559
rect 29635 96513 29681 96559
rect 29759 96513 29805 96559
rect 29883 96513 29929 96559
rect 30007 96513 30053 96559
rect 30131 96513 30177 96559
rect 30255 96513 30301 96559
rect 30379 96513 30425 96559
rect 30503 96513 30549 96559
rect 30627 96513 30673 96559
rect 30751 96513 30797 96559
rect 30875 96513 30921 96559
rect 30999 96513 31045 96559
rect 31123 96513 31169 96559
rect 31247 96513 31293 96559
rect 31371 96513 31417 96559
rect 31495 96513 31541 96559
rect 31619 96513 31665 96559
rect 31743 96513 31789 96559
rect 31867 96513 31913 96559
rect 31991 96513 32037 96559
rect 32115 96513 32161 96559
rect 32239 96513 32285 96559
rect 32363 96513 32409 96559
rect 32487 96513 32533 96559
rect 32611 96513 32657 96559
rect 32735 96513 32781 96559
rect 32859 96513 32905 96559
rect 32983 96513 33029 96559
rect 33107 96513 33153 96559
rect 33231 96513 33277 96559
rect 33355 96513 33401 96559
rect 33479 96513 33525 96559
rect 33603 96513 33649 96559
rect 33727 96513 33773 96559
rect 33851 96513 33897 96559
rect 33975 96513 34021 96559
rect 34099 96513 34145 96559
rect 34223 96513 34269 96559
rect 34347 96513 34393 96559
rect 34471 96513 34517 96559
rect 34595 96513 34641 96559
rect 34719 96513 34765 96559
rect 34843 96513 34889 96559
rect 34967 96513 35013 96559
rect 35091 96513 35137 96559
rect 35215 96513 35261 96559
rect 35339 96513 35385 96559
rect 35463 96513 35509 96559
rect 35587 96513 35633 96559
rect 35711 96513 35757 96559
rect 35835 96513 35881 96559
rect 35959 96513 36005 96559
rect 36083 96513 36129 96559
rect 36207 96513 36253 96559
rect 36331 96513 36377 96559
rect 36455 96513 36501 96559
rect 36579 96513 36625 96559
rect 36703 96513 36749 96559
rect 36827 96513 36873 96559
rect 36951 96513 36997 96559
rect 37075 96513 37121 96559
rect 37199 96513 37245 96559
rect 37323 96513 37369 96559
rect 37447 96513 37493 96559
rect 37571 96513 37617 96559
rect 37695 96513 37741 96559
rect 37819 96513 37865 96559
rect 37943 96513 37989 96559
rect 38067 96513 38113 96559
rect 38191 96513 38237 96559
rect 38315 96513 38361 96559
rect 38439 96513 38485 96559
rect 38563 96513 38609 96559
rect 38687 96513 38733 96559
rect 38811 96513 38857 96559
rect 38935 96513 38981 96559
rect 39059 96513 39105 96559
rect 39183 96513 39229 96559
rect 39307 96513 39353 96559
rect 39431 96513 39477 96559
rect 39555 96513 39601 96559
rect 39679 96513 39725 96559
rect 39803 96513 39849 96559
rect 39927 96513 39973 96559
rect 40051 96513 40097 96559
rect 40175 96513 40221 96559
rect 40299 96513 40345 96559
rect 40423 96513 40469 96559
rect 40547 96513 40593 96559
rect 40671 96513 40717 96559
rect 40795 96513 40841 96559
rect 40919 96513 40965 96559
rect 41043 96513 41089 96559
rect 41167 96513 41213 96559
rect 41291 96513 41337 96559
rect 41415 96513 41461 96559
rect 41539 96513 41585 96559
rect 41663 96513 41709 96559
rect 41787 96513 41833 96559
rect 41911 96513 41957 96559
rect 42035 96513 42081 96559
rect 42159 96513 42205 96559
rect 42283 96513 42329 96559
rect 42407 96513 42453 96559
rect 42531 96513 42577 96559
rect 42655 96513 42701 96559
rect 42779 96513 42825 96559
rect 42903 96513 42949 96559
rect 43027 96513 43073 96559
rect 43151 96513 43197 96559
rect 43275 96513 43321 96559
rect 43399 96513 43445 96559
rect 43523 96513 43569 96559
rect 43647 96513 43693 96559
rect 43771 96513 43817 96559
rect 43895 96513 43941 96559
rect 44019 96513 44065 96559
rect 44143 96513 44189 96559
rect 44267 96513 44313 96559
rect 44391 96513 44437 96559
rect 44515 96513 44561 96559
rect 44639 96513 44685 96559
rect 44763 96513 44809 96559
rect 44887 96513 44933 96559
rect 45011 96513 45057 96559
rect 45135 96513 45181 96559
rect 45259 96513 45305 96559
rect 45383 96513 45429 96559
rect 45507 96513 45553 96559
rect 45631 96513 45677 96559
rect 45755 96513 45801 96559
rect 45879 96513 45925 96559
rect 46003 96513 46049 96559
rect 46127 96513 46173 96559
rect 46251 96513 46297 96559
rect 46375 96513 46421 96559
rect 46499 96513 46545 96559
rect 46623 96513 46669 96559
rect 46747 96513 46793 96559
rect 46871 96513 46917 96559
rect 46995 96513 47041 96559
rect 47119 96513 47165 96559
rect 47243 96513 47289 96559
rect 47367 96513 47413 96559
rect 47491 96513 47537 96559
rect 47615 96513 47661 96559
rect 47739 96513 47785 96559
rect 47863 96513 47909 96559
rect 47987 96513 48033 96559
rect 48111 96513 48157 96559
rect 48235 96513 48281 96559
rect 48359 96513 48405 96559
rect 48483 96513 48529 96559
rect 48607 96513 48653 96559
rect 48731 96513 48777 96559
rect 48855 96513 48901 96559
rect 48979 96513 49025 96559
rect 49103 96513 49149 96559
rect 49227 96513 49273 96559
rect 49351 96513 49397 96559
rect 49475 96513 49521 96559
rect 49599 96513 49645 96559
rect 49723 96513 49769 96559
rect 49847 96513 49893 96559
rect 49971 96513 50017 96559
rect 50095 96513 50141 96559
rect 50219 96513 50265 96559
rect 50343 96513 50389 96559
rect 50467 96513 50513 96559
rect 50591 96513 50637 96559
rect 50715 96513 50761 96559
rect 50839 96513 50885 96559
rect 50963 96513 51009 96559
rect 51087 96513 51133 96559
rect 51211 96513 51257 96559
rect 51335 96513 51381 96559
rect 51459 96513 51505 96559
rect 51583 96513 51629 96559
rect 51707 96513 51753 96559
rect 51831 96513 51877 96559
rect 51955 96513 52001 96559
rect 52079 96513 52125 96559
rect 52203 96513 52249 96559
rect 52327 96513 52373 96559
rect 52451 96513 52497 96559
rect 52575 96513 52621 96559
rect 52699 96513 52745 96559
rect 52823 96513 52869 96559
rect 52947 96513 52993 96559
rect 53071 96513 53117 96559
rect 53195 96513 53241 96559
rect 53319 96513 53365 96559
rect 53443 96513 53489 96559
rect 53567 96513 53613 96559
rect 53691 96513 53737 96559
rect 53815 96513 53861 96559
rect 53939 96513 53985 96559
rect 54063 96513 54109 96559
rect 54187 96513 54233 96559
rect 54311 96513 54357 96559
rect 54435 96513 54481 96559
rect 54559 96513 54605 96559
rect 54683 96513 54729 96559
rect 54807 96513 54853 96559
rect 54931 96513 54977 96559
rect 55055 96513 55101 96559
rect 55179 96513 55225 96559
rect 55303 96513 55349 96559
rect 55427 96513 55473 96559
rect 55551 96513 55597 96559
rect 55675 96513 55721 96559
rect 55799 96513 55845 96559
rect 55923 96513 55969 96559
rect 56047 96513 56093 96559
rect 56171 96513 56217 96559
rect 56295 96513 56341 96559
rect 56419 96513 56465 96559
rect 56543 96513 56589 96559
rect 56667 96513 56713 96559
rect 56791 96513 56837 96559
rect 56915 96513 56961 96559
rect 57039 96513 57085 96559
rect 57163 96513 57209 96559
rect 57287 96513 57333 96559
rect 57411 96513 57457 96559
rect 57535 96513 57581 96559
rect 57659 96513 57705 96559
rect 57783 96513 57829 96559
rect 57907 96513 57953 96559
rect 58031 96513 58077 96559
rect 58155 96513 58201 96559
rect 58279 96513 58325 96559
rect 58403 96513 58449 96559
rect 58527 96513 58573 96559
rect 58651 96513 58697 96559
rect 58775 96513 58821 96559
rect 58899 96513 58945 96559
rect 59023 96513 59069 96559
rect 59147 96513 59193 96559
rect 59271 96513 59317 96559
rect 59395 96513 59441 96559
rect 59519 96513 59565 96559
rect 59643 96513 59689 96559
rect 59767 96513 59813 96559
rect 59891 96513 59937 96559
rect 60015 96513 60061 96559
rect 60139 96513 60185 96559
rect 60263 96513 60309 96559
rect 60387 96513 60433 96559
rect 60511 96513 60557 96559
rect 60635 96513 60681 96559
rect 60759 96513 60805 96559
rect 60883 96513 60929 96559
rect 61007 96513 61053 96559
rect 61131 96513 61177 96559
rect 61255 96513 61301 96559
rect 61379 96513 61425 96559
rect 61503 96513 61549 96559
rect 61627 96513 61673 96559
rect 61751 96513 61797 96559
rect 61875 96513 61921 96559
rect 61999 96513 62045 96559
rect 62123 96513 62169 96559
rect 62247 96513 62293 96559
rect 62371 96513 62417 96559
rect 62495 96513 62541 96559
rect 62619 96513 62665 96559
rect 62743 96513 62789 96559
rect 62867 96513 62913 96559
rect 62991 96513 63037 96559
rect 63115 96513 63161 96559
rect 63239 96513 63285 96559
rect 63363 96513 63409 96559
rect 63487 96513 63533 96559
rect 63611 96513 63657 96559
rect 63735 96513 63781 96559
rect 63859 96513 63905 96559
rect 63983 96513 64029 96559
rect 64107 96513 64153 96559
rect 64231 96513 64277 96559
rect 64355 96513 64401 96559
rect 64479 96513 64525 96559
rect 64603 96513 64649 96559
rect 64727 96513 64773 96559
rect 64851 96513 64897 96559
rect 64975 96513 65021 96559
rect 65099 96513 65145 96559
rect 65223 96513 65269 96559
rect 65347 96513 65393 96559
rect 65471 96513 65517 96559
rect 65595 96513 65641 96559
rect 65719 96513 65765 96559
rect 65843 96513 65889 96559
rect 65967 96513 66013 96559
rect 66091 96513 66137 96559
rect 66215 96513 66261 96559
rect 66339 96513 66385 96559
rect 66463 96513 66509 96559
rect 66587 96513 66633 96559
rect 66711 96513 66757 96559
rect 66835 96513 66881 96559
rect 66959 96513 67005 96559
rect 67083 96513 67129 96559
rect 67207 96513 67253 96559
rect 67331 96513 67377 96559
rect 67455 96513 67501 96559
rect 67579 96513 67625 96559
rect 67703 96513 67749 96559
rect 67827 96513 67873 96559
rect 67951 96513 67997 96559
rect 68075 96513 68121 96559
rect 68199 96513 68245 96559
rect 68323 96513 68369 96559
rect 68447 96513 68493 96559
rect 68571 96513 68617 96559
rect 68695 96513 68741 96559
rect 68819 96513 68865 96559
rect 68943 96513 68989 96559
rect 69067 96513 69113 96559
rect 69191 96513 69237 96559
rect 69315 96513 69361 96559
rect 69439 96513 69485 96559
rect 69563 96513 69609 96559
rect 69687 96513 69733 96559
rect 69811 96513 69857 96559
rect 69935 96513 69981 96559
rect 70059 96513 70105 96559
rect 70183 96513 70229 96559
rect 70307 96513 70353 96559
rect 70431 96513 70477 96559
rect 70555 96513 70601 96559
rect 70679 96513 70725 96559
rect 70803 96513 70849 96559
rect 70927 96513 70973 96559
rect 71051 96513 71097 96559
rect 71175 96513 71221 96559
rect 71299 96513 71345 96559
rect 71423 96513 71469 96559
rect 71547 96513 71593 96559
rect 71671 96513 71717 96559
rect 71795 96513 71841 96559
rect 71919 96513 71965 96559
rect 72043 96513 72089 96559
rect 72167 96513 72213 96559
rect 72291 96513 72337 96559
rect 72415 96513 72461 96559
rect 72539 96513 72585 96559
rect 72663 96513 72709 96559
rect 72787 96513 72833 96559
rect 72911 96513 72957 96559
rect 73035 96513 73081 96559
rect 73159 96513 73205 96559
rect 73283 96513 73329 96559
rect 73407 96513 73453 96559
rect 73531 96513 73577 96559
rect 73655 96513 73701 96559
rect 73779 96513 73825 96559
rect 73903 96513 73949 96559
rect 74027 96513 74073 96559
rect 74151 96513 74197 96559
rect 74275 96513 74321 96559
rect 74399 96513 74445 96559
rect 74523 96513 74569 96559
rect 74647 96513 74693 96559
rect 74771 96513 74817 96559
rect 74895 96513 74941 96559
rect 75019 96513 75065 96559
rect 75143 96513 75189 96559
rect 75267 96513 75313 96559
rect 75391 96513 75437 96559
rect 75515 96513 75561 96559
rect 75639 96513 75685 96559
rect 75763 96513 75809 96559
rect 75887 96513 75933 96559
rect 76011 96513 76057 96559
rect 76135 96513 76181 96559
rect 76259 96513 76305 96559
rect 76383 96513 76429 96559
rect 76507 96513 76553 96559
rect 76631 96513 76677 96559
rect 76755 96513 76801 96559
rect 76879 96513 76925 96559
rect 77003 96513 77049 96559
rect 77127 96513 77173 96559
rect 77251 96513 77297 96559
rect 77375 96513 77421 96559
rect 77499 96513 77545 96559
rect 77623 96513 77669 96559
rect 77747 96513 77793 96559
rect 77871 96513 77917 96559
rect 77995 96513 78041 96559
rect 78119 96513 78165 96559
rect 78243 96513 78289 96559
rect 78367 96513 78413 96559
rect 78491 96513 78537 96559
rect 78615 96513 78661 96559
rect 78739 96513 78785 96559
rect 78863 96513 78909 96559
rect 78987 96513 79033 96559
rect 79111 96513 79157 96559
rect 79235 96513 79281 96559
rect 79359 96513 79405 96559
rect 79483 96513 79529 96559
rect 79607 96513 79653 96559
rect 79731 96513 79777 96559
rect 79855 96513 79901 96559
rect 79979 96513 80025 96559
rect 80103 96513 80149 96559
rect 80227 96513 80273 96559
rect 80351 96513 80397 96559
rect 80475 96513 80521 96559
rect 80599 96513 80645 96559
rect 80723 96513 80769 96559
rect 80847 96513 80893 96559
rect 80971 96513 81017 96559
rect 81095 96513 81141 96559
rect 81219 96513 81265 96559
rect 81343 96513 81389 96559
rect 81467 96513 81513 96559
rect 81591 96513 81637 96559
rect 81715 96513 81761 96559
rect 81839 96513 81885 96559
rect 81963 96513 82009 96559
rect 82087 96513 82133 96559
rect 82211 96513 82257 96559
rect 82335 96513 82381 96559
rect 82459 96513 82505 96559
rect 82583 96513 82629 96559
rect 82707 96513 82753 96559
rect 82831 96513 82877 96559
rect 82955 96513 83001 96559
rect 83079 96513 83125 96559
rect 83203 96513 83249 96559
rect 83327 96513 83373 96559
rect 83451 96513 83497 96559
rect 83575 96513 83621 96559
rect 83699 96513 83745 96559
rect 83823 96513 83869 96559
rect 83947 96513 83993 96559
rect 84071 96513 84117 96559
rect 84195 96513 84241 96559
rect 84319 96513 84365 96559
rect 84443 96513 84489 96559
rect 84567 96513 84613 96559
rect 84691 96513 84737 96559
rect 84815 96513 84861 96559
rect 84939 96513 84985 96559
rect 85063 96513 85109 96559
rect 85187 96513 85233 96559
rect 85311 96513 85357 96559
rect 85435 96513 85481 96559
rect 85559 96513 85605 96559
rect 85683 96513 85729 96559
rect 85807 96513 85853 96559
rect 85931 96513 85977 96559
rect 371 96389 417 96435
rect 495 96389 541 96435
rect 619 96389 665 96435
rect 743 96389 789 96435
rect 867 96389 913 96435
rect 991 96389 1037 96435
rect 1115 96389 1161 96435
rect 1239 96389 1285 96435
rect 1363 96389 1409 96435
rect 1487 96389 1533 96435
rect 1611 96389 1657 96435
rect 1735 96389 1781 96435
rect 1859 96389 1905 96435
rect 1983 96389 2029 96435
rect 2107 96389 2153 96435
rect 2231 96389 2277 96435
rect 2355 96389 2401 96435
rect 2479 96389 2525 96435
rect 2603 96389 2649 96435
rect 2727 96389 2773 96435
rect 2851 96389 2897 96435
rect 2975 96389 3021 96435
rect 3099 96389 3145 96435
rect 3223 96389 3269 96435
rect 3347 96389 3393 96435
rect 3471 96389 3517 96435
rect 3595 96389 3641 96435
rect 3719 96389 3765 96435
rect 3843 96389 3889 96435
rect 3967 96389 4013 96435
rect 4091 96389 4137 96435
rect 4215 96389 4261 96435
rect 4339 96389 4385 96435
rect 4463 96389 4509 96435
rect 4587 96389 4633 96435
rect 4711 96389 4757 96435
rect 4835 96389 4881 96435
rect 4959 96389 5005 96435
rect 5083 96389 5129 96435
rect 5207 96389 5253 96435
rect 5331 96389 5377 96435
rect 5455 96389 5501 96435
rect 5579 96389 5625 96435
rect 5703 96389 5749 96435
rect 5827 96389 5873 96435
rect 5951 96389 5997 96435
rect 6075 96389 6121 96435
rect 6199 96389 6245 96435
rect 6323 96389 6369 96435
rect 6447 96389 6493 96435
rect 6571 96389 6617 96435
rect 6695 96389 6741 96435
rect 6819 96389 6865 96435
rect 6943 96389 6989 96435
rect 7067 96389 7113 96435
rect 7191 96389 7237 96435
rect 7315 96389 7361 96435
rect 7439 96389 7485 96435
rect 7563 96389 7609 96435
rect 7687 96389 7733 96435
rect 7811 96389 7857 96435
rect 7935 96389 7981 96435
rect 8059 96389 8105 96435
rect 8183 96389 8229 96435
rect 8307 96389 8353 96435
rect 8431 96389 8477 96435
rect 8555 96389 8601 96435
rect 8679 96389 8725 96435
rect 8803 96389 8849 96435
rect 8927 96389 8973 96435
rect 9051 96389 9097 96435
rect 9175 96389 9221 96435
rect 9299 96389 9345 96435
rect 9423 96389 9469 96435
rect 9547 96389 9593 96435
rect 9671 96389 9717 96435
rect 9795 96389 9841 96435
rect 9919 96389 9965 96435
rect 10043 96389 10089 96435
rect 10167 96389 10213 96435
rect 10291 96389 10337 96435
rect 10415 96389 10461 96435
rect 10539 96389 10585 96435
rect 10663 96389 10709 96435
rect 10787 96389 10833 96435
rect 10911 96389 10957 96435
rect 11035 96389 11081 96435
rect 11159 96389 11205 96435
rect 11283 96389 11329 96435
rect 11407 96389 11453 96435
rect 11531 96389 11577 96435
rect 11655 96389 11701 96435
rect 11779 96389 11825 96435
rect 11903 96389 11949 96435
rect 12027 96389 12073 96435
rect 12151 96389 12197 96435
rect 12275 96389 12321 96435
rect 12399 96389 12445 96435
rect 12523 96389 12569 96435
rect 12647 96389 12693 96435
rect 12771 96389 12817 96435
rect 12895 96389 12941 96435
rect 13019 96389 13065 96435
rect 13143 96389 13189 96435
rect 13267 96389 13313 96435
rect 13391 96389 13437 96435
rect 13515 96389 13561 96435
rect 13639 96389 13685 96435
rect 13763 96389 13809 96435
rect 13887 96389 13933 96435
rect 14011 96389 14057 96435
rect 14135 96389 14181 96435
rect 14259 96389 14305 96435
rect 14383 96389 14429 96435
rect 14507 96389 14553 96435
rect 14631 96389 14677 96435
rect 14755 96389 14801 96435
rect 14879 96389 14925 96435
rect 15003 96389 15049 96435
rect 15127 96389 15173 96435
rect 15251 96389 15297 96435
rect 15375 96389 15421 96435
rect 15499 96389 15545 96435
rect 15623 96389 15669 96435
rect 15747 96389 15793 96435
rect 15871 96389 15917 96435
rect 15995 96389 16041 96435
rect 16119 96389 16165 96435
rect 16243 96389 16289 96435
rect 16367 96389 16413 96435
rect 16491 96389 16537 96435
rect 16615 96389 16661 96435
rect 16739 96389 16785 96435
rect 16863 96389 16909 96435
rect 16987 96389 17033 96435
rect 17111 96389 17157 96435
rect 17235 96389 17281 96435
rect 17359 96389 17405 96435
rect 17483 96389 17529 96435
rect 17607 96389 17653 96435
rect 17731 96389 17777 96435
rect 17855 96389 17901 96435
rect 17979 96389 18025 96435
rect 18103 96389 18149 96435
rect 18227 96389 18273 96435
rect 18351 96389 18397 96435
rect 18475 96389 18521 96435
rect 18599 96389 18645 96435
rect 18723 96389 18769 96435
rect 18847 96389 18893 96435
rect 18971 96389 19017 96435
rect 19095 96389 19141 96435
rect 19219 96389 19265 96435
rect 19343 96389 19389 96435
rect 19467 96389 19513 96435
rect 19591 96389 19637 96435
rect 19715 96389 19761 96435
rect 19839 96389 19885 96435
rect 19963 96389 20009 96435
rect 20087 96389 20133 96435
rect 20211 96389 20257 96435
rect 20335 96389 20381 96435
rect 20459 96389 20505 96435
rect 20583 96389 20629 96435
rect 20707 96389 20753 96435
rect 20831 96389 20877 96435
rect 20955 96389 21001 96435
rect 21079 96389 21125 96435
rect 21203 96389 21249 96435
rect 21327 96389 21373 96435
rect 21451 96389 21497 96435
rect 21575 96389 21621 96435
rect 21699 96389 21745 96435
rect 21823 96389 21869 96435
rect 21947 96389 21993 96435
rect 22071 96389 22117 96435
rect 22195 96389 22241 96435
rect 22319 96389 22365 96435
rect 22443 96389 22489 96435
rect 22567 96389 22613 96435
rect 22691 96389 22737 96435
rect 22815 96389 22861 96435
rect 22939 96389 22985 96435
rect 23063 96389 23109 96435
rect 23187 96389 23233 96435
rect 23311 96389 23357 96435
rect 23435 96389 23481 96435
rect 23559 96389 23605 96435
rect 23683 96389 23729 96435
rect 23807 96389 23853 96435
rect 23931 96389 23977 96435
rect 24055 96389 24101 96435
rect 24179 96389 24225 96435
rect 24303 96389 24349 96435
rect 24427 96389 24473 96435
rect 24551 96389 24597 96435
rect 24675 96389 24721 96435
rect 24799 96389 24845 96435
rect 24923 96389 24969 96435
rect 25047 96389 25093 96435
rect 25171 96389 25217 96435
rect 25295 96389 25341 96435
rect 25419 96389 25465 96435
rect 25543 96389 25589 96435
rect 25667 96389 25713 96435
rect 25791 96389 25837 96435
rect 25915 96389 25961 96435
rect 26039 96389 26085 96435
rect 26163 96389 26209 96435
rect 26287 96389 26333 96435
rect 26411 96389 26457 96435
rect 26535 96389 26581 96435
rect 26659 96389 26705 96435
rect 26783 96389 26829 96435
rect 26907 96389 26953 96435
rect 27031 96389 27077 96435
rect 27155 96389 27201 96435
rect 27279 96389 27325 96435
rect 27403 96389 27449 96435
rect 27527 96389 27573 96435
rect 27651 96389 27697 96435
rect 27775 96389 27821 96435
rect 27899 96389 27945 96435
rect 28023 96389 28069 96435
rect 28147 96389 28193 96435
rect 28271 96389 28317 96435
rect 28395 96389 28441 96435
rect 28519 96389 28565 96435
rect 28643 96389 28689 96435
rect 28767 96389 28813 96435
rect 28891 96389 28937 96435
rect 29015 96389 29061 96435
rect 29139 96389 29185 96435
rect 29263 96389 29309 96435
rect 29387 96389 29433 96435
rect 29511 96389 29557 96435
rect 29635 96389 29681 96435
rect 29759 96389 29805 96435
rect 29883 96389 29929 96435
rect 30007 96389 30053 96435
rect 30131 96389 30177 96435
rect 30255 96389 30301 96435
rect 30379 96389 30425 96435
rect 30503 96389 30549 96435
rect 30627 96389 30673 96435
rect 30751 96389 30797 96435
rect 30875 96389 30921 96435
rect 30999 96389 31045 96435
rect 31123 96389 31169 96435
rect 31247 96389 31293 96435
rect 31371 96389 31417 96435
rect 31495 96389 31541 96435
rect 31619 96389 31665 96435
rect 31743 96389 31789 96435
rect 31867 96389 31913 96435
rect 31991 96389 32037 96435
rect 32115 96389 32161 96435
rect 32239 96389 32285 96435
rect 32363 96389 32409 96435
rect 32487 96389 32533 96435
rect 32611 96389 32657 96435
rect 32735 96389 32781 96435
rect 32859 96389 32905 96435
rect 32983 96389 33029 96435
rect 33107 96389 33153 96435
rect 33231 96389 33277 96435
rect 33355 96389 33401 96435
rect 33479 96389 33525 96435
rect 33603 96389 33649 96435
rect 33727 96389 33773 96435
rect 33851 96389 33897 96435
rect 33975 96389 34021 96435
rect 34099 96389 34145 96435
rect 34223 96389 34269 96435
rect 34347 96389 34393 96435
rect 34471 96389 34517 96435
rect 34595 96389 34641 96435
rect 34719 96389 34765 96435
rect 34843 96389 34889 96435
rect 34967 96389 35013 96435
rect 35091 96389 35137 96435
rect 35215 96389 35261 96435
rect 35339 96389 35385 96435
rect 35463 96389 35509 96435
rect 35587 96389 35633 96435
rect 35711 96389 35757 96435
rect 35835 96389 35881 96435
rect 35959 96389 36005 96435
rect 36083 96389 36129 96435
rect 36207 96389 36253 96435
rect 36331 96389 36377 96435
rect 36455 96389 36501 96435
rect 36579 96389 36625 96435
rect 36703 96389 36749 96435
rect 36827 96389 36873 96435
rect 36951 96389 36997 96435
rect 37075 96389 37121 96435
rect 37199 96389 37245 96435
rect 37323 96389 37369 96435
rect 37447 96389 37493 96435
rect 37571 96389 37617 96435
rect 37695 96389 37741 96435
rect 37819 96389 37865 96435
rect 37943 96389 37989 96435
rect 38067 96389 38113 96435
rect 38191 96389 38237 96435
rect 38315 96389 38361 96435
rect 38439 96389 38485 96435
rect 38563 96389 38609 96435
rect 38687 96389 38733 96435
rect 38811 96389 38857 96435
rect 38935 96389 38981 96435
rect 39059 96389 39105 96435
rect 39183 96389 39229 96435
rect 39307 96389 39353 96435
rect 39431 96389 39477 96435
rect 39555 96389 39601 96435
rect 39679 96389 39725 96435
rect 39803 96389 39849 96435
rect 39927 96389 39973 96435
rect 40051 96389 40097 96435
rect 40175 96389 40221 96435
rect 40299 96389 40345 96435
rect 40423 96389 40469 96435
rect 40547 96389 40593 96435
rect 40671 96389 40717 96435
rect 40795 96389 40841 96435
rect 40919 96389 40965 96435
rect 41043 96389 41089 96435
rect 41167 96389 41213 96435
rect 41291 96389 41337 96435
rect 41415 96389 41461 96435
rect 41539 96389 41585 96435
rect 41663 96389 41709 96435
rect 41787 96389 41833 96435
rect 41911 96389 41957 96435
rect 42035 96389 42081 96435
rect 42159 96389 42205 96435
rect 42283 96389 42329 96435
rect 42407 96389 42453 96435
rect 42531 96389 42577 96435
rect 42655 96389 42701 96435
rect 42779 96389 42825 96435
rect 42903 96389 42949 96435
rect 43027 96389 43073 96435
rect 43151 96389 43197 96435
rect 43275 96389 43321 96435
rect 43399 96389 43445 96435
rect 43523 96389 43569 96435
rect 43647 96389 43693 96435
rect 43771 96389 43817 96435
rect 43895 96389 43941 96435
rect 44019 96389 44065 96435
rect 44143 96389 44189 96435
rect 44267 96389 44313 96435
rect 44391 96389 44437 96435
rect 44515 96389 44561 96435
rect 44639 96389 44685 96435
rect 44763 96389 44809 96435
rect 44887 96389 44933 96435
rect 45011 96389 45057 96435
rect 45135 96389 45181 96435
rect 45259 96389 45305 96435
rect 45383 96389 45429 96435
rect 45507 96389 45553 96435
rect 45631 96389 45677 96435
rect 45755 96389 45801 96435
rect 45879 96389 45925 96435
rect 46003 96389 46049 96435
rect 46127 96389 46173 96435
rect 46251 96389 46297 96435
rect 46375 96389 46421 96435
rect 46499 96389 46545 96435
rect 46623 96389 46669 96435
rect 46747 96389 46793 96435
rect 46871 96389 46917 96435
rect 46995 96389 47041 96435
rect 47119 96389 47165 96435
rect 47243 96389 47289 96435
rect 47367 96389 47413 96435
rect 47491 96389 47537 96435
rect 47615 96389 47661 96435
rect 47739 96389 47785 96435
rect 47863 96389 47909 96435
rect 47987 96389 48033 96435
rect 48111 96389 48157 96435
rect 48235 96389 48281 96435
rect 48359 96389 48405 96435
rect 48483 96389 48529 96435
rect 48607 96389 48653 96435
rect 48731 96389 48777 96435
rect 48855 96389 48901 96435
rect 48979 96389 49025 96435
rect 49103 96389 49149 96435
rect 49227 96389 49273 96435
rect 49351 96389 49397 96435
rect 49475 96389 49521 96435
rect 49599 96389 49645 96435
rect 49723 96389 49769 96435
rect 49847 96389 49893 96435
rect 49971 96389 50017 96435
rect 50095 96389 50141 96435
rect 50219 96389 50265 96435
rect 50343 96389 50389 96435
rect 50467 96389 50513 96435
rect 50591 96389 50637 96435
rect 50715 96389 50761 96435
rect 50839 96389 50885 96435
rect 50963 96389 51009 96435
rect 51087 96389 51133 96435
rect 51211 96389 51257 96435
rect 51335 96389 51381 96435
rect 51459 96389 51505 96435
rect 51583 96389 51629 96435
rect 51707 96389 51753 96435
rect 51831 96389 51877 96435
rect 51955 96389 52001 96435
rect 52079 96389 52125 96435
rect 52203 96389 52249 96435
rect 52327 96389 52373 96435
rect 52451 96389 52497 96435
rect 52575 96389 52621 96435
rect 52699 96389 52745 96435
rect 52823 96389 52869 96435
rect 52947 96389 52993 96435
rect 53071 96389 53117 96435
rect 53195 96389 53241 96435
rect 53319 96389 53365 96435
rect 53443 96389 53489 96435
rect 53567 96389 53613 96435
rect 53691 96389 53737 96435
rect 53815 96389 53861 96435
rect 53939 96389 53985 96435
rect 54063 96389 54109 96435
rect 54187 96389 54233 96435
rect 54311 96389 54357 96435
rect 54435 96389 54481 96435
rect 54559 96389 54605 96435
rect 54683 96389 54729 96435
rect 54807 96389 54853 96435
rect 54931 96389 54977 96435
rect 55055 96389 55101 96435
rect 55179 96389 55225 96435
rect 55303 96389 55349 96435
rect 55427 96389 55473 96435
rect 55551 96389 55597 96435
rect 55675 96389 55721 96435
rect 55799 96389 55845 96435
rect 55923 96389 55969 96435
rect 56047 96389 56093 96435
rect 56171 96389 56217 96435
rect 56295 96389 56341 96435
rect 56419 96389 56465 96435
rect 56543 96389 56589 96435
rect 56667 96389 56713 96435
rect 56791 96389 56837 96435
rect 56915 96389 56961 96435
rect 57039 96389 57085 96435
rect 57163 96389 57209 96435
rect 57287 96389 57333 96435
rect 57411 96389 57457 96435
rect 57535 96389 57581 96435
rect 57659 96389 57705 96435
rect 57783 96389 57829 96435
rect 57907 96389 57953 96435
rect 58031 96389 58077 96435
rect 58155 96389 58201 96435
rect 58279 96389 58325 96435
rect 58403 96389 58449 96435
rect 58527 96389 58573 96435
rect 58651 96389 58697 96435
rect 58775 96389 58821 96435
rect 58899 96389 58945 96435
rect 59023 96389 59069 96435
rect 59147 96389 59193 96435
rect 59271 96389 59317 96435
rect 59395 96389 59441 96435
rect 59519 96389 59565 96435
rect 59643 96389 59689 96435
rect 59767 96389 59813 96435
rect 59891 96389 59937 96435
rect 60015 96389 60061 96435
rect 60139 96389 60185 96435
rect 60263 96389 60309 96435
rect 60387 96389 60433 96435
rect 60511 96389 60557 96435
rect 60635 96389 60681 96435
rect 60759 96389 60805 96435
rect 60883 96389 60929 96435
rect 61007 96389 61053 96435
rect 61131 96389 61177 96435
rect 61255 96389 61301 96435
rect 61379 96389 61425 96435
rect 61503 96389 61549 96435
rect 61627 96389 61673 96435
rect 61751 96389 61797 96435
rect 61875 96389 61921 96435
rect 61999 96389 62045 96435
rect 62123 96389 62169 96435
rect 62247 96389 62293 96435
rect 62371 96389 62417 96435
rect 62495 96389 62541 96435
rect 62619 96389 62665 96435
rect 62743 96389 62789 96435
rect 62867 96389 62913 96435
rect 62991 96389 63037 96435
rect 63115 96389 63161 96435
rect 63239 96389 63285 96435
rect 63363 96389 63409 96435
rect 63487 96389 63533 96435
rect 63611 96389 63657 96435
rect 63735 96389 63781 96435
rect 63859 96389 63905 96435
rect 63983 96389 64029 96435
rect 64107 96389 64153 96435
rect 64231 96389 64277 96435
rect 64355 96389 64401 96435
rect 64479 96389 64525 96435
rect 64603 96389 64649 96435
rect 64727 96389 64773 96435
rect 64851 96389 64897 96435
rect 64975 96389 65021 96435
rect 65099 96389 65145 96435
rect 65223 96389 65269 96435
rect 65347 96389 65393 96435
rect 65471 96389 65517 96435
rect 65595 96389 65641 96435
rect 65719 96389 65765 96435
rect 65843 96389 65889 96435
rect 65967 96389 66013 96435
rect 66091 96389 66137 96435
rect 66215 96389 66261 96435
rect 66339 96389 66385 96435
rect 66463 96389 66509 96435
rect 66587 96389 66633 96435
rect 66711 96389 66757 96435
rect 66835 96389 66881 96435
rect 66959 96389 67005 96435
rect 67083 96389 67129 96435
rect 67207 96389 67253 96435
rect 67331 96389 67377 96435
rect 67455 96389 67501 96435
rect 67579 96389 67625 96435
rect 67703 96389 67749 96435
rect 67827 96389 67873 96435
rect 67951 96389 67997 96435
rect 68075 96389 68121 96435
rect 68199 96389 68245 96435
rect 68323 96389 68369 96435
rect 68447 96389 68493 96435
rect 68571 96389 68617 96435
rect 68695 96389 68741 96435
rect 68819 96389 68865 96435
rect 68943 96389 68989 96435
rect 69067 96389 69113 96435
rect 69191 96389 69237 96435
rect 69315 96389 69361 96435
rect 69439 96389 69485 96435
rect 69563 96389 69609 96435
rect 69687 96389 69733 96435
rect 69811 96389 69857 96435
rect 69935 96389 69981 96435
rect 70059 96389 70105 96435
rect 70183 96389 70229 96435
rect 70307 96389 70353 96435
rect 70431 96389 70477 96435
rect 70555 96389 70601 96435
rect 70679 96389 70725 96435
rect 70803 96389 70849 96435
rect 70927 96389 70973 96435
rect 71051 96389 71097 96435
rect 71175 96389 71221 96435
rect 71299 96389 71345 96435
rect 71423 96389 71469 96435
rect 71547 96389 71593 96435
rect 71671 96389 71717 96435
rect 71795 96389 71841 96435
rect 71919 96389 71965 96435
rect 72043 96389 72089 96435
rect 72167 96389 72213 96435
rect 72291 96389 72337 96435
rect 72415 96389 72461 96435
rect 72539 96389 72585 96435
rect 72663 96389 72709 96435
rect 72787 96389 72833 96435
rect 72911 96389 72957 96435
rect 73035 96389 73081 96435
rect 73159 96389 73205 96435
rect 73283 96389 73329 96435
rect 73407 96389 73453 96435
rect 73531 96389 73577 96435
rect 73655 96389 73701 96435
rect 73779 96389 73825 96435
rect 73903 96389 73949 96435
rect 74027 96389 74073 96435
rect 74151 96389 74197 96435
rect 74275 96389 74321 96435
rect 74399 96389 74445 96435
rect 74523 96389 74569 96435
rect 74647 96389 74693 96435
rect 74771 96389 74817 96435
rect 74895 96389 74941 96435
rect 75019 96389 75065 96435
rect 75143 96389 75189 96435
rect 75267 96389 75313 96435
rect 75391 96389 75437 96435
rect 75515 96389 75561 96435
rect 75639 96389 75685 96435
rect 75763 96389 75809 96435
rect 75887 96389 75933 96435
rect 76011 96389 76057 96435
rect 76135 96389 76181 96435
rect 76259 96389 76305 96435
rect 76383 96389 76429 96435
rect 76507 96389 76553 96435
rect 76631 96389 76677 96435
rect 76755 96389 76801 96435
rect 76879 96389 76925 96435
rect 77003 96389 77049 96435
rect 77127 96389 77173 96435
rect 77251 96389 77297 96435
rect 77375 96389 77421 96435
rect 77499 96389 77545 96435
rect 77623 96389 77669 96435
rect 77747 96389 77793 96435
rect 77871 96389 77917 96435
rect 77995 96389 78041 96435
rect 78119 96389 78165 96435
rect 78243 96389 78289 96435
rect 78367 96389 78413 96435
rect 78491 96389 78537 96435
rect 78615 96389 78661 96435
rect 78739 96389 78785 96435
rect 78863 96389 78909 96435
rect 78987 96389 79033 96435
rect 79111 96389 79157 96435
rect 79235 96389 79281 96435
rect 79359 96389 79405 96435
rect 79483 96389 79529 96435
rect 79607 96389 79653 96435
rect 79731 96389 79777 96435
rect 79855 96389 79901 96435
rect 79979 96389 80025 96435
rect 80103 96389 80149 96435
rect 80227 96389 80273 96435
rect 80351 96389 80397 96435
rect 80475 96389 80521 96435
rect 80599 96389 80645 96435
rect 80723 96389 80769 96435
rect 80847 96389 80893 96435
rect 80971 96389 81017 96435
rect 81095 96389 81141 96435
rect 81219 96389 81265 96435
rect 81343 96389 81389 96435
rect 81467 96389 81513 96435
rect 81591 96389 81637 96435
rect 81715 96389 81761 96435
rect 81839 96389 81885 96435
rect 81963 96389 82009 96435
rect 82087 96389 82133 96435
rect 82211 96389 82257 96435
rect 82335 96389 82381 96435
rect 82459 96389 82505 96435
rect 82583 96389 82629 96435
rect 82707 96389 82753 96435
rect 82831 96389 82877 96435
rect 82955 96389 83001 96435
rect 83079 96389 83125 96435
rect 83203 96389 83249 96435
rect 83327 96389 83373 96435
rect 83451 96389 83497 96435
rect 83575 96389 83621 96435
rect 83699 96389 83745 96435
rect 83823 96389 83869 96435
rect 83947 96389 83993 96435
rect 84071 96389 84117 96435
rect 84195 96389 84241 96435
rect 84319 96389 84365 96435
rect 84443 96389 84489 96435
rect 84567 96389 84613 96435
rect 84691 96389 84737 96435
rect 84815 96389 84861 96435
rect 84939 96389 84985 96435
rect 85063 96389 85109 96435
rect 85187 96389 85233 96435
rect 85311 96389 85357 96435
rect 85435 96389 85481 96435
rect 85559 96389 85605 96435
rect 85683 96389 85729 96435
rect 85807 96389 85853 96435
rect 85931 96389 85977 96435
rect 371 96265 417 96311
rect 495 96265 541 96311
rect 619 96265 665 96311
rect 743 96265 789 96311
rect 867 96265 913 96311
rect 991 96265 1037 96311
rect 1115 96265 1161 96311
rect 1239 96265 1285 96311
rect 1363 96265 1409 96311
rect 1487 96265 1533 96311
rect 1611 96265 1657 96311
rect 1735 96265 1781 96311
rect 1859 96265 1905 96311
rect 1983 96265 2029 96311
rect 2107 96265 2153 96311
rect 2231 96265 2277 96311
rect 2355 96265 2401 96311
rect 2479 96265 2525 96311
rect 2603 96265 2649 96311
rect 2727 96265 2773 96311
rect 2851 96265 2897 96311
rect 2975 96265 3021 96311
rect 3099 96265 3145 96311
rect 3223 96265 3269 96311
rect 3347 96265 3393 96311
rect 3471 96265 3517 96311
rect 3595 96265 3641 96311
rect 3719 96265 3765 96311
rect 3843 96265 3889 96311
rect 3967 96265 4013 96311
rect 4091 96265 4137 96311
rect 4215 96265 4261 96311
rect 4339 96265 4385 96311
rect 4463 96265 4509 96311
rect 4587 96265 4633 96311
rect 4711 96265 4757 96311
rect 4835 96265 4881 96311
rect 4959 96265 5005 96311
rect 5083 96265 5129 96311
rect 5207 96265 5253 96311
rect 5331 96265 5377 96311
rect 5455 96265 5501 96311
rect 5579 96265 5625 96311
rect 5703 96265 5749 96311
rect 5827 96265 5873 96311
rect 5951 96265 5997 96311
rect 6075 96265 6121 96311
rect 6199 96265 6245 96311
rect 6323 96265 6369 96311
rect 6447 96265 6493 96311
rect 6571 96265 6617 96311
rect 6695 96265 6741 96311
rect 6819 96265 6865 96311
rect 6943 96265 6989 96311
rect 7067 96265 7113 96311
rect 7191 96265 7237 96311
rect 7315 96265 7361 96311
rect 7439 96265 7485 96311
rect 7563 96265 7609 96311
rect 7687 96265 7733 96311
rect 7811 96265 7857 96311
rect 7935 96265 7981 96311
rect 8059 96265 8105 96311
rect 8183 96265 8229 96311
rect 8307 96265 8353 96311
rect 8431 96265 8477 96311
rect 8555 96265 8601 96311
rect 8679 96265 8725 96311
rect 8803 96265 8849 96311
rect 8927 96265 8973 96311
rect 9051 96265 9097 96311
rect 9175 96265 9221 96311
rect 9299 96265 9345 96311
rect 9423 96265 9469 96311
rect 9547 96265 9593 96311
rect 9671 96265 9717 96311
rect 9795 96265 9841 96311
rect 9919 96265 9965 96311
rect 10043 96265 10089 96311
rect 10167 96265 10213 96311
rect 10291 96265 10337 96311
rect 10415 96265 10461 96311
rect 10539 96265 10585 96311
rect 10663 96265 10709 96311
rect 10787 96265 10833 96311
rect 10911 96265 10957 96311
rect 11035 96265 11081 96311
rect 11159 96265 11205 96311
rect 11283 96265 11329 96311
rect 11407 96265 11453 96311
rect 11531 96265 11577 96311
rect 11655 96265 11701 96311
rect 11779 96265 11825 96311
rect 11903 96265 11949 96311
rect 12027 96265 12073 96311
rect 12151 96265 12197 96311
rect 12275 96265 12321 96311
rect 12399 96265 12445 96311
rect 12523 96265 12569 96311
rect 12647 96265 12693 96311
rect 12771 96265 12817 96311
rect 12895 96265 12941 96311
rect 13019 96265 13065 96311
rect 13143 96265 13189 96311
rect 13267 96265 13313 96311
rect 13391 96265 13437 96311
rect 13515 96265 13561 96311
rect 13639 96265 13685 96311
rect 13763 96265 13809 96311
rect 13887 96265 13933 96311
rect 14011 96265 14057 96311
rect 14135 96265 14181 96311
rect 14259 96265 14305 96311
rect 14383 96265 14429 96311
rect 14507 96265 14553 96311
rect 14631 96265 14677 96311
rect 14755 96265 14801 96311
rect 14879 96265 14925 96311
rect 15003 96265 15049 96311
rect 15127 96265 15173 96311
rect 15251 96265 15297 96311
rect 15375 96265 15421 96311
rect 15499 96265 15545 96311
rect 15623 96265 15669 96311
rect 15747 96265 15793 96311
rect 15871 96265 15917 96311
rect 15995 96265 16041 96311
rect 16119 96265 16165 96311
rect 16243 96265 16289 96311
rect 16367 96265 16413 96311
rect 16491 96265 16537 96311
rect 16615 96265 16661 96311
rect 16739 96265 16785 96311
rect 16863 96265 16909 96311
rect 16987 96265 17033 96311
rect 17111 96265 17157 96311
rect 17235 96265 17281 96311
rect 17359 96265 17405 96311
rect 17483 96265 17529 96311
rect 17607 96265 17653 96311
rect 17731 96265 17777 96311
rect 17855 96265 17901 96311
rect 17979 96265 18025 96311
rect 18103 96265 18149 96311
rect 18227 96265 18273 96311
rect 18351 96265 18397 96311
rect 18475 96265 18521 96311
rect 18599 96265 18645 96311
rect 18723 96265 18769 96311
rect 18847 96265 18893 96311
rect 18971 96265 19017 96311
rect 19095 96265 19141 96311
rect 19219 96265 19265 96311
rect 19343 96265 19389 96311
rect 19467 96265 19513 96311
rect 19591 96265 19637 96311
rect 19715 96265 19761 96311
rect 19839 96265 19885 96311
rect 19963 96265 20009 96311
rect 20087 96265 20133 96311
rect 20211 96265 20257 96311
rect 20335 96265 20381 96311
rect 20459 96265 20505 96311
rect 20583 96265 20629 96311
rect 20707 96265 20753 96311
rect 20831 96265 20877 96311
rect 20955 96265 21001 96311
rect 21079 96265 21125 96311
rect 21203 96265 21249 96311
rect 21327 96265 21373 96311
rect 21451 96265 21497 96311
rect 21575 96265 21621 96311
rect 21699 96265 21745 96311
rect 21823 96265 21869 96311
rect 21947 96265 21993 96311
rect 22071 96265 22117 96311
rect 22195 96265 22241 96311
rect 22319 96265 22365 96311
rect 22443 96265 22489 96311
rect 22567 96265 22613 96311
rect 22691 96265 22737 96311
rect 22815 96265 22861 96311
rect 22939 96265 22985 96311
rect 23063 96265 23109 96311
rect 23187 96265 23233 96311
rect 23311 96265 23357 96311
rect 23435 96265 23481 96311
rect 23559 96265 23605 96311
rect 23683 96265 23729 96311
rect 23807 96265 23853 96311
rect 23931 96265 23977 96311
rect 24055 96265 24101 96311
rect 24179 96265 24225 96311
rect 24303 96265 24349 96311
rect 24427 96265 24473 96311
rect 24551 96265 24597 96311
rect 24675 96265 24721 96311
rect 24799 96265 24845 96311
rect 24923 96265 24969 96311
rect 25047 96265 25093 96311
rect 25171 96265 25217 96311
rect 25295 96265 25341 96311
rect 25419 96265 25465 96311
rect 25543 96265 25589 96311
rect 25667 96265 25713 96311
rect 25791 96265 25837 96311
rect 25915 96265 25961 96311
rect 26039 96265 26085 96311
rect 26163 96265 26209 96311
rect 26287 96265 26333 96311
rect 26411 96265 26457 96311
rect 26535 96265 26581 96311
rect 26659 96265 26705 96311
rect 26783 96265 26829 96311
rect 26907 96265 26953 96311
rect 27031 96265 27077 96311
rect 27155 96265 27201 96311
rect 27279 96265 27325 96311
rect 27403 96265 27449 96311
rect 27527 96265 27573 96311
rect 27651 96265 27697 96311
rect 27775 96265 27821 96311
rect 27899 96265 27945 96311
rect 28023 96265 28069 96311
rect 28147 96265 28193 96311
rect 28271 96265 28317 96311
rect 28395 96265 28441 96311
rect 28519 96265 28565 96311
rect 28643 96265 28689 96311
rect 28767 96265 28813 96311
rect 28891 96265 28937 96311
rect 29015 96265 29061 96311
rect 29139 96265 29185 96311
rect 29263 96265 29309 96311
rect 29387 96265 29433 96311
rect 29511 96265 29557 96311
rect 29635 96265 29681 96311
rect 29759 96265 29805 96311
rect 29883 96265 29929 96311
rect 30007 96265 30053 96311
rect 30131 96265 30177 96311
rect 30255 96265 30301 96311
rect 30379 96265 30425 96311
rect 30503 96265 30549 96311
rect 30627 96265 30673 96311
rect 30751 96265 30797 96311
rect 30875 96265 30921 96311
rect 30999 96265 31045 96311
rect 31123 96265 31169 96311
rect 31247 96265 31293 96311
rect 31371 96265 31417 96311
rect 31495 96265 31541 96311
rect 31619 96265 31665 96311
rect 31743 96265 31789 96311
rect 31867 96265 31913 96311
rect 31991 96265 32037 96311
rect 32115 96265 32161 96311
rect 32239 96265 32285 96311
rect 32363 96265 32409 96311
rect 32487 96265 32533 96311
rect 32611 96265 32657 96311
rect 32735 96265 32781 96311
rect 32859 96265 32905 96311
rect 32983 96265 33029 96311
rect 33107 96265 33153 96311
rect 33231 96265 33277 96311
rect 33355 96265 33401 96311
rect 33479 96265 33525 96311
rect 33603 96265 33649 96311
rect 33727 96265 33773 96311
rect 33851 96265 33897 96311
rect 33975 96265 34021 96311
rect 34099 96265 34145 96311
rect 34223 96265 34269 96311
rect 34347 96265 34393 96311
rect 34471 96265 34517 96311
rect 34595 96265 34641 96311
rect 34719 96265 34765 96311
rect 34843 96265 34889 96311
rect 34967 96265 35013 96311
rect 35091 96265 35137 96311
rect 35215 96265 35261 96311
rect 35339 96265 35385 96311
rect 35463 96265 35509 96311
rect 35587 96265 35633 96311
rect 35711 96265 35757 96311
rect 35835 96265 35881 96311
rect 35959 96265 36005 96311
rect 36083 96265 36129 96311
rect 36207 96265 36253 96311
rect 36331 96265 36377 96311
rect 36455 96265 36501 96311
rect 36579 96265 36625 96311
rect 36703 96265 36749 96311
rect 36827 96265 36873 96311
rect 36951 96265 36997 96311
rect 37075 96265 37121 96311
rect 37199 96265 37245 96311
rect 37323 96265 37369 96311
rect 37447 96265 37493 96311
rect 37571 96265 37617 96311
rect 37695 96265 37741 96311
rect 37819 96265 37865 96311
rect 37943 96265 37989 96311
rect 38067 96265 38113 96311
rect 38191 96265 38237 96311
rect 38315 96265 38361 96311
rect 38439 96265 38485 96311
rect 38563 96265 38609 96311
rect 38687 96265 38733 96311
rect 38811 96265 38857 96311
rect 38935 96265 38981 96311
rect 39059 96265 39105 96311
rect 39183 96265 39229 96311
rect 39307 96265 39353 96311
rect 39431 96265 39477 96311
rect 39555 96265 39601 96311
rect 39679 96265 39725 96311
rect 39803 96265 39849 96311
rect 39927 96265 39973 96311
rect 40051 96265 40097 96311
rect 40175 96265 40221 96311
rect 40299 96265 40345 96311
rect 40423 96265 40469 96311
rect 40547 96265 40593 96311
rect 40671 96265 40717 96311
rect 40795 96265 40841 96311
rect 40919 96265 40965 96311
rect 41043 96265 41089 96311
rect 41167 96265 41213 96311
rect 41291 96265 41337 96311
rect 41415 96265 41461 96311
rect 41539 96265 41585 96311
rect 41663 96265 41709 96311
rect 41787 96265 41833 96311
rect 41911 96265 41957 96311
rect 42035 96265 42081 96311
rect 42159 96265 42205 96311
rect 42283 96265 42329 96311
rect 42407 96265 42453 96311
rect 42531 96265 42577 96311
rect 42655 96265 42701 96311
rect 42779 96265 42825 96311
rect 42903 96265 42949 96311
rect 43027 96265 43073 96311
rect 43151 96265 43197 96311
rect 43275 96265 43321 96311
rect 43399 96265 43445 96311
rect 43523 96265 43569 96311
rect 43647 96265 43693 96311
rect 43771 96265 43817 96311
rect 43895 96265 43941 96311
rect 44019 96265 44065 96311
rect 44143 96265 44189 96311
rect 44267 96265 44313 96311
rect 44391 96265 44437 96311
rect 44515 96265 44561 96311
rect 44639 96265 44685 96311
rect 44763 96265 44809 96311
rect 44887 96265 44933 96311
rect 45011 96265 45057 96311
rect 45135 96265 45181 96311
rect 45259 96265 45305 96311
rect 45383 96265 45429 96311
rect 45507 96265 45553 96311
rect 45631 96265 45677 96311
rect 45755 96265 45801 96311
rect 45879 96265 45925 96311
rect 46003 96265 46049 96311
rect 46127 96265 46173 96311
rect 46251 96265 46297 96311
rect 46375 96265 46421 96311
rect 46499 96265 46545 96311
rect 46623 96265 46669 96311
rect 46747 96265 46793 96311
rect 46871 96265 46917 96311
rect 46995 96265 47041 96311
rect 47119 96265 47165 96311
rect 47243 96265 47289 96311
rect 47367 96265 47413 96311
rect 47491 96265 47537 96311
rect 47615 96265 47661 96311
rect 47739 96265 47785 96311
rect 47863 96265 47909 96311
rect 47987 96265 48033 96311
rect 48111 96265 48157 96311
rect 48235 96265 48281 96311
rect 48359 96265 48405 96311
rect 48483 96265 48529 96311
rect 48607 96265 48653 96311
rect 48731 96265 48777 96311
rect 48855 96265 48901 96311
rect 48979 96265 49025 96311
rect 49103 96265 49149 96311
rect 49227 96265 49273 96311
rect 49351 96265 49397 96311
rect 49475 96265 49521 96311
rect 49599 96265 49645 96311
rect 49723 96265 49769 96311
rect 49847 96265 49893 96311
rect 49971 96265 50017 96311
rect 50095 96265 50141 96311
rect 50219 96265 50265 96311
rect 50343 96265 50389 96311
rect 50467 96265 50513 96311
rect 50591 96265 50637 96311
rect 50715 96265 50761 96311
rect 50839 96265 50885 96311
rect 50963 96265 51009 96311
rect 51087 96265 51133 96311
rect 51211 96265 51257 96311
rect 51335 96265 51381 96311
rect 51459 96265 51505 96311
rect 51583 96265 51629 96311
rect 51707 96265 51753 96311
rect 51831 96265 51877 96311
rect 51955 96265 52001 96311
rect 52079 96265 52125 96311
rect 52203 96265 52249 96311
rect 52327 96265 52373 96311
rect 52451 96265 52497 96311
rect 52575 96265 52621 96311
rect 52699 96265 52745 96311
rect 52823 96265 52869 96311
rect 52947 96265 52993 96311
rect 53071 96265 53117 96311
rect 53195 96265 53241 96311
rect 53319 96265 53365 96311
rect 53443 96265 53489 96311
rect 53567 96265 53613 96311
rect 53691 96265 53737 96311
rect 53815 96265 53861 96311
rect 53939 96265 53985 96311
rect 54063 96265 54109 96311
rect 54187 96265 54233 96311
rect 54311 96265 54357 96311
rect 54435 96265 54481 96311
rect 54559 96265 54605 96311
rect 54683 96265 54729 96311
rect 54807 96265 54853 96311
rect 54931 96265 54977 96311
rect 55055 96265 55101 96311
rect 55179 96265 55225 96311
rect 55303 96265 55349 96311
rect 55427 96265 55473 96311
rect 55551 96265 55597 96311
rect 55675 96265 55721 96311
rect 55799 96265 55845 96311
rect 55923 96265 55969 96311
rect 56047 96265 56093 96311
rect 56171 96265 56217 96311
rect 56295 96265 56341 96311
rect 56419 96265 56465 96311
rect 56543 96265 56589 96311
rect 56667 96265 56713 96311
rect 56791 96265 56837 96311
rect 56915 96265 56961 96311
rect 57039 96265 57085 96311
rect 57163 96265 57209 96311
rect 57287 96265 57333 96311
rect 57411 96265 57457 96311
rect 57535 96265 57581 96311
rect 57659 96265 57705 96311
rect 57783 96265 57829 96311
rect 57907 96265 57953 96311
rect 58031 96265 58077 96311
rect 58155 96265 58201 96311
rect 58279 96265 58325 96311
rect 58403 96265 58449 96311
rect 58527 96265 58573 96311
rect 58651 96265 58697 96311
rect 58775 96265 58821 96311
rect 58899 96265 58945 96311
rect 59023 96265 59069 96311
rect 59147 96265 59193 96311
rect 59271 96265 59317 96311
rect 59395 96265 59441 96311
rect 59519 96265 59565 96311
rect 59643 96265 59689 96311
rect 59767 96265 59813 96311
rect 59891 96265 59937 96311
rect 60015 96265 60061 96311
rect 60139 96265 60185 96311
rect 60263 96265 60309 96311
rect 60387 96265 60433 96311
rect 60511 96265 60557 96311
rect 60635 96265 60681 96311
rect 60759 96265 60805 96311
rect 60883 96265 60929 96311
rect 61007 96265 61053 96311
rect 61131 96265 61177 96311
rect 61255 96265 61301 96311
rect 61379 96265 61425 96311
rect 61503 96265 61549 96311
rect 61627 96265 61673 96311
rect 61751 96265 61797 96311
rect 61875 96265 61921 96311
rect 61999 96265 62045 96311
rect 62123 96265 62169 96311
rect 62247 96265 62293 96311
rect 62371 96265 62417 96311
rect 62495 96265 62541 96311
rect 62619 96265 62665 96311
rect 62743 96265 62789 96311
rect 62867 96265 62913 96311
rect 62991 96265 63037 96311
rect 63115 96265 63161 96311
rect 63239 96265 63285 96311
rect 63363 96265 63409 96311
rect 63487 96265 63533 96311
rect 63611 96265 63657 96311
rect 63735 96265 63781 96311
rect 63859 96265 63905 96311
rect 63983 96265 64029 96311
rect 64107 96265 64153 96311
rect 64231 96265 64277 96311
rect 64355 96265 64401 96311
rect 64479 96265 64525 96311
rect 64603 96265 64649 96311
rect 64727 96265 64773 96311
rect 64851 96265 64897 96311
rect 64975 96265 65021 96311
rect 65099 96265 65145 96311
rect 65223 96265 65269 96311
rect 65347 96265 65393 96311
rect 65471 96265 65517 96311
rect 65595 96265 65641 96311
rect 65719 96265 65765 96311
rect 65843 96265 65889 96311
rect 65967 96265 66013 96311
rect 66091 96265 66137 96311
rect 66215 96265 66261 96311
rect 66339 96265 66385 96311
rect 66463 96265 66509 96311
rect 66587 96265 66633 96311
rect 66711 96265 66757 96311
rect 66835 96265 66881 96311
rect 66959 96265 67005 96311
rect 67083 96265 67129 96311
rect 67207 96265 67253 96311
rect 67331 96265 67377 96311
rect 67455 96265 67501 96311
rect 67579 96265 67625 96311
rect 67703 96265 67749 96311
rect 67827 96265 67873 96311
rect 67951 96265 67997 96311
rect 68075 96265 68121 96311
rect 68199 96265 68245 96311
rect 68323 96265 68369 96311
rect 68447 96265 68493 96311
rect 68571 96265 68617 96311
rect 68695 96265 68741 96311
rect 68819 96265 68865 96311
rect 68943 96265 68989 96311
rect 69067 96265 69113 96311
rect 69191 96265 69237 96311
rect 69315 96265 69361 96311
rect 69439 96265 69485 96311
rect 69563 96265 69609 96311
rect 69687 96265 69733 96311
rect 69811 96265 69857 96311
rect 69935 96265 69981 96311
rect 70059 96265 70105 96311
rect 70183 96265 70229 96311
rect 70307 96265 70353 96311
rect 70431 96265 70477 96311
rect 70555 96265 70601 96311
rect 70679 96265 70725 96311
rect 70803 96265 70849 96311
rect 70927 96265 70973 96311
rect 71051 96265 71097 96311
rect 71175 96265 71221 96311
rect 71299 96265 71345 96311
rect 71423 96265 71469 96311
rect 71547 96265 71593 96311
rect 71671 96265 71717 96311
rect 71795 96265 71841 96311
rect 71919 96265 71965 96311
rect 72043 96265 72089 96311
rect 72167 96265 72213 96311
rect 72291 96265 72337 96311
rect 72415 96265 72461 96311
rect 72539 96265 72585 96311
rect 72663 96265 72709 96311
rect 72787 96265 72833 96311
rect 72911 96265 72957 96311
rect 73035 96265 73081 96311
rect 73159 96265 73205 96311
rect 73283 96265 73329 96311
rect 73407 96265 73453 96311
rect 73531 96265 73577 96311
rect 73655 96265 73701 96311
rect 73779 96265 73825 96311
rect 73903 96265 73949 96311
rect 74027 96265 74073 96311
rect 74151 96265 74197 96311
rect 74275 96265 74321 96311
rect 74399 96265 74445 96311
rect 74523 96265 74569 96311
rect 74647 96265 74693 96311
rect 74771 96265 74817 96311
rect 74895 96265 74941 96311
rect 75019 96265 75065 96311
rect 75143 96265 75189 96311
rect 75267 96265 75313 96311
rect 75391 96265 75437 96311
rect 75515 96265 75561 96311
rect 75639 96265 75685 96311
rect 75763 96265 75809 96311
rect 75887 96265 75933 96311
rect 76011 96265 76057 96311
rect 76135 96265 76181 96311
rect 76259 96265 76305 96311
rect 76383 96265 76429 96311
rect 76507 96265 76553 96311
rect 76631 96265 76677 96311
rect 76755 96265 76801 96311
rect 76879 96265 76925 96311
rect 77003 96265 77049 96311
rect 77127 96265 77173 96311
rect 77251 96265 77297 96311
rect 77375 96265 77421 96311
rect 77499 96265 77545 96311
rect 77623 96265 77669 96311
rect 77747 96265 77793 96311
rect 77871 96265 77917 96311
rect 77995 96265 78041 96311
rect 78119 96265 78165 96311
rect 78243 96265 78289 96311
rect 78367 96265 78413 96311
rect 78491 96265 78537 96311
rect 78615 96265 78661 96311
rect 78739 96265 78785 96311
rect 78863 96265 78909 96311
rect 78987 96265 79033 96311
rect 79111 96265 79157 96311
rect 79235 96265 79281 96311
rect 79359 96265 79405 96311
rect 79483 96265 79529 96311
rect 79607 96265 79653 96311
rect 79731 96265 79777 96311
rect 79855 96265 79901 96311
rect 79979 96265 80025 96311
rect 80103 96265 80149 96311
rect 80227 96265 80273 96311
rect 80351 96265 80397 96311
rect 80475 96265 80521 96311
rect 80599 96265 80645 96311
rect 80723 96265 80769 96311
rect 80847 96265 80893 96311
rect 80971 96265 81017 96311
rect 81095 96265 81141 96311
rect 81219 96265 81265 96311
rect 81343 96265 81389 96311
rect 81467 96265 81513 96311
rect 81591 96265 81637 96311
rect 81715 96265 81761 96311
rect 81839 96265 81885 96311
rect 81963 96265 82009 96311
rect 82087 96265 82133 96311
rect 82211 96265 82257 96311
rect 82335 96265 82381 96311
rect 82459 96265 82505 96311
rect 82583 96265 82629 96311
rect 82707 96265 82753 96311
rect 82831 96265 82877 96311
rect 82955 96265 83001 96311
rect 83079 96265 83125 96311
rect 83203 96265 83249 96311
rect 83327 96265 83373 96311
rect 83451 96265 83497 96311
rect 83575 96265 83621 96311
rect 83699 96265 83745 96311
rect 83823 96265 83869 96311
rect 83947 96265 83993 96311
rect 84071 96265 84117 96311
rect 84195 96265 84241 96311
rect 84319 96265 84365 96311
rect 84443 96265 84489 96311
rect 84567 96265 84613 96311
rect 84691 96265 84737 96311
rect 84815 96265 84861 96311
rect 84939 96265 84985 96311
rect 85063 96265 85109 96311
rect 85187 96265 85233 96311
rect 85311 96265 85357 96311
rect 85435 96265 85481 96311
rect 85559 96265 85605 96311
rect 85683 96265 85729 96311
rect 85807 96265 85853 96311
rect 85931 96265 85977 96311
rect 371 1117 717 96163
rect 27398 1117 27744 96163
rect 27822 35996 28668 96142
rect 56382 35996 57228 96142
rect 27822 34174 57168 34620
rect 28639 3860 28685 3906
rect 28755 3860 28801 3906
rect 28871 3860 28917 3906
rect 28987 3860 29033 3906
rect 29103 3860 29149 3906
rect 29219 3860 29265 3906
rect 29335 3860 29381 3906
rect 29451 3860 29497 3906
rect 29567 3860 29613 3906
rect 29683 3860 29729 3906
rect 29799 3860 29845 3906
rect 29915 3860 29961 3906
rect 30031 3860 30077 3906
rect 30147 3860 30193 3906
rect 30263 3860 30309 3906
rect 30379 3860 30425 3906
rect 30495 3860 30541 3906
rect 30611 3860 30657 3906
rect 30727 3860 30773 3906
rect 30843 3860 30889 3906
rect 30959 3860 31005 3906
rect 31075 3860 31121 3906
rect 31191 3860 31237 3906
rect 31307 3860 31353 3906
rect 31423 3860 31469 3906
rect 31539 3860 31585 3906
rect 31655 3860 31701 3906
rect 31771 3860 31817 3906
rect 31887 3860 31933 3906
rect 32003 3860 32049 3906
rect 32119 3860 32165 3906
rect 32235 3860 32281 3906
rect 32351 3860 32397 3906
rect 32467 3860 32513 3906
rect 32583 3860 32629 3906
rect 32699 3860 32745 3906
rect 32815 3860 32861 3906
rect 32931 3860 32977 3906
rect 33047 3860 33093 3906
rect 33163 3860 33209 3906
rect 33279 3860 33325 3906
rect 33395 3860 33441 3906
rect 33511 3860 33557 3906
rect 33627 3860 33673 3906
rect 33743 3860 33789 3906
rect 33859 3860 33905 3906
rect 33975 3860 34021 3906
rect 34091 3860 34137 3906
rect 34207 3860 34253 3906
rect 34323 3860 34369 3906
rect 34439 3860 34485 3906
rect 34555 3860 34601 3906
rect 34671 3860 34717 3906
rect 34787 3860 34833 3906
rect 34903 3860 34949 3906
rect 35019 3860 35065 3906
rect 35135 3860 35181 3906
rect 35251 3860 35297 3906
rect 35367 3860 35413 3906
rect 35483 3860 35529 3906
rect 35599 3860 35645 3906
rect 35715 3860 35761 3906
rect 35831 3860 35877 3906
rect 35947 3860 35993 3906
rect 36063 3860 36109 3906
rect 36179 3860 36225 3906
rect 36295 3860 36341 3906
rect 36411 3860 36457 3906
rect 36527 3860 36573 3906
rect 36643 3860 36689 3906
rect 36759 3860 36805 3906
rect 36875 3860 36921 3906
rect 36991 3860 37037 3906
rect 37107 3860 37153 3906
rect 37223 3860 37269 3906
rect 37339 3860 37385 3906
rect 37455 3860 37501 3906
rect 37571 3860 37617 3906
rect 37687 3860 37733 3906
rect 37803 3860 37849 3906
rect 37919 3860 37965 3906
rect 38035 3860 38081 3906
rect 38151 3860 38197 3906
rect 38267 3860 38313 3906
rect 38383 3860 38429 3906
rect 38499 3860 38545 3906
rect 38615 3860 38661 3906
rect 38731 3860 38777 3906
rect 38847 3860 38893 3906
rect 38963 3860 39009 3906
rect 39079 3860 39125 3906
rect 39195 3860 39241 3906
rect 39311 3860 39357 3906
rect 39427 3860 39473 3906
rect 39543 3860 39589 3906
rect 39659 3860 39705 3906
rect 39775 3860 39821 3906
rect 39891 3860 39937 3906
rect 40007 3860 40053 3906
rect 40123 3860 40169 3906
rect 28639 3744 28685 3790
rect 28755 3744 28801 3790
rect 28871 3744 28917 3790
rect 28987 3744 29033 3790
rect 29103 3744 29149 3790
rect 29219 3744 29265 3790
rect 29335 3744 29381 3790
rect 29451 3744 29497 3790
rect 29567 3744 29613 3790
rect 29683 3744 29729 3790
rect 29799 3744 29845 3790
rect 29915 3744 29961 3790
rect 30031 3744 30077 3790
rect 30147 3744 30193 3790
rect 30263 3744 30309 3790
rect 30379 3744 30425 3790
rect 30495 3744 30541 3790
rect 30611 3744 30657 3790
rect 30727 3744 30773 3790
rect 30843 3744 30889 3790
rect 30959 3744 31005 3790
rect 31075 3744 31121 3790
rect 31191 3744 31237 3790
rect 31307 3744 31353 3790
rect 31423 3744 31469 3790
rect 31539 3744 31585 3790
rect 31655 3744 31701 3790
rect 31771 3744 31817 3790
rect 31887 3744 31933 3790
rect 32003 3744 32049 3790
rect 32119 3744 32165 3790
rect 32235 3744 32281 3790
rect 32351 3744 32397 3790
rect 32467 3744 32513 3790
rect 32583 3744 32629 3790
rect 32699 3744 32745 3790
rect 32815 3744 32861 3790
rect 32931 3744 32977 3790
rect 33047 3744 33093 3790
rect 33163 3744 33209 3790
rect 33279 3744 33325 3790
rect 33395 3744 33441 3790
rect 33511 3744 33557 3790
rect 33627 3744 33673 3790
rect 33743 3744 33789 3790
rect 33859 3744 33905 3790
rect 33975 3744 34021 3790
rect 34091 3744 34137 3790
rect 34207 3744 34253 3790
rect 34323 3744 34369 3790
rect 34439 3744 34485 3790
rect 34555 3744 34601 3790
rect 34671 3744 34717 3790
rect 34787 3744 34833 3790
rect 34903 3744 34949 3790
rect 35019 3744 35065 3790
rect 35135 3744 35181 3790
rect 35251 3744 35297 3790
rect 35367 3744 35413 3790
rect 35483 3744 35529 3790
rect 35599 3744 35645 3790
rect 35715 3744 35761 3790
rect 35831 3744 35877 3790
rect 35947 3744 35993 3790
rect 36063 3744 36109 3790
rect 36179 3744 36225 3790
rect 36295 3744 36341 3790
rect 36411 3744 36457 3790
rect 36527 3744 36573 3790
rect 36643 3744 36689 3790
rect 36759 3744 36805 3790
rect 36875 3744 36921 3790
rect 36991 3744 37037 3790
rect 37107 3744 37153 3790
rect 37223 3744 37269 3790
rect 37339 3744 37385 3790
rect 37455 3744 37501 3790
rect 37571 3744 37617 3790
rect 37687 3744 37733 3790
rect 37803 3744 37849 3790
rect 37919 3744 37965 3790
rect 38035 3744 38081 3790
rect 38151 3744 38197 3790
rect 38267 3744 38313 3790
rect 38383 3744 38429 3790
rect 38499 3744 38545 3790
rect 38615 3744 38661 3790
rect 38731 3744 38777 3790
rect 38847 3744 38893 3790
rect 38963 3744 39009 3790
rect 39079 3744 39125 3790
rect 39195 3744 39241 3790
rect 39311 3744 39357 3790
rect 39427 3744 39473 3790
rect 39543 3744 39589 3790
rect 39659 3744 39705 3790
rect 39775 3744 39821 3790
rect 39891 3744 39937 3790
rect 40007 3744 40053 3790
rect 40123 3744 40169 3790
rect 28639 3628 28685 3674
rect 28755 3628 28801 3674
rect 28871 3628 28917 3674
rect 28987 3628 29033 3674
rect 29103 3628 29149 3674
rect 29219 3628 29265 3674
rect 29335 3628 29381 3674
rect 29451 3628 29497 3674
rect 29567 3628 29613 3674
rect 29683 3628 29729 3674
rect 29799 3628 29845 3674
rect 29915 3628 29961 3674
rect 30031 3628 30077 3674
rect 30147 3628 30193 3674
rect 30263 3628 30309 3674
rect 30379 3628 30425 3674
rect 30495 3628 30541 3674
rect 30611 3628 30657 3674
rect 30727 3628 30773 3674
rect 30843 3628 30889 3674
rect 30959 3628 31005 3674
rect 31075 3628 31121 3674
rect 31191 3628 31237 3674
rect 31307 3628 31353 3674
rect 31423 3628 31469 3674
rect 31539 3628 31585 3674
rect 31655 3628 31701 3674
rect 31771 3628 31817 3674
rect 31887 3628 31933 3674
rect 32003 3628 32049 3674
rect 32119 3628 32165 3674
rect 32235 3628 32281 3674
rect 32351 3628 32397 3674
rect 32467 3628 32513 3674
rect 32583 3628 32629 3674
rect 32699 3628 32745 3674
rect 32815 3628 32861 3674
rect 32931 3628 32977 3674
rect 33047 3628 33093 3674
rect 33163 3628 33209 3674
rect 33279 3628 33325 3674
rect 33395 3628 33441 3674
rect 33511 3628 33557 3674
rect 33627 3628 33673 3674
rect 33743 3628 33789 3674
rect 33859 3628 33905 3674
rect 33975 3628 34021 3674
rect 34091 3628 34137 3674
rect 34207 3628 34253 3674
rect 34323 3628 34369 3674
rect 34439 3628 34485 3674
rect 34555 3628 34601 3674
rect 34671 3628 34717 3674
rect 34787 3628 34833 3674
rect 34903 3628 34949 3674
rect 35019 3628 35065 3674
rect 35135 3628 35181 3674
rect 35251 3628 35297 3674
rect 35367 3628 35413 3674
rect 35483 3628 35529 3674
rect 35599 3628 35645 3674
rect 35715 3628 35761 3674
rect 35831 3628 35877 3674
rect 35947 3628 35993 3674
rect 36063 3628 36109 3674
rect 36179 3628 36225 3674
rect 36295 3628 36341 3674
rect 36411 3628 36457 3674
rect 36527 3628 36573 3674
rect 36643 3628 36689 3674
rect 36759 3628 36805 3674
rect 36875 3628 36921 3674
rect 36991 3628 37037 3674
rect 37107 3628 37153 3674
rect 37223 3628 37269 3674
rect 37339 3628 37385 3674
rect 37455 3628 37501 3674
rect 37571 3628 37617 3674
rect 37687 3628 37733 3674
rect 37803 3628 37849 3674
rect 37919 3628 37965 3674
rect 38035 3628 38081 3674
rect 38151 3628 38197 3674
rect 38267 3628 38313 3674
rect 38383 3628 38429 3674
rect 38499 3628 38545 3674
rect 38615 3628 38661 3674
rect 38731 3628 38777 3674
rect 38847 3628 38893 3674
rect 38963 3628 39009 3674
rect 39079 3628 39125 3674
rect 39195 3628 39241 3674
rect 39311 3628 39357 3674
rect 39427 3628 39473 3674
rect 39543 3628 39589 3674
rect 39659 3628 39705 3674
rect 39775 3628 39821 3674
rect 39891 3628 39937 3674
rect 40007 3628 40053 3674
rect 40123 3628 40169 3674
rect 28639 3512 28685 3558
rect 28755 3512 28801 3558
rect 28871 3512 28917 3558
rect 28987 3512 29033 3558
rect 29103 3512 29149 3558
rect 29219 3512 29265 3558
rect 29335 3512 29381 3558
rect 29451 3512 29497 3558
rect 29567 3512 29613 3558
rect 29683 3512 29729 3558
rect 29799 3512 29845 3558
rect 29915 3512 29961 3558
rect 30031 3512 30077 3558
rect 30147 3512 30193 3558
rect 30263 3512 30309 3558
rect 30379 3512 30425 3558
rect 30495 3512 30541 3558
rect 30611 3512 30657 3558
rect 30727 3512 30773 3558
rect 30843 3512 30889 3558
rect 30959 3512 31005 3558
rect 31075 3512 31121 3558
rect 31191 3512 31237 3558
rect 31307 3512 31353 3558
rect 31423 3512 31469 3558
rect 31539 3512 31585 3558
rect 31655 3512 31701 3558
rect 31771 3512 31817 3558
rect 31887 3512 31933 3558
rect 32003 3512 32049 3558
rect 32119 3512 32165 3558
rect 32235 3512 32281 3558
rect 32351 3512 32397 3558
rect 32467 3512 32513 3558
rect 32583 3512 32629 3558
rect 32699 3512 32745 3558
rect 32815 3512 32861 3558
rect 32931 3512 32977 3558
rect 33047 3512 33093 3558
rect 33163 3512 33209 3558
rect 33279 3512 33325 3558
rect 33395 3512 33441 3558
rect 33511 3512 33557 3558
rect 33627 3512 33673 3558
rect 33743 3512 33789 3558
rect 33859 3512 33905 3558
rect 33975 3512 34021 3558
rect 34091 3512 34137 3558
rect 34207 3512 34253 3558
rect 34323 3512 34369 3558
rect 34439 3512 34485 3558
rect 34555 3512 34601 3558
rect 34671 3512 34717 3558
rect 34787 3512 34833 3558
rect 34903 3512 34949 3558
rect 35019 3512 35065 3558
rect 35135 3512 35181 3558
rect 35251 3512 35297 3558
rect 35367 3512 35413 3558
rect 35483 3512 35529 3558
rect 35599 3512 35645 3558
rect 35715 3512 35761 3558
rect 35831 3512 35877 3558
rect 35947 3512 35993 3558
rect 36063 3512 36109 3558
rect 36179 3512 36225 3558
rect 36295 3512 36341 3558
rect 36411 3512 36457 3558
rect 36527 3512 36573 3558
rect 36643 3512 36689 3558
rect 36759 3512 36805 3558
rect 36875 3512 36921 3558
rect 36991 3512 37037 3558
rect 37107 3512 37153 3558
rect 37223 3512 37269 3558
rect 37339 3512 37385 3558
rect 37455 3512 37501 3558
rect 37571 3512 37617 3558
rect 37687 3512 37733 3558
rect 37803 3512 37849 3558
rect 37919 3512 37965 3558
rect 38035 3512 38081 3558
rect 38151 3512 38197 3558
rect 38267 3512 38313 3558
rect 38383 3512 38429 3558
rect 38499 3512 38545 3558
rect 38615 3512 38661 3558
rect 38731 3512 38777 3558
rect 38847 3512 38893 3558
rect 38963 3512 39009 3558
rect 39079 3512 39125 3558
rect 39195 3512 39241 3558
rect 39311 3512 39357 3558
rect 39427 3512 39473 3558
rect 39543 3512 39589 3558
rect 39659 3512 39705 3558
rect 39775 3512 39821 3558
rect 39891 3512 39937 3558
rect 40007 3512 40053 3558
rect 40123 3512 40169 3558
rect 28639 3396 28685 3442
rect 28755 3396 28801 3442
rect 28871 3396 28917 3442
rect 28987 3396 29033 3442
rect 29103 3396 29149 3442
rect 29219 3396 29265 3442
rect 29335 3396 29381 3442
rect 29451 3396 29497 3442
rect 29567 3396 29613 3442
rect 29683 3396 29729 3442
rect 29799 3396 29845 3442
rect 29915 3396 29961 3442
rect 30031 3396 30077 3442
rect 30147 3396 30193 3442
rect 30263 3396 30309 3442
rect 30379 3396 30425 3442
rect 30495 3396 30541 3442
rect 30611 3396 30657 3442
rect 30727 3396 30773 3442
rect 30843 3396 30889 3442
rect 30959 3396 31005 3442
rect 31075 3396 31121 3442
rect 31191 3396 31237 3442
rect 31307 3396 31353 3442
rect 31423 3396 31469 3442
rect 31539 3396 31585 3442
rect 31655 3396 31701 3442
rect 31771 3396 31817 3442
rect 31887 3396 31933 3442
rect 32003 3396 32049 3442
rect 32119 3396 32165 3442
rect 32235 3396 32281 3442
rect 32351 3396 32397 3442
rect 32467 3396 32513 3442
rect 32583 3396 32629 3442
rect 32699 3396 32745 3442
rect 32815 3396 32861 3442
rect 32931 3396 32977 3442
rect 33047 3396 33093 3442
rect 33163 3396 33209 3442
rect 33279 3396 33325 3442
rect 33395 3396 33441 3442
rect 33511 3396 33557 3442
rect 33627 3396 33673 3442
rect 33743 3396 33789 3442
rect 33859 3396 33905 3442
rect 33975 3396 34021 3442
rect 34091 3396 34137 3442
rect 34207 3396 34253 3442
rect 34323 3396 34369 3442
rect 34439 3396 34485 3442
rect 34555 3396 34601 3442
rect 34671 3396 34717 3442
rect 34787 3396 34833 3442
rect 34903 3396 34949 3442
rect 35019 3396 35065 3442
rect 35135 3396 35181 3442
rect 35251 3396 35297 3442
rect 35367 3396 35413 3442
rect 35483 3396 35529 3442
rect 35599 3396 35645 3442
rect 35715 3396 35761 3442
rect 35831 3396 35877 3442
rect 35947 3396 35993 3442
rect 36063 3396 36109 3442
rect 36179 3396 36225 3442
rect 36295 3396 36341 3442
rect 36411 3396 36457 3442
rect 36527 3396 36573 3442
rect 36643 3396 36689 3442
rect 36759 3396 36805 3442
rect 36875 3396 36921 3442
rect 36991 3396 37037 3442
rect 37107 3396 37153 3442
rect 37223 3396 37269 3442
rect 37339 3396 37385 3442
rect 37455 3396 37501 3442
rect 37571 3396 37617 3442
rect 37687 3396 37733 3442
rect 37803 3396 37849 3442
rect 37919 3396 37965 3442
rect 38035 3396 38081 3442
rect 38151 3396 38197 3442
rect 38267 3396 38313 3442
rect 38383 3396 38429 3442
rect 38499 3396 38545 3442
rect 38615 3396 38661 3442
rect 38731 3396 38777 3442
rect 38847 3396 38893 3442
rect 38963 3396 39009 3442
rect 39079 3396 39125 3442
rect 39195 3396 39241 3442
rect 39311 3396 39357 3442
rect 39427 3396 39473 3442
rect 39543 3396 39589 3442
rect 39659 3396 39705 3442
rect 39775 3396 39821 3442
rect 39891 3396 39937 3442
rect 40007 3396 40053 3442
rect 40123 3396 40169 3442
rect 28639 3280 28685 3326
rect 28755 3280 28801 3326
rect 28871 3280 28917 3326
rect 28987 3280 29033 3326
rect 29103 3280 29149 3326
rect 29219 3280 29265 3326
rect 29335 3280 29381 3326
rect 29451 3280 29497 3326
rect 29567 3280 29613 3326
rect 29683 3280 29729 3326
rect 29799 3280 29845 3326
rect 29915 3280 29961 3326
rect 30031 3280 30077 3326
rect 30147 3280 30193 3326
rect 30263 3280 30309 3326
rect 30379 3280 30425 3326
rect 30495 3280 30541 3326
rect 30611 3280 30657 3326
rect 30727 3280 30773 3326
rect 30843 3280 30889 3326
rect 30959 3280 31005 3326
rect 31075 3280 31121 3326
rect 31191 3280 31237 3326
rect 31307 3280 31353 3326
rect 31423 3280 31469 3326
rect 31539 3280 31585 3326
rect 31655 3280 31701 3326
rect 31771 3280 31817 3326
rect 31887 3280 31933 3326
rect 32003 3280 32049 3326
rect 32119 3280 32165 3326
rect 32235 3280 32281 3326
rect 32351 3280 32397 3326
rect 32467 3280 32513 3326
rect 32583 3280 32629 3326
rect 32699 3280 32745 3326
rect 32815 3280 32861 3326
rect 32931 3280 32977 3326
rect 33047 3280 33093 3326
rect 33163 3280 33209 3326
rect 33279 3280 33325 3326
rect 33395 3280 33441 3326
rect 33511 3280 33557 3326
rect 33627 3280 33673 3326
rect 33743 3280 33789 3326
rect 33859 3280 33905 3326
rect 33975 3280 34021 3326
rect 34091 3280 34137 3326
rect 34207 3280 34253 3326
rect 34323 3280 34369 3326
rect 34439 3280 34485 3326
rect 34555 3280 34601 3326
rect 34671 3280 34717 3326
rect 34787 3280 34833 3326
rect 34903 3280 34949 3326
rect 35019 3280 35065 3326
rect 35135 3280 35181 3326
rect 35251 3280 35297 3326
rect 35367 3280 35413 3326
rect 35483 3280 35529 3326
rect 35599 3280 35645 3326
rect 35715 3280 35761 3326
rect 35831 3280 35877 3326
rect 35947 3280 35993 3326
rect 36063 3280 36109 3326
rect 36179 3280 36225 3326
rect 36295 3280 36341 3326
rect 36411 3280 36457 3326
rect 36527 3280 36573 3326
rect 36643 3280 36689 3326
rect 36759 3280 36805 3326
rect 36875 3280 36921 3326
rect 36991 3280 37037 3326
rect 37107 3280 37153 3326
rect 37223 3280 37269 3326
rect 37339 3280 37385 3326
rect 37455 3280 37501 3326
rect 37571 3280 37617 3326
rect 37687 3280 37733 3326
rect 37803 3280 37849 3326
rect 37919 3280 37965 3326
rect 38035 3280 38081 3326
rect 38151 3280 38197 3326
rect 38267 3280 38313 3326
rect 38383 3280 38429 3326
rect 38499 3280 38545 3326
rect 38615 3280 38661 3326
rect 38731 3280 38777 3326
rect 38847 3280 38893 3326
rect 38963 3280 39009 3326
rect 39079 3280 39125 3326
rect 39195 3280 39241 3326
rect 39311 3280 39357 3326
rect 39427 3280 39473 3326
rect 39543 3280 39589 3326
rect 39659 3280 39705 3326
rect 39775 3280 39821 3326
rect 39891 3280 39937 3326
rect 40007 3280 40053 3326
rect 40123 3280 40169 3326
rect 28639 3164 28685 3210
rect 28755 3164 28801 3210
rect 28871 3164 28917 3210
rect 28987 3164 29033 3210
rect 29103 3164 29149 3210
rect 29219 3164 29265 3210
rect 29335 3164 29381 3210
rect 29451 3164 29497 3210
rect 29567 3164 29613 3210
rect 29683 3164 29729 3210
rect 29799 3164 29845 3210
rect 29915 3164 29961 3210
rect 30031 3164 30077 3210
rect 30147 3164 30193 3210
rect 30263 3164 30309 3210
rect 30379 3164 30425 3210
rect 30495 3164 30541 3210
rect 30611 3164 30657 3210
rect 30727 3164 30773 3210
rect 30843 3164 30889 3210
rect 30959 3164 31005 3210
rect 31075 3164 31121 3210
rect 31191 3164 31237 3210
rect 31307 3164 31353 3210
rect 31423 3164 31469 3210
rect 31539 3164 31585 3210
rect 31655 3164 31701 3210
rect 31771 3164 31817 3210
rect 31887 3164 31933 3210
rect 32003 3164 32049 3210
rect 32119 3164 32165 3210
rect 32235 3164 32281 3210
rect 32351 3164 32397 3210
rect 32467 3164 32513 3210
rect 32583 3164 32629 3210
rect 32699 3164 32745 3210
rect 32815 3164 32861 3210
rect 32931 3164 32977 3210
rect 33047 3164 33093 3210
rect 33163 3164 33209 3210
rect 33279 3164 33325 3210
rect 33395 3164 33441 3210
rect 33511 3164 33557 3210
rect 33627 3164 33673 3210
rect 33743 3164 33789 3210
rect 33859 3164 33905 3210
rect 33975 3164 34021 3210
rect 34091 3164 34137 3210
rect 34207 3164 34253 3210
rect 34323 3164 34369 3210
rect 34439 3164 34485 3210
rect 34555 3164 34601 3210
rect 34671 3164 34717 3210
rect 34787 3164 34833 3210
rect 34903 3164 34949 3210
rect 35019 3164 35065 3210
rect 35135 3164 35181 3210
rect 35251 3164 35297 3210
rect 35367 3164 35413 3210
rect 35483 3164 35529 3210
rect 35599 3164 35645 3210
rect 35715 3164 35761 3210
rect 35831 3164 35877 3210
rect 35947 3164 35993 3210
rect 36063 3164 36109 3210
rect 36179 3164 36225 3210
rect 36295 3164 36341 3210
rect 36411 3164 36457 3210
rect 36527 3164 36573 3210
rect 36643 3164 36689 3210
rect 36759 3164 36805 3210
rect 36875 3164 36921 3210
rect 36991 3164 37037 3210
rect 37107 3164 37153 3210
rect 37223 3164 37269 3210
rect 37339 3164 37385 3210
rect 37455 3164 37501 3210
rect 37571 3164 37617 3210
rect 37687 3164 37733 3210
rect 37803 3164 37849 3210
rect 37919 3164 37965 3210
rect 38035 3164 38081 3210
rect 38151 3164 38197 3210
rect 38267 3164 38313 3210
rect 38383 3164 38429 3210
rect 38499 3164 38545 3210
rect 38615 3164 38661 3210
rect 38731 3164 38777 3210
rect 38847 3164 38893 3210
rect 38963 3164 39009 3210
rect 39079 3164 39125 3210
rect 39195 3164 39241 3210
rect 39311 3164 39357 3210
rect 39427 3164 39473 3210
rect 39543 3164 39589 3210
rect 39659 3164 39705 3210
rect 39775 3164 39821 3210
rect 39891 3164 39937 3210
rect 40007 3164 40053 3210
rect 40123 3164 40169 3210
rect 28639 3048 28685 3094
rect 28755 3048 28801 3094
rect 28871 3048 28917 3094
rect 28987 3048 29033 3094
rect 29103 3048 29149 3094
rect 29219 3048 29265 3094
rect 29335 3048 29381 3094
rect 29451 3048 29497 3094
rect 29567 3048 29613 3094
rect 29683 3048 29729 3094
rect 29799 3048 29845 3094
rect 29915 3048 29961 3094
rect 30031 3048 30077 3094
rect 30147 3048 30193 3094
rect 30263 3048 30309 3094
rect 30379 3048 30425 3094
rect 30495 3048 30541 3094
rect 30611 3048 30657 3094
rect 30727 3048 30773 3094
rect 30843 3048 30889 3094
rect 30959 3048 31005 3094
rect 31075 3048 31121 3094
rect 31191 3048 31237 3094
rect 31307 3048 31353 3094
rect 31423 3048 31469 3094
rect 31539 3048 31585 3094
rect 31655 3048 31701 3094
rect 31771 3048 31817 3094
rect 31887 3048 31933 3094
rect 32003 3048 32049 3094
rect 32119 3048 32165 3094
rect 32235 3048 32281 3094
rect 32351 3048 32397 3094
rect 32467 3048 32513 3094
rect 32583 3048 32629 3094
rect 32699 3048 32745 3094
rect 32815 3048 32861 3094
rect 32931 3048 32977 3094
rect 33047 3048 33093 3094
rect 33163 3048 33209 3094
rect 33279 3048 33325 3094
rect 33395 3048 33441 3094
rect 33511 3048 33557 3094
rect 33627 3048 33673 3094
rect 33743 3048 33789 3094
rect 33859 3048 33905 3094
rect 33975 3048 34021 3094
rect 34091 3048 34137 3094
rect 34207 3048 34253 3094
rect 34323 3048 34369 3094
rect 34439 3048 34485 3094
rect 34555 3048 34601 3094
rect 34671 3048 34717 3094
rect 34787 3048 34833 3094
rect 34903 3048 34949 3094
rect 35019 3048 35065 3094
rect 35135 3048 35181 3094
rect 35251 3048 35297 3094
rect 35367 3048 35413 3094
rect 35483 3048 35529 3094
rect 35599 3048 35645 3094
rect 35715 3048 35761 3094
rect 35831 3048 35877 3094
rect 35947 3048 35993 3094
rect 36063 3048 36109 3094
rect 36179 3048 36225 3094
rect 36295 3048 36341 3094
rect 36411 3048 36457 3094
rect 36527 3048 36573 3094
rect 36643 3048 36689 3094
rect 36759 3048 36805 3094
rect 36875 3048 36921 3094
rect 36991 3048 37037 3094
rect 37107 3048 37153 3094
rect 37223 3048 37269 3094
rect 37339 3048 37385 3094
rect 37455 3048 37501 3094
rect 37571 3048 37617 3094
rect 37687 3048 37733 3094
rect 37803 3048 37849 3094
rect 37919 3048 37965 3094
rect 38035 3048 38081 3094
rect 38151 3048 38197 3094
rect 38267 3048 38313 3094
rect 38383 3048 38429 3094
rect 38499 3048 38545 3094
rect 38615 3048 38661 3094
rect 38731 3048 38777 3094
rect 38847 3048 38893 3094
rect 38963 3048 39009 3094
rect 39079 3048 39125 3094
rect 39195 3048 39241 3094
rect 39311 3048 39357 3094
rect 39427 3048 39473 3094
rect 39543 3048 39589 3094
rect 39659 3048 39705 3094
rect 39775 3048 39821 3094
rect 39891 3048 39937 3094
rect 40007 3048 40053 3094
rect 40123 3048 40169 3094
rect 28639 2932 28685 2978
rect 28755 2932 28801 2978
rect 28871 2932 28917 2978
rect 28987 2932 29033 2978
rect 29103 2932 29149 2978
rect 29219 2932 29265 2978
rect 29335 2932 29381 2978
rect 29451 2932 29497 2978
rect 29567 2932 29613 2978
rect 29683 2932 29729 2978
rect 29799 2932 29845 2978
rect 29915 2932 29961 2978
rect 30031 2932 30077 2978
rect 30147 2932 30193 2978
rect 30263 2932 30309 2978
rect 30379 2932 30425 2978
rect 30495 2932 30541 2978
rect 30611 2932 30657 2978
rect 30727 2932 30773 2978
rect 30843 2932 30889 2978
rect 30959 2932 31005 2978
rect 31075 2932 31121 2978
rect 31191 2932 31237 2978
rect 31307 2932 31353 2978
rect 31423 2932 31469 2978
rect 31539 2932 31585 2978
rect 31655 2932 31701 2978
rect 31771 2932 31817 2978
rect 31887 2932 31933 2978
rect 32003 2932 32049 2978
rect 32119 2932 32165 2978
rect 32235 2932 32281 2978
rect 32351 2932 32397 2978
rect 32467 2932 32513 2978
rect 32583 2932 32629 2978
rect 32699 2932 32745 2978
rect 32815 2932 32861 2978
rect 32931 2932 32977 2978
rect 33047 2932 33093 2978
rect 33163 2932 33209 2978
rect 33279 2932 33325 2978
rect 33395 2932 33441 2978
rect 33511 2932 33557 2978
rect 33627 2932 33673 2978
rect 33743 2932 33789 2978
rect 33859 2932 33905 2978
rect 33975 2932 34021 2978
rect 34091 2932 34137 2978
rect 34207 2932 34253 2978
rect 34323 2932 34369 2978
rect 34439 2932 34485 2978
rect 34555 2932 34601 2978
rect 34671 2932 34717 2978
rect 34787 2932 34833 2978
rect 34903 2932 34949 2978
rect 35019 2932 35065 2978
rect 35135 2932 35181 2978
rect 35251 2932 35297 2978
rect 35367 2932 35413 2978
rect 35483 2932 35529 2978
rect 35599 2932 35645 2978
rect 35715 2932 35761 2978
rect 35831 2932 35877 2978
rect 35947 2932 35993 2978
rect 36063 2932 36109 2978
rect 36179 2932 36225 2978
rect 36295 2932 36341 2978
rect 36411 2932 36457 2978
rect 36527 2932 36573 2978
rect 36643 2932 36689 2978
rect 36759 2932 36805 2978
rect 36875 2932 36921 2978
rect 36991 2932 37037 2978
rect 37107 2932 37153 2978
rect 37223 2932 37269 2978
rect 37339 2932 37385 2978
rect 37455 2932 37501 2978
rect 37571 2932 37617 2978
rect 37687 2932 37733 2978
rect 37803 2932 37849 2978
rect 37919 2932 37965 2978
rect 38035 2932 38081 2978
rect 38151 2932 38197 2978
rect 38267 2932 38313 2978
rect 38383 2932 38429 2978
rect 38499 2932 38545 2978
rect 38615 2932 38661 2978
rect 38731 2932 38777 2978
rect 38847 2932 38893 2978
rect 38963 2932 39009 2978
rect 39079 2932 39125 2978
rect 39195 2932 39241 2978
rect 39311 2932 39357 2978
rect 39427 2932 39473 2978
rect 39543 2932 39589 2978
rect 39659 2932 39705 2978
rect 39775 2932 39821 2978
rect 39891 2932 39937 2978
rect 40007 2932 40053 2978
rect 40123 2932 40169 2978
rect 28639 2816 28685 2862
rect 28755 2816 28801 2862
rect 28871 2816 28917 2862
rect 28987 2816 29033 2862
rect 29103 2816 29149 2862
rect 29219 2816 29265 2862
rect 29335 2816 29381 2862
rect 29451 2816 29497 2862
rect 29567 2816 29613 2862
rect 29683 2816 29729 2862
rect 29799 2816 29845 2862
rect 29915 2816 29961 2862
rect 30031 2816 30077 2862
rect 30147 2816 30193 2862
rect 30263 2816 30309 2862
rect 30379 2816 30425 2862
rect 30495 2816 30541 2862
rect 30611 2816 30657 2862
rect 30727 2816 30773 2862
rect 30843 2816 30889 2862
rect 30959 2816 31005 2862
rect 31075 2816 31121 2862
rect 31191 2816 31237 2862
rect 31307 2816 31353 2862
rect 31423 2816 31469 2862
rect 31539 2816 31585 2862
rect 31655 2816 31701 2862
rect 31771 2816 31817 2862
rect 31887 2816 31933 2862
rect 32003 2816 32049 2862
rect 32119 2816 32165 2862
rect 32235 2816 32281 2862
rect 32351 2816 32397 2862
rect 32467 2816 32513 2862
rect 32583 2816 32629 2862
rect 32699 2816 32745 2862
rect 32815 2816 32861 2862
rect 32931 2816 32977 2862
rect 33047 2816 33093 2862
rect 33163 2816 33209 2862
rect 33279 2816 33325 2862
rect 33395 2816 33441 2862
rect 33511 2816 33557 2862
rect 33627 2816 33673 2862
rect 33743 2816 33789 2862
rect 33859 2816 33905 2862
rect 33975 2816 34021 2862
rect 34091 2816 34137 2862
rect 34207 2816 34253 2862
rect 34323 2816 34369 2862
rect 34439 2816 34485 2862
rect 34555 2816 34601 2862
rect 34671 2816 34717 2862
rect 34787 2816 34833 2862
rect 34903 2816 34949 2862
rect 35019 2816 35065 2862
rect 35135 2816 35181 2862
rect 35251 2816 35297 2862
rect 35367 2816 35413 2862
rect 35483 2816 35529 2862
rect 35599 2816 35645 2862
rect 35715 2816 35761 2862
rect 35831 2816 35877 2862
rect 35947 2816 35993 2862
rect 36063 2816 36109 2862
rect 36179 2816 36225 2862
rect 36295 2816 36341 2862
rect 36411 2816 36457 2862
rect 36527 2816 36573 2862
rect 36643 2816 36689 2862
rect 36759 2816 36805 2862
rect 36875 2816 36921 2862
rect 36991 2816 37037 2862
rect 37107 2816 37153 2862
rect 37223 2816 37269 2862
rect 37339 2816 37385 2862
rect 37455 2816 37501 2862
rect 37571 2816 37617 2862
rect 37687 2816 37733 2862
rect 37803 2816 37849 2862
rect 37919 2816 37965 2862
rect 38035 2816 38081 2862
rect 38151 2816 38197 2862
rect 38267 2816 38313 2862
rect 38383 2816 38429 2862
rect 38499 2816 38545 2862
rect 38615 2816 38661 2862
rect 38731 2816 38777 2862
rect 38847 2816 38893 2862
rect 38963 2816 39009 2862
rect 39079 2816 39125 2862
rect 39195 2816 39241 2862
rect 39311 2816 39357 2862
rect 39427 2816 39473 2862
rect 39543 2816 39589 2862
rect 39659 2816 39705 2862
rect 39775 2816 39821 2862
rect 39891 2816 39937 2862
rect 40007 2816 40053 2862
rect 40123 2816 40169 2862
rect 28639 2700 28685 2746
rect 28755 2700 28801 2746
rect 28871 2700 28917 2746
rect 28987 2700 29033 2746
rect 29103 2700 29149 2746
rect 29219 2700 29265 2746
rect 29335 2700 29381 2746
rect 29451 2700 29497 2746
rect 29567 2700 29613 2746
rect 29683 2700 29729 2746
rect 29799 2700 29845 2746
rect 29915 2700 29961 2746
rect 30031 2700 30077 2746
rect 30147 2700 30193 2746
rect 30263 2700 30309 2746
rect 30379 2700 30425 2746
rect 30495 2700 30541 2746
rect 30611 2700 30657 2746
rect 30727 2700 30773 2746
rect 30843 2700 30889 2746
rect 30959 2700 31005 2746
rect 31075 2700 31121 2746
rect 31191 2700 31237 2746
rect 31307 2700 31353 2746
rect 31423 2700 31469 2746
rect 31539 2700 31585 2746
rect 31655 2700 31701 2746
rect 31771 2700 31817 2746
rect 31887 2700 31933 2746
rect 32003 2700 32049 2746
rect 32119 2700 32165 2746
rect 32235 2700 32281 2746
rect 32351 2700 32397 2746
rect 32467 2700 32513 2746
rect 32583 2700 32629 2746
rect 32699 2700 32745 2746
rect 32815 2700 32861 2746
rect 32931 2700 32977 2746
rect 33047 2700 33093 2746
rect 33163 2700 33209 2746
rect 33279 2700 33325 2746
rect 33395 2700 33441 2746
rect 33511 2700 33557 2746
rect 33627 2700 33673 2746
rect 33743 2700 33789 2746
rect 33859 2700 33905 2746
rect 33975 2700 34021 2746
rect 34091 2700 34137 2746
rect 34207 2700 34253 2746
rect 34323 2700 34369 2746
rect 34439 2700 34485 2746
rect 34555 2700 34601 2746
rect 34671 2700 34717 2746
rect 34787 2700 34833 2746
rect 34903 2700 34949 2746
rect 35019 2700 35065 2746
rect 35135 2700 35181 2746
rect 35251 2700 35297 2746
rect 35367 2700 35413 2746
rect 35483 2700 35529 2746
rect 35599 2700 35645 2746
rect 35715 2700 35761 2746
rect 35831 2700 35877 2746
rect 35947 2700 35993 2746
rect 36063 2700 36109 2746
rect 36179 2700 36225 2746
rect 36295 2700 36341 2746
rect 36411 2700 36457 2746
rect 36527 2700 36573 2746
rect 36643 2700 36689 2746
rect 36759 2700 36805 2746
rect 36875 2700 36921 2746
rect 36991 2700 37037 2746
rect 37107 2700 37153 2746
rect 37223 2700 37269 2746
rect 37339 2700 37385 2746
rect 37455 2700 37501 2746
rect 37571 2700 37617 2746
rect 37687 2700 37733 2746
rect 37803 2700 37849 2746
rect 37919 2700 37965 2746
rect 38035 2700 38081 2746
rect 38151 2700 38197 2746
rect 38267 2700 38313 2746
rect 38383 2700 38429 2746
rect 38499 2700 38545 2746
rect 38615 2700 38661 2746
rect 38731 2700 38777 2746
rect 38847 2700 38893 2746
rect 38963 2700 39009 2746
rect 39079 2700 39125 2746
rect 39195 2700 39241 2746
rect 39311 2700 39357 2746
rect 39427 2700 39473 2746
rect 39543 2700 39589 2746
rect 39659 2700 39705 2746
rect 39775 2700 39821 2746
rect 39891 2700 39937 2746
rect 40007 2700 40053 2746
rect 40123 2700 40169 2746
rect 28639 2584 28685 2630
rect 28755 2584 28801 2630
rect 28871 2584 28917 2630
rect 28987 2584 29033 2630
rect 29103 2584 29149 2630
rect 29219 2584 29265 2630
rect 29335 2584 29381 2630
rect 29451 2584 29497 2630
rect 29567 2584 29613 2630
rect 29683 2584 29729 2630
rect 29799 2584 29845 2630
rect 29915 2584 29961 2630
rect 30031 2584 30077 2630
rect 30147 2584 30193 2630
rect 30263 2584 30309 2630
rect 30379 2584 30425 2630
rect 30495 2584 30541 2630
rect 30611 2584 30657 2630
rect 30727 2584 30773 2630
rect 30843 2584 30889 2630
rect 30959 2584 31005 2630
rect 31075 2584 31121 2630
rect 31191 2584 31237 2630
rect 31307 2584 31353 2630
rect 31423 2584 31469 2630
rect 31539 2584 31585 2630
rect 31655 2584 31701 2630
rect 31771 2584 31817 2630
rect 31887 2584 31933 2630
rect 32003 2584 32049 2630
rect 32119 2584 32165 2630
rect 32235 2584 32281 2630
rect 32351 2584 32397 2630
rect 32467 2584 32513 2630
rect 32583 2584 32629 2630
rect 32699 2584 32745 2630
rect 32815 2584 32861 2630
rect 32931 2584 32977 2630
rect 33047 2584 33093 2630
rect 33163 2584 33209 2630
rect 33279 2584 33325 2630
rect 33395 2584 33441 2630
rect 33511 2584 33557 2630
rect 33627 2584 33673 2630
rect 33743 2584 33789 2630
rect 33859 2584 33905 2630
rect 33975 2584 34021 2630
rect 34091 2584 34137 2630
rect 34207 2584 34253 2630
rect 34323 2584 34369 2630
rect 34439 2584 34485 2630
rect 34555 2584 34601 2630
rect 34671 2584 34717 2630
rect 34787 2584 34833 2630
rect 34903 2584 34949 2630
rect 35019 2584 35065 2630
rect 35135 2584 35181 2630
rect 35251 2584 35297 2630
rect 35367 2584 35413 2630
rect 35483 2584 35529 2630
rect 35599 2584 35645 2630
rect 35715 2584 35761 2630
rect 35831 2584 35877 2630
rect 35947 2584 35993 2630
rect 36063 2584 36109 2630
rect 36179 2584 36225 2630
rect 36295 2584 36341 2630
rect 36411 2584 36457 2630
rect 36527 2584 36573 2630
rect 36643 2584 36689 2630
rect 36759 2584 36805 2630
rect 36875 2584 36921 2630
rect 36991 2584 37037 2630
rect 37107 2584 37153 2630
rect 37223 2584 37269 2630
rect 37339 2584 37385 2630
rect 37455 2584 37501 2630
rect 37571 2584 37617 2630
rect 37687 2584 37733 2630
rect 37803 2584 37849 2630
rect 37919 2584 37965 2630
rect 38035 2584 38081 2630
rect 38151 2584 38197 2630
rect 38267 2584 38313 2630
rect 38383 2584 38429 2630
rect 38499 2584 38545 2630
rect 38615 2584 38661 2630
rect 38731 2584 38777 2630
rect 38847 2584 38893 2630
rect 38963 2584 39009 2630
rect 39079 2584 39125 2630
rect 39195 2584 39241 2630
rect 39311 2584 39357 2630
rect 39427 2584 39473 2630
rect 39543 2584 39589 2630
rect 39659 2584 39705 2630
rect 39775 2584 39821 2630
rect 39891 2584 39937 2630
rect 40007 2584 40053 2630
rect 40123 2584 40169 2630
rect 28639 2468 28685 2514
rect 28755 2468 28801 2514
rect 28871 2468 28917 2514
rect 28987 2468 29033 2514
rect 29103 2468 29149 2514
rect 29219 2468 29265 2514
rect 29335 2468 29381 2514
rect 29451 2468 29497 2514
rect 29567 2468 29613 2514
rect 29683 2468 29729 2514
rect 29799 2468 29845 2514
rect 29915 2468 29961 2514
rect 30031 2468 30077 2514
rect 30147 2468 30193 2514
rect 30263 2468 30309 2514
rect 30379 2468 30425 2514
rect 30495 2468 30541 2514
rect 30611 2468 30657 2514
rect 30727 2468 30773 2514
rect 30843 2468 30889 2514
rect 30959 2468 31005 2514
rect 31075 2468 31121 2514
rect 31191 2468 31237 2514
rect 31307 2468 31353 2514
rect 31423 2468 31469 2514
rect 31539 2468 31585 2514
rect 31655 2468 31701 2514
rect 31771 2468 31817 2514
rect 31887 2468 31933 2514
rect 32003 2468 32049 2514
rect 32119 2468 32165 2514
rect 32235 2468 32281 2514
rect 32351 2468 32397 2514
rect 32467 2468 32513 2514
rect 32583 2468 32629 2514
rect 32699 2468 32745 2514
rect 32815 2468 32861 2514
rect 32931 2468 32977 2514
rect 33047 2468 33093 2514
rect 33163 2468 33209 2514
rect 33279 2468 33325 2514
rect 33395 2468 33441 2514
rect 33511 2468 33557 2514
rect 33627 2468 33673 2514
rect 33743 2468 33789 2514
rect 33859 2468 33905 2514
rect 33975 2468 34021 2514
rect 34091 2468 34137 2514
rect 34207 2468 34253 2514
rect 34323 2468 34369 2514
rect 34439 2468 34485 2514
rect 34555 2468 34601 2514
rect 34671 2468 34717 2514
rect 34787 2468 34833 2514
rect 34903 2468 34949 2514
rect 35019 2468 35065 2514
rect 35135 2468 35181 2514
rect 35251 2468 35297 2514
rect 35367 2468 35413 2514
rect 35483 2468 35529 2514
rect 35599 2468 35645 2514
rect 35715 2468 35761 2514
rect 35831 2468 35877 2514
rect 35947 2468 35993 2514
rect 36063 2468 36109 2514
rect 36179 2468 36225 2514
rect 36295 2468 36341 2514
rect 36411 2468 36457 2514
rect 36527 2468 36573 2514
rect 36643 2468 36689 2514
rect 36759 2468 36805 2514
rect 36875 2468 36921 2514
rect 36991 2468 37037 2514
rect 37107 2468 37153 2514
rect 37223 2468 37269 2514
rect 37339 2468 37385 2514
rect 37455 2468 37501 2514
rect 37571 2468 37617 2514
rect 37687 2468 37733 2514
rect 37803 2468 37849 2514
rect 37919 2468 37965 2514
rect 38035 2468 38081 2514
rect 38151 2468 38197 2514
rect 38267 2468 38313 2514
rect 38383 2468 38429 2514
rect 38499 2468 38545 2514
rect 38615 2468 38661 2514
rect 38731 2468 38777 2514
rect 38847 2468 38893 2514
rect 38963 2468 39009 2514
rect 39079 2468 39125 2514
rect 39195 2468 39241 2514
rect 39311 2468 39357 2514
rect 39427 2468 39473 2514
rect 39543 2468 39589 2514
rect 39659 2468 39705 2514
rect 39775 2468 39821 2514
rect 39891 2468 39937 2514
rect 40007 2468 40053 2514
rect 40123 2468 40169 2514
rect 28639 2352 28685 2398
rect 28755 2352 28801 2398
rect 28871 2352 28917 2398
rect 28987 2352 29033 2398
rect 29103 2352 29149 2398
rect 29219 2352 29265 2398
rect 29335 2352 29381 2398
rect 29451 2352 29497 2398
rect 29567 2352 29613 2398
rect 29683 2352 29729 2398
rect 29799 2352 29845 2398
rect 29915 2352 29961 2398
rect 30031 2352 30077 2398
rect 30147 2352 30193 2398
rect 30263 2352 30309 2398
rect 30379 2352 30425 2398
rect 30495 2352 30541 2398
rect 30611 2352 30657 2398
rect 30727 2352 30773 2398
rect 30843 2352 30889 2398
rect 30959 2352 31005 2398
rect 31075 2352 31121 2398
rect 31191 2352 31237 2398
rect 31307 2352 31353 2398
rect 31423 2352 31469 2398
rect 31539 2352 31585 2398
rect 31655 2352 31701 2398
rect 31771 2352 31817 2398
rect 31887 2352 31933 2398
rect 32003 2352 32049 2398
rect 32119 2352 32165 2398
rect 32235 2352 32281 2398
rect 32351 2352 32397 2398
rect 32467 2352 32513 2398
rect 32583 2352 32629 2398
rect 32699 2352 32745 2398
rect 32815 2352 32861 2398
rect 32931 2352 32977 2398
rect 33047 2352 33093 2398
rect 33163 2352 33209 2398
rect 33279 2352 33325 2398
rect 33395 2352 33441 2398
rect 33511 2352 33557 2398
rect 33627 2352 33673 2398
rect 33743 2352 33789 2398
rect 33859 2352 33905 2398
rect 33975 2352 34021 2398
rect 34091 2352 34137 2398
rect 34207 2352 34253 2398
rect 34323 2352 34369 2398
rect 34439 2352 34485 2398
rect 34555 2352 34601 2398
rect 34671 2352 34717 2398
rect 34787 2352 34833 2398
rect 34903 2352 34949 2398
rect 35019 2352 35065 2398
rect 35135 2352 35181 2398
rect 35251 2352 35297 2398
rect 35367 2352 35413 2398
rect 35483 2352 35529 2398
rect 35599 2352 35645 2398
rect 35715 2352 35761 2398
rect 35831 2352 35877 2398
rect 35947 2352 35993 2398
rect 36063 2352 36109 2398
rect 36179 2352 36225 2398
rect 36295 2352 36341 2398
rect 36411 2352 36457 2398
rect 36527 2352 36573 2398
rect 36643 2352 36689 2398
rect 36759 2352 36805 2398
rect 36875 2352 36921 2398
rect 36991 2352 37037 2398
rect 37107 2352 37153 2398
rect 37223 2352 37269 2398
rect 37339 2352 37385 2398
rect 37455 2352 37501 2398
rect 37571 2352 37617 2398
rect 37687 2352 37733 2398
rect 37803 2352 37849 2398
rect 37919 2352 37965 2398
rect 38035 2352 38081 2398
rect 38151 2352 38197 2398
rect 38267 2352 38313 2398
rect 38383 2352 38429 2398
rect 38499 2352 38545 2398
rect 38615 2352 38661 2398
rect 38731 2352 38777 2398
rect 38847 2352 38893 2398
rect 38963 2352 39009 2398
rect 39079 2352 39125 2398
rect 39195 2352 39241 2398
rect 39311 2352 39357 2398
rect 39427 2352 39473 2398
rect 39543 2352 39589 2398
rect 39659 2352 39705 2398
rect 39775 2352 39821 2398
rect 39891 2352 39937 2398
rect 40007 2352 40053 2398
rect 40123 2352 40169 2398
rect 28639 2236 28685 2282
rect 28755 2236 28801 2282
rect 28871 2236 28917 2282
rect 28987 2236 29033 2282
rect 29103 2236 29149 2282
rect 29219 2236 29265 2282
rect 29335 2236 29381 2282
rect 29451 2236 29497 2282
rect 29567 2236 29613 2282
rect 29683 2236 29729 2282
rect 29799 2236 29845 2282
rect 29915 2236 29961 2282
rect 30031 2236 30077 2282
rect 30147 2236 30193 2282
rect 30263 2236 30309 2282
rect 30379 2236 30425 2282
rect 30495 2236 30541 2282
rect 30611 2236 30657 2282
rect 30727 2236 30773 2282
rect 30843 2236 30889 2282
rect 30959 2236 31005 2282
rect 31075 2236 31121 2282
rect 31191 2236 31237 2282
rect 31307 2236 31353 2282
rect 31423 2236 31469 2282
rect 31539 2236 31585 2282
rect 31655 2236 31701 2282
rect 31771 2236 31817 2282
rect 31887 2236 31933 2282
rect 32003 2236 32049 2282
rect 32119 2236 32165 2282
rect 32235 2236 32281 2282
rect 32351 2236 32397 2282
rect 32467 2236 32513 2282
rect 32583 2236 32629 2282
rect 32699 2236 32745 2282
rect 32815 2236 32861 2282
rect 32931 2236 32977 2282
rect 33047 2236 33093 2282
rect 33163 2236 33209 2282
rect 33279 2236 33325 2282
rect 33395 2236 33441 2282
rect 33511 2236 33557 2282
rect 33627 2236 33673 2282
rect 33743 2236 33789 2282
rect 33859 2236 33905 2282
rect 33975 2236 34021 2282
rect 34091 2236 34137 2282
rect 34207 2236 34253 2282
rect 34323 2236 34369 2282
rect 34439 2236 34485 2282
rect 34555 2236 34601 2282
rect 34671 2236 34717 2282
rect 34787 2236 34833 2282
rect 34903 2236 34949 2282
rect 35019 2236 35065 2282
rect 35135 2236 35181 2282
rect 35251 2236 35297 2282
rect 35367 2236 35413 2282
rect 35483 2236 35529 2282
rect 35599 2236 35645 2282
rect 35715 2236 35761 2282
rect 35831 2236 35877 2282
rect 35947 2236 35993 2282
rect 36063 2236 36109 2282
rect 36179 2236 36225 2282
rect 36295 2236 36341 2282
rect 36411 2236 36457 2282
rect 36527 2236 36573 2282
rect 36643 2236 36689 2282
rect 36759 2236 36805 2282
rect 36875 2236 36921 2282
rect 36991 2236 37037 2282
rect 37107 2236 37153 2282
rect 37223 2236 37269 2282
rect 37339 2236 37385 2282
rect 37455 2236 37501 2282
rect 37571 2236 37617 2282
rect 37687 2236 37733 2282
rect 37803 2236 37849 2282
rect 37919 2236 37965 2282
rect 38035 2236 38081 2282
rect 38151 2236 38197 2282
rect 38267 2236 38313 2282
rect 38383 2236 38429 2282
rect 38499 2236 38545 2282
rect 38615 2236 38661 2282
rect 38731 2236 38777 2282
rect 38847 2236 38893 2282
rect 38963 2236 39009 2282
rect 39079 2236 39125 2282
rect 39195 2236 39241 2282
rect 39311 2236 39357 2282
rect 39427 2236 39473 2282
rect 39543 2236 39589 2282
rect 39659 2236 39705 2282
rect 39775 2236 39821 2282
rect 39891 2236 39937 2282
rect 40007 2236 40053 2282
rect 40123 2236 40169 2282
rect 28639 2120 28685 2166
rect 28755 2120 28801 2166
rect 28871 2120 28917 2166
rect 28987 2120 29033 2166
rect 29103 2120 29149 2166
rect 29219 2120 29265 2166
rect 29335 2120 29381 2166
rect 29451 2120 29497 2166
rect 29567 2120 29613 2166
rect 29683 2120 29729 2166
rect 29799 2120 29845 2166
rect 29915 2120 29961 2166
rect 30031 2120 30077 2166
rect 30147 2120 30193 2166
rect 30263 2120 30309 2166
rect 30379 2120 30425 2166
rect 30495 2120 30541 2166
rect 30611 2120 30657 2166
rect 30727 2120 30773 2166
rect 30843 2120 30889 2166
rect 30959 2120 31005 2166
rect 31075 2120 31121 2166
rect 31191 2120 31237 2166
rect 31307 2120 31353 2166
rect 31423 2120 31469 2166
rect 31539 2120 31585 2166
rect 31655 2120 31701 2166
rect 31771 2120 31817 2166
rect 31887 2120 31933 2166
rect 32003 2120 32049 2166
rect 32119 2120 32165 2166
rect 32235 2120 32281 2166
rect 32351 2120 32397 2166
rect 32467 2120 32513 2166
rect 32583 2120 32629 2166
rect 32699 2120 32745 2166
rect 32815 2120 32861 2166
rect 32931 2120 32977 2166
rect 33047 2120 33093 2166
rect 33163 2120 33209 2166
rect 33279 2120 33325 2166
rect 33395 2120 33441 2166
rect 33511 2120 33557 2166
rect 33627 2120 33673 2166
rect 33743 2120 33789 2166
rect 33859 2120 33905 2166
rect 33975 2120 34021 2166
rect 34091 2120 34137 2166
rect 34207 2120 34253 2166
rect 34323 2120 34369 2166
rect 34439 2120 34485 2166
rect 34555 2120 34601 2166
rect 34671 2120 34717 2166
rect 34787 2120 34833 2166
rect 34903 2120 34949 2166
rect 35019 2120 35065 2166
rect 35135 2120 35181 2166
rect 35251 2120 35297 2166
rect 35367 2120 35413 2166
rect 35483 2120 35529 2166
rect 35599 2120 35645 2166
rect 35715 2120 35761 2166
rect 35831 2120 35877 2166
rect 35947 2120 35993 2166
rect 36063 2120 36109 2166
rect 36179 2120 36225 2166
rect 36295 2120 36341 2166
rect 36411 2120 36457 2166
rect 36527 2120 36573 2166
rect 36643 2120 36689 2166
rect 36759 2120 36805 2166
rect 36875 2120 36921 2166
rect 36991 2120 37037 2166
rect 37107 2120 37153 2166
rect 37223 2120 37269 2166
rect 37339 2120 37385 2166
rect 37455 2120 37501 2166
rect 37571 2120 37617 2166
rect 37687 2120 37733 2166
rect 37803 2120 37849 2166
rect 37919 2120 37965 2166
rect 38035 2120 38081 2166
rect 38151 2120 38197 2166
rect 38267 2120 38313 2166
rect 38383 2120 38429 2166
rect 38499 2120 38545 2166
rect 38615 2120 38661 2166
rect 38731 2120 38777 2166
rect 38847 2120 38893 2166
rect 38963 2120 39009 2166
rect 39079 2120 39125 2166
rect 39195 2120 39241 2166
rect 39311 2120 39357 2166
rect 39427 2120 39473 2166
rect 39543 2120 39589 2166
rect 39659 2120 39705 2166
rect 39775 2120 39821 2166
rect 39891 2120 39937 2166
rect 40007 2120 40053 2166
rect 40123 2120 40169 2166
rect 28639 2004 28685 2050
rect 28755 2004 28801 2050
rect 28871 2004 28917 2050
rect 28987 2004 29033 2050
rect 29103 2004 29149 2050
rect 29219 2004 29265 2050
rect 29335 2004 29381 2050
rect 29451 2004 29497 2050
rect 29567 2004 29613 2050
rect 29683 2004 29729 2050
rect 29799 2004 29845 2050
rect 29915 2004 29961 2050
rect 30031 2004 30077 2050
rect 30147 2004 30193 2050
rect 30263 2004 30309 2050
rect 30379 2004 30425 2050
rect 30495 2004 30541 2050
rect 30611 2004 30657 2050
rect 30727 2004 30773 2050
rect 30843 2004 30889 2050
rect 30959 2004 31005 2050
rect 31075 2004 31121 2050
rect 31191 2004 31237 2050
rect 31307 2004 31353 2050
rect 31423 2004 31469 2050
rect 31539 2004 31585 2050
rect 31655 2004 31701 2050
rect 31771 2004 31817 2050
rect 31887 2004 31933 2050
rect 32003 2004 32049 2050
rect 32119 2004 32165 2050
rect 32235 2004 32281 2050
rect 32351 2004 32397 2050
rect 32467 2004 32513 2050
rect 32583 2004 32629 2050
rect 32699 2004 32745 2050
rect 32815 2004 32861 2050
rect 32931 2004 32977 2050
rect 33047 2004 33093 2050
rect 33163 2004 33209 2050
rect 33279 2004 33325 2050
rect 33395 2004 33441 2050
rect 33511 2004 33557 2050
rect 33627 2004 33673 2050
rect 33743 2004 33789 2050
rect 33859 2004 33905 2050
rect 33975 2004 34021 2050
rect 34091 2004 34137 2050
rect 34207 2004 34253 2050
rect 34323 2004 34369 2050
rect 34439 2004 34485 2050
rect 34555 2004 34601 2050
rect 34671 2004 34717 2050
rect 34787 2004 34833 2050
rect 34903 2004 34949 2050
rect 35019 2004 35065 2050
rect 35135 2004 35181 2050
rect 35251 2004 35297 2050
rect 35367 2004 35413 2050
rect 35483 2004 35529 2050
rect 35599 2004 35645 2050
rect 35715 2004 35761 2050
rect 35831 2004 35877 2050
rect 35947 2004 35993 2050
rect 36063 2004 36109 2050
rect 36179 2004 36225 2050
rect 36295 2004 36341 2050
rect 36411 2004 36457 2050
rect 36527 2004 36573 2050
rect 36643 2004 36689 2050
rect 36759 2004 36805 2050
rect 36875 2004 36921 2050
rect 36991 2004 37037 2050
rect 37107 2004 37153 2050
rect 37223 2004 37269 2050
rect 37339 2004 37385 2050
rect 37455 2004 37501 2050
rect 37571 2004 37617 2050
rect 37687 2004 37733 2050
rect 37803 2004 37849 2050
rect 37919 2004 37965 2050
rect 38035 2004 38081 2050
rect 38151 2004 38197 2050
rect 38267 2004 38313 2050
rect 38383 2004 38429 2050
rect 38499 2004 38545 2050
rect 38615 2004 38661 2050
rect 38731 2004 38777 2050
rect 38847 2004 38893 2050
rect 38963 2004 39009 2050
rect 39079 2004 39125 2050
rect 39195 2004 39241 2050
rect 39311 2004 39357 2050
rect 39427 2004 39473 2050
rect 39543 2004 39589 2050
rect 39659 2004 39705 2050
rect 39775 2004 39821 2050
rect 39891 2004 39937 2050
rect 40007 2004 40053 2050
rect 40123 2004 40169 2050
rect 28639 1888 28685 1934
rect 28755 1888 28801 1934
rect 28871 1888 28917 1934
rect 28987 1888 29033 1934
rect 29103 1888 29149 1934
rect 29219 1888 29265 1934
rect 29335 1888 29381 1934
rect 29451 1888 29497 1934
rect 29567 1888 29613 1934
rect 29683 1888 29729 1934
rect 29799 1888 29845 1934
rect 29915 1888 29961 1934
rect 30031 1888 30077 1934
rect 30147 1888 30193 1934
rect 30263 1888 30309 1934
rect 30379 1888 30425 1934
rect 30495 1888 30541 1934
rect 30611 1888 30657 1934
rect 30727 1888 30773 1934
rect 30843 1888 30889 1934
rect 30959 1888 31005 1934
rect 31075 1888 31121 1934
rect 31191 1888 31237 1934
rect 31307 1888 31353 1934
rect 31423 1888 31469 1934
rect 31539 1888 31585 1934
rect 31655 1888 31701 1934
rect 31771 1888 31817 1934
rect 31887 1888 31933 1934
rect 32003 1888 32049 1934
rect 32119 1888 32165 1934
rect 32235 1888 32281 1934
rect 32351 1888 32397 1934
rect 32467 1888 32513 1934
rect 32583 1888 32629 1934
rect 32699 1888 32745 1934
rect 32815 1888 32861 1934
rect 32931 1888 32977 1934
rect 33047 1888 33093 1934
rect 33163 1888 33209 1934
rect 33279 1888 33325 1934
rect 33395 1888 33441 1934
rect 33511 1888 33557 1934
rect 33627 1888 33673 1934
rect 33743 1888 33789 1934
rect 33859 1888 33905 1934
rect 33975 1888 34021 1934
rect 34091 1888 34137 1934
rect 34207 1888 34253 1934
rect 34323 1888 34369 1934
rect 34439 1888 34485 1934
rect 34555 1888 34601 1934
rect 34671 1888 34717 1934
rect 34787 1888 34833 1934
rect 34903 1888 34949 1934
rect 35019 1888 35065 1934
rect 35135 1888 35181 1934
rect 35251 1888 35297 1934
rect 35367 1888 35413 1934
rect 35483 1888 35529 1934
rect 35599 1888 35645 1934
rect 35715 1888 35761 1934
rect 35831 1888 35877 1934
rect 35947 1888 35993 1934
rect 36063 1888 36109 1934
rect 36179 1888 36225 1934
rect 36295 1888 36341 1934
rect 36411 1888 36457 1934
rect 36527 1888 36573 1934
rect 36643 1888 36689 1934
rect 36759 1888 36805 1934
rect 36875 1888 36921 1934
rect 36991 1888 37037 1934
rect 37107 1888 37153 1934
rect 37223 1888 37269 1934
rect 37339 1888 37385 1934
rect 37455 1888 37501 1934
rect 37571 1888 37617 1934
rect 37687 1888 37733 1934
rect 37803 1888 37849 1934
rect 37919 1888 37965 1934
rect 38035 1888 38081 1934
rect 38151 1888 38197 1934
rect 38267 1888 38313 1934
rect 38383 1888 38429 1934
rect 38499 1888 38545 1934
rect 38615 1888 38661 1934
rect 38731 1888 38777 1934
rect 38847 1888 38893 1934
rect 38963 1888 39009 1934
rect 39079 1888 39125 1934
rect 39195 1888 39241 1934
rect 39311 1888 39357 1934
rect 39427 1888 39473 1934
rect 39543 1888 39589 1934
rect 39659 1888 39705 1934
rect 39775 1888 39821 1934
rect 39891 1888 39937 1934
rect 40007 1888 40053 1934
rect 40123 1888 40169 1934
rect 28639 1772 28685 1818
rect 28755 1772 28801 1818
rect 28871 1772 28917 1818
rect 28987 1772 29033 1818
rect 29103 1772 29149 1818
rect 29219 1772 29265 1818
rect 29335 1772 29381 1818
rect 29451 1772 29497 1818
rect 29567 1772 29613 1818
rect 29683 1772 29729 1818
rect 29799 1772 29845 1818
rect 29915 1772 29961 1818
rect 30031 1772 30077 1818
rect 30147 1772 30193 1818
rect 30263 1772 30309 1818
rect 30379 1772 30425 1818
rect 30495 1772 30541 1818
rect 30611 1772 30657 1818
rect 30727 1772 30773 1818
rect 30843 1772 30889 1818
rect 30959 1772 31005 1818
rect 31075 1772 31121 1818
rect 31191 1772 31237 1818
rect 31307 1772 31353 1818
rect 31423 1772 31469 1818
rect 31539 1772 31585 1818
rect 31655 1772 31701 1818
rect 31771 1772 31817 1818
rect 31887 1772 31933 1818
rect 32003 1772 32049 1818
rect 32119 1772 32165 1818
rect 32235 1772 32281 1818
rect 32351 1772 32397 1818
rect 32467 1772 32513 1818
rect 32583 1772 32629 1818
rect 32699 1772 32745 1818
rect 32815 1772 32861 1818
rect 32931 1772 32977 1818
rect 33047 1772 33093 1818
rect 33163 1772 33209 1818
rect 33279 1772 33325 1818
rect 33395 1772 33441 1818
rect 33511 1772 33557 1818
rect 33627 1772 33673 1818
rect 33743 1772 33789 1818
rect 33859 1772 33905 1818
rect 33975 1772 34021 1818
rect 34091 1772 34137 1818
rect 34207 1772 34253 1818
rect 34323 1772 34369 1818
rect 34439 1772 34485 1818
rect 34555 1772 34601 1818
rect 34671 1772 34717 1818
rect 34787 1772 34833 1818
rect 34903 1772 34949 1818
rect 35019 1772 35065 1818
rect 35135 1772 35181 1818
rect 35251 1772 35297 1818
rect 35367 1772 35413 1818
rect 35483 1772 35529 1818
rect 35599 1772 35645 1818
rect 35715 1772 35761 1818
rect 35831 1772 35877 1818
rect 35947 1772 35993 1818
rect 36063 1772 36109 1818
rect 36179 1772 36225 1818
rect 36295 1772 36341 1818
rect 36411 1772 36457 1818
rect 36527 1772 36573 1818
rect 36643 1772 36689 1818
rect 36759 1772 36805 1818
rect 36875 1772 36921 1818
rect 36991 1772 37037 1818
rect 37107 1772 37153 1818
rect 37223 1772 37269 1818
rect 37339 1772 37385 1818
rect 37455 1772 37501 1818
rect 37571 1772 37617 1818
rect 37687 1772 37733 1818
rect 37803 1772 37849 1818
rect 37919 1772 37965 1818
rect 38035 1772 38081 1818
rect 38151 1772 38197 1818
rect 38267 1772 38313 1818
rect 38383 1772 38429 1818
rect 38499 1772 38545 1818
rect 38615 1772 38661 1818
rect 38731 1772 38777 1818
rect 38847 1772 38893 1818
rect 38963 1772 39009 1818
rect 39079 1772 39125 1818
rect 39195 1772 39241 1818
rect 39311 1772 39357 1818
rect 39427 1772 39473 1818
rect 39543 1772 39589 1818
rect 39659 1772 39705 1818
rect 39775 1772 39821 1818
rect 39891 1772 39937 1818
rect 40007 1772 40053 1818
rect 40123 1772 40169 1818
rect 28639 1656 28685 1702
rect 28755 1656 28801 1702
rect 28871 1656 28917 1702
rect 28987 1656 29033 1702
rect 29103 1656 29149 1702
rect 29219 1656 29265 1702
rect 29335 1656 29381 1702
rect 29451 1656 29497 1702
rect 29567 1656 29613 1702
rect 29683 1656 29729 1702
rect 29799 1656 29845 1702
rect 29915 1656 29961 1702
rect 30031 1656 30077 1702
rect 30147 1656 30193 1702
rect 30263 1656 30309 1702
rect 30379 1656 30425 1702
rect 30495 1656 30541 1702
rect 30611 1656 30657 1702
rect 30727 1656 30773 1702
rect 30843 1656 30889 1702
rect 30959 1656 31005 1702
rect 31075 1656 31121 1702
rect 31191 1656 31237 1702
rect 31307 1656 31353 1702
rect 31423 1656 31469 1702
rect 31539 1656 31585 1702
rect 31655 1656 31701 1702
rect 31771 1656 31817 1702
rect 31887 1656 31933 1702
rect 32003 1656 32049 1702
rect 32119 1656 32165 1702
rect 32235 1656 32281 1702
rect 32351 1656 32397 1702
rect 32467 1656 32513 1702
rect 32583 1656 32629 1702
rect 32699 1656 32745 1702
rect 32815 1656 32861 1702
rect 32931 1656 32977 1702
rect 33047 1656 33093 1702
rect 33163 1656 33209 1702
rect 33279 1656 33325 1702
rect 33395 1656 33441 1702
rect 33511 1656 33557 1702
rect 33627 1656 33673 1702
rect 33743 1656 33789 1702
rect 33859 1656 33905 1702
rect 33975 1656 34021 1702
rect 34091 1656 34137 1702
rect 34207 1656 34253 1702
rect 34323 1656 34369 1702
rect 34439 1656 34485 1702
rect 34555 1656 34601 1702
rect 34671 1656 34717 1702
rect 34787 1656 34833 1702
rect 34903 1656 34949 1702
rect 35019 1656 35065 1702
rect 35135 1656 35181 1702
rect 35251 1656 35297 1702
rect 35367 1656 35413 1702
rect 35483 1656 35529 1702
rect 35599 1656 35645 1702
rect 35715 1656 35761 1702
rect 35831 1656 35877 1702
rect 35947 1656 35993 1702
rect 36063 1656 36109 1702
rect 36179 1656 36225 1702
rect 36295 1656 36341 1702
rect 36411 1656 36457 1702
rect 36527 1656 36573 1702
rect 36643 1656 36689 1702
rect 36759 1656 36805 1702
rect 36875 1656 36921 1702
rect 36991 1656 37037 1702
rect 37107 1656 37153 1702
rect 37223 1656 37269 1702
rect 37339 1656 37385 1702
rect 37455 1656 37501 1702
rect 37571 1656 37617 1702
rect 37687 1656 37733 1702
rect 37803 1656 37849 1702
rect 37919 1656 37965 1702
rect 38035 1656 38081 1702
rect 38151 1656 38197 1702
rect 38267 1656 38313 1702
rect 38383 1656 38429 1702
rect 38499 1656 38545 1702
rect 38615 1656 38661 1702
rect 38731 1656 38777 1702
rect 38847 1656 38893 1702
rect 38963 1656 39009 1702
rect 39079 1656 39125 1702
rect 39195 1656 39241 1702
rect 39311 1656 39357 1702
rect 39427 1656 39473 1702
rect 39543 1656 39589 1702
rect 39659 1656 39705 1702
rect 39775 1656 39821 1702
rect 39891 1656 39937 1702
rect 40007 1656 40053 1702
rect 40123 1656 40169 1702
rect 50845 3860 50891 3906
rect 50961 3860 51007 3906
rect 51077 3860 51123 3906
rect 51193 3860 51239 3906
rect 51309 3860 51355 3906
rect 51425 3860 51471 3906
rect 51541 3860 51587 3906
rect 51657 3860 51703 3906
rect 51773 3860 51819 3906
rect 51889 3860 51935 3906
rect 52005 3860 52051 3906
rect 52121 3860 52167 3906
rect 52237 3860 52283 3906
rect 52353 3860 52399 3906
rect 52469 3860 52515 3906
rect 52585 3860 52631 3906
rect 52701 3860 52747 3906
rect 52817 3860 52863 3906
rect 52933 3860 52979 3906
rect 53049 3860 53095 3906
rect 53165 3860 53211 3906
rect 53281 3860 53327 3906
rect 53397 3860 53443 3906
rect 53513 3860 53559 3906
rect 53629 3860 53675 3906
rect 53745 3860 53791 3906
rect 53861 3860 53907 3906
rect 53977 3860 54023 3906
rect 54093 3860 54139 3906
rect 54209 3860 54255 3906
rect 54325 3860 54371 3906
rect 54441 3860 54487 3906
rect 54557 3860 54603 3906
rect 54673 3860 54719 3906
rect 54789 3860 54835 3906
rect 54905 3860 54951 3906
rect 55021 3860 55067 3906
rect 55137 3860 55183 3906
rect 55253 3860 55299 3906
rect 55369 3860 55415 3906
rect 55485 3860 55531 3906
rect 55601 3860 55647 3906
rect 55717 3860 55763 3906
rect 55833 3860 55879 3906
rect 55949 3860 55995 3906
rect 56065 3860 56111 3906
rect 56181 3860 56227 3906
rect 56297 3860 56343 3906
rect 56413 3860 56459 3906
rect 56529 3860 56575 3906
rect 50845 3744 50891 3790
rect 50961 3744 51007 3790
rect 51077 3744 51123 3790
rect 51193 3744 51239 3790
rect 51309 3744 51355 3790
rect 51425 3744 51471 3790
rect 51541 3744 51587 3790
rect 51657 3744 51703 3790
rect 51773 3744 51819 3790
rect 51889 3744 51935 3790
rect 52005 3744 52051 3790
rect 52121 3744 52167 3790
rect 52237 3744 52283 3790
rect 52353 3744 52399 3790
rect 52469 3744 52515 3790
rect 52585 3744 52631 3790
rect 52701 3744 52747 3790
rect 52817 3744 52863 3790
rect 52933 3744 52979 3790
rect 53049 3744 53095 3790
rect 53165 3744 53211 3790
rect 53281 3744 53327 3790
rect 53397 3744 53443 3790
rect 53513 3744 53559 3790
rect 53629 3744 53675 3790
rect 53745 3744 53791 3790
rect 53861 3744 53907 3790
rect 53977 3744 54023 3790
rect 54093 3744 54139 3790
rect 54209 3744 54255 3790
rect 54325 3744 54371 3790
rect 54441 3744 54487 3790
rect 54557 3744 54603 3790
rect 54673 3744 54719 3790
rect 54789 3744 54835 3790
rect 54905 3744 54951 3790
rect 55021 3744 55067 3790
rect 55137 3744 55183 3790
rect 55253 3744 55299 3790
rect 55369 3744 55415 3790
rect 55485 3744 55531 3790
rect 55601 3744 55647 3790
rect 55717 3744 55763 3790
rect 55833 3744 55879 3790
rect 55949 3744 55995 3790
rect 56065 3744 56111 3790
rect 56181 3744 56227 3790
rect 56297 3744 56343 3790
rect 56413 3744 56459 3790
rect 56529 3744 56575 3790
rect 50845 3628 50891 3674
rect 50961 3628 51007 3674
rect 51077 3628 51123 3674
rect 51193 3628 51239 3674
rect 51309 3628 51355 3674
rect 51425 3628 51471 3674
rect 51541 3628 51587 3674
rect 51657 3628 51703 3674
rect 51773 3628 51819 3674
rect 51889 3628 51935 3674
rect 52005 3628 52051 3674
rect 52121 3628 52167 3674
rect 52237 3628 52283 3674
rect 52353 3628 52399 3674
rect 52469 3628 52515 3674
rect 52585 3628 52631 3674
rect 52701 3628 52747 3674
rect 52817 3628 52863 3674
rect 52933 3628 52979 3674
rect 53049 3628 53095 3674
rect 53165 3628 53211 3674
rect 53281 3628 53327 3674
rect 53397 3628 53443 3674
rect 53513 3628 53559 3674
rect 53629 3628 53675 3674
rect 53745 3628 53791 3674
rect 53861 3628 53907 3674
rect 53977 3628 54023 3674
rect 54093 3628 54139 3674
rect 54209 3628 54255 3674
rect 54325 3628 54371 3674
rect 54441 3628 54487 3674
rect 54557 3628 54603 3674
rect 54673 3628 54719 3674
rect 54789 3628 54835 3674
rect 54905 3628 54951 3674
rect 55021 3628 55067 3674
rect 55137 3628 55183 3674
rect 55253 3628 55299 3674
rect 55369 3628 55415 3674
rect 55485 3628 55531 3674
rect 55601 3628 55647 3674
rect 55717 3628 55763 3674
rect 55833 3628 55879 3674
rect 55949 3628 55995 3674
rect 56065 3628 56111 3674
rect 56181 3628 56227 3674
rect 56297 3628 56343 3674
rect 56413 3628 56459 3674
rect 56529 3628 56575 3674
rect 50845 3512 50891 3558
rect 50961 3512 51007 3558
rect 51077 3512 51123 3558
rect 51193 3512 51239 3558
rect 51309 3512 51355 3558
rect 51425 3512 51471 3558
rect 51541 3512 51587 3558
rect 51657 3512 51703 3558
rect 51773 3512 51819 3558
rect 51889 3512 51935 3558
rect 52005 3512 52051 3558
rect 52121 3512 52167 3558
rect 52237 3512 52283 3558
rect 52353 3512 52399 3558
rect 52469 3512 52515 3558
rect 52585 3512 52631 3558
rect 52701 3512 52747 3558
rect 52817 3512 52863 3558
rect 52933 3512 52979 3558
rect 53049 3512 53095 3558
rect 53165 3512 53211 3558
rect 53281 3512 53327 3558
rect 53397 3512 53443 3558
rect 53513 3512 53559 3558
rect 53629 3512 53675 3558
rect 53745 3512 53791 3558
rect 53861 3512 53907 3558
rect 53977 3512 54023 3558
rect 54093 3512 54139 3558
rect 54209 3512 54255 3558
rect 54325 3512 54371 3558
rect 54441 3512 54487 3558
rect 54557 3512 54603 3558
rect 54673 3512 54719 3558
rect 54789 3512 54835 3558
rect 54905 3512 54951 3558
rect 55021 3512 55067 3558
rect 55137 3512 55183 3558
rect 55253 3512 55299 3558
rect 55369 3512 55415 3558
rect 55485 3512 55531 3558
rect 55601 3512 55647 3558
rect 55717 3512 55763 3558
rect 55833 3512 55879 3558
rect 55949 3512 55995 3558
rect 56065 3512 56111 3558
rect 56181 3512 56227 3558
rect 56297 3512 56343 3558
rect 56413 3512 56459 3558
rect 56529 3512 56575 3558
rect 50845 3396 50891 3442
rect 50961 3396 51007 3442
rect 51077 3396 51123 3442
rect 51193 3396 51239 3442
rect 51309 3396 51355 3442
rect 51425 3396 51471 3442
rect 51541 3396 51587 3442
rect 51657 3396 51703 3442
rect 51773 3396 51819 3442
rect 51889 3396 51935 3442
rect 52005 3396 52051 3442
rect 52121 3396 52167 3442
rect 52237 3396 52283 3442
rect 52353 3396 52399 3442
rect 52469 3396 52515 3442
rect 52585 3396 52631 3442
rect 52701 3396 52747 3442
rect 52817 3396 52863 3442
rect 52933 3396 52979 3442
rect 53049 3396 53095 3442
rect 53165 3396 53211 3442
rect 53281 3396 53327 3442
rect 53397 3396 53443 3442
rect 53513 3396 53559 3442
rect 53629 3396 53675 3442
rect 53745 3396 53791 3442
rect 53861 3396 53907 3442
rect 53977 3396 54023 3442
rect 54093 3396 54139 3442
rect 54209 3396 54255 3442
rect 54325 3396 54371 3442
rect 54441 3396 54487 3442
rect 54557 3396 54603 3442
rect 54673 3396 54719 3442
rect 54789 3396 54835 3442
rect 54905 3396 54951 3442
rect 55021 3396 55067 3442
rect 55137 3396 55183 3442
rect 55253 3396 55299 3442
rect 55369 3396 55415 3442
rect 55485 3396 55531 3442
rect 55601 3396 55647 3442
rect 55717 3396 55763 3442
rect 55833 3396 55879 3442
rect 55949 3396 55995 3442
rect 56065 3396 56111 3442
rect 56181 3396 56227 3442
rect 56297 3396 56343 3442
rect 56413 3396 56459 3442
rect 56529 3396 56575 3442
rect 50845 3280 50891 3326
rect 50961 3280 51007 3326
rect 51077 3280 51123 3326
rect 51193 3280 51239 3326
rect 51309 3280 51355 3326
rect 51425 3280 51471 3326
rect 51541 3280 51587 3326
rect 51657 3280 51703 3326
rect 51773 3280 51819 3326
rect 51889 3280 51935 3326
rect 52005 3280 52051 3326
rect 52121 3280 52167 3326
rect 52237 3280 52283 3326
rect 52353 3280 52399 3326
rect 52469 3280 52515 3326
rect 52585 3280 52631 3326
rect 52701 3280 52747 3326
rect 52817 3280 52863 3326
rect 52933 3280 52979 3326
rect 53049 3280 53095 3326
rect 53165 3280 53211 3326
rect 53281 3280 53327 3326
rect 53397 3280 53443 3326
rect 53513 3280 53559 3326
rect 53629 3280 53675 3326
rect 53745 3280 53791 3326
rect 53861 3280 53907 3326
rect 53977 3280 54023 3326
rect 54093 3280 54139 3326
rect 54209 3280 54255 3326
rect 54325 3280 54371 3326
rect 54441 3280 54487 3326
rect 54557 3280 54603 3326
rect 54673 3280 54719 3326
rect 54789 3280 54835 3326
rect 54905 3280 54951 3326
rect 55021 3280 55067 3326
rect 55137 3280 55183 3326
rect 55253 3280 55299 3326
rect 55369 3280 55415 3326
rect 55485 3280 55531 3326
rect 55601 3280 55647 3326
rect 55717 3280 55763 3326
rect 55833 3280 55879 3326
rect 55949 3280 55995 3326
rect 56065 3280 56111 3326
rect 56181 3280 56227 3326
rect 56297 3280 56343 3326
rect 56413 3280 56459 3326
rect 56529 3280 56575 3326
rect 50845 3164 50891 3210
rect 50961 3164 51007 3210
rect 51077 3164 51123 3210
rect 51193 3164 51239 3210
rect 51309 3164 51355 3210
rect 51425 3164 51471 3210
rect 51541 3164 51587 3210
rect 51657 3164 51703 3210
rect 51773 3164 51819 3210
rect 51889 3164 51935 3210
rect 52005 3164 52051 3210
rect 52121 3164 52167 3210
rect 52237 3164 52283 3210
rect 52353 3164 52399 3210
rect 52469 3164 52515 3210
rect 52585 3164 52631 3210
rect 52701 3164 52747 3210
rect 52817 3164 52863 3210
rect 52933 3164 52979 3210
rect 53049 3164 53095 3210
rect 53165 3164 53211 3210
rect 53281 3164 53327 3210
rect 53397 3164 53443 3210
rect 53513 3164 53559 3210
rect 53629 3164 53675 3210
rect 53745 3164 53791 3210
rect 53861 3164 53907 3210
rect 53977 3164 54023 3210
rect 54093 3164 54139 3210
rect 54209 3164 54255 3210
rect 54325 3164 54371 3210
rect 54441 3164 54487 3210
rect 54557 3164 54603 3210
rect 54673 3164 54719 3210
rect 54789 3164 54835 3210
rect 54905 3164 54951 3210
rect 55021 3164 55067 3210
rect 55137 3164 55183 3210
rect 55253 3164 55299 3210
rect 55369 3164 55415 3210
rect 55485 3164 55531 3210
rect 55601 3164 55647 3210
rect 55717 3164 55763 3210
rect 55833 3164 55879 3210
rect 55949 3164 55995 3210
rect 56065 3164 56111 3210
rect 56181 3164 56227 3210
rect 56297 3164 56343 3210
rect 56413 3164 56459 3210
rect 56529 3164 56575 3210
rect 50845 3048 50891 3094
rect 50961 3048 51007 3094
rect 51077 3048 51123 3094
rect 51193 3048 51239 3094
rect 51309 3048 51355 3094
rect 51425 3048 51471 3094
rect 51541 3048 51587 3094
rect 51657 3048 51703 3094
rect 51773 3048 51819 3094
rect 51889 3048 51935 3094
rect 52005 3048 52051 3094
rect 52121 3048 52167 3094
rect 52237 3048 52283 3094
rect 52353 3048 52399 3094
rect 52469 3048 52515 3094
rect 52585 3048 52631 3094
rect 52701 3048 52747 3094
rect 52817 3048 52863 3094
rect 52933 3048 52979 3094
rect 53049 3048 53095 3094
rect 53165 3048 53211 3094
rect 53281 3048 53327 3094
rect 53397 3048 53443 3094
rect 53513 3048 53559 3094
rect 53629 3048 53675 3094
rect 53745 3048 53791 3094
rect 53861 3048 53907 3094
rect 53977 3048 54023 3094
rect 54093 3048 54139 3094
rect 54209 3048 54255 3094
rect 54325 3048 54371 3094
rect 54441 3048 54487 3094
rect 54557 3048 54603 3094
rect 54673 3048 54719 3094
rect 54789 3048 54835 3094
rect 54905 3048 54951 3094
rect 55021 3048 55067 3094
rect 55137 3048 55183 3094
rect 55253 3048 55299 3094
rect 55369 3048 55415 3094
rect 55485 3048 55531 3094
rect 55601 3048 55647 3094
rect 55717 3048 55763 3094
rect 55833 3048 55879 3094
rect 55949 3048 55995 3094
rect 56065 3048 56111 3094
rect 56181 3048 56227 3094
rect 56297 3048 56343 3094
rect 56413 3048 56459 3094
rect 56529 3048 56575 3094
rect 50845 2932 50891 2978
rect 50961 2932 51007 2978
rect 51077 2932 51123 2978
rect 51193 2932 51239 2978
rect 51309 2932 51355 2978
rect 51425 2932 51471 2978
rect 51541 2932 51587 2978
rect 51657 2932 51703 2978
rect 51773 2932 51819 2978
rect 51889 2932 51935 2978
rect 52005 2932 52051 2978
rect 52121 2932 52167 2978
rect 52237 2932 52283 2978
rect 52353 2932 52399 2978
rect 52469 2932 52515 2978
rect 52585 2932 52631 2978
rect 52701 2932 52747 2978
rect 52817 2932 52863 2978
rect 52933 2932 52979 2978
rect 53049 2932 53095 2978
rect 53165 2932 53211 2978
rect 53281 2932 53327 2978
rect 53397 2932 53443 2978
rect 53513 2932 53559 2978
rect 53629 2932 53675 2978
rect 53745 2932 53791 2978
rect 53861 2932 53907 2978
rect 53977 2932 54023 2978
rect 54093 2932 54139 2978
rect 54209 2932 54255 2978
rect 54325 2932 54371 2978
rect 54441 2932 54487 2978
rect 54557 2932 54603 2978
rect 54673 2932 54719 2978
rect 54789 2932 54835 2978
rect 54905 2932 54951 2978
rect 55021 2932 55067 2978
rect 55137 2932 55183 2978
rect 55253 2932 55299 2978
rect 55369 2932 55415 2978
rect 55485 2932 55531 2978
rect 55601 2932 55647 2978
rect 55717 2932 55763 2978
rect 55833 2932 55879 2978
rect 55949 2932 55995 2978
rect 56065 2932 56111 2978
rect 56181 2932 56227 2978
rect 56297 2932 56343 2978
rect 56413 2932 56459 2978
rect 56529 2932 56575 2978
rect 50845 2816 50891 2862
rect 50961 2816 51007 2862
rect 51077 2816 51123 2862
rect 51193 2816 51239 2862
rect 51309 2816 51355 2862
rect 51425 2816 51471 2862
rect 51541 2816 51587 2862
rect 51657 2816 51703 2862
rect 51773 2816 51819 2862
rect 51889 2816 51935 2862
rect 52005 2816 52051 2862
rect 52121 2816 52167 2862
rect 52237 2816 52283 2862
rect 52353 2816 52399 2862
rect 52469 2816 52515 2862
rect 52585 2816 52631 2862
rect 52701 2816 52747 2862
rect 52817 2816 52863 2862
rect 52933 2816 52979 2862
rect 53049 2816 53095 2862
rect 53165 2816 53211 2862
rect 53281 2816 53327 2862
rect 53397 2816 53443 2862
rect 53513 2816 53559 2862
rect 53629 2816 53675 2862
rect 53745 2816 53791 2862
rect 53861 2816 53907 2862
rect 53977 2816 54023 2862
rect 54093 2816 54139 2862
rect 54209 2816 54255 2862
rect 54325 2816 54371 2862
rect 54441 2816 54487 2862
rect 54557 2816 54603 2862
rect 54673 2816 54719 2862
rect 54789 2816 54835 2862
rect 54905 2816 54951 2862
rect 55021 2816 55067 2862
rect 55137 2816 55183 2862
rect 55253 2816 55299 2862
rect 55369 2816 55415 2862
rect 55485 2816 55531 2862
rect 55601 2816 55647 2862
rect 55717 2816 55763 2862
rect 55833 2816 55879 2862
rect 55949 2816 55995 2862
rect 56065 2816 56111 2862
rect 56181 2816 56227 2862
rect 56297 2816 56343 2862
rect 56413 2816 56459 2862
rect 56529 2816 56575 2862
rect 50845 2700 50891 2746
rect 50961 2700 51007 2746
rect 51077 2700 51123 2746
rect 51193 2700 51239 2746
rect 51309 2700 51355 2746
rect 51425 2700 51471 2746
rect 51541 2700 51587 2746
rect 51657 2700 51703 2746
rect 51773 2700 51819 2746
rect 51889 2700 51935 2746
rect 52005 2700 52051 2746
rect 52121 2700 52167 2746
rect 52237 2700 52283 2746
rect 52353 2700 52399 2746
rect 52469 2700 52515 2746
rect 52585 2700 52631 2746
rect 52701 2700 52747 2746
rect 52817 2700 52863 2746
rect 52933 2700 52979 2746
rect 53049 2700 53095 2746
rect 53165 2700 53211 2746
rect 53281 2700 53327 2746
rect 53397 2700 53443 2746
rect 53513 2700 53559 2746
rect 53629 2700 53675 2746
rect 53745 2700 53791 2746
rect 53861 2700 53907 2746
rect 53977 2700 54023 2746
rect 54093 2700 54139 2746
rect 54209 2700 54255 2746
rect 54325 2700 54371 2746
rect 54441 2700 54487 2746
rect 54557 2700 54603 2746
rect 54673 2700 54719 2746
rect 54789 2700 54835 2746
rect 54905 2700 54951 2746
rect 55021 2700 55067 2746
rect 55137 2700 55183 2746
rect 55253 2700 55299 2746
rect 55369 2700 55415 2746
rect 55485 2700 55531 2746
rect 55601 2700 55647 2746
rect 55717 2700 55763 2746
rect 55833 2700 55879 2746
rect 55949 2700 55995 2746
rect 56065 2700 56111 2746
rect 56181 2700 56227 2746
rect 56297 2700 56343 2746
rect 56413 2700 56459 2746
rect 56529 2700 56575 2746
rect 50845 2584 50891 2630
rect 50961 2584 51007 2630
rect 51077 2584 51123 2630
rect 51193 2584 51239 2630
rect 51309 2584 51355 2630
rect 51425 2584 51471 2630
rect 51541 2584 51587 2630
rect 51657 2584 51703 2630
rect 51773 2584 51819 2630
rect 51889 2584 51935 2630
rect 52005 2584 52051 2630
rect 52121 2584 52167 2630
rect 52237 2584 52283 2630
rect 52353 2584 52399 2630
rect 52469 2584 52515 2630
rect 52585 2584 52631 2630
rect 52701 2584 52747 2630
rect 52817 2584 52863 2630
rect 52933 2584 52979 2630
rect 53049 2584 53095 2630
rect 53165 2584 53211 2630
rect 53281 2584 53327 2630
rect 53397 2584 53443 2630
rect 53513 2584 53559 2630
rect 53629 2584 53675 2630
rect 53745 2584 53791 2630
rect 53861 2584 53907 2630
rect 53977 2584 54023 2630
rect 54093 2584 54139 2630
rect 54209 2584 54255 2630
rect 54325 2584 54371 2630
rect 54441 2584 54487 2630
rect 54557 2584 54603 2630
rect 54673 2584 54719 2630
rect 54789 2584 54835 2630
rect 54905 2584 54951 2630
rect 55021 2584 55067 2630
rect 55137 2584 55183 2630
rect 55253 2584 55299 2630
rect 55369 2584 55415 2630
rect 55485 2584 55531 2630
rect 55601 2584 55647 2630
rect 55717 2584 55763 2630
rect 55833 2584 55879 2630
rect 55949 2584 55995 2630
rect 56065 2584 56111 2630
rect 56181 2584 56227 2630
rect 56297 2584 56343 2630
rect 56413 2584 56459 2630
rect 56529 2584 56575 2630
rect 50845 2468 50891 2514
rect 50961 2468 51007 2514
rect 51077 2468 51123 2514
rect 51193 2468 51239 2514
rect 51309 2468 51355 2514
rect 51425 2468 51471 2514
rect 51541 2468 51587 2514
rect 51657 2468 51703 2514
rect 51773 2468 51819 2514
rect 51889 2468 51935 2514
rect 52005 2468 52051 2514
rect 52121 2468 52167 2514
rect 52237 2468 52283 2514
rect 52353 2468 52399 2514
rect 52469 2468 52515 2514
rect 52585 2468 52631 2514
rect 52701 2468 52747 2514
rect 52817 2468 52863 2514
rect 52933 2468 52979 2514
rect 53049 2468 53095 2514
rect 53165 2468 53211 2514
rect 53281 2468 53327 2514
rect 53397 2468 53443 2514
rect 53513 2468 53559 2514
rect 53629 2468 53675 2514
rect 53745 2468 53791 2514
rect 53861 2468 53907 2514
rect 53977 2468 54023 2514
rect 54093 2468 54139 2514
rect 54209 2468 54255 2514
rect 54325 2468 54371 2514
rect 54441 2468 54487 2514
rect 54557 2468 54603 2514
rect 54673 2468 54719 2514
rect 54789 2468 54835 2514
rect 54905 2468 54951 2514
rect 55021 2468 55067 2514
rect 55137 2468 55183 2514
rect 55253 2468 55299 2514
rect 55369 2468 55415 2514
rect 55485 2468 55531 2514
rect 55601 2468 55647 2514
rect 55717 2468 55763 2514
rect 55833 2468 55879 2514
rect 55949 2468 55995 2514
rect 56065 2468 56111 2514
rect 56181 2468 56227 2514
rect 56297 2468 56343 2514
rect 56413 2468 56459 2514
rect 56529 2468 56575 2514
rect 50845 2352 50891 2398
rect 50961 2352 51007 2398
rect 51077 2352 51123 2398
rect 51193 2352 51239 2398
rect 51309 2352 51355 2398
rect 51425 2352 51471 2398
rect 51541 2352 51587 2398
rect 51657 2352 51703 2398
rect 51773 2352 51819 2398
rect 51889 2352 51935 2398
rect 52005 2352 52051 2398
rect 52121 2352 52167 2398
rect 52237 2352 52283 2398
rect 52353 2352 52399 2398
rect 52469 2352 52515 2398
rect 52585 2352 52631 2398
rect 52701 2352 52747 2398
rect 52817 2352 52863 2398
rect 52933 2352 52979 2398
rect 53049 2352 53095 2398
rect 53165 2352 53211 2398
rect 53281 2352 53327 2398
rect 53397 2352 53443 2398
rect 53513 2352 53559 2398
rect 53629 2352 53675 2398
rect 53745 2352 53791 2398
rect 53861 2352 53907 2398
rect 53977 2352 54023 2398
rect 54093 2352 54139 2398
rect 54209 2352 54255 2398
rect 54325 2352 54371 2398
rect 54441 2352 54487 2398
rect 54557 2352 54603 2398
rect 54673 2352 54719 2398
rect 54789 2352 54835 2398
rect 54905 2352 54951 2398
rect 55021 2352 55067 2398
rect 55137 2352 55183 2398
rect 55253 2352 55299 2398
rect 55369 2352 55415 2398
rect 55485 2352 55531 2398
rect 55601 2352 55647 2398
rect 55717 2352 55763 2398
rect 55833 2352 55879 2398
rect 55949 2352 55995 2398
rect 56065 2352 56111 2398
rect 56181 2352 56227 2398
rect 56297 2352 56343 2398
rect 56413 2352 56459 2398
rect 56529 2352 56575 2398
rect 50845 2236 50891 2282
rect 50961 2236 51007 2282
rect 51077 2236 51123 2282
rect 51193 2236 51239 2282
rect 51309 2236 51355 2282
rect 51425 2236 51471 2282
rect 51541 2236 51587 2282
rect 51657 2236 51703 2282
rect 51773 2236 51819 2282
rect 51889 2236 51935 2282
rect 52005 2236 52051 2282
rect 52121 2236 52167 2282
rect 52237 2236 52283 2282
rect 52353 2236 52399 2282
rect 52469 2236 52515 2282
rect 52585 2236 52631 2282
rect 52701 2236 52747 2282
rect 52817 2236 52863 2282
rect 52933 2236 52979 2282
rect 53049 2236 53095 2282
rect 53165 2236 53211 2282
rect 53281 2236 53327 2282
rect 53397 2236 53443 2282
rect 53513 2236 53559 2282
rect 53629 2236 53675 2282
rect 53745 2236 53791 2282
rect 53861 2236 53907 2282
rect 53977 2236 54023 2282
rect 54093 2236 54139 2282
rect 54209 2236 54255 2282
rect 54325 2236 54371 2282
rect 54441 2236 54487 2282
rect 54557 2236 54603 2282
rect 54673 2236 54719 2282
rect 54789 2236 54835 2282
rect 54905 2236 54951 2282
rect 55021 2236 55067 2282
rect 55137 2236 55183 2282
rect 55253 2236 55299 2282
rect 55369 2236 55415 2282
rect 55485 2236 55531 2282
rect 55601 2236 55647 2282
rect 55717 2236 55763 2282
rect 55833 2236 55879 2282
rect 55949 2236 55995 2282
rect 56065 2236 56111 2282
rect 56181 2236 56227 2282
rect 56297 2236 56343 2282
rect 56413 2236 56459 2282
rect 56529 2236 56575 2282
rect 50845 2120 50891 2166
rect 50961 2120 51007 2166
rect 51077 2120 51123 2166
rect 51193 2120 51239 2166
rect 51309 2120 51355 2166
rect 51425 2120 51471 2166
rect 51541 2120 51587 2166
rect 51657 2120 51703 2166
rect 51773 2120 51819 2166
rect 51889 2120 51935 2166
rect 52005 2120 52051 2166
rect 52121 2120 52167 2166
rect 52237 2120 52283 2166
rect 52353 2120 52399 2166
rect 52469 2120 52515 2166
rect 52585 2120 52631 2166
rect 52701 2120 52747 2166
rect 52817 2120 52863 2166
rect 52933 2120 52979 2166
rect 53049 2120 53095 2166
rect 53165 2120 53211 2166
rect 53281 2120 53327 2166
rect 53397 2120 53443 2166
rect 53513 2120 53559 2166
rect 53629 2120 53675 2166
rect 53745 2120 53791 2166
rect 53861 2120 53907 2166
rect 53977 2120 54023 2166
rect 54093 2120 54139 2166
rect 54209 2120 54255 2166
rect 54325 2120 54371 2166
rect 54441 2120 54487 2166
rect 54557 2120 54603 2166
rect 54673 2120 54719 2166
rect 54789 2120 54835 2166
rect 54905 2120 54951 2166
rect 55021 2120 55067 2166
rect 55137 2120 55183 2166
rect 55253 2120 55299 2166
rect 55369 2120 55415 2166
rect 55485 2120 55531 2166
rect 55601 2120 55647 2166
rect 55717 2120 55763 2166
rect 55833 2120 55879 2166
rect 55949 2120 55995 2166
rect 56065 2120 56111 2166
rect 56181 2120 56227 2166
rect 56297 2120 56343 2166
rect 56413 2120 56459 2166
rect 56529 2120 56575 2166
rect 50845 2004 50891 2050
rect 50961 2004 51007 2050
rect 51077 2004 51123 2050
rect 51193 2004 51239 2050
rect 51309 2004 51355 2050
rect 51425 2004 51471 2050
rect 51541 2004 51587 2050
rect 51657 2004 51703 2050
rect 51773 2004 51819 2050
rect 51889 2004 51935 2050
rect 52005 2004 52051 2050
rect 52121 2004 52167 2050
rect 52237 2004 52283 2050
rect 52353 2004 52399 2050
rect 52469 2004 52515 2050
rect 52585 2004 52631 2050
rect 52701 2004 52747 2050
rect 52817 2004 52863 2050
rect 52933 2004 52979 2050
rect 53049 2004 53095 2050
rect 53165 2004 53211 2050
rect 53281 2004 53327 2050
rect 53397 2004 53443 2050
rect 53513 2004 53559 2050
rect 53629 2004 53675 2050
rect 53745 2004 53791 2050
rect 53861 2004 53907 2050
rect 53977 2004 54023 2050
rect 54093 2004 54139 2050
rect 54209 2004 54255 2050
rect 54325 2004 54371 2050
rect 54441 2004 54487 2050
rect 54557 2004 54603 2050
rect 54673 2004 54719 2050
rect 54789 2004 54835 2050
rect 54905 2004 54951 2050
rect 55021 2004 55067 2050
rect 55137 2004 55183 2050
rect 55253 2004 55299 2050
rect 55369 2004 55415 2050
rect 55485 2004 55531 2050
rect 55601 2004 55647 2050
rect 55717 2004 55763 2050
rect 55833 2004 55879 2050
rect 55949 2004 55995 2050
rect 56065 2004 56111 2050
rect 56181 2004 56227 2050
rect 56297 2004 56343 2050
rect 56413 2004 56459 2050
rect 56529 2004 56575 2050
rect 50845 1888 50891 1934
rect 50961 1888 51007 1934
rect 51077 1888 51123 1934
rect 51193 1888 51239 1934
rect 51309 1888 51355 1934
rect 51425 1888 51471 1934
rect 51541 1888 51587 1934
rect 51657 1888 51703 1934
rect 51773 1888 51819 1934
rect 51889 1888 51935 1934
rect 52005 1888 52051 1934
rect 52121 1888 52167 1934
rect 52237 1888 52283 1934
rect 52353 1888 52399 1934
rect 52469 1888 52515 1934
rect 52585 1888 52631 1934
rect 52701 1888 52747 1934
rect 52817 1888 52863 1934
rect 52933 1888 52979 1934
rect 53049 1888 53095 1934
rect 53165 1888 53211 1934
rect 53281 1888 53327 1934
rect 53397 1888 53443 1934
rect 53513 1888 53559 1934
rect 53629 1888 53675 1934
rect 53745 1888 53791 1934
rect 53861 1888 53907 1934
rect 53977 1888 54023 1934
rect 54093 1888 54139 1934
rect 54209 1888 54255 1934
rect 54325 1888 54371 1934
rect 54441 1888 54487 1934
rect 54557 1888 54603 1934
rect 54673 1888 54719 1934
rect 54789 1888 54835 1934
rect 54905 1888 54951 1934
rect 55021 1888 55067 1934
rect 55137 1888 55183 1934
rect 55253 1888 55299 1934
rect 55369 1888 55415 1934
rect 55485 1888 55531 1934
rect 55601 1888 55647 1934
rect 55717 1888 55763 1934
rect 55833 1888 55879 1934
rect 55949 1888 55995 1934
rect 56065 1888 56111 1934
rect 56181 1888 56227 1934
rect 56297 1888 56343 1934
rect 56413 1888 56459 1934
rect 56529 1888 56575 1934
rect 50845 1772 50891 1818
rect 50961 1772 51007 1818
rect 51077 1772 51123 1818
rect 51193 1772 51239 1818
rect 51309 1772 51355 1818
rect 51425 1772 51471 1818
rect 51541 1772 51587 1818
rect 51657 1772 51703 1818
rect 51773 1772 51819 1818
rect 51889 1772 51935 1818
rect 52005 1772 52051 1818
rect 52121 1772 52167 1818
rect 52237 1772 52283 1818
rect 52353 1772 52399 1818
rect 52469 1772 52515 1818
rect 52585 1772 52631 1818
rect 52701 1772 52747 1818
rect 52817 1772 52863 1818
rect 52933 1772 52979 1818
rect 53049 1772 53095 1818
rect 53165 1772 53211 1818
rect 53281 1772 53327 1818
rect 53397 1772 53443 1818
rect 53513 1772 53559 1818
rect 53629 1772 53675 1818
rect 53745 1772 53791 1818
rect 53861 1772 53907 1818
rect 53977 1772 54023 1818
rect 54093 1772 54139 1818
rect 54209 1772 54255 1818
rect 54325 1772 54371 1818
rect 54441 1772 54487 1818
rect 54557 1772 54603 1818
rect 54673 1772 54719 1818
rect 54789 1772 54835 1818
rect 54905 1772 54951 1818
rect 55021 1772 55067 1818
rect 55137 1772 55183 1818
rect 55253 1772 55299 1818
rect 55369 1772 55415 1818
rect 55485 1772 55531 1818
rect 55601 1772 55647 1818
rect 55717 1772 55763 1818
rect 55833 1772 55879 1818
rect 55949 1772 55995 1818
rect 56065 1772 56111 1818
rect 56181 1772 56227 1818
rect 56297 1772 56343 1818
rect 56413 1772 56459 1818
rect 56529 1772 56575 1818
rect 50845 1656 50891 1702
rect 50961 1656 51007 1702
rect 51077 1656 51123 1702
rect 51193 1656 51239 1702
rect 51309 1656 51355 1702
rect 51425 1656 51471 1702
rect 51541 1656 51587 1702
rect 51657 1656 51703 1702
rect 51773 1656 51819 1702
rect 51889 1656 51935 1702
rect 52005 1656 52051 1702
rect 52121 1656 52167 1702
rect 52237 1656 52283 1702
rect 52353 1656 52399 1702
rect 52469 1656 52515 1702
rect 52585 1656 52631 1702
rect 52701 1656 52747 1702
rect 52817 1656 52863 1702
rect 52933 1656 52979 1702
rect 53049 1656 53095 1702
rect 53165 1656 53211 1702
rect 53281 1656 53327 1702
rect 53397 1656 53443 1702
rect 53513 1656 53559 1702
rect 53629 1656 53675 1702
rect 53745 1656 53791 1702
rect 53861 1656 53907 1702
rect 53977 1656 54023 1702
rect 54093 1656 54139 1702
rect 54209 1656 54255 1702
rect 54325 1656 54371 1702
rect 54441 1656 54487 1702
rect 54557 1656 54603 1702
rect 54673 1656 54719 1702
rect 54789 1656 54835 1702
rect 54905 1656 54951 1702
rect 55021 1656 55067 1702
rect 55137 1656 55183 1702
rect 55253 1656 55299 1702
rect 55369 1656 55415 1702
rect 55485 1656 55531 1702
rect 55601 1656 55647 1702
rect 55717 1656 55763 1702
rect 55833 1656 55879 1702
rect 55949 1656 55995 1702
rect 56065 1656 56111 1702
rect 56181 1656 56227 1702
rect 56297 1656 56343 1702
rect 56413 1656 56459 1702
rect 56529 1656 56575 1702
rect 57306 1117 57652 96163
rect 85733 1117 86079 96163
rect 371 969 417 1015
rect 495 969 541 1015
rect 619 969 665 1015
rect 743 969 789 1015
rect 867 969 913 1015
rect 991 969 1037 1015
rect 1115 969 1161 1015
rect 1239 969 1285 1015
rect 1363 969 1409 1015
rect 1487 969 1533 1015
rect 1611 969 1657 1015
rect 1735 969 1781 1015
rect 1859 969 1905 1015
rect 1983 969 2029 1015
rect 2107 969 2153 1015
rect 2231 969 2277 1015
rect 2355 969 2401 1015
rect 2479 969 2525 1015
rect 2603 969 2649 1015
rect 2727 969 2773 1015
rect 2851 969 2897 1015
rect 2975 969 3021 1015
rect 3099 969 3145 1015
rect 3223 969 3269 1015
rect 3347 969 3393 1015
rect 3471 969 3517 1015
rect 3595 969 3641 1015
rect 3719 969 3765 1015
rect 3843 969 3889 1015
rect 3967 969 4013 1015
rect 4091 969 4137 1015
rect 4215 969 4261 1015
rect 4339 969 4385 1015
rect 4463 969 4509 1015
rect 4587 969 4633 1015
rect 4711 969 4757 1015
rect 4835 969 4881 1015
rect 4959 969 5005 1015
rect 5083 969 5129 1015
rect 5207 969 5253 1015
rect 5331 969 5377 1015
rect 5455 969 5501 1015
rect 5579 969 5625 1015
rect 5703 969 5749 1015
rect 5827 969 5873 1015
rect 5951 969 5997 1015
rect 6075 969 6121 1015
rect 6199 969 6245 1015
rect 6323 969 6369 1015
rect 6447 969 6493 1015
rect 6571 969 6617 1015
rect 6695 969 6741 1015
rect 6819 969 6865 1015
rect 6943 969 6989 1015
rect 7067 969 7113 1015
rect 7191 969 7237 1015
rect 7315 969 7361 1015
rect 7439 969 7485 1015
rect 7563 969 7609 1015
rect 7687 969 7733 1015
rect 7811 969 7857 1015
rect 7935 969 7981 1015
rect 8059 969 8105 1015
rect 8183 969 8229 1015
rect 8307 969 8353 1015
rect 8431 969 8477 1015
rect 8555 969 8601 1015
rect 8679 969 8725 1015
rect 8803 969 8849 1015
rect 8927 969 8973 1015
rect 9051 969 9097 1015
rect 9175 969 9221 1015
rect 9299 969 9345 1015
rect 9423 969 9469 1015
rect 9547 969 9593 1015
rect 9671 969 9717 1015
rect 9795 969 9841 1015
rect 9919 969 9965 1015
rect 10043 969 10089 1015
rect 10167 969 10213 1015
rect 10291 969 10337 1015
rect 10415 969 10461 1015
rect 10539 969 10585 1015
rect 10663 969 10709 1015
rect 10787 969 10833 1015
rect 10911 969 10957 1015
rect 11035 969 11081 1015
rect 11159 969 11205 1015
rect 11283 969 11329 1015
rect 11407 969 11453 1015
rect 11531 969 11577 1015
rect 11655 969 11701 1015
rect 11779 969 11825 1015
rect 11903 969 11949 1015
rect 12027 969 12073 1015
rect 12151 969 12197 1015
rect 12275 969 12321 1015
rect 12399 969 12445 1015
rect 12523 969 12569 1015
rect 12647 969 12693 1015
rect 12771 969 12817 1015
rect 12895 969 12941 1015
rect 13019 969 13065 1015
rect 13143 969 13189 1015
rect 13267 969 13313 1015
rect 13391 969 13437 1015
rect 13515 969 13561 1015
rect 13639 969 13685 1015
rect 13763 969 13809 1015
rect 13887 969 13933 1015
rect 14011 969 14057 1015
rect 14135 969 14181 1015
rect 14259 969 14305 1015
rect 14383 969 14429 1015
rect 14507 969 14553 1015
rect 14631 969 14677 1015
rect 14755 969 14801 1015
rect 14879 969 14925 1015
rect 15003 969 15049 1015
rect 15127 969 15173 1015
rect 15251 969 15297 1015
rect 15375 969 15421 1015
rect 15499 969 15545 1015
rect 15623 969 15669 1015
rect 15747 969 15793 1015
rect 15871 969 15917 1015
rect 15995 969 16041 1015
rect 16119 969 16165 1015
rect 16243 969 16289 1015
rect 16367 969 16413 1015
rect 16491 969 16537 1015
rect 16615 969 16661 1015
rect 16739 969 16785 1015
rect 16863 969 16909 1015
rect 16987 969 17033 1015
rect 17111 969 17157 1015
rect 17235 969 17281 1015
rect 17359 969 17405 1015
rect 17483 969 17529 1015
rect 17607 969 17653 1015
rect 17731 969 17777 1015
rect 17855 969 17901 1015
rect 17979 969 18025 1015
rect 18103 969 18149 1015
rect 18227 969 18273 1015
rect 18351 969 18397 1015
rect 18475 969 18521 1015
rect 18599 969 18645 1015
rect 18723 969 18769 1015
rect 18847 969 18893 1015
rect 18971 969 19017 1015
rect 19095 969 19141 1015
rect 19219 969 19265 1015
rect 19343 969 19389 1015
rect 19467 969 19513 1015
rect 19591 969 19637 1015
rect 19715 969 19761 1015
rect 19839 969 19885 1015
rect 19963 969 20009 1015
rect 20087 969 20133 1015
rect 20211 969 20257 1015
rect 20335 969 20381 1015
rect 20459 969 20505 1015
rect 20583 969 20629 1015
rect 20707 969 20753 1015
rect 20831 969 20877 1015
rect 20955 969 21001 1015
rect 21079 969 21125 1015
rect 21203 969 21249 1015
rect 21327 969 21373 1015
rect 21451 969 21497 1015
rect 21575 969 21621 1015
rect 21699 969 21745 1015
rect 21823 969 21869 1015
rect 21947 969 21993 1015
rect 22071 969 22117 1015
rect 22195 969 22241 1015
rect 22319 969 22365 1015
rect 22443 969 22489 1015
rect 22567 969 22613 1015
rect 22691 969 22737 1015
rect 22815 969 22861 1015
rect 22939 969 22985 1015
rect 23063 969 23109 1015
rect 23187 969 23233 1015
rect 23311 969 23357 1015
rect 23435 969 23481 1015
rect 23559 969 23605 1015
rect 23683 969 23729 1015
rect 23807 969 23853 1015
rect 23931 969 23977 1015
rect 24055 969 24101 1015
rect 24179 969 24225 1015
rect 24303 969 24349 1015
rect 24427 969 24473 1015
rect 24551 969 24597 1015
rect 24675 969 24721 1015
rect 24799 969 24845 1015
rect 24923 969 24969 1015
rect 25047 969 25093 1015
rect 25171 969 25217 1015
rect 25295 969 25341 1015
rect 25419 969 25465 1015
rect 25543 969 25589 1015
rect 25667 969 25713 1015
rect 25791 969 25837 1015
rect 25915 969 25961 1015
rect 26039 969 26085 1015
rect 26163 969 26209 1015
rect 26287 969 26333 1015
rect 26411 969 26457 1015
rect 26535 969 26581 1015
rect 26659 969 26705 1015
rect 26783 969 26829 1015
rect 26907 969 26953 1015
rect 27031 969 27077 1015
rect 27155 969 27201 1015
rect 27279 969 27325 1015
rect 27403 969 27449 1015
rect 27527 969 27573 1015
rect 27651 969 27697 1015
rect 27775 969 27821 1015
rect 27899 969 27945 1015
rect 28023 969 28069 1015
rect 28147 969 28193 1015
rect 28271 969 28317 1015
rect 28395 969 28441 1015
rect 28519 969 28565 1015
rect 28643 969 28689 1015
rect 28767 969 28813 1015
rect 28891 969 28937 1015
rect 29015 969 29061 1015
rect 29139 969 29185 1015
rect 29263 969 29309 1015
rect 29387 969 29433 1015
rect 29511 969 29557 1015
rect 29635 969 29681 1015
rect 29759 969 29805 1015
rect 29883 969 29929 1015
rect 30007 969 30053 1015
rect 30131 969 30177 1015
rect 30255 969 30301 1015
rect 30379 969 30425 1015
rect 30503 969 30549 1015
rect 30627 969 30673 1015
rect 30751 969 30797 1015
rect 30875 969 30921 1015
rect 30999 969 31045 1015
rect 31123 969 31169 1015
rect 31247 969 31293 1015
rect 31371 969 31417 1015
rect 31495 969 31541 1015
rect 31619 969 31665 1015
rect 31743 969 31789 1015
rect 31867 969 31913 1015
rect 31991 969 32037 1015
rect 32115 969 32161 1015
rect 32239 969 32285 1015
rect 32363 969 32409 1015
rect 32487 969 32533 1015
rect 32611 969 32657 1015
rect 32735 969 32781 1015
rect 32859 969 32905 1015
rect 32983 969 33029 1015
rect 33107 969 33153 1015
rect 33231 969 33277 1015
rect 33355 969 33401 1015
rect 33479 969 33525 1015
rect 33603 969 33649 1015
rect 33727 969 33773 1015
rect 33851 969 33897 1015
rect 33975 969 34021 1015
rect 34099 969 34145 1015
rect 34223 969 34269 1015
rect 34347 969 34393 1015
rect 34471 969 34517 1015
rect 34595 969 34641 1015
rect 34719 969 34765 1015
rect 34843 969 34889 1015
rect 34967 969 35013 1015
rect 35091 969 35137 1015
rect 35215 969 35261 1015
rect 35339 969 35385 1015
rect 35463 969 35509 1015
rect 35587 969 35633 1015
rect 35711 969 35757 1015
rect 35835 969 35881 1015
rect 35959 969 36005 1015
rect 36083 969 36129 1015
rect 36207 969 36253 1015
rect 36331 969 36377 1015
rect 36455 969 36501 1015
rect 36579 969 36625 1015
rect 36703 969 36749 1015
rect 36827 969 36873 1015
rect 36951 969 36997 1015
rect 37075 969 37121 1015
rect 37199 969 37245 1015
rect 37323 969 37369 1015
rect 37447 969 37493 1015
rect 37571 969 37617 1015
rect 37695 969 37741 1015
rect 37819 969 37865 1015
rect 37943 969 37989 1015
rect 38067 969 38113 1015
rect 38191 969 38237 1015
rect 38315 969 38361 1015
rect 38439 969 38485 1015
rect 38563 969 38609 1015
rect 38687 969 38733 1015
rect 38811 969 38857 1015
rect 38935 969 38981 1015
rect 39059 969 39105 1015
rect 39183 969 39229 1015
rect 39307 969 39353 1015
rect 39431 969 39477 1015
rect 39555 969 39601 1015
rect 39679 969 39725 1015
rect 39803 969 39849 1015
rect 39927 969 39973 1015
rect 40051 969 40097 1015
rect 40175 969 40221 1015
rect 40299 969 40345 1015
rect 40423 969 40469 1015
rect 40547 969 40593 1015
rect 40671 969 40717 1015
rect 40795 969 40841 1015
rect 40919 969 40965 1015
rect 41043 969 41089 1015
rect 41167 969 41213 1015
rect 41291 969 41337 1015
rect 41415 969 41461 1015
rect 41539 969 41585 1015
rect 41663 969 41709 1015
rect 41787 969 41833 1015
rect 41911 969 41957 1015
rect 42035 969 42081 1015
rect 42159 969 42205 1015
rect 42283 969 42329 1015
rect 42407 969 42453 1015
rect 42531 969 42577 1015
rect 42655 969 42701 1015
rect 42779 969 42825 1015
rect 42903 969 42949 1015
rect 43027 969 43073 1015
rect 43151 969 43197 1015
rect 43275 969 43321 1015
rect 43399 969 43445 1015
rect 43523 969 43569 1015
rect 43647 969 43693 1015
rect 43771 969 43817 1015
rect 43895 969 43941 1015
rect 44019 969 44065 1015
rect 44143 969 44189 1015
rect 44267 969 44313 1015
rect 44391 969 44437 1015
rect 44515 969 44561 1015
rect 44639 969 44685 1015
rect 44763 969 44809 1015
rect 44887 969 44933 1015
rect 45011 969 45057 1015
rect 45135 969 45181 1015
rect 45259 969 45305 1015
rect 45383 969 45429 1015
rect 45507 969 45553 1015
rect 45631 969 45677 1015
rect 45755 969 45801 1015
rect 45879 969 45925 1015
rect 46003 969 46049 1015
rect 46127 969 46173 1015
rect 46251 969 46297 1015
rect 46375 969 46421 1015
rect 46499 969 46545 1015
rect 46623 969 46669 1015
rect 46747 969 46793 1015
rect 46871 969 46917 1015
rect 46995 969 47041 1015
rect 47119 969 47165 1015
rect 47243 969 47289 1015
rect 47367 969 47413 1015
rect 47491 969 47537 1015
rect 47615 969 47661 1015
rect 47739 969 47785 1015
rect 47863 969 47909 1015
rect 47987 969 48033 1015
rect 48111 969 48157 1015
rect 48235 969 48281 1015
rect 48359 969 48405 1015
rect 48483 969 48529 1015
rect 48607 969 48653 1015
rect 48731 969 48777 1015
rect 48855 969 48901 1015
rect 48979 969 49025 1015
rect 49103 969 49149 1015
rect 49227 969 49273 1015
rect 49351 969 49397 1015
rect 49475 969 49521 1015
rect 49599 969 49645 1015
rect 49723 969 49769 1015
rect 49847 969 49893 1015
rect 49971 969 50017 1015
rect 50095 969 50141 1015
rect 50219 969 50265 1015
rect 50343 969 50389 1015
rect 50467 969 50513 1015
rect 50591 969 50637 1015
rect 50715 969 50761 1015
rect 50839 969 50885 1015
rect 50963 969 51009 1015
rect 51087 969 51133 1015
rect 51211 969 51257 1015
rect 51335 969 51381 1015
rect 51459 969 51505 1015
rect 51583 969 51629 1015
rect 51707 969 51753 1015
rect 51831 969 51877 1015
rect 51955 969 52001 1015
rect 52079 969 52125 1015
rect 52203 969 52249 1015
rect 52327 969 52373 1015
rect 52451 969 52497 1015
rect 52575 969 52621 1015
rect 52699 969 52745 1015
rect 52823 969 52869 1015
rect 52947 969 52993 1015
rect 53071 969 53117 1015
rect 53195 969 53241 1015
rect 53319 969 53365 1015
rect 53443 969 53489 1015
rect 53567 969 53613 1015
rect 53691 969 53737 1015
rect 53815 969 53861 1015
rect 53939 969 53985 1015
rect 54063 969 54109 1015
rect 54187 969 54233 1015
rect 54311 969 54357 1015
rect 54435 969 54481 1015
rect 54559 969 54605 1015
rect 54683 969 54729 1015
rect 54807 969 54853 1015
rect 54931 969 54977 1015
rect 55055 969 55101 1015
rect 55179 969 55225 1015
rect 55303 969 55349 1015
rect 55427 969 55473 1015
rect 55551 969 55597 1015
rect 55675 969 55721 1015
rect 55799 969 55845 1015
rect 55923 969 55969 1015
rect 56047 969 56093 1015
rect 56171 969 56217 1015
rect 56295 969 56341 1015
rect 56419 969 56465 1015
rect 56543 969 56589 1015
rect 56667 969 56713 1015
rect 56791 969 56837 1015
rect 56915 969 56961 1015
rect 57039 969 57085 1015
rect 57163 969 57209 1015
rect 57287 969 57333 1015
rect 57411 969 57457 1015
rect 57535 969 57581 1015
rect 57659 969 57705 1015
rect 57783 969 57829 1015
rect 57907 969 57953 1015
rect 58031 969 58077 1015
rect 58155 969 58201 1015
rect 58279 969 58325 1015
rect 58403 969 58449 1015
rect 58527 969 58573 1015
rect 58651 969 58697 1015
rect 58775 969 58821 1015
rect 58899 969 58945 1015
rect 59023 969 59069 1015
rect 59147 969 59193 1015
rect 59271 969 59317 1015
rect 59395 969 59441 1015
rect 59519 969 59565 1015
rect 59643 969 59689 1015
rect 59767 969 59813 1015
rect 59891 969 59937 1015
rect 60015 969 60061 1015
rect 60139 969 60185 1015
rect 60263 969 60309 1015
rect 60387 969 60433 1015
rect 60511 969 60557 1015
rect 60635 969 60681 1015
rect 60759 969 60805 1015
rect 60883 969 60929 1015
rect 61007 969 61053 1015
rect 61131 969 61177 1015
rect 61255 969 61301 1015
rect 61379 969 61425 1015
rect 61503 969 61549 1015
rect 61627 969 61673 1015
rect 61751 969 61797 1015
rect 61875 969 61921 1015
rect 61999 969 62045 1015
rect 62123 969 62169 1015
rect 62247 969 62293 1015
rect 62371 969 62417 1015
rect 62495 969 62541 1015
rect 62619 969 62665 1015
rect 62743 969 62789 1015
rect 62867 969 62913 1015
rect 62991 969 63037 1015
rect 63115 969 63161 1015
rect 63239 969 63285 1015
rect 63363 969 63409 1015
rect 63487 969 63533 1015
rect 63611 969 63657 1015
rect 63735 969 63781 1015
rect 63859 969 63905 1015
rect 63983 969 64029 1015
rect 64107 969 64153 1015
rect 64231 969 64277 1015
rect 64355 969 64401 1015
rect 64479 969 64525 1015
rect 64603 969 64649 1015
rect 64727 969 64773 1015
rect 64851 969 64897 1015
rect 64975 969 65021 1015
rect 65099 969 65145 1015
rect 65223 969 65269 1015
rect 65347 969 65393 1015
rect 65471 969 65517 1015
rect 65595 969 65641 1015
rect 65719 969 65765 1015
rect 65843 969 65889 1015
rect 65967 969 66013 1015
rect 66091 969 66137 1015
rect 66215 969 66261 1015
rect 66339 969 66385 1015
rect 66463 969 66509 1015
rect 66587 969 66633 1015
rect 66711 969 66757 1015
rect 66835 969 66881 1015
rect 66959 969 67005 1015
rect 67083 969 67129 1015
rect 67207 969 67253 1015
rect 67331 969 67377 1015
rect 67455 969 67501 1015
rect 67579 969 67625 1015
rect 67703 969 67749 1015
rect 67827 969 67873 1015
rect 67951 969 67997 1015
rect 68075 969 68121 1015
rect 68199 969 68245 1015
rect 68323 969 68369 1015
rect 68447 969 68493 1015
rect 68571 969 68617 1015
rect 68695 969 68741 1015
rect 68819 969 68865 1015
rect 68943 969 68989 1015
rect 69067 969 69113 1015
rect 69191 969 69237 1015
rect 69315 969 69361 1015
rect 69439 969 69485 1015
rect 69563 969 69609 1015
rect 69687 969 69733 1015
rect 69811 969 69857 1015
rect 69935 969 69981 1015
rect 70059 969 70105 1015
rect 70183 969 70229 1015
rect 70307 969 70353 1015
rect 70431 969 70477 1015
rect 70555 969 70601 1015
rect 70679 969 70725 1015
rect 70803 969 70849 1015
rect 70927 969 70973 1015
rect 71051 969 71097 1015
rect 71175 969 71221 1015
rect 71299 969 71345 1015
rect 71423 969 71469 1015
rect 71547 969 71593 1015
rect 71671 969 71717 1015
rect 71795 969 71841 1015
rect 71919 969 71965 1015
rect 72043 969 72089 1015
rect 72167 969 72213 1015
rect 72291 969 72337 1015
rect 72415 969 72461 1015
rect 72539 969 72585 1015
rect 72663 969 72709 1015
rect 72787 969 72833 1015
rect 72911 969 72957 1015
rect 73035 969 73081 1015
rect 73159 969 73205 1015
rect 73283 969 73329 1015
rect 73407 969 73453 1015
rect 73531 969 73577 1015
rect 73655 969 73701 1015
rect 73779 969 73825 1015
rect 73903 969 73949 1015
rect 74027 969 74073 1015
rect 74151 969 74197 1015
rect 74275 969 74321 1015
rect 74399 969 74445 1015
rect 74523 969 74569 1015
rect 74647 969 74693 1015
rect 74771 969 74817 1015
rect 74895 969 74941 1015
rect 75019 969 75065 1015
rect 75143 969 75189 1015
rect 75267 969 75313 1015
rect 75391 969 75437 1015
rect 75515 969 75561 1015
rect 75639 969 75685 1015
rect 75763 969 75809 1015
rect 75887 969 75933 1015
rect 76011 969 76057 1015
rect 76135 969 76181 1015
rect 76259 969 76305 1015
rect 76383 969 76429 1015
rect 76507 969 76553 1015
rect 76631 969 76677 1015
rect 76755 969 76801 1015
rect 76879 969 76925 1015
rect 77003 969 77049 1015
rect 77127 969 77173 1015
rect 77251 969 77297 1015
rect 77375 969 77421 1015
rect 77499 969 77545 1015
rect 77623 969 77669 1015
rect 77747 969 77793 1015
rect 77871 969 77917 1015
rect 77995 969 78041 1015
rect 78119 969 78165 1015
rect 78243 969 78289 1015
rect 78367 969 78413 1015
rect 78491 969 78537 1015
rect 78615 969 78661 1015
rect 78739 969 78785 1015
rect 78863 969 78909 1015
rect 78987 969 79033 1015
rect 79111 969 79157 1015
rect 79235 969 79281 1015
rect 79359 969 79405 1015
rect 79483 969 79529 1015
rect 79607 969 79653 1015
rect 79731 969 79777 1015
rect 79855 969 79901 1015
rect 79979 969 80025 1015
rect 80103 969 80149 1015
rect 80227 969 80273 1015
rect 80351 969 80397 1015
rect 80475 969 80521 1015
rect 80599 969 80645 1015
rect 80723 969 80769 1015
rect 80847 969 80893 1015
rect 80971 969 81017 1015
rect 81095 969 81141 1015
rect 81219 969 81265 1015
rect 81343 969 81389 1015
rect 81467 969 81513 1015
rect 81591 969 81637 1015
rect 81715 969 81761 1015
rect 81839 969 81885 1015
rect 81963 969 82009 1015
rect 82087 969 82133 1015
rect 82211 969 82257 1015
rect 82335 969 82381 1015
rect 82459 969 82505 1015
rect 82583 969 82629 1015
rect 82707 969 82753 1015
rect 82831 969 82877 1015
rect 82955 969 83001 1015
rect 83079 969 83125 1015
rect 83203 969 83249 1015
rect 83327 969 83373 1015
rect 83451 969 83497 1015
rect 83575 969 83621 1015
rect 83699 969 83745 1015
rect 83823 969 83869 1015
rect 83947 969 83993 1015
rect 84071 969 84117 1015
rect 84195 969 84241 1015
rect 84319 969 84365 1015
rect 84443 969 84489 1015
rect 84567 969 84613 1015
rect 84691 969 84737 1015
rect 84815 969 84861 1015
rect 84939 969 84985 1015
rect 85063 969 85109 1015
rect 85187 969 85233 1015
rect 85311 969 85357 1015
rect 85435 969 85481 1015
rect 85559 969 85605 1015
rect 85683 969 85729 1015
rect 85807 969 85853 1015
rect 85931 969 85977 1015
rect 371 845 417 891
rect 495 845 541 891
rect 619 845 665 891
rect 743 845 789 891
rect 867 845 913 891
rect 991 845 1037 891
rect 1115 845 1161 891
rect 1239 845 1285 891
rect 1363 845 1409 891
rect 1487 845 1533 891
rect 1611 845 1657 891
rect 1735 845 1781 891
rect 1859 845 1905 891
rect 1983 845 2029 891
rect 2107 845 2153 891
rect 2231 845 2277 891
rect 2355 845 2401 891
rect 2479 845 2525 891
rect 2603 845 2649 891
rect 2727 845 2773 891
rect 2851 845 2897 891
rect 2975 845 3021 891
rect 3099 845 3145 891
rect 3223 845 3269 891
rect 3347 845 3393 891
rect 3471 845 3517 891
rect 3595 845 3641 891
rect 3719 845 3765 891
rect 3843 845 3889 891
rect 3967 845 4013 891
rect 4091 845 4137 891
rect 4215 845 4261 891
rect 4339 845 4385 891
rect 4463 845 4509 891
rect 4587 845 4633 891
rect 4711 845 4757 891
rect 4835 845 4881 891
rect 4959 845 5005 891
rect 5083 845 5129 891
rect 5207 845 5253 891
rect 5331 845 5377 891
rect 5455 845 5501 891
rect 5579 845 5625 891
rect 5703 845 5749 891
rect 5827 845 5873 891
rect 5951 845 5997 891
rect 6075 845 6121 891
rect 6199 845 6245 891
rect 6323 845 6369 891
rect 6447 845 6493 891
rect 6571 845 6617 891
rect 6695 845 6741 891
rect 6819 845 6865 891
rect 6943 845 6989 891
rect 7067 845 7113 891
rect 7191 845 7237 891
rect 7315 845 7361 891
rect 7439 845 7485 891
rect 7563 845 7609 891
rect 7687 845 7733 891
rect 7811 845 7857 891
rect 7935 845 7981 891
rect 8059 845 8105 891
rect 8183 845 8229 891
rect 8307 845 8353 891
rect 8431 845 8477 891
rect 8555 845 8601 891
rect 8679 845 8725 891
rect 8803 845 8849 891
rect 8927 845 8973 891
rect 9051 845 9097 891
rect 9175 845 9221 891
rect 9299 845 9345 891
rect 9423 845 9469 891
rect 9547 845 9593 891
rect 9671 845 9717 891
rect 9795 845 9841 891
rect 9919 845 9965 891
rect 10043 845 10089 891
rect 10167 845 10213 891
rect 10291 845 10337 891
rect 10415 845 10461 891
rect 10539 845 10585 891
rect 10663 845 10709 891
rect 10787 845 10833 891
rect 10911 845 10957 891
rect 11035 845 11081 891
rect 11159 845 11205 891
rect 11283 845 11329 891
rect 11407 845 11453 891
rect 11531 845 11577 891
rect 11655 845 11701 891
rect 11779 845 11825 891
rect 11903 845 11949 891
rect 12027 845 12073 891
rect 12151 845 12197 891
rect 12275 845 12321 891
rect 12399 845 12445 891
rect 12523 845 12569 891
rect 12647 845 12693 891
rect 12771 845 12817 891
rect 12895 845 12941 891
rect 13019 845 13065 891
rect 13143 845 13189 891
rect 13267 845 13313 891
rect 13391 845 13437 891
rect 13515 845 13561 891
rect 13639 845 13685 891
rect 13763 845 13809 891
rect 13887 845 13933 891
rect 14011 845 14057 891
rect 14135 845 14181 891
rect 14259 845 14305 891
rect 14383 845 14429 891
rect 14507 845 14553 891
rect 14631 845 14677 891
rect 14755 845 14801 891
rect 14879 845 14925 891
rect 15003 845 15049 891
rect 15127 845 15173 891
rect 15251 845 15297 891
rect 15375 845 15421 891
rect 15499 845 15545 891
rect 15623 845 15669 891
rect 15747 845 15793 891
rect 15871 845 15917 891
rect 15995 845 16041 891
rect 16119 845 16165 891
rect 16243 845 16289 891
rect 16367 845 16413 891
rect 16491 845 16537 891
rect 16615 845 16661 891
rect 16739 845 16785 891
rect 16863 845 16909 891
rect 16987 845 17033 891
rect 17111 845 17157 891
rect 17235 845 17281 891
rect 17359 845 17405 891
rect 17483 845 17529 891
rect 17607 845 17653 891
rect 17731 845 17777 891
rect 17855 845 17901 891
rect 17979 845 18025 891
rect 18103 845 18149 891
rect 18227 845 18273 891
rect 18351 845 18397 891
rect 18475 845 18521 891
rect 18599 845 18645 891
rect 18723 845 18769 891
rect 18847 845 18893 891
rect 18971 845 19017 891
rect 19095 845 19141 891
rect 19219 845 19265 891
rect 19343 845 19389 891
rect 19467 845 19513 891
rect 19591 845 19637 891
rect 19715 845 19761 891
rect 19839 845 19885 891
rect 19963 845 20009 891
rect 20087 845 20133 891
rect 20211 845 20257 891
rect 20335 845 20381 891
rect 20459 845 20505 891
rect 20583 845 20629 891
rect 20707 845 20753 891
rect 20831 845 20877 891
rect 20955 845 21001 891
rect 21079 845 21125 891
rect 21203 845 21249 891
rect 21327 845 21373 891
rect 21451 845 21497 891
rect 21575 845 21621 891
rect 21699 845 21745 891
rect 21823 845 21869 891
rect 21947 845 21993 891
rect 22071 845 22117 891
rect 22195 845 22241 891
rect 22319 845 22365 891
rect 22443 845 22489 891
rect 22567 845 22613 891
rect 22691 845 22737 891
rect 22815 845 22861 891
rect 22939 845 22985 891
rect 23063 845 23109 891
rect 23187 845 23233 891
rect 23311 845 23357 891
rect 23435 845 23481 891
rect 23559 845 23605 891
rect 23683 845 23729 891
rect 23807 845 23853 891
rect 23931 845 23977 891
rect 24055 845 24101 891
rect 24179 845 24225 891
rect 24303 845 24349 891
rect 24427 845 24473 891
rect 24551 845 24597 891
rect 24675 845 24721 891
rect 24799 845 24845 891
rect 24923 845 24969 891
rect 25047 845 25093 891
rect 25171 845 25217 891
rect 25295 845 25341 891
rect 25419 845 25465 891
rect 25543 845 25589 891
rect 25667 845 25713 891
rect 25791 845 25837 891
rect 25915 845 25961 891
rect 26039 845 26085 891
rect 26163 845 26209 891
rect 26287 845 26333 891
rect 26411 845 26457 891
rect 26535 845 26581 891
rect 26659 845 26705 891
rect 26783 845 26829 891
rect 26907 845 26953 891
rect 27031 845 27077 891
rect 27155 845 27201 891
rect 27279 845 27325 891
rect 27403 845 27449 891
rect 27527 845 27573 891
rect 27651 845 27697 891
rect 27775 845 27821 891
rect 27899 845 27945 891
rect 28023 845 28069 891
rect 28147 845 28193 891
rect 28271 845 28317 891
rect 28395 845 28441 891
rect 28519 845 28565 891
rect 28643 845 28689 891
rect 28767 845 28813 891
rect 28891 845 28937 891
rect 29015 845 29061 891
rect 29139 845 29185 891
rect 29263 845 29309 891
rect 29387 845 29433 891
rect 29511 845 29557 891
rect 29635 845 29681 891
rect 29759 845 29805 891
rect 29883 845 29929 891
rect 30007 845 30053 891
rect 30131 845 30177 891
rect 30255 845 30301 891
rect 30379 845 30425 891
rect 30503 845 30549 891
rect 30627 845 30673 891
rect 30751 845 30797 891
rect 30875 845 30921 891
rect 30999 845 31045 891
rect 31123 845 31169 891
rect 31247 845 31293 891
rect 31371 845 31417 891
rect 31495 845 31541 891
rect 31619 845 31665 891
rect 31743 845 31789 891
rect 31867 845 31913 891
rect 31991 845 32037 891
rect 32115 845 32161 891
rect 32239 845 32285 891
rect 32363 845 32409 891
rect 32487 845 32533 891
rect 32611 845 32657 891
rect 32735 845 32781 891
rect 32859 845 32905 891
rect 32983 845 33029 891
rect 33107 845 33153 891
rect 33231 845 33277 891
rect 33355 845 33401 891
rect 33479 845 33525 891
rect 33603 845 33649 891
rect 33727 845 33773 891
rect 33851 845 33897 891
rect 33975 845 34021 891
rect 34099 845 34145 891
rect 34223 845 34269 891
rect 34347 845 34393 891
rect 34471 845 34517 891
rect 34595 845 34641 891
rect 34719 845 34765 891
rect 34843 845 34889 891
rect 34967 845 35013 891
rect 35091 845 35137 891
rect 35215 845 35261 891
rect 35339 845 35385 891
rect 35463 845 35509 891
rect 35587 845 35633 891
rect 35711 845 35757 891
rect 35835 845 35881 891
rect 35959 845 36005 891
rect 36083 845 36129 891
rect 36207 845 36253 891
rect 36331 845 36377 891
rect 36455 845 36501 891
rect 36579 845 36625 891
rect 36703 845 36749 891
rect 36827 845 36873 891
rect 36951 845 36997 891
rect 37075 845 37121 891
rect 37199 845 37245 891
rect 37323 845 37369 891
rect 37447 845 37493 891
rect 37571 845 37617 891
rect 37695 845 37741 891
rect 37819 845 37865 891
rect 37943 845 37989 891
rect 38067 845 38113 891
rect 38191 845 38237 891
rect 38315 845 38361 891
rect 38439 845 38485 891
rect 38563 845 38609 891
rect 38687 845 38733 891
rect 38811 845 38857 891
rect 38935 845 38981 891
rect 39059 845 39105 891
rect 39183 845 39229 891
rect 39307 845 39353 891
rect 39431 845 39477 891
rect 39555 845 39601 891
rect 39679 845 39725 891
rect 39803 845 39849 891
rect 39927 845 39973 891
rect 40051 845 40097 891
rect 40175 845 40221 891
rect 40299 845 40345 891
rect 40423 845 40469 891
rect 40547 845 40593 891
rect 40671 845 40717 891
rect 40795 845 40841 891
rect 40919 845 40965 891
rect 41043 845 41089 891
rect 41167 845 41213 891
rect 41291 845 41337 891
rect 41415 845 41461 891
rect 41539 845 41585 891
rect 41663 845 41709 891
rect 41787 845 41833 891
rect 41911 845 41957 891
rect 42035 845 42081 891
rect 42159 845 42205 891
rect 42283 845 42329 891
rect 42407 845 42453 891
rect 42531 845 42577 891
rect 42655 845 42701 891
rect 42779 845 42825 891
rect 42903 845 42949 891
rect 43027 845 43073 891
rect 43151 845 43197 891
rect 43275 845 43321 891
rect 43399 845 43445 891
rect 43523 845 43569 891
rect 43647 845 43693 891
rect 43771 845 43817 891
rect 43895 845 43941 891
rect 44019 845 44065 891
rect 44143 845 44189 891
rect 44267 845 44313 891
rect 44391 845 44437 891
rect 44515 845 44561 891
rect 44639 845 44685 891
rect 44763 845 44809 891
rect 44887 845 44933 891
rect 45011 845 45057 891
rect 45135 845 45181 891
rect 45259 845 45305 891
rect 45383 845 45429 891
rect 45507 845 45553 891
rect 45631 845 45677 891
rect 45755 845 45801 891
rect 45879 845 45925 891
rect 46003 845 46049 891
rect 46127 845 46173 891
rect 46251 845 46297 891
rect 46375 845 46421 891
rect 46499 845 46545 891
rect 46623 845 46669 891
rect 46747 845 46793 891
rect 46871 845 46917 891
rect 46995 845 47041 891
rect 47119 845 47165 891
rect 47243 845 47289 891
rect 47367 845 47413 891
rect 47491 845 47537 891
rect 47615 845 47661 891
rect 47739 845 47785 891
rect 47863 845 47909 891
rect 47987 845 48033 891
rect 48111 845 48157 891
rect 48235 845 48281 891
rect 48359 845 48405 891
rect 48483 845 48529 891
rect 48607 845 48653 891
rect 48731 845 48777 891
rect 48855 845 48901 891
rect 48979 845 49025 891
rect 49103 845 49149 891
rect 49227 845 49273 891
rect 49351 845 49397 891
rect 49475 845 49521 891
rect 49599 845 49645 891
rect 49723 845 49769 891
rect 49847 845 49893 891
rect 49971 845 50017 891
rect 50095 845 50141 891
rect 50219 845 50265 891
rect 50343 845 50389 891
rect 50467 845 50513 891
rect 50591 845 50637 891
rect 50715 845 50761 891
rect 50839 845 50885 891
rect 50963 845 51009 891
rect 51087 845 51133 891
rect 51211 845 51257 891
rect 51335 845 51381 891
rect 51459 845 51505 891
rect 51583 845 51629 891
rect 51707 845 51753 891
rect 51831 845 51877 891
rect 51955 845 52001 891
rect 52079 845 52125 891
rect 52203 845 52249 891
rect 52327 845 52373 891
rect 52451 845 52497 891
rect 52575 845 52621 891
rect 52699 845 52745 891
rect 52823 845 52869 891
rect 52947 845 52993 891
rect 53071 845 53117 891
rect 53195 845 53241 891
rect 53319 845 53365 891
rect 53443 845 53489 891
rect 53567 845 53613 891
rect 53691 845 53737 891
rect 53815 845 53861 891
rect 53939 845 53985 891
rect 54063 845 54109 891
rect 54187 845 54233 891
rect 54311 845 54357 891
rect 54435 845 54481 891
rect 54559 845 54605 891
rect 54683 845 54729 891
rect 54807 845 54853 891
rect 54931 845 54977 891
rect 55055 845 55101 891
rect 55179 845 55225 891
rect 55303 845 55349 891
rect 55427 845 55473 891
rect 55551 845 55597 891
rect 55675 845 55721 891
rect 55799 845 55845 891
rect 55923 845 55969 891
rect 56047 845 56093 891
rect 56171 845 56217 891
rect 56295 845 56341 891
rect 56419 845 56465 891
rect 56543 845 56589 891
rect 56667 845 56713 891
rect 56791 845 56837 891
rect 56915 845 56961 891
rect 57039 845 57085 891
rect 57163 845 57209 891
rect 57287 845 57333 891
rect 57411 845 57457 891
rect 57535 845 57581 891
rect 57659 845 57705 891
rect 57783 845 57829 891
rect 57907 845 57953 891
rect 58031 845 58077 891
rect 58155 845 58201 891
rect 58279 845 58325 891
rect 58403 845 58449 891
rect 58527 845 58573 891
rect 58651 845 58697 891
rect 58775 845 58821 891
rect 58899 845 58945 891
rect 59023 845 59069 891
rect 59147 845 59193 891
rect 59271 845 59317 891
rect 59395 845 59441 891
rect 59519 845 59565 891
rect 59643 845 59689 891
rect 59767 845 59813 891
rect 59891 845 59937 891
rect 60015 845 60061 891
rect 60139 845 60185 891
rect 60263 845 60309 891
rect 60387 845 60433 891
rect 60511 845 60557 891
rect 60635 845 60681 891
rect 60759 845 60805 891
rect 60883 845 60929 891
rect 61007 845 61053 891
rect 61131 845 61177 891
rect 61255 845 61301 891
rect 61379 845 61425 891
rect 61503 845 61549 891
rect 61627 845 61673 891
rect 61751 845 61797 891
rect 61875 845 61921 891
rect 61999 845 62045 891
rect 62123 845 62169 891
rect 62247 845 62293 891
rect 62371 845 62417 891
rect 62495 845 62541 891
rect 62619 845 62665 891
rect 62743 845 62789 891
rect 62867 845 62913 891
rect 62991 845 63037 891
rect 63115 845 63161 891
rect 63239 845 63285 891
rect 63363 845 63409 891
rect 63487 845 63533 891
rect 63611 845 63657 891
rect 63735 845 63781 891
rect 63859 845 63905 891
rect 63983 845 64029 891
rect 64107 845 64153 891
rect 64231 845 64277 891
rect 64355 845 64401 891
rect 64479 845 64525 891
rect 64603 845 64649 891
rect 64727 845 64773 891
rect 64851 845 64897 891
rect 64975 845 65021 891
rect 65099 845 65145 891
rect 65223 845 65269 891
rect 65347 845 65393 891
rect 65471 845 65517 891
rect 65595 845 65641 891
rect 65719 845 65765 891
rect 65843 845 65889 891
rect 65967 845 66013 891
rect 66091 845 66137 891
rect 66215 845 66261 891
rect 66339 845 66385 891
rect 66463 845 66509 891
rect 66587 845 66633 891
rect 66711 845 66757 891
rect 66835 845 66881 891
rect 66959 845 67005 891
rect 67083 845 67129 891
rect 67207 845 67253 891
rect 67331 845 67377 891
rect 67455 845 67501 891
rect 67579 845 67625 891
rect 67703 845 67749 891
rect 67827 845 67873 891
rect 67951 845 67997 891
rect 68075 845 68121 891
rect 68199 845 68245 891
rect 68323 845 68369 891
rect 68447 845 68493 891
rect 68571 845 68617 891
rect 68695 845 68741 891
rect 68819 845 68865 891
rect 68943 845 68989 891
rect 69067 845 69113 891
rect 69191 845 69237 891
rect 69315 845 69361 891
rect 69439 845 69485 891
rect 69563 845 69609 891
rect 69687 845 69733 891
rect 69811 845 69857 891
rect 69935 845 69981 891
rect 70059 845 70105 891
rect 70183 845 70229 891
rect 70307 845 70353 891
rect 70431 845 70477 891
rect 70555 845 70601 891
rect 70679 845 70725 891
rect 70803 845 70849 891
rect 70927 845 70973 891
rect 71051 845 71097 891
rect 71175 845 71221 891
rect 71299 845 71345 891
rect 71423 845 71469 891
rect 71547 845 71593 891
rect 71671 845 71717 891
rect 71795 845 71841 891
rect 71919 845 71965 891
rect 72043 845 72089 891
rect 72167 845 72213 891
rect 72291 845 72337 891
rect 72415 845 72461 891
rect 72539 845 72585 891
rect 72663 845 72709 891
rect 72787 845 72833 891
rect 72911 845 72957 891
rect 73035 845 73081 891
rect 73159 845 73205 891
rect 73283 845 73329 891
rect 73407 845 73453 891
rect 73531 845 73577 891
rect 73655 845 73701 891
rect 73779 845 73825 891
rect 73903 845 73949 891
rect 74027 845 74073 891
rect 74151 845 74197 891
rect 74275 845 74321 891
rect 74399 845 74445 891
rect 74523 845 74569 891
rect 74647 845 74693 891
rect 74771 845 74817 891
rect 74895 845 74941 891
rect 75019 845 75065 891
rect 75143 845 75189 891
rect 75267 845 75313 891
rect 75391 845 75437 891
rect 75515 845 75561 891
rect 75639 845 75685 891
rect 75763 845 75809 891
rect 75887 845 75933 891
rect 76011 845 76057 891
rect 76135 845 76181 891
rect 76259 845 76305 891
rect 76383 845 76429 891
rect 76507 845 76553 891
rect 76631 845 76677 891
rect 76755 845 76801 891
rect 76879 845 76925 891
rect 77003 845 77049 891
rect 77127 845 77173 891
rect 77251 845 77297 891
rect 77375 845 77421 891
rect 77499 845 77545 891
rect 77623 845 77669 891
rect 77747 845 77793 891
rect 77871 845 77917 891
rect 77995 845 78041 891
rect 78119 845 78165 891
rect 78243 845 78289 891
rect 78367 845 78413 891
rect 78491 845 78537 891
rect 78615 845 78661 891
rect 78739 845 78785 891
rect 78863 845 78909 891
rect 78987 845 79033 891
rect 79111 845 79157 891
rect 79235 845 79281 891
rect 79359 845 79405 891
rect 79483 845 79529 891
rect 79607 845 79653 891
rect 79731 845 79777 891
rect 79855 845 79901 891
rect 79979 845 80025 891
rect 80103 845 80149 891
rect 80227 845 80273 891
rect 80351 845 80397 891
rect 80475 845 80521 891
rect 80599 845 80645 891
rect 80723 845 80769 891
rect 80847 845 80893 891
rect 80971 845 81017 891
rect 81095 845 81141 891
rect 81219 845 81265 891
rect 81343 845 81389 891
rect 81467 845 81513 891
rect 81591 845 81637 891
rect 81715 845 81761 891
rect 81839 845 81885 891
rect 81963 845 82009 891
rect 82087 845 82133 891
rect 82211 845 82257 891
rect 82335 845 82381 891
rect 82459 845 82505 891
rect 82583 845 82629 891
rect 82707 845 82753 891
rect 82831 845 82877 891
rect 82955 845 83001 891
rect 83079 845 83125 891
rect 83203 845 83249 891
rect 83327 845 83373 891
rect 83451 845 83497 891
rect 83575 845 83621 891
rect 83699 845 83745 891
rect 83823 845 83869 891
rect 83947 845 83993 891
rect 84071 845 84117 891
rect 84195 845 84241 891
rect 84319 845 84365 891
rect 84443 845 84489 891
rect 84567 845 84613 891
rect 84691 845 84737 891
rect 84815 845 84861 891
rect 84939 845 84985 891
rect 85063 845 85109 891
rect 85187 845 85233 891
rect 85311 845 85357 891
rect 85435 845 85481 891
rect 85559 845 85605 891
rect 85683 845 85729 891
rect 85807 845 85853 891
rect 85931 845 85977 891
rect 371 721 417 767
rect 495 721 541 767
rect 619 721 665 767
rect 743 721 789 767
rect 867 721 913 767
rect 991 721 1037 767
rect 1115 721 1161 767
rect 1239 721 1285 767
rect 1363 721 1409 767
rect 1487 721 1533 767
rect 1611 721 1657 767
rect 1735 721 1781 767
rect 1859 721 1905 767
rect 1983 721 2029 767
rect 2107 721 2153 767
rect 2231 721 2277 767
rect 2355 721 2401 767
rect 2479 721 2525 767
rect 2603 721 2649 767
rect 2727 721 2773 767
rect 2851 721 2897 767
rect 2975 721 3021 767
rect 3099 721 3145 767
rect 3223 721 3269 767
rect 3347 721 3393 767
rect 3471 721 3517 767
rect 3595 721 3641 767
rect 3719 721 3765 767
rect 3843 721 3889 767
rect 3967 721 4013 767
rect 4091 721 4137 767
rect 4215 721 4261 767
rect 4339 721 4385 767
rect 4463 721 4509 767
rect 4587 721 4633 767
rect 4711 721 4757 767
rect 4835 721 4881 767
rect 4959 721 5005 767
rect 5083 721 5129 767
rect 5207 721 5253 767
rect 5331 721 5377 767
rect 5455 721 5501 767
rect 5579 721 5625 767
rect 5703 721 5749 767
rect 5827 721 5873 767
rect 5951 721 5997 767
rect 6075 721 6121 767
rect 6199 721 6245 767
rect 6323 721 6369 767
rect 6447 721 6493 767
rect 6571 721 6617 767
rect 6695 721 6741 767
rect 6819 721 6865 767
rect 6943 721 6989 767
rect 7067 721 7113 767
rect 7191 721 7237 767
rect 7315 721 7361 767
rect 7439 721 7485 767
rect 7563 721 7609 767
rect 7687 721 7733 767
rect 7811 721 7857 767
rect 7935 721 7981 767
rect 8059 721 8105 767
rect 8183 721 8229 767
rect 8307 721 8353 767
rect 8431 721 8477 767
rect 8555 721 8601 767
rect 8679 721 8725 767
rect 8803 721 8849 767
rect 8927 721 8973 767
rect 9051 721 9097 767
rect 9175 721 9221 767
rect 9299 721 9345 767
rect 9423 721 9469 767
rect 9547 721 9593 767
rect 9671 721 9717 767
rect 9795 721 9841 767
rect 9919 721 9965 767
rect 10043 721 10089 767
rect 10167 721 10213 767
rect 10291 721 10337 767
rect 10415 721 10461 767
rect 10539 721 10585 767
rect 10663 721 10709 767
rect 10787 721 10833 767
rect 10911 721 10957 767
rect 11035 721 11081 767
rect 11159 721 11205 767
rect 11283 721 11329 767
rect 11407 721 11453 767
rect 11531 721 11577 767
rect 11655 721 11701 767
rect 11779 721 11825 767
rect 11903 721 11949 767
rect 12027 721 12073 767
rect 12151 721 12197 767
rect 12275 721 12321 767
rect 12399 721 12445 767
rect 12523 721 12569 767
rect 12647 721 12693 767
rect 12771 721 12817 767
rect 12895 721 12941 767
rect 13019 721 13065 767
rect 13143 721 13189 767
rect 13267 721 13313 767
rect 13391 721 13437 767
rect 13515 721 13561 767
rect 13639 721 13685 767
rect 13763 721 13809 767
rect 13887 721 13933 767
rect 14011 721 14057 767
rect 14135 721 14181 767
rect 14259 721 14305 767
rect 14383 721 14429 767
rect 14507 721 14553 767
rect 14631 721 14677 767
rect 14755 721 14801 767
rect 14879 721 14925 767
rect 15003 721 15049 767
rect 15127 721 15173 767
rect 15251 721 15297 767
rect 15375 721 15421 767
rect 15499 721 15545 767
rect 15623 721 15669 767
rect 15747 721 15793 767
rect 15871 721 15917 767
rect 15995 721 16041 767
rect 16119 721 16165 767
rect 16243 721 16289 767
rect 16367 721 16413 767
rect 16491 721 16537 767
rect 16615 721 16661 767
rect 16739 721 16785 767
rect 16863 721 16909 767
rect 16987 721 17033 767
rect 17111 721 17157 767
rect 17235 721 17281 767
rect 17359 721 17405 767
rect 17483 721 17529 767
rect 17607 721 17653 767
rect 17731 721 17777 767
rect 17855 721 17901 767
rect 17979 721 18025 767
rect 18103 721 18149 767
rect 18227 721 18273 767
rect 18351 721 18397 767
rect 18475 721 18521 767
rect 18599 721 18645 767
rect 18723 721 18769 767
rect 18847 721 18893 767
rect 18971 721 19017 767
rect 19095 721 19141 767
rect 19219 721 19265 767
rect 19343 721 19389 767
rect 19467 721 19513 767
rect 19591 721 19637 767
rect 19715 721 19761 767
rect 19839 721 19885 767
rect 19963 721 20009 767
rect 20087 721 20133 767
rect 20211 721 20257 767
rect 20335 721 20381 767
rect 20459 721 20505 767
rect 20583 721 20629 767
rect 20707 721 20753 767
rect 20831 721 20877 767
rect 20955 721 21001 767
rect 21079 721 21125 767
rect 21203 721 21249 767
rect 21327 721 21373 767
rect 21451 721 21497 767
rect 21575 721 21621 767
rect 21699 721 21745 767
rect 21823 721 21869 767
rect 21947 721 21993 767
rect 22071 721 22117 767
rect 22195 721 22241 767
rect 22319 721 22365 767
rect 22443 721 22489 767
rect 22567 721 22613 767
rect 22691 721 22737 767
rect 22815 721 22861 767
rect 22939 721 22985 767
rect 23063 721 23109 767
rect 23187 721 23233 767
rect 23311 721 23357 767
rect 23435 721 23481 767
rect 23559 721 23605 767
rect 23683 721 23729 767
rect 23807 721 23853 767
rect 23931 721 23977 767
rect 24055 721 24101 767
rect 24179 721 24225 767
rect 24303 721 24349 767
rect 24427 721 24473 767
rect 24551 721 24597 767
rect 24675 721 24721 767
rect 24799 721 24845 767
rect 24923 721 24969 767
rect 25047 721 25093 767
rect 25171 721 25217 767
rect 25295 721 25341 767
rect 25419 721 25465 767
rect 25543 721 25589 767
rect 25667 721 25713 767
rect 25791 721 25837 767
rect 25915 721 25961 767
rect 26039 721 26085 767
rect 26163 721 26209 767
rect 26287 721 26333 767
rect 26411 721 26457 767
rect 26535 721 26581 767
rect 26659 721 26705 767
rect 26783 721 26829 767
rect 26907 721 26953 767
rect 27031 721 27077 767
rect 27155 721 27201 767
rect 27279 721 27325 767
rect 27403 721 27449 767
rect 27527 721 27573 767
rect 27651 721 27697 767
rect 27775 721 27821 767
rect 27899 721 27945 767
rect 28023 721 28069 767
rect 28147 721 28193 767
rect 28271 721 28317 767
rect 28395 721 28441 767
rect 28519 721 28565 767
rect 28643 721 28689 767
rect 28767 721 28813 767
rect 28891 721 28937 767
rect 29015 721 29061 767
rect 29139 721 29185 767
rect 29263 721 29309 767
rect 29387 721 29433 767
rect 29511 721 29557 767
rect 29635 721 29681 767
rect 29759 721 29805 767
rect 29883 721 29929 767
rect 30007 721 30053 767
rect 30131 721 30177 767
rect 30255 721 30301 767
rect 30379 721 30425 767
rect 30503 721 30549 767
rect 30627 721 30673 767
rect 30751 721 30797 767
rect 30875 721 30921 767
rect 30999 721 31045 767
rect 31123 721 31169 767
rect 31247 721 31293 767
rect 31371 721 31417 767
rect 31495 721 31541 767
rect 31619 721 31665 767
rect 31743 721 31789 767
rect 31867 721 31913 767
rect 31991 721 32037 767
rect 32115 721 32161 767
rect 32239 721 32285 767
rect 32363 721 32409 767
rect 32487 721 32533 767
rect 32611 721 32657 767
rect 32735 721 32781 767
rect 32859 721 32905 767
rect 32983 721 33029 767
rect 33107 721 33153 767
rect 33231 721 33277 767
rect 33355 721 33401 767
rect 33479 721 33525 767
rect 33603 721 33649 767
rect 33727 721 33773 767
rect 33851 721 33897 767
rect 33975 721 34021 767
rect 34099 721 34145 767
rect 34223 721 34269 767
rect 34347 721 34393 767
rect 34471 721 34517 767
rect 34595 721 34641 767
rect 34719 721 34765 767
rect 34843 721 34889 767
rect 34967 721 35013 767
rect 35091 721 35137 767
rect 35215 721 35261 767
rect 35339 721 35385 767
rect 35463 721 35509 767
rect 35587 721 35633 767
rect 35711 721 35757 767
rect 35835 721 35881 767
rect 35959 721 36005 767
rect 36083 721 36129 767
rect 36207 721 36253 767
rect 36331 721 36377 767
rect 36455 721 36501 767
rect 36579 721 36625 767
rect 36703 721 36749 767
rect 36827 721 36873 767
rect 36951 721 36997 767
rect 37075 721 37121 767
rect 37199 721 37245 767
rect 37323 721 37369 767
rect 37447 721 37493 767
rect 37571 721 37617 767
rect 37695 721 37741 767
rect 37819 721 37865 767
rect 37943 721 37989 767
rect 38067 721 38113 767
rect 38191 721 38237 767
rect 38315 721 38361 767
rect 38439 721 38485 767
rect 38563 721 38609 767
rect 38687 721 38733 767
rect 38811 721 38857 767
rect 38935 721 38981 767
rect 39059 721 39105 767
rect 39183 721 39229 767
rect 39307 721 39353 767
rect 39431 721 39477 767
rect 39555 721 39601 767
rect 39679 721 39725 767
rect 39803 721 39849 767
rect 39927 721 39973 767
rect 40051 721 40097 767
rect 40175 721 40221 767
rect 40299 721 40345 767
rect 40423 721 40469 767
rect 40547 721 40593 767
rect 40671 721 40717 767
rect 40795 721 40841 767
rect 40919 721 40965 767
rect 41043 721 41089 767
rect 41167 721 41213 767
rect 41291 721 41337 767
rect 41415 721 41461 767
rect 41539 721 41585 767
rect 41663 721 41709 767
rect 41787 721 41833 767
rect 41911 721 41957 767
rect 42035 721 42081 767
rect 42159 721 42205 767
rect 42283 721 42329 767
rect 42407 721 42453 767
rect 42531 721 42577 767
rect 42655 721 42701 767
rect 42779 721 42825 767
rect 42903 721 42949 767
rect 43027 721 43073 767
rect 43151 721 43197 767
rect 43275 721 43321 767
rect 43399 721 43445 767
rect 43523 721 43569 767
rect 43647 721 43693 767
rect 43771 721 43817 767
rect 43895 721 43941 767
rect 44019 721 44065 767
rect 44143 721 44189 767
rect 44267 721 44313 767
rect 44391 721 44437 767
rect 44515 721 44561 767
rect 44639 721 44685 767
rect 44763 721 44809 767
rect 44887 721 44933 767
rect 45011 721 45057 767
rect 45135 721 45181 767
rect 45259 721 45305 767
rect 45383 721 45429 767
rect 45507 721 45553 767
rect 45631 721 45677 767
rect 45755 721 45801 767
rect 45879 721 45925 767
rect 46003 721 46049 767
rect 46127 721 46173 767
rect 46251 721 46297 767
rect 46375 721 46421 767
rect 46499 721 46545 767
rect 46623 721 46669 767
rect 46747 721 46793 767
rect 46871 721 46917 767
rect 46995 721 47041 767
rect 47119 721 47165 767
rect 47243 721 47289 767
rect 47367 721 47413 767
rect 47491 721 47537 767
rect 47615 721 47661 767
rect 47739 721 47785 767
rect 47863 721 47909 767
rect 47987 721 48033 767
rect 48111 721 48157 767
rect 48235 721 48281 767
rect 48359 721 48405 767
rect 48483 721 48529 767
rect 48607 721 48653 767
rect 48731 721 48777 767
rect 48855 721 48901 767
rect 48979 721 49025 767
rect 49103 721 49149 767
rect 49227 721 49273 767
rect 49351 721 49397 767
rect 49475 721 49521 767
rect 49599 721 49645 767
rect 49723 721 49769 767
rect 49847 721 49893 767
rect 49971 721 50017 767
rect 50095 721 50141 767
rect 50219 721 50265 767
rect 50343 721 50389 767
rect 50467 721 50513 767
rect 50591 721 50637 767
rect 50715 721 50761 767
rect 50839 721 50885 767
rect 50963 721 51009 767
rect 51087 721 51133 767
rect 51211 721 51257 767
rect 51335 721 51381 767
rect 51459 721 51505 767
rect 51583 721 51629 767
rect 51707 721 51753 767
rect 51831 721 51877 767
rect 51955 721 52001 767
rect 52079 721 52125 767
rect 52203 721 52249 767
rect 52327 721 52373 767
rect 52451 721 52497 767
rect 52575 721 52621 767
rect 52699 721 52745 767
rect 52823 721 52869 767
rect 52947 721 52993 767
rect 53071 721 53117 767
rect 53195 721 53241 767
rect 53319 721 53365 767
rect 53443 721 53489 767
rect 53567 721 53613 767
rect 53691 721 53737 767
rect 53815 721 53861 767
rect 53939 721 53985 767
rect 54063 721 54109 767
rect 54187 721 54233 767
rect 54311 721 54357 767
rect 54435 721 54481 767
rect 54559 721 54605 767
rect 54683 721 54729 767
rect 54807 721 54853 767
rect 54931 721 54977 767
rect 55055 721 55101 767
rect 55179 721 55225 767
rect 55303 721 55349 767
rect 55427 721 55473 767
rect 55551 721 55597 767
rect 55675 721 55721 767
rect 55799 721 55845 767
rect 55923 721 55969 767
rect 56047 721 56093 767
rect 56171 721 56217 767
rect 56295 721 56341 767
rect 56419 721 56465 767
rect 56543 721 56589 767
rect 56667 721 56713 767
rect 56791 721 56837 767
rect 56915 721 56961 767
rect 57039 721 57085 767
rect 57163 721 57209 767
rect 57287 721 57333 767
rect 57411 721 57457 767
rect 57535 721 57581 767
rect 57659 721 57705 767
rect 57783 721 57829 767
rect 57907 721 57953 767
rect 58031 721 58077 767
rect 58155 721 58201 767
rect 58279 721 58325 767
rect 58403 721 58449 767
rect 58527 721 58573 767
rect 58651 721 58697 767
rect 58775 721 58821 767
rect 58899 721 58945 767
rect 59023 721 59069 767
rect 59147 721 59193 767
rect 59271 721 59317 767
rect 59395 721 59441 767
rect 59519 721 59565 767
rect 59643 721 59689 767
rect 59767 721 59813 767
rect 59891 721 59937 767
rect 60015 721 60061 767
rect 60139 721 60185 767
rect 60263 721 60309 767
rect 60387 721 60433 767
rect 60511 721 60557 767
rect 60635 721 60681 767
rect 60759 721 60805 767
rect 60883 721 60929 767
rect 61007 721 61053 767
rect 61131 721 61177 767
rect 61255 721 61301 767
rect 61379 721 61425 767
rect 61503 721 61549 767
rect 61627 721 61673 767
rect 61751 721 61797 767
rect 61875 721 61921 767
rect 61999 721 62045 767
rect 62123 721 62169 767
rect 62247 721 62293 767
rect 62371 721 62417 767
rect 62495 721 62541 767
rect 62619 721 62665 767
rect 62743 721 62789 767
rect 62867 721 62913 767
rect 62991 721 63037 767
rect 63115 721 63161 767
rect 63239 721 63285 767
rect 63363 721 63409 767
rect 63487 721 63533 767
rect 63611 721 63657 767
rect 63735 721 63781 767
rect 63859 721 63905 767
rect 63983 721 64029 767
rect 64107 721 64153 767
rect 64231 721 64277 767
rect 64355 721 64401 767
rect 64479 721 64525 767
rect 64603 721 64649 767
rect 64727 721 64773 767
rect 64851 721 64897 767
rect 64975 721 65021 767
rect 65099 721 65145 767
rect 65223 721 65269 767
rect 65347 721 65393 767
rect 65471 721 65517 767
rect 65595 721 65641 767
rect 65719 721 65765 767
rect 65843 721 65889 767
rect 65967 721 66013 767
rect 66091 721 66137 767
rect 66215 721 66261 767
rect 66339 721 66385 767
rect 66463 721 66509 767
rect 66587 721 66633 767
rect 66711 721 66757 767
rect 66835 721 66881 767
rect 66959 721 67005 767
rect 67083 721 67129 767
rect 67207 721 67253 767
rect 67331 721 67377 767
rect 67455 721 67501 767
rect 67579 721 67625 767
rect 67703 721 67749 767
rect 67827 721 67873 767
rect 67951 721 67997 767
rect 68075 721 68121 767
rect 68199 721 68245 767
rect 68323 721 68369 767
rect 68447 721 68493 767
rect 68571 721 68617 767
rect 68695 721 68741 767
rect 68819 721 68865 767
rect 68943 721 68989 767
rect 69067 721 69113 767
rect 69191 721 69237 767
rect 69315 721 69361 767
rect 69439 721 69485 767
rect 69563 721 69609 767
rect 69687 721 69733 767
rect 69811 721 69857 767
rect 69935 721 69981 767
rect 70059 721 70105 767
rect 70183 721 70229 767
rect 70307 721 70353 767
rect 70431 721 70477 767
rect 70555 721 70601 767
rect 70679 721 70725 767
rect 70803 721 70849 767
rect 70927 721 70973 767
rect 71051 721 71097 767
rect 71175 721 71221 767
rect 71299 721 71345 767
rect 71423 721 71469 767
rect 71547 721 71593 767
rect 71671 721 71717 767
rect 71795 721 71841 767
rect 71919 721 71965 767
rect 72043 721 72089 767
rect 72167 721 72213 767
rect 72291 721 72337 767
rect 72415 721 72461 767
rect 72539 721 72585 767
rect 72663 721 72709 767
rect 72787 721 72833 767
rect 72911 721 72957 767
rect 73035 721 73081 767
rect 73159 721 73205 767
rect 73283 721 73329 767
rect 73407 721 73453 767
rect 73531 721 73577 767
rect 73655 721 73701 767
rect 73779 721 73825 767
rect 73903 721 73949 767
rect 74027 721 74073 767
rect 74151 721 74197 767
rect 74275 721 74321 767
rect 74399 721 74445 767
rect 74523 721 74569 767
rect 74647 721 74693 767
rect 74771 721 74817 767
rect 74895 721 74941 767
rect 75019 721 75065 767
rect 75143 721 75189 767
rect 75267 721 75313 767
rect 75391 721 75437 767
rect 75515 721 75561 767
rect 75639 721 75685 767
rect 75763 721 75809 767
rect 75887 721 75933 767
rect 76011 721 76057 767
rect 76135 721 76181 767
rect 76259 721 76305 767
rect 76383 721 76429 767
rect 76507 721 76553 767
rect 76631 721 76677 767
rect 76755 721 76801 767
rect 76879 721 76925 767
rect 77003 721 77049 767
rect 77127 721 77173 767
rect 77251 721 77297 767
rect 77375 721 77421 767
rect 77499 721 77545 767
rect 77623 721 77669 767
rect 77747 721 77793 767
rect 77871 721 77917 767
rect 77995 721 78041 767
rect 78119 721 78165 767
rect 78243 721 78289 767
rect 78367 721 78413 767
rect 78491 721 78537 767
rect 78615 721 78661 767
rect 78739 721 78785 767
rect 78863 721 78909 767
rect 78987 721 79033 767
rect 79111 721 79157 767
rect 79235 721 79281 767
rect 79359 721 79405 767
rect 79483 721 79529 767
rect 79607 721 79653 767
rect 79731 721 79777 767
rect 79855 721 79901 767
rect 79979 721 80025 767
rect 80103 721 80149 767
rect 80227 721 80273 767
rect 80351 721 80397 767
rect 80475 721 80521 767
rect 80599 721 80645 767
rect 80723 721 80769 767
rect 80847 721 80893 767
rect 80971 721 81017 767
rect 81095 721 81141 767
rect 81219 721 81265 767
rect 81343 721 81389 767
rect 81467 721 81513 767
rect 81591 721 81637 767
rect 81715 721 81761 767
rect 81839 721 81885 767
rect 81963 721 82009 767
rect 82087 721 82133 767
rect 82211 721 82257 767
rect 82335 721 82381 767
rect 82459 721 82505 767
rect 82583 721 82629 767
rect 82707 721 82753 767
rect 82831 721 82877 767
rect 82955 721 83001 767
rect 83079 721 83125 767
rect 83203 721 83249 767
rect 83327 721 83373 767
rect 83451 721 83497 767
rect 83575 721 83621 767
rect 83699 721 83745 767
rect 83823 721 83869 767
rect 83947 721 83993 767
rect 84071 721 84117 767
rect 84195 721 84241 767
rect 84319 721 84365 767
rect 84443 721 84489 767
rect 84567 721 84613 767
rect 84691 721 84737 767
rect 84815 721 84861 767
rect 84939 721 84985 767
rect 85063 721 85109 767
rect 85187 721 85233 767
rect 85311 721 85357 767
rect 85435 721 85481 767
rect 85559 721 85605 767
rect 85683 721 85729 767
rect 85807 721 85853 767
rect 85931 721 85977 767
rect 371 597 417 643
rect 495 597 541 643
rect 619 597 665 643
rect 743 597 789 643
rect 867 597 913 643
rect 991 597 1037 643
rect 1115 597 1161 643
rect 1239 597 1285 643
rect 1363 597 1409 643
rect 1487 597 1533 643
rect 1611 597 1657 643
rect 1735 597 1781 643
rect 1859 597 1905 643
rect 1983 597 2029 643
rect 2107 597 2153 643
rect 2231 597 2277 643
rect 2355 597 2401 643
rect 2479 597 2525 643
rect 2603 597 2649 643
rect 2727 597 2773 643
rect 2851 597 2897 643
rect 2975 597 3021 643
rect 3099 597 3145 643
rect 3223 597 3269 643
rect 3347 597 3393 643
rect 3471 597 3517 643
rect 3595 597 3641 643
rect 3719 597 3765 643
rect 3843 597 3889 643
rect 3967 597 4013 643
rect 4091 597 4137 643
rect 4215 597 4261 643
rect 4339 597 4385 643
rect 4463 597 4509 643
rect 4587 597 4633 643
rect 4711 597 4757 643
rect 4835 597 4881 643
rect 4959 597 5005 643
rect 5083 597 5129 643
rect 5207 597 5253 643
rect 5331 597 5377 643
rect 5455 597 5501 643
rect 5579 597 5625 643
rect 5703 597 5749 643
rect 5827 597 5873 643
rect 5951 597 5997 643
rect 6075 597 6121 643
rect 6199 597 6245 643
rect 6323 597 6369 643
rect 6447 597 6493 643
rect 6571 597 6617 643
rect 6695 597 6741 643
rect 6819 597 6865 643
rect 6943 597 6989 643
rect 7067 597 7113 643
rect 7191 597 7237 643
rect 7315 597 7361 643
rect 7439 597 7485 643
rect 7563 597 7609 643
rect 7687 597 7733 643
rect 7811 597 7857 643
rect 7935 597 7981 643
rect 8059 597 8105 643
rect 8183 597 8229 643
rect 8307 597 8353 643
rect 8431 597 8477 643
rect 8555 597 8601 643
rect 8679 597 8725 643
rect 8803 597 8849 643
rect 8927 597 8973 643
rect 9051 597 9097 643
rect 9175 597 9221 643
rect 9299 597 9345 643
rect 9423 597 9469 643
rect 9547 597 9593 643
rect 9671 597 9717 643
rect 9795 597 9841 643
rect 9919 597 9965 643
rect 10043 597 10089 643
rect 10167 597 10213 643
rect 10291 597 10337 643
rect 10415 597 10461 643
rect 10539 597 10585 643
rect 10663 597 10709 643
rect 10787 597 10833 643
rect 10911 597 10957 643
rect 11035 597 11081 643
rect 11159 597 11205 643
rect 11283 597 11329 643
rect 11407 597 11453 643
rect 11531 597 11577 643
rect 11655 597 11701 643
rect 11779 597 11825 643
rect 11903 597 11949 643
rect 12027 597 12073 643
rect 12151 597 12197 643
rect 12275 597 12321 643
rect 12399 597 12445 643
rect 12523 597 12569 643
rect 12647 597 12693 643
rect 12771 597 12817 643
rect 12895 597 12941 643
rect 13019 597 13065 643
rect 13143 597 13189 643
rect 13267 597 13313 643
rect 13391 597 13437 643
rect 13515 597 13561 643
rect 13639 597 13685 643
rect 13763 597 13809 643
rect 13887 597 13933 643
rect 14011 597 14057 643
rect 14135 597 14181 643
rect 14259 597 14305 643
rect 14383 597 14429 643
rect 14507 597 14553 643
rect 14631 597 14677 643
rect 14755 597 14801 643
rect 14879 597 14925 643
rect 15003 597 15049 643
rect 15127 597 15173 643
rect 15251 597 15297 643
rect 15375 597 15421 643
rect 15499 597 15545 643
rect 15623 597 15669 643
rect 15747 597 15793 643
rect 15871 597 15917 643
rect 15995 597 16041 643
rect 16119 597 16165 643
rect 16243 597 16289 643
rect 16367 597 16413 643
rect 16491 597 16537 643
rect 16615 597 16661 643
rect 16739 597 16785 643
rect 16863 597 16909 643
rect 16987 597 17033 643
rect 17111 597 17157 643
rect 17235 597 17281 643
rect 17359 597 17405 643
rect 17483 597 17529 643
rect 17607 597 17653 643
rect 17731 597 17777 643
rect 17855 597 17901 643
rect 17979 597 18025 643
rect 18103 597 18149 643
rect 18227 597 18273 643
rect 18351 597 18397 643
rect 18475 597 18521 643
rect 18599 597 18645 643
rect 18723 597 18769 643
rect 18847 597 18893 643
rect 18971 597 19017 643
rect 19095 597 19141 643
rect 19219 597 19265 643
rect 19343 597 19389 643
rect 19467 597 19513 643
rect 19591 597 19637 643
rect 19715 597 19761 643
rect 19839 597 19885 643
rect 19963 597 20009 643
rect 20087 597 20133 643
rect 20211 597 20257 643
rect 20335 597 20381 643
rect 20459 597 20505 643
rect 20583 597 20629 643
rect 20707 597 20753 643
rect 20831 597 20877 643
rect 20955 597 21001 643
rect 21079 597 21125 643
rect 21203 597 21249 643
rect 21327 597 21373 643
rect 21451 597 21497 643
rect 21575 597 21621 643
rect 21699 597 21745 643
rect 21823 597 21869 643
rect 21947 597 21993 643
rect 22071 597 22117 643
rect 22195 597 22241 643
rect 22319 597 22365 643
rect 22443 597 22489 643
rect 22567 597 22613 643
rect 22691 597 22737 643
rect 22815 597 22861 643
rect 22939 597 22985 643
rect 23063 597 23109 643
rect 23187 597 23233 643
rect 23311 597 23357 643
rect 23435 597 23481 643
rect 23559 597 23605 643
rect 23683 597 23729 643
rect 23807 597 23853 643
rect 23931 597 23977 643
rect 24055 597 24101 643
rect 24179 597 24225 643
rect 24303 597 24349 643
rect 24427 597 24473 643
rect 24551 597 24597 643
rect 24675 597 24721 643
rect 24799 597 24845 643
rect 24923 597 24969 643
rect 25047 597 25093 643
rect 25171 597 25217 643
rect 25295 597 25341 643
rect 25419 597 25465 643
rect 25543 597 25589 643
rect 25667 597 25713 643
rect 25791 597 25837 643
rect 25915 597 25961 643
rect 26039 597 26085 643
rect 26163 597 26209 643
rect 26287 597 26333 643
rect 26411 597 26457 643
rect 26535 597 26581 643
rect 26659 597 26705 643
rect 26783 597 26829 643
rect 26907 597 26953 643
rect 27031 597 27077 643
rect 27155 597 27201 643
rect 27279 597 27325 643
rect 27403 597 27449 643
rect 27527 597 27573 643
rect 27651 597 27697 643
rect 27775 597 27821 643
rect 27899 597 27945 643
rect 28023 597 28069 643
rect 28147 597 28193 643
rect 28271 597 28317 643
rect 28395 597 28441 643
rect 28519 597 28565 643
rect 28643 597 28689 643
rect 28767 597 28813 643
rect 28891 597 28937 643
rect 29015 597 29061 643
rect 29139 597 29185 643
rect 29263 597 29309 643
rect 29387 597 29433 643
rect 29511 597 29557 643
rect 29635 597 29681 643
rect 29759 597 29805 643
rect 29883 597 29929 643
rect 30007 597 30053 643
rect 30131 597 30177 643
rect 30255 597 30301 643
rect 30379 597 30425 643
rect 30503 597 30549 643
rect 30627 597 30673 643
rect 30751 597 30797 643
rect 30875 597 30921 643
rect 30999 597 31045 643
rect 31123 597 31169 643
rect 31247 597 31293 643
rect 31371 597 31417 643
rect 31495 597 31541 643
rect 31619 597 31665 643
rect 31743 597 31789 643
rect 31867 597 31913 643
rect 31991 597 32037 643
rect 32115 597 32161 643
rect 32239 597 32285 643
rect 32363 597 32409 643
rect 32487 597 32533 643
rect 32611 597 32657 643
rect 32735 597 32781 643
rect 32859 597 32905 643
rect 32983 597 33029 643
rect 33107 597 33153 643
rect 33231 597 33277 643
rect 33355 597 33401 643
rect 33479 597 33525 643
rect 33603 597 33649 643
rect 33727 597 33773 643
rect 33851 597 33897 643
rect 33975 597 34021 643
rect 34099 597 34145 643
rect 34223 597 34269 643
rect 34347 597 34393 643
rect 34471 597 34517 643
rect 34595 597 34641 643
rect 34719 597 34765 643
rect 34843 597 34889 643
rect 34967 597 35013 643
rect 35091 597 35137 643
rect 35215 597 35261 643
rect 35339 597 35385 643
rect 35463 597 35509 643
rect 35587 597 35633 643
rect 35711 597 35757 643
rect 35835 597 35881 643
rect 35959 597 36005 643
rect 36083 597 36129 643
rect 36207 597 36253 643
rect 36331 597 36377 643
rect 36455 597 36501 643
rect 36579 597 36625 643
rect 36703 597 36749 643
rect 36827 597 36873 643
rect 36951 597 36997 643
rect 37075 597 37121 643
rect 37199 597 37245 643
rect 37323 597 37369 643
rect 37447 597 37493 643
rect 37571 597 37617 643
rect 37695 597 37741 643
rect 37819 597 37865 643
rect 37943 597 37989 643
rect 38067 597 38113 643
rect 38191 597 38237 643
rect 38315 597 38361 643
rect 38439 597 38485 643
rect 38563 597 38609 643
rect 38687 597 38733 643
rect 38811 597 38857 643
rect 38935 597 38981 643
rect 39059 597 39105 643
rect 39183 597 39229 643
rect 39307 597 39353 643
rect 39431 597 39477 643
rect 39555 597 39601 643
rect 39679 597 39725 643
rect 39803 597 39849 643
rect 39927 597 39973 643
rect 40051 597 40097 643
rect 40175 597 40221 643
rect 40299 597 40345 643
rect 40423 597 40469 643
rect 40547 597 40593 643
rect 40671 597 40717 643
rect 40795 597 40841 643
rect 40919 597 40965 643
rect 41043 597 41089 643
rect 41167 597 41213 643
rect 41291 597 41337 643
rect 41415 597 41461 643
rect 41539 597 41585 643
rect 41663 597 41709 643
rect 41787 597 41833 643
rect 41911 597 41957 643
rect 42035 597 42081 643
rect 42159 597 42205 643
rect 42283 597 42329 643
rect 42407 597 42453 643
rect 42531 597 42577 643
rect 42655 597 42701 643
rect 42779 597 42825 643
rect 42903 597 42949 643
rect 43027 597 43073 643
rect 43151 597 43197 643
rect 43275 597 43321 643
rect 43399 597 43445 643
rect 43523 597 43569 643
rect 43647 597 43693 643
rect 43771 597 43817 643
rect 43895 597 43941 643
rect 44019 597 44065 643
rect 44143 597 44189 643
rect 44267 597 44313 643
rect 44391 597 44437 643
rect 44515 597 44561 643
rect 44639 597 44685 643
rect 44763 597 44809 643
rect 44887 597 44933 643
rect 45011 597 45057 643
rect 45135 597 45181 643
rect 45259 597 45305 643
rect 45383 597 45429 643
rect 45507 597 45553 643
rect 45631 597 45677 643
rect 45755 597 45801 643
rect 45879 597 45925 643
rect 46003 597 46049 643
rect 46127 597 46173 643
rect 46251 597 46297 643
rect 46375 597 46421 643
rect 46499 597 46545 643
rect 46623 597 46669 643
rect 46747 597 46793 643
rect 46871 597 46917 643
rect 46995 597 47041 643
rect 47119 597 47165 643
rect 47243 597 47289 643
rect 47367 597 47413 643
rect 47491 597 47537 643
rect 47615 597 47661 643
rect 47739 597 47785 643
rect 47863 597 47909 643
rect 47987 597 48033 643
rect 48111 597 48157 643
rect 48235 597 48281 643
rect 48359 597 48405 643
rect 48483 597 48529 643
rect 48607 597 48653 643
rect 48731 597 48777 643
rect 48855 597 48901 643
rect 48979 597 49025 643
rect 49103 597 49149 643
rect 49227 597 49273 643
rect 49351 597 49397 643
rect 49475 597 49521 643
rect 49599 597 49645 643
rect 49723 597 49769 643
rect 49847 597 49893 643
rect 49971 597 50017 643
rect 50095 597 50141 643
rect 50219 597 50265 643
rect 50343 597 50389 643
rect 50467 597 50513 643
rect 50591 597 50637 643
rect 50715 597 50761 643
rect 50839 597 50885 643
rect 50963 597 51009 643
rect 51087 597 51133 643
rect 51211 597 51257 643
rect 51335 597 51381 643
rect 51459 597 51505 643
rect 51583 597 51629 643
rect 51707 597 51753 643
rect 51831 597 51877 643
rect 51955 597 52001 643
rect 52079 597 52125 643
rect 52203 597 52249 643
rect 52327 597 52373 643
rect 52451 597 52497 643
rect 52575 597 52621 643
rect 52699 597 52745 643
rect 52823 597 52869 643
rect 52947 597 52993 643
rect 53071 597 53117 643
rect 53195 597 53241 643
rect 53319 597 53365 643
rect 53443 597 53489 643
rect 53567 597 53613 643
rect 53691 597 53737 643
rect 53815 597 53861 643
rect 53939 597 53985 643
rect 54063 597 54109 643
rect 54187 597 54233 643
rect 54311 597 54357 643
rect 54435 597 54481 643
rect 54559 597 54605 643
rect 54683 597 54729 643
rect 54807 597 54853 643
rect 54931 597 54977 643
rect 55055 597 55101 643
rect 55179 597 55225 643
rect 55303 597 55349 643
rect 55427 597 55473 643
rect 55551 597 55597 643
rect 55675 597 55721 643
rect 55799 597 55845 643
rect 55923 597 55969 643
rect 56047 597 56093 643
rect 56171 597 56217 643
rect 56295 597 56341 643
rect 56419 597 56465 643
rect 56543 597 56589 643
rect 56667 597 56713 643
rect 56791 597 56837 643
rect 56915 597 56961 643
rect 57039 597 57085 643
rect 57163 597 57209 643
rect 57287 597 57333 643
rect 57411 597 57457 643
rect 57535 597 57581 643
rect 57659 597 57705 643
rect 57783 597 57829 643
rect 57907 597 57953 643
rect 58031 597 58077 643
rect 58155 597 58201 643
rect 58279 597 58325 643
rect 58403 597 58449 643
rect 58527 597 58573 643
rect 58651 597 58697 643
rect 58775 597 58821 643
rect 58899 597 58945 643
rect 59023 597 59069 643
rect 59147 597 59193 643
rect 59271 597 59317 643
rect 59395 597 59441 643
rect 59519 597 59565 643
rect 59643 597 59689 643
rect 59767 597 59813 643
rect 59891 597 59937 643
rect 60015 597 60061 643
rect 60139 597 60185 643
rect 60263 597 60309 643
rect 60387 597 60433 643
rect 60511 597 60557 643
rect 60635 597 60681 643
rect 60759 597 60805 643
rect 60883 597 60929 643
rect 61007 597 61053 643
rect 61131 597 61177 643
rect 61255 597 61301 643
rect 61379 597 61425 643
rect 61503 597 61549 643
rect 61627 597 61673 643
rect 61751 597 61797 643
rect 61875 597 61921 643
rect 61999 597 62045 643
rect 62123 597 62169 643
rect 62247 597 62293 643
rect 62371 597 62417 643
rect 62495 597 62541 643
rect 62619 597 62665 643
rect 62743 597 62789 643
rect 62867 597 62913 643
rect 62991 597 63037 643
rect 63115 597 63161 643
rect 63239 597 63285 643
rect 63363 597 63409 643
rect 63487 597 63533 643
rect 63611 597 63657 643
rect 63735 597 63781 643
rect 63859 597 63905 643
rect 63983 597 64029 643
rect 64107 597 64153 643
rect 64231 597 64277 643
rect 64355 597 64401 643
rect 64479 597 64525 643
rect 64603 597 64649 643
rect 64727 597 64773 643
rect 64851 597 64897 643
rect 64975 597 65021 643
rect 65099 597 65145 643
rect 65223 597 65269 643
rect 65347 597 65393 643
rect 65471 597 65517 643
rect 65595 597 65641 643
rect 65719 597 65765 643
rect 65843 597 65889 643
rect 65967 597 66013 643
rect 66091 597 66137 643
rect 66215 597 66261 643
rect 66339 597 66385 643
rect 66463 597 66509 643
rect 66587 597 66633 643
rect 66711 597 66757 643
rect 66835 597 66881 643
rect 66959 597 67005 643
rect 67083 597 67129 643
rect 67207 597 67253 643
rect 67331 597 67377 643
rect 67455 597 67501 643
rect 67579 597 67625 643
rect 67703 597 67749 643
rect 67827 597 67873 643
rect 67951 597 67997 643
rect 68075 597 68121 643
rect 68199 597 68245 643
rect 68323 597 68369 643
rect 68447 597 68493 643
rect 68571 597 68617 643
rect 68695 597 68741 643
rect 68819 597 68865 643
rect 68943 597 68989 643
rect 69067 597 69113 643
rect 69191 597 69237 643
rect 69315 597 69361 643
rect 69439 597 69485 643
rect 69563 597 69609 643
rect 69687 597 69733 643
rect 69811 597 69857 643
rect 69935 597 69981 643
rect 70059 597 70105 643
rect 70183 597 70229 643
rect 70307 597 70353 643
rect 70431 597 70477 643
rect 70555 597 70601 643
rect 70679 597 70725 643
rect 70803 597 70849 643
rect 70927 597 70973 643
rect 71051 597 71097 643
rect 71175 597 71221 643
rect 71299 597 71345 643
rect 71423 597 71469 643
rect 71547 597 71593 643
rect 71671 597 71717 643
rect 71795 597 71841 643
rect 71919 597 71965 643
rect 72043 597 72089 643
rect 72167 597 72213 643
rect 72291 597 72337 643
rect 72415 597 72461 643
rect 72539 597 72585 643
rect 72663 597 72709 643
rect 72787 597 72833 643
rect 72911 597 72957 643
rect 73035 597 73081 643
rect 73159 597 73205 643
rect 73283 597 73329 643
rect 73407 597 73453 643
rect 73531 597 73577 643
rect 73655 597 73701 643
rect 73779 597 73825 643
rect 73903 597 73949 643
rect 74027 597 74073 643
rect 74151 597 74197 643
rect 74275 597 74321 643
rect 74399 597 74445 643
rect 74523 597 74569 643
rect 74647 597 74693 643
rect 74771 597 74817 643
rect 74895 597 74941 643
rect 75019 597 75065 643
rect 75143 597 75189 643
rect 75267 597 75313 643
rect 75391 597 75437 643
rect 75515 597 75561 643
rect 75639 597 75685 643
rect 75763 597 75809 643
rect 75887 597 75933 643
rect 76011 597 76057 643
rect 76135 597 76181 643
rect 76259 597 76305 643
rect 76383 597 76429 643
rect 76507 597 76553 643
rect 76631 597 76677 643
rect 76755 597 76801 643
rect 76879 597 76925 643
rect 77003 597 77049 643
rect 77127 597 77173 643
rect 77251 597 77297 643
rect 77375 597 77421 643
rect 77499 597 77545 643
rect 77623 597 77669 643
rect 77747 597 77793 643
rect 77871 597 77917 643
rect 77995 597 78041 643
rect 78119 597 78165 643
rect 78243 597 78289 643
rect 78367 597 78413 643
rect 78491 597 78537 643
rect 78615 597 78661 643
rect 78739 597 78785 643
rect 78863 597 78909 643
rect 78987 597 79033 643
rect 79111 597 79157 643
rect 79235 597 79281 643
rect 79359 597 79405 643
rect 79483 597 79529 643
rect 79607 597 79653 643
rect 79731 597 79777 643
rect 79855 597 79901 643
rect 79979 597 80025 643
rect 80103 597 80149 643
rect 80227 597 80273 643
rect 80351 597 80397 643
rect 80475 597 80521 643
rect 80599 597 80645 643
rect 80723 597 80769 643
rect 80847 597 80893 643
rect 80971 597 81017 643
rect 81095 597 81141 643
rect 81219 597 81265 643
rect 81343 597 81389 643
rect 81467 597 81513 643
rect 81591 597 81637 643
rect 81715 597 81761 643
rect 81839 597 81885 643
rect 81963 597 82009 643
rect 82087 597 82133 643
rect 82211 597 82257 643
rect 82335 597 82381 643
rect 82459 597 82505 643
rect 82583 597 82629 643
rect 82707 597 82753 643
rect 82831 597 82877 643
rect 82955 597 83001 643
rect 83079 597 83125 643
rect 83203 597 83249 643
rect 83327 597 83373 643
rect 83451 597 83497 643
rect 83575 597 83621 643
rect 83699 597 83745 643
rect 83823 597 83869 643
rect 83947 597 83993 643
rect 84071 597 84117 643
rect 84195 597 84241 643
rect 84319 597 84365 643
rect 84443 597 84489 643
rect 84567 597 84613 643
rect 84691 597 84737 643
rect 84815 597 84861 643
rect 84939 597 84985 643
rect 85063 597 85109 643
rect 85187 597 85233 643
rect 85311 597 85357 643
rect 85435 597 85481 643
rect 85559 597 85605 643
rect 85683 597 85729 643
rect 85807 597 85853 643
rect 85931 597 85977 643
<< metal1 >>
rect 282 96683 86090 96694
rect 282 96637 371 96683
rect 417 96637 495 96683
rect 541 96637 619 96683
rect 665 96637 743 96683
rect 789 96637 867 96683
rect 913 96637 991 96683
rect 1037 96637 1115 96683
rect 1161 96637 1239 96683
rect 1285 96637 1363 96683
rect 1409 96637 1487 96683
rect 1533 96637 1611 96683
rect 1657 96637 1735 96683
rect 1781 96637 1859 96683
rect 1905 96637 1983 96683
rect 2029 96637 2107 96683
rect 2153 96637 2231 96683
rect 2277 96637 2355 96683
rect 2401 96637 2479 96683
rect 2525 96637 2603 96683
rect 2649 96637 2727 96683
rect 2773 96637 2851 96683
rect 2897 96637 2975 96683
rect 3021 96637 3099 96683
rect 3145 96637 3223 96683
rect 3269 96637 3347 96683
rect 3393 96637 3471 96683
rect 3517 96637 3595 96683
rect 3641 96637 3719 96683
rect 3765 96637 3843 96683
rect 3889 96637 3967 96683
rect 4013 96637 4091 96683
rect 4137 96637 4215 96683
rect 4261 96637 4339 96683
rect 4385 96637 4463 96683
rect 4509 96637 4587 96683
rect 4633 96637 4711 96683
rect 4757 96637 4835 96683
rect 4881 96637 4959 96683
rect 5005 96637 5083 96683
rect 5129 96637 5207 96683
rect 5253 96637 5331 96683
rect 5377 96637 5455 96683
rect 5501 96637 5579 96683
rect 5625 96637 5703 96683
rect 5749 96637 5827 96683
rect 5873 96637 5951 96683
rect 5997 96637 6075 96683
rect 6121 96637 6199 96683
rect 6245 96637 6323 96683
rect 6369 96637 6447 96683
rect 6493 96637 6571 96683
rect 6617 96637 6695 96683
rect 6741 96637 6819 96683
rect 6865 96637 6943 96683
rect 6989 96637 7067 96683
rect 7113 96637 7191 96683
rect 7237 96637 7315 96683
rect 7361 96637 7439 96683
rect 7485 96637 7563 96683
rect 7609 96637 7687 96683
rect 7733 96637 7811 96683
rect 7857 96637 7935 96683
rect 7981 96637 8059 96683
rect 8105 96637 8183 96683
rect 8229 96637 8307 96683
rect 8353 96637 8431 96683
rect 8477 96637 8555 96683
rect 8601 96637 8679 96683
rect 8725 96637 8803 96683
rect 8849 96637 8927 96683
rect 8973 96637 9051 96683
rect 9097 96637 9175 96683
rect 9221 96637 9299 96683
rect 9345 96637 9423 96683
rect 9469 96637 9547 96683
rect 9593 96637 9671 96683
rect 9717 96637 9795 96683
rect 9841 96637 9919 96683
rect 9965 96637 10043 96683
rect 10089 96637 10167 96683
rect 10213 96637 10291 96683
rect 10337 96637 10415 96683
rect 10461 96637 10539 96683
rect 10585 96637 10663 96683
rect 10709 96637 10787 96683
rect 10833 96637 10911 96683
rect 10957 96637 11035 96683
rect 11081 96637 11159 96683
rect 11205 96637 11283 96683
rect 11329 96637 11407 96683
rect 11453 96637 11531 96683
rect 11577 96637 11655 96683
rect 11701 96637 11779 96683
rect 11825 96637 11903 96683
rect 11949 96637 12027 96683
rect 12073 96637 12151 96683
rect 12197 96637 12275 96683
rect 12321 96637 12399 96683
rect 12445 96637 12523 96683
rect 12569 96637 12647 96683
rect 12693 96637 12771 96683
rect 12817 96637 12895 96683
rect 12941 96637 13019 96683
rect 13065 96637 13143 96683
rect 13189 96637 13267 96683
rect 13313 96637 13391 96683
rect 13437 96637 13515 96683
rect 13561 96637 13639 96683
rect 13685 96637 13763 96683
rect 13809 96637 13887 96683
rect 13933 96637 14011 96683
rect 14057 96637 14135 96683
rect 14181 96637 14259 96683
rect 14305 96637 14383 96683
rect 14429 96637 14507 96683
rect 14553 96637 14631 96683
rect 14677 96637 14755 96683
rect 14801 96637 14879 96683
rect 14925 96637 15003 96683
rect 15049 96637 15127 96683
rect 15173 96637 15251 96683
rect 15297 96637 15375 96683
rect 15421 96637 15499 96683
rect 15545 96637 15623 96683
rect 15669 96637 15747 96683
rect 15793 96637 15871 96683
rect 15917 96637 15995 96683
rect 16041 96637 16119 96683
rect 16165 96637 16243 96683
rect 16289 96637 16367 96683
rect 16413 96637 16491 96683
rect 16537 96637 16615 96683
rect 16661 96637 16739 96683
rect 16785 96637 16863 96683
rect 16909 96637 16987 96683
rect 17033 96637 17111 96683
rect 17157 96637 17235 96683
rect 17281 96637 17359 96683
rect 17405 96637 17483 96683
rect 17529 96637 17607 96683
rect 17653 96637 17731 96683
rect 17777 96637 17855 96683
rect 17901 96637 17979 96683
rect 18025 96637 18103 96683
rect 18149 96637 18227 96683
rect 18273 96637 18351 96683
rect 18397 96637 18475 96683
rect 18521 96637 18599 96683
rect 18645 96637 18723 96683
rect 18769 96637 18847 96683
rect 18893 96637 18971 96683
rect 19017 96637 19095 96683
rect 19141 96637 19219 96683
rect 19265 96637 19343 96683
rect 19389 96637 19467 96683
rect 19513 96637 19591 96683
rect 19637 96637 19715 96683
rect 19761 96637 19839 96683
rect 19885 96637 19963 96683
rect 20009 96637 20087 96683
rect 20133 96637 20211 96683
rect 20257 96637 20335 96683
rect 20381 96637 20459 96683
rect 20505 96637 20583 96683
rect 20629 96637 20707 96683
rect 20753 96637 20831 96683
rect 20877 96637 20955 96683
rect 21001 96637 21079 96683
rect 21125 96637 21203 96683
rect 21249 96637 21327 96683
rect 21373 96637 21451 96683
rect 21497 96637 21575 96683
rect 21621 96637 21699 96683
rect 21745 96637 21823 96683
rect 21869 96637 21947 96683
rect 21993 96637 22071 96683
rect 22117 96637 22195 96683
rect 22241 96637 22319 96683
rect 22365 96637 22443 96683
rect 22489 96637 22567 96683
rect 22613 96637 22691 96683
rect 22737 96637 22815 96683
rect 22861 96637 22939 96683
rect 22985 96637 23063 96683
rect 23109 96637 23187 96683
rect 23233 96637 23311 96683
rect 23357 96637 23435 96683
rect 23481 96637 23559 96683
rect 23605 96637 23683 96683
rect 23729 96637 23807 96683
rect 23853 96637 23931 96683
rect 23977 96637 24055 96683
rect 24101 96637 24179 96683
rect 24225 96637 24303 96683
rect 24349 96637 24427 96683
rect 24473 96637 24551 96683
rect 24597 96637 24675 96683
rect 24721 96637 24799 96683
rect 24845 96637 24923 96683
rect 24969 96637 25047 96683
rect 25093 96637 25171 96683
rect 25217 96637 25295 96683
rect 25341 96637 25419 96683
rect 25465 96637 25543 96683
rect 25589 96637 25667 96683
rect 25713 96637 25791 96683
rect 25837 96637 25915 96683
rect 25961 96637 26039 96683
rect 26085 96637 26163 96683
rect 26209 96637 26287 96683
rect 26333 96637 26411 96683
rect 26457 96637 26535 96683
rect 26581 96637 26659 96683
rect 26705 96637 26783 96683
rect 26829 96637 26907 96683
rect 26953 96637 27031 96683
rect 27077 96637 27155 96683
rect 27201 96637 27279 96683
rect 27325 96637 27403 96683
rect 27449 96637 27527 96683
rect 27573 96637 27651 96683
rect 27697 96637 27775 96683
rect 27821 96637 27899 96683
rect 27945 96637 28023 96683
rect 28069 96637 28147 96683
rect 28193 96637 28271 96683
rect 28317 96637 28395 96683
rect 28441 96637 28519 96683
rect 28565 96637 28643 96683
rect 28689 96637 28767 96683
rect 28813 96637 28891 96683
rect 28937 96637 29015 96683
rect 29061 96637 29139 96683
rect 29185 96637 29263 96683
rect 29309 96637 29387 96683
rect 29433 96637 29511 96683
rect 29557 96637 29635 96683
rect 29681 96637 29759 96683
rect 29805 96637 29883 96683
rect 29929 96637 30007 96683
rect 30053 96637 30131 96683
rect 30177 96637 30255 96683
rect 30301 96637 30379 96683
rect 30425 96637 30503 96683
rect 30549 96637 30627 96683
rect 30673 96637 30751 96683
rect 30797 96637 30875 96683
rect 30921 96637 30999 96683
rect 31045 96637 31123 96683
rect 31169 96637 31247 96683
rect 31293 96637 31371 96683
rect 31417 96637 31495 96683
rect 31541 96637 31619 96683
rect 31665 96637 31743 96683
rect 31789 96637 31867 96683
rect 31913 96637 31991 96683
rect 32037 96637 32115 96683
rect 32161 96637 32239 96683
rect 32285 96637 32363 96683
rect 32409 96637 32487 96683
rect 32533 96637 32611 96683
rect 32657 96637 32735 96683
rect 32781 96637 32859 96683
rect 32905 96637 32983 96683
rect 33029 96637 33107 96683
rect 33153 96637 33231 96683
rect 33277 96637 33355 96683
rect 33401 96637 33479 96683
rect 33525 96637 33603 96683
rect 33649 96637 33727 96683
rect 33773 96637 33851 96683
rect 33897 96637 33975 96683
rect 34021 96637 34099 96683
rect 34145 96637 34223 96683
rect 34269 96637 34347 96683
rect 34393 96637 34471 96683
rect 34517 96637 34595 96683
rect 34641 96637 34719 96683
rect 34765 96637 34843 96683
rect 34889 96637 34967 96683
rect 35013 96637 35091 96683
rect 35137 96637 35215 96683
rect 35261 96637 35339 96683
rect 35385 96637 35463 96683
rect 35509 96637 35587 96683
rect 35633 96637 35711 96683
rect 35757 96637 35835 96683
rect 35881 96637 35959 96683
rect 36005 96637 36083 96683
rect 36129 96637 36207 96683
rect 36253 96637 36331 96683
rect 36377 96637 36455 96683
rect 36501 96637 36579 96683
rect 36625 96637 36703 96683
rect 36749 96637 36827 96683
rect 36873 96637 36951 96683
rect 36997 96637 37075 96683
rect 37121 96637 37199 96683
rect 37245 96637 37323 96683
rect 37369 96637 37447 96683
rect 37493 96637 37571 96683
rect 37617 96637 37695 96683
rect 37741 96637 37819 96683
rect 37865 96637 37943 96683
rect 37989 96637 38067 96683
rect 38113 96637 38191 96683
rect 38237 96637 38315 96683
rect 38361 96637 38439 96683
rect 38485 96637 38563 96683
rect 38609 96637 38687 96683
rect 38733 96637 38811 96683
rect 38857 96637 38935 96683
rect 38981 96637 39059 96683
rect 39105 96637 39183 96683
rect 39229 96637 39307 96683
rect 39353 96637 39431 96683
rect 39477 96637 39555 96683
rect 39601 96637 39679 96683
rect 39725 96637 39803 96683
rect 39849 96637 39927 96683
rect 39973 96637 40051 96683
rect 40097 96637 40175 96683
rect 40221 96637 40299 96683
rect 40345 96637 40423 96683
rect 40469 96637 40547 96683
rect 40593 96637 40671 96683
rect 40717 96637 40795 96683
rect 40841 96637 40919 96683
rect 40965 96637 41043 96683
rect 41089 96637 41167 96683
rect 41213 96637 41291 96683
rect 41337 96637 41415 96683
rect 41461 96637 41539 96683
rect 41585 96637 41663 96683
rect 41709 96637 41787 96683
rect 41833 96637 41911 96683
rect 41957 96637 42035 96683
rect 42081 96637 42159 96683
rect 42205 96637 42283 96683
rect 42329 96637 42407 96683
rect 42453 96637 42531 96683
rect 42577 96637 42655 96683
rect 42701 96637 42779 96683
rect 42825 96637 42903 96683
rect 42949 96637 43027 96683
rect 43073 96637 43151 96683
rect 43197 96637 43275 96683
rect 43321 96637 43399 96683
rect 43445 96637 43523 96683
rect 43569 96637 43647 96683
rect 43693 96637 43771 96683
rect 43817 96637 43895 96683
rect 43941 96637 44019 96683
rect 44065 96637 44143 96683
rect 44189 96637 44267 96683
rect 44313 96637 44391 96683
rect 44437 96637 44515 96683
rect 44561 96637 44639 96683
rect 44685 96637 44763 96683
rect 44809 96637 44887 96683
rect 44933 96637 45011 96683
rect 45057 96637 45135 96683
rect 45181 96637 45259 96683
rect 45305 96637 45383 96683
rect 45429 96637 45507 96683
rect 45553 96637 45631 96683
rect 45677 96637 45755 96683
rect 45801 96637 45879 96683
rect 45925 96637 46003 96683
rect 46049 96637 46127 96683
rect 46173 96637 46251 96683
rect 46297 96637 46375 96683
rect 46421 96637 46499 96683
rect 46545 96637 46623 96683
rect 46669 96637 46747 96683
rect 46793 96637 46871 96683
rect 46917 96637 46995 96683
rect 47041 96637 47119 96683
rect 47165 96637 47243 96683
rect 47289 96637 47367 96683
rect 47413 96637 47491 96683
rect 47537 96637 47615 96683
rect 47661 96637 47739 96683
rect 47785 96637 47863 96683
rect 47909 96637 47987 96683
rect 48033 96637 48111 96683
rect 48157 96637 48235 96683
rect 48281 96637 48359 96683
rect 48405 96637 48483 96683
rect 48529 96637 48607 96683
rect 48653 96637 48731 96683
rect 48777 96637 48855 96683
rect 48901 96637 48979 96683
rect 49025 96637 49103 96683
rect 49149 96637 49227 96683
rect 49273 96637 49351 96683
rect 49397 96637 49475 96683
rect 49521 96637 49599 96683
rect 49645 96637 49723 96683
rect 49769 96637 49847 96683
rect 49893 96637 49971 96683
rect 50017 96637 50095 96683
rect 50141 96637 50219 96683
rect 50265 96637 50343 96683
rect 50389 96637 50467 96683
rect 50513 96637 50591 96683
rect 50637 96637 50715 96683
rect 50761 96637 50839 96683
rect 50885 96637 50963 96683
rect 51009 96637 51087 96683
rect 51133 96637 51211 96683
rect 51257 96637 51335 96683
rect 51381 96637 51459 96683
rect 51505 96637 51583 96683
rect 51629 96637 51707 96683
rect 51753 96637 51831 96683
rect 51877 96637 51955 96683
rect 52001 96637 52079 96683
rect 52125 96637 52203 96683
rect 52249 96637 52327 96683
rect 52373 96637 52451 96683
rect 52497 96637 52575 96683
rect 52621 96637 52699 96683
rect 52745 96637 52823 96683
rect 52869 96637 52947 96683
rect 52993 96637 53071 96683
rect 53117 96637 53195 96683
rect 53241 96637 53319 96683
rect 53365 96637 53443 96683
rect 53489 96637 53567 96683
rect 53613 96637 53691 96683
rect 53737 96637 53815 96683
rect 53861 96637 53939 96683
rect 53985 96637 54063 96683
rect 54109 96637 54187 96683
rect 54233 96637 54311 96683
rect 54357 96637 54435 96683
rect 54481 96637 54559 96683
rect 54605 96637 54683 96683
rect 54729 96637 54807 96683
rect 54853 96637 54931 96683
rect 54977 96637 55055 96683
rect 55101 96637 55179 96683
rect 55225 96637 55303 96683
rect 55349 96637 55427 96683
rect 55473 96637 55551 96683
rect 55597 96637 55675 96683
rect 55721 96637 55799 96683
rect 55845 96637 55923 96683
rect 55969 96637 56047 96683
rect 56093 96637 56171 96683
rect 56217 96637 56295 96683
rect 56341 96637 56419 96683
rect 56465 96637 56543 96683
rect 56589 96637 56667 96683
rect 56713 96637 56791 96683
rect 56837 96637 56915 96683
rect 56961 96637 57039 96683
rect 57085 96637 57163 96683
rect 57209 96637 57287 96683
rect 57333 96637 57411 96683
rect 57457 96637 57535 96683
rect 57581 96637 57659 96683
rect 57705 96637 57783 96683
rect 57829 96637 57907 96683
rect 57953 96637 58031 96683
rect 58077 96637 58155 96683
rect 58201 96637 58279 96683
rect 58325 96637 58403 96683
rect 58449 96637 58527 96683
rect 58573 96637 58651 96683
rect 58697 96637 58775 96683
rect 58821 96637 58899 96683
rect 58945 96637 59023 96683
rect 59069 96637 59147 96683
rect 59193 96637 59271 96683
rect 59317 96637 59395 96683
rect 59441 96637 59519 96683
rect 59565 96637 59643 96683
rect 59689 96637 59767 96683
rect 59813 96637 59891 96683
rect 59937 96637 60015 96683
rect 60061 96637 60139 96683
rect 60185 96637 60263 96683
rect 60309 96637 60387 96683
rect 60433 96637 60511 96683
rect 60557 96637 60635 96683
rect 60681 96637 60759 96683
rect 60805 96637 60883 96683
rect 60929 96637 61007 96683
rect 61053 96637 61131 96683
rect 61177 96637 61255 96683
rect 61301 96637 61379 96683
rect 61425 96637 61503 96683
rect 61549 96637 61627 96683
rect 61673 96637 61751 96683
rect 61797 96637 61875 96683
rect 61921 96637 61999 96683
rect 62045 96637 62123 96683
rect 62169 96637 62247 96683
rect 62293 96637 62371 96683
rect 62417 96637 62495 96683
rect 62541 96637 62619 96683
rect 62665 96637 62743 96683
rect 62789 96637 62867 96683
rect 62913 96637 62991 96683
rect 63037 96637 63115 96683
rect 63161 96637 63239 96683
rect 63285 96637 63363 96683
rect 63409 96637 63487 96683
rect 63533 96637 63611 96683
rect 63657 96637 63735 96683
rect 63781 96637 63859 96683
rect 63905 96637 63983 96683
rect 64029 96637 64107 96683
rect 64153 96637 64231 96683
rect 64277 96637 64355 96683
rect 64401 96637 64479 96683
rect 64525 96637 64603 96683
rect 64649 96637 64727 96683
rect 64773 96637 64851 96683
rect 64897 96637 64975 96683
rect 65021 96637 65099 96683
rect 65145 96637 65223 96683
rect 65269 96637 65347 96683
rect 65393 96637 65471 96683
rect 65517 96637 65595 96683
rect 65641 96637 65719 96683
rect 65765 96637 65843 96683
rect 65889 96637 65967 96683
rect 66013 96637 66091 96683
rect 66137 96637 66215 96683
rect 66261 96637 66339 96683
rect 66385 96637 66463 96683
rect 66509 96637 66587 96683
rect 66633 96637 66711 96683
rect 66757 96637 66835 96683
rect 66881 96637 66959 96683
rect 67005 96637 67083 96683
rect 67129 96637 67207 96683
rect 67253 96637 67331 96683
rect 67377 96637 67455 96683
rect 67501 96637 67579 96683
rect 67625 96637 67703 96683
rect 67749 96637 67827 96683
rect 67873 96637 67951 96683
rect 67997 96637 68075 96683
rect 68121 96637 68199 96683
rect 68245 96637 68323 96683
rect 68369 96637 68447 96683
rect 68493 96637 68571 96683
rect 68617 96637 68695 96683
rect 68741 96637 68819 96683
rect 68865 96637 68943 96683
rect 68989 96637 69067 96683
rect 69113 96637 69191 96683
rect 69237 96637 69315 96683
rect 69361 96637 69439 96683
rect 69485 96637 69563 96683
rect 69609 96637 69687 96683
rect 69733 96637 69811 96683
rect 69857 96637 69935 96683
rect 69981 96637 70059 96683
rect 70105 96637 70183 96683
rect 70229 96637 70307 96683
rect 70353 96637 70431 96683
rect 70477 96637 70555 96683
rect 70601 96637 70679 96683
rect 70725 96637 70803 96683
rect 70849 96637 70927 96683
rect 70973 96637 71051 96683
rect 71097 96637 71175 96683
rect 71221 96637 71299 96683
rect 71345 96637 71423 96683
rect 71469 96637 71547 96683
rect 71593 96637 71671 96683
rect 71717 96637 71795 96683
rect 71841 96637 71919 96683
rect 71965 96637 72043 96683
rect 72089 96637 72167 96683
rect 72213 96637 72291 96683
rect 72337 96637 72415 96683
rect 72461 96637 72539 96683
rect 72585 96637 72663 96683
rect 72709 96637 72787 96683
rect 72833 96637 72911 96683
rect 72957 96637 73035 96683
rect 73081 96637 73159 96683
rect 73205 96637 73283 96683
rect 73329 96637 73407 96683
rect 73453 96637 73531 96683
rect 73577 96637 73655 96683
rect 73701 96637 73779 96683
rect 73825 96637 73903 96683
rect 73949 96637 74027 96683
rect 74073 96637 74151 96683
rect 74197 96637 74275 96683
rect 74321 96637 74399 96683
rect 74445 96637 74523 96683
rect 74569 96637 74647 96683
rect 74693 96637 74771 96683
rect 74817 96637 74895 96683
rect 74941 96637 75019 96683
rect 75065 96637 75143 96683
rect 75189 96637 75267 96683
rect 75313 96637 75391 96683
rect 75437 96637 75515 96683
rect 75561 96637 75639 96683
rect 75685 96637 75763 96683
rect 75809 96637 75887 96683
rect 75933 96637 76011 96683
rect 76057 96637 76135 96683
rect 76181 96637 76259 96683
rect 76305 96637 76383 96683
rect 76429 96637 76507 96683
rect 76553 96637 76631 96683
rect 76677 96637 76755 96683
rect 76801 96637 76879 96683
rect 76925 96637 77003 96683
rect 77049 96637 77127 96683
rect 77173 96637 77251 96683
rect 77297 96637 77375 96683
rect 77421 96637 77499 96683
rect 77545 96637 77623 96683
rect 77669 96637 77747 96683
rect 77793 96637 77871 96683
rect 77917 96637 77995 96683
rect 78041 96637 78119 96683
rect 78165 96637 78243 96683
rect 78289 96637 78367 96683
rect 78413 96637 78491 96683
rect 78537 96637 78615 96683
rect 78661 96637 78739 96683
rect 78785 96637 78863 96683
rect 78909 96637 78987 96683
rect 79033 96637 79111 96683
rect 79157 96637 79235 96683
rect 79281 96637 79359 96683
rect 79405 96637 79483 96683
rect 79529 96637 79607 96683
rect 79653 96637 79731 96683
rect 79777 96637 79855 96683
rect 79901 96637 79979 96683
rect 80025 96637 80103 96683
rect 80149 96637 80227 96683
rect 80273 96637 80351 96683
rect 80397 96637 80475 96683
rect 80521 96637 80599 96683
rect 80645 96637 80723 96683
rect 80769 96637 80847 96683
rect 80893 96637 80971 96683
rect 81017 96637 81095 96683
rect 81141 96637 81219 96683
rect 81265 96637 81343 96683
rect 81389 96637 81467 96683
rect 81513 96637 81591 96683
rect 81637 96637 81715 96683
rect 81761 96637 81839 96683
rect 81885 96637 81963 96683
rect 82009 96637 82087 96683
rect 82133 96637 82211 96683
rect 82257 96637 82335 96683
rect 82381 96637 82459 96683
rect 82505 96637 82583 96683
rect 82629 96637 82707 96683
rect 82753 96637 82831 96683
rect 82877 96637 82955 96683
rect 83001 96637 83079 96683
rect 83125 96637 83203 96683
rect 83249 96637 83327 96683
rect 83373 96637 83451 96683
rect 83497 96637 83575 96683
rect 83621 96637 83699 96683
rect 83745 96637 83823 96683
rect 83869 96637 83947 96683
rect 83993 96637 84071 96683
rect 84117 96637 84195 96683
rect 84241 96637 84319 96683
rect 84365 96637 84443 96683
rect 84489 96637 84567 96683
rect 84613 96637 84691 96683
rect 84737 96637 84815 96683
rect 84861 96637 84939 96683
rect 84985 96637 85063 96683
rect 85109 96637 85187 96683
rect 85233 96637 85311 96683
rect 85357 96637 85435 96683
rect 85481 96637 85559 96683
rect 85605 96637 85683 96683
rect 85729 96637 85807 96683
rect 85853 96637 85931 96683
rect 85977 96637 86090 96683
rect 282 96559 86090 96637
rect 282 96513 371 96559
rect 417 96513 495 96559
rect 541 96513 619 96559
rect 665 96513 743 96559
rect 789 96513 867 96559
rect 913 96513 991 96559
rect 1037 96513 1115 96559
rect 1161 96513 1239 96559
rect 1285 96513 1363 96559
rect 1409 96513 1487 96559
rect 1533 96513 1611 96559
rect 1657 96513 1735 96559
rect 1781 96513 1859 96559
rect 1905 96513 1983 96559
rect 2029 96513 2107 96559
rect 2153 96513 2231 96559
rect 2277 96513 2355 96559
rect 2401 96513 2479 96559
rect 2525 96513 2603 96559
rect 2649 96513 2727 96559
rect 2773 96513 2851 96559
rect 2897 96513 2975 96559
rect 3021 96513 3099 96559
rect 3145 96513 3223 96559
rect 3269 96513 3347 96559
rect 3393 96513 3471 96559
rect 3517 96513 3595 96559
rect 3641 96513 3719 96559
rect 3765 96513 3843 96559
rect 3889 96513 3967 96559
rect 4013 96513 4091 96559
rect 4137 96513 4215 96559
rect 4261 96513 4339 96559
rect 4385 96513 4463 96559
rect 4509 96513 4587 96559
rect 4633 96513 4711 96559
rect 4757 96513 4835 96559
rect 4881 96513 4959 96559
rect 5005 96513 5083 96559
rect 5129 96513 5207 96559
rect 5253 96513 5331 96559
rect 5377 96513 5455 96559
rect 5501 96513 5579 96559
rect 5625 96513 5703 96559
rect 5749 96513 5827 96559
rect 5873 96513 5951 96559
rect 5997 96513 6075 96559
rect 6121 96513 6199 96559
rect 6245 96513 6323 96559
rect 6369 96513 6447 96559
rect 6493 96513 6571 96559
rect 6617 96513 6695 96559
rect 6741 96513 6819 96559
rect 6865 96513 6943 96559
rect 6989 96513 7067 96559
rect 7113 96513 7191 96559
rect 7237 96513 7315 96559
rect 7361 96513 7439 96559
rect 7485 96513 7563 96559
rect 7609 96513 7687 96559
rect 7733 96513 7811 96559
rect 7857 96513 7935 96559
rect 7981 96513 8059 96559
rect 8105 96513 8183 96559
rect 8229 96513 8307 96559
rect 8353 96513 8431 96559
rect 8477 96513 8555 96559
rect 8601 96513 8679 96559
rect 8725 96513 8803 96559
rect 8849 96513 8927 96559
rect 8973 96513 9051 96559
rect 9097 96513 9175 96559
rect 9221 96513 9299 96559
rect 9345 96513 9423 96559
rect 9469 96513 9547 96559
rect 9593 96513 9671 96559
rect 9717 96513 9795 96559
rect 9841 96513 9919 96559
rect 9965 96513 10043 96559
rect 10089 96513 10167 96559
rect 10213 96513 10291 96559
rect 10337 96513 10415 96559
rect 10461 96513 10539 96559
rect 10585 96513 10663 96559
rect 10709 96513 10787 96559
rect 10833 96513 10911 96559
rect 10957 96513 11035 96559
rect 11081 96513 11159 96559
rect 11205 96513 11283 96559
rect 11329 96513 11407 96559
rect 11453 96513 11531 96559
rect 11577 96513 11655 96559
rect 11701 96513 11779 96559
rect 11825 96513 11903 96559
rect 11949 96513 12027 96559
rect 12073 96513 12151 96559
rect 12197 96513 12275 96559
rect 12321 96513 12399 96559
rect 12445 96513 12523 96559
rect 12569 96513 12647 96559
rect 12693 96513 12771 96559
rect 12817 96513 12895 96559
rect 12941 96513 13019 96559
rect 13065 96513 13143 96559
rect 13189 96513 13267 96559
rect 13313 96513 13391 96559
rect 13437 96513 13515 96559
rect 13561 96513 13639 96559
rect 13685 96513 13763 96559
rect 13809 96513 13887 96559
rect 13933 96513 14011 96559
rect 14057 96513 14135 96559
rect 14181 96513 14259 96559
rect 14305 96513 14383 96559
rect 14429 96513 14507 96559
rect 14553 96513 14631 96559
rect 14677 96513 14755 96559
rect 14801 96513 14879 96559
rect 14925 96513 15003 96559
rect 15049 96513 15127 96559
rect 15173 96513 15251 96559
rect 15297 96513 15375 96559
rect 15421 96513 15499 96559
rect 15545 96513 15623 96559
rect 15669 96513 15747 96559
rect 15793 96513 15871 96559
rect 15917 96513 15995 96559
rect 16041 96513 16119 96559
rect 16165 96513 16243 96559
rect 16289 96513 16367 96559
rect 16413 96513 16491 96559
rect 16537 96513 16615 96559
rect 16661 96513 16739 96559
rect 16785 96513 16863 96559
rect 16909 96513 16987 96559
rect 17033 96513 17111 96559
rect 17157 96513 17235 96559
rect 17281 96513 17359 96559
rect 17405 96513 17483 96559
rect 17529 96513 17607 96559
rect 17653 96513 17731 96559
rect 17777 96513 17855 96559
rect 17901 96513 17979 96559
rect 18025 96513 18103 96559
rect 18149 96513 18227 96559
rect 18273 96513 18351 96559
rect 18397 96513 18475 96559
rect 18521 96513 18599 96559
rect 18645 96513 18723 96559
rect 18769 96513 18847 96559
rect 18893 96513 18971 96559
rect 19017 96513 19095 96559
rect 19141 96513 19219 96559
rect 19265 96513 19343 96559
rect 19389 96513 19467 96559
rect 19513 96513 19591 96559
rect 19637 96513 19715 96559
rect 19761 96513 19839 96559
rect 19885 96513 19963 96559
rect 20009 96513 20087 96559
rect 20133 96513 20211 96559
rect 20257 96513 20335 96559
rect 20381 96513 20459 96559
rect 20505 96513 20583 96559
rect 20629 96513 20707 96559
rect 20753 96513 20831 96559
rect 20877 96513 20955 96559
rect 21001 96513 21079 96559
rect 21125 96513 21203 96559
rect 21249 96513 21327 96559
rect 21373 96513 21451 96559
rect 21497 96513 21575 96559
rect 21621 96513 21699 96559
rect 21745 96513 21823 96559
rect 21869 96513 21947 96559
rect 21993 96513 22071 96559
rect 22117 96513 22195 96559
rect 22241 96513 22319 96559
rect 22365 96513 22443 96559
rect 22489 96513 22567 96559
rect 22613 96513 22691 96559
rect 22737 96513 22815 96559
rect 22861 96513 22939 96559
rect 22985 96513 23063 96559
rect 23109 96513 23187 96559
rect 23233 96513 23311 96559
rect 23357 96513 23435 96559
rect 23481 96513 23559 96559
rect 23605 96513 23683 96559
rect 23729 96513 23807 96559
rect 23853 96513 23931 96559
rect 23977 96513 24055 96559
rect 24101 96513 24179 96559
rect 24225 96513 24303 96559
rect 24349 96513 24427 96559
rect 24473 96513 24551 96559
rect 24597 96513 24675 96559
rect 24721 96513 24799 96559
rect 24845 96513 24923 96559
rect 24969 96513 25047 96559
rect 25093 96513 25171 96559
rect 25217 96513 25295 96559
rect 25341 96513 25419 96559
rect 25465 96513 25543 96559
rect 25589 96513 25667 96559
rect 25713 96513 25791 96559
rect 25837 96513 25915 96559
rect 25961 96513 26039 96559
rect 26085 96513 26163 96559
rect 26209 96513 26287 96559
rect 26333 96513 26411 96559
rect 26457 96513 26535 96559
rect 26581 96513 26659 96559
rect 26705 96513 26783 96559
rect 26829 96513 26907 96559
rect 26953 96513 27031 96559
rect 27077 96513 27155 96559
rect 27201 96513 27279 96559
rect 27325 96513 27403 96559
rect 27449 96513 27527 96559
rect 27573 96513 27651 96559
rect 27697 96513 27775 96559
rect 27821 96513 27899 96559
rect 27945 96513 28023 96559
rect 28069 96513 28147 96559
rect 28193 96513 28271 96559
rect 28317 96513 28395 96559
rect 28441 96513 28519 96559
rect 28565 96513 28643 96559
rect 28689 96513 28767 96559
rect 28813 96513 28891 96559
rect 28937 96513 29015 96559
rect 29061 96513 29139 96559
rect 29185 96513 29263 96559
rect 29309 96513 29387 96559
rect 29433 96513 29511 96559
rect 29557 96513 29635 96559
rect 29681 96513 29759 96559
rect 29805 96513 29883 96559
rect 29929 96513 30007 96559
rect 30053 96513 30131 96559
rect 30177 96513 30255 96559
rect 30301 96513 30379 96559
rect 30425 96513 30503 96559
rect 30549 96513 30627 96559
rect 30673 96513 30751 96559
rect 30797 96513 30875 96559
rect 30921 96513 30999 96559
rect 31045 96513 31123 96559
rect 31169 96513 31247 96559
rect 31293 96513 31371 96559
rect 31417 96513 31495 96559
rect 31541 96513 31619 96559
rect 31665 96513 31743 96559
rect 31789 96513 31867 96559
rect 31913 96513 31991 96559
rect 32037 96513 32115 96559
rect 32161 96513 32239 96559
rect 32285 96513 32363 96559
rect 32409 96513 32487 96559
rect 32533 96513 32611 96559
rect 32657 96513 32735 96559
rect 32781 96513 32859 96559
rect 32905 96513 32983 96559
rect 33029 96513 33107 96559
rect 33153 96513 33231 96559
rect 33277 96513 33355 96559
rect 33401 96513 33479 96559
rect 33525 96513 33603 96559
rect 33649 96513 33727 96559
rect 33773 96513 33851 96559
rect 33897 96513 33975 96559
rect 34021 96513 34099 96559
rect 34145 96513 34223 96559
rect 34269 96513 34347 96559
rect 34393 96513 34471 96559
rect 34517 96513 34595 96559
rect 34641 96513 34719 96559
rect 34765 96513 34843 96559
rect 34889 96513 34967 96559
rect 35013 96513 35091 96559
rect 35137 96513 35215 96559
rect 35261 96513 35339 96559
rect 35385 96513 35463 96559
rect 35509 96513 35587 96559
rect 35633 96513 35711 96559
rect 35757 96513 35835 96559
rect 35881 96513 35959 96559
rect 36005 96513 36083 96559
rect 36129 96513 36207 96559
rect 36253 96513 36331 96559
rect 36377 96513 36455 96559
rect 36501 96513 36579 96559
rect 36625 96513 36703 96559
rect 36749 96513 36827 96559
rect 36873 96513 36951 96559
rect 36997 96513 37075 96559
rect 37121 96513 37199 96559
rect 37245 96513 37323 96559
rect 37369 96513 37447 96559
rect 37493 96513 37571 96559
rect 37617 96513 37695 96559
rect 37741 96513 37819 96559
rect 37865 96513 37943 96559
rect 37989 96513 38067 96559
rect 38113 96513 38191 96559
rect 38237 96513 38315 96559
rect 38361 96513 38439 96559
rect 38485 96513 38563 96559
rect 38609 96513 38687 96559
rect 38733 96513 38811 96559
rect 38857 96513 38935 96559
rect 38981 96513 39059 96559
rect 39105 96513 39183 96559
rect 39229 96513 39307 96559
rect 39353 96513 39431 96559
rect 39477 96513 39555 96559
rect 39601 96513 39679 96559
rect 39725 96513 39803 96559
rect 39849 96513 39927 96559
rect 39973 96513 40051 96559
rect 40097 96513 40175 96559
rect 40221 96513 40299 96559
rect 40345 96513 40423 96559
rect 40469 96513 40547 96559
rect 40593 96513 40671 96559
rect 40717 96513 40795 96559
rect 40841 96513 40919 96559
rect 40965 96513 41043 96559
rect 41089 96513 41167 96559
rect 41213 96513 41291 96559
rect 41337 96513 41415 96559
rect 41461 96513 41539 96559
rect 41585 96513 41663 96559
rect 41709 96513 41787 96559
rect 41833 96513 41911 96559
rect 41957 96513 42035 96559
rect 42081 96513 42159 96559
rect 42205 96513 42283 96559
rect 42329 96513 42407 96559
rect 42453 96513 42531 96559
rect 42577 96513 42655 96559
rect 42701 96513 42779 96559
rect 42825 96513 42903 96559
rect 42949 96513 43027 96559
rect 43073 96513 43151 96559
rect 43197 96513 43275 96559
rect 43321 96513 43399 96559
rect 43445 96513 43523 96559
rect 43569 96513 43647 96559
rect 43693 96513 43771 96559
rect 43817 96513 43895 96559
rect 43941 96513 44019 96559
rect 44065 96513 44143 96559
rect 44189 96513 44267 96559
rect 44313 96513 44391 96559
rect 44437 96513 44515 96559
rect 44561 96513 44639 96559
rect 44685 96513 44763 96559
rect 44809 96513 44887 96559
rect 44933 96513 45011 96559
rect 45057 96513 45135 96559
rect 45181 96513 45259 96559
rect 45305 96513 45383 96559
rect 45429 96513 45507 96559
rect 45553 96513 45631 96559
rect 45677 96513 45755 96559
rect 45801 96513 45879 96559
rect 45925 96513 46003 96559
rect 46049 96513 46127 96559
rect 46173 96513 46251 96559
rect 46297 96513 46375 96559
rect 46421 96513 46499 96559
rect 46545 96513 46623 96559
rect 46669 96513 46747 96559
rect 46793 96513 46871 96559
rect 46917 96513 46995 96559
rect 47041 96513 47119 96559
rect 47165 96513 47243 96559
rect 47289 96513 47367 96559
rect 47413 96513 47491 96559
rect 47537 96513 47615 96559
rect 47661 96513 47739 96559
rect 47785 96513 47863 96559
rect 47909 96513 47987 96559
rect 48033 96513 48111 96559
rect 48157 96513 48235 96559
rect 48281 96513 48359 96559
rect 48405 96513 48483 96559
rect 48529 96513 48607 96559
rect 48653 96513 48731 96559
rect 48777 96513 48855 96559
rect 48901 96513 48979 96559
rect 49025 96513 49103 96559
rect 49149 96513 49227 96559
rect 49273 96513 49351 96559
rect 49397 96513 49475 96559
rect 49521 96513 49599 96559
rect 49645 96513 49723 96559
rect 49769 96513 49847 96559
rect 49893 96513 49971 96559
rect 50017 96513 50095 96559
rect 50141 96513 50219 96559
rect 50265 96513 50343 96559
rect 50389 96513 50467 96559
rect 50513 96513 50591 96559
rect 50637 96513 50715 96559
rect 50761 96513 50839 96559
rect 50885 96513 50963 96559
rect 51009 96513 51087 96559
rect 51133 96513 51211 96559
rect 51257 96513 51335 96559
rect 51381 96513 51459 96559
rect 51505 96513 51583 96559
rect 51629 96513 51707 96559
rect 51753 96513 51831 96559
rect 51877 96513 51955 96559
rect 52001 96513 52079 96559
rect 52125 96513 52203 96559
rect 52249 96513 52327 96559
rect 52373 96513 52451 96559
rect 52497 96513 52575 96559
rect 52621 96513 52699 96559
rect 52745 96513 52823 96559
rect 52869 96513 52947 96559
rect 52993 96513 53071 96559
rect 53117 96513 53195 96559
rect 53241 96513 53319 96559
rect 53365 96513 53443 96559
rect 53489 96513 53567 96559
rect 53613 96513 53691 96559
rect 53737 96513 53815 96559
rect 53861 96513 53939 96559
rect 53985 96513 54063 96559
rect 54109 96513 54187 96559
rect 54233 96513 54311 96559
rect 54357 96513 54435 96559
rect 54481 96513 54559 96559
rect 54605 96513 54683 96559
rect 54729 96513 54807 96559
rect 54853 96513 54931 96559
rect 54977 96513 55055 96559
rect 55101 96513 55179 96559
rect 55225 96513 55303 96559
rect 55349 96513 55427 96559
rect 55473 96513 55551 96559
rect 55597 96513 55675 96559
rect 55721 96513 55799 96559
rect 55845 96513 55923 96559
rect 55969 96513 56047 96559
rect 56093 96513 56171 96559
rect 56217 96513 56295 96559
rect 56341 96513 56419 96559
rect 56465 96513 56543 96559
rect 56589 96513 56667 96559
rect 56713 96513 56791 96559
rect 56837 96513 56915 96559
rect 56961 96513 57039 96559
rect 57085 96513 57163 96559
rect 57209 96513 57287 96559
rect 57333 96513 57411 96559
rect 57457 96513 57535 96559
rect 57581 96513 57659 96559
rect 57705 96513 57783 96559
rect 57829 96513 57907 96559
rect 57953 96513 58031 96559
rect 58077 96513 58155 96559
rect 58201 96513 58279 96559
rect 58325 96513 58403 96559
rect 58449 96513 58527 96559
rect 58573 96513 58651 96559
rect 58697 96513 58775 96559
rect 58821 96513 58899 96559
rect 58945 96513 59023 96559
rect 59069 96513 59147 96559
rect 59193 96513 59271 96559
rect 59317 96513 59395 96559
rect 59441 96513 59519 96559
rect 59565 96513 59643 96559
rect 59689 96513 59767 96559
rect 59813 96513 59891 96559
rect 59937 96513 60015 96559
rect 60061 96513 60139 96559
rect 60185 96513 60263 96559
rect 60309 96513 60387 96559
rect 60433 96513 60511 96559
rect 60557 96513 60635 96559
rect 60681 96513 60759 96559
rect 60805 96513 60883 96559
rect 60929 96513 61007 96559
rect 61053 96513 61131 96559
rect 61177 96513 61255 96559
rect 61301 96513 61379 96559
rect 61425 96513 61503 96559
rect 61549 96513 61627 96559
rect 61673 96513 61751 96559
rect 61797 96513 61875 96559
rect 61921 96513 61999 96559
rect 62045 96513 62123 96559
rect 62169 96513 62247 96559
rect 62293 96513 62371 96559
rect 62417 96513 62495 96559
rect 62541 96513 62619 96559
rect 62665 96513 62743 96559
rect 62789 96513 62867 96559
rect 62913 96513 62991 96559
rect 63037 96513 63115 96559
rect 63161 96513 63239 96559
rect 63285 96513 63363 96559
rect 63409 96513 63487 96559
rect 63533 96513 63611 96559
rect 63657 96513 63735 96559
rect 63781 96513 63859 96559
rect 63905 96513 63983 96559
rect 64029 96513 64107 96559
rect 64153 96513 64231 96559
rect 64277 96513 64355 96559
rect 64401 96513 64479 96559
rect 64525 96513 64603 96559
rect 64649 96513 64727 96559
rect 64773 96513 64851 96559
rect 64897 96513 64975 96559
rect 65021 96513 65099 96559
rect 65145 96513 65223 96559
rect 65269 96513 65347 96559
rect 65393 96513 65471 96559
rect 65517 96513 65595 96559
rect 65641 96513 65719 96559
rect 65765 96513 65843 96559
rect 65889 96513 65967 96559
rect 66013 96513 66091 96559
rect 66137 96513 66215 96559
rect 66261 96513 66339 96559
rect 66385 96513 66463 96559
rect 66509 96513 66587 96559
rect 66633 96513 66711 96559
rect 66757 96513 66835 96559
rect 66881 96513 66959 96559
rect 67005 96513 67083 96559
rect 67129 96513 67207 96559
rect 67253 96513 67331 96559
rect 67377 96513 67455 96559
rect 67501 96513 67579 96559
rect 67625 96513 67703 96559
rect 67749 96513 67827 96559
rect 67873 96513 67951 96559
rect 67997 96513 68075 96559
rect 68121 96513 68199 96559
rect 68245 96513 68323 96559
rect 68369 96513 68447 96559
rect 68493 96513 68571 96559
rect 68617 96513 68695 96559
rect 68741 96513 68819 96559
rect 68865 96513 68943 96559
rect 68989 96513 69067 96559
rect 69113 96513 69191 96559
rect 69237 96513 69315 96559
rect 69361 96513 69439 96559
rect 69485 96513 69563 96559
rect 69609 96513 69687 96559
rect 69733 96513 69811 96559
rect 69857 96513 69935 96559
rect 69981 96513 70059 96559
rect 70105 96513 70183 96559
rect 70229 96513 70307 96559
rect 70353 96513 70431 96559
rect 70477 96513 70555 96559
rect 70601 96513 70679 96559
rect 70725 96513 70803 96559
rect 70849 96513 70927 96559
rect 70973 96513 71051 96559
rect 71097 96513 71175 96559
rect 71221 96513 71299 96559
rect 71345 96513 71423 96559
rect 71469 96513 71547 96559
rect 71593 96513 71671 96559
rect 71717 96513 71795 96559
rect 71841 96513 71919 96559
rect 71965 96513 72043 96559
rect 72089 96513 72167 96559
rect 72213 96513 72291 96559
rect 72337 96513 72415 96559
rect 72461 96513 72539 96559
rect 72585 96513 72663 96559
rect 72709 96513 72787 96559
rect 72833 96513 72911 96559
rect 72957 96513 73035 96559
rect 73081 96513 73159 96559
rect 73205 96513 73283 96559
rect 73329 96513 73407 96559
rect 73453 96513 73531 96559
rect 73577 96513 73655 96559
rect 73701 96513 73779 96559
rect 73825 96513 73903 96559
rect 73949 96513 74027 96559
rect 74073 96513 74151 96559
rect 74197 96513 74275 96559
rect 74321 96513 74399 96559
rect 74445 96513 74523 96559
rect 74569 96513 74647 96559
rect 74693 96513 74771 96559
rect 74817 96513 74895 96559
rect 74941 96513 75019 96559
rect 75065 96513 75143 96559
rect 75189 96513 75267 96559
rect 75313 96513 75391 96559
rect 75437 96513 75515 96559
rect 75561 96513 75639 96559
rect 75685 96513 75763 96559
rect 75809 96513 75887 96559
rect 75933 96513 76011 96559
rect 76057 96513 76135 96559
rect 76181 96513 76259 96559
rect 76305 96513 76383 96559
rect 76429 96513 76507 96559
rect 76553 96513 76631 96559
rect 76677 96513 76755 96559
rect 76801 96513 76879 96559
rect 76925 96513 77003 96559
rect 77049 96513 77127 96559
rect 77173 96513 77251 96559
rect 77297 96513 77375 96559
rect 77421 96513 77499 96559
rect 77545 96513 77623 96559
rect 77669 96513 77747 96559
rect 77793 96513 77871 96559
rect 77917 96513 77995 96559
rect 78041 96513 78119 96559
rect 78165 96513 78243 96559
rect 78289 96513 78367 96559
rect 78413 96513 78491 96559
rect 78537 96513 78615 96559
rect 78661 96513 78739 96559
rect 78785 96513 78863 96559
rect 78909 96513 78987 96559
rect 79033 96513 79111 96559
rect 79157 96513 79235 96559
rect 79281 96513 79359 96559
rect 79405 96513 79483 96559
rect 79529 96513 79607 96559
rect 79653 96513 79731 96559
rect 79777 96513 79855 96559
rect 79901 96513 79979 96559
rect 80025 96513 80103 96559
rect 80149 96513 80227 96559
rect 80273 96513 80351 96559
rect 80397 96513 80475 96559
rect 80521 96513 80599 96559
rect 80645 96513 80723 96559
rect 80769 96513 80847 96559
rect 80893 96513 80971 96559
rect 81017 96513 81095 96559
rect 81141 96513 81219 96559
rect 81265 96513 81343 96559
rect 81389 96513 81467 96559
rect 81513 96513 81591 96559
rect 81637 96513 81715 96559
rect 81761 96513 81839 96559
rect 81885 96513 81963 96559
rect 82009 96513 82087 96559
rect 82133 96513 82211 96559
rect 82257 96513 82335 96559
rect 82381 96513 82459 96559
rect 82505 96513 82583 96559
rect 82629 96513 82707 96559
rect 82753 96513 82831 96559
rect 82877 96513 82955 96559
rect 83001 96513 83079 96559
rect 83125 96513 83203 96559
rect 83249 96513 83327 96559
rect 83373 96513 83451 96559
rect 83497 96513 83575 96559
rect 83621 96513 83699 96559
rect 83745 96513 83823 96559
rect 83869 96513 83947 96559
rect 83993 96513 84071 96559
rect 84117 96513 84195 96559
rect 84241 96513 84319 96559
rect 84365 96513 84443 96559
rect 84489 96513 84567 96559
rect 84613 96513 84691 96559
rect 84737 96513 84815 96559
rect 84861 96513 84939 96559
rect 84985 96513 85063 96559
rect 85109 96513 85187 96559
rect 85233 96513 85311 96559
rect 85357 96513 85435 96559
rect 85481 96513 85559 96559
rect 85605 96513 85683 96559
rect 85729 96513 85807 96559
rect 85853 96513 85931 96559
rect 85977 96513 86090 96559
rect 282 96435 86090 96513
rect 282 96389 371 96435
rect 417 96389 495 96435
rect 541 96389 619 96435
rect 665 96389 743 96435
rect 789 96389 867 96435
rect 913 96389 991 96435
rect 1037 96389 1115 96435
rect 1161 96389 1239 96435
rect 1285 96389 1363 96435
rect 1409 96389 1487 96435
rect 1533 96389 1611 96435
rect 1657 96389 1735 96435
rect 1781 96389 1859 96435
rect 1905 96389 1983 96435
rect 2029 96389 2107 96435
rect 2153 96389 2231 96435
rect 2277 96389 2355 96435
rect 2401 96389 2479 96435
rect 2525 96389 2603 96435
rect 2649 96389 2727 96435
rect 2773 96389 2851 96435
rect 2897 96389 2975 96435
rect 3021 96389 3099 96435
rect 3145 96389 3223 96435
rect 3269 96389 3347 96435
rect 3393 96389 3471 96435
rect 3517 96389 3595 96435
rect 3641 96389 3719 96435
rect 3765 96389 3843 96435
rect 3889 96389 3967 96435
rect 4013 96389 4091 96435
rect 4137 96389 4215 96435
rect 4261 96389 4339 96435
rect 4385 96389 4463 96435
rect 4509 96389 4587 96435
rect 4633 96389 4711 96435
rect 4757 96389 4835 96435
rect 4881 96389 4959 96435
rect 5005 96389 5083 96435
rect 5129 96389 5207 96435
rect 5253 96389 5331 96435
rect 5377 96389 5455 96435
rect 5501 96389 5579 96435
rect 5625 96389 5703 96435
rect 5749 96389 5827 96435
rect 5873 96389 5951 96435
rect 5997 96389 6075 96435
rect 6121 96389 6199 96435
rect 6245 96389 6323 96435
rect 6369 96389 6447 96435
rect 6493 96389 6571 96435
rect 6617 96389 6695 96435
rect 6741 96389 6819 96435
rect 6865 96389 6943 96435
rect 6989 96389 7067 96435
rect 7113 96389 7191 96435
rect 7237 96389 7315 96435
rect 7361 96389 7439 96435
rect 7485 96389 7563 96435
rect 7609 96389 7687 96435
rect 7733 96389 7811 96435
rect 7857 96389 7935 96435
rect 7981 96389 8059 96435
rect 8105 96389 8183 96435
rect 8229 96389 8307 96435
rect 8353 96389 8431 96435
rect 8477 96389 8555 96435
rect 8601 96389 8679 96435
rect 8725 96389 8803 96435
rect 8849 96389 8927 96435
rect 8973 96389 9051 96435
rect 9097 96389 9175 96435
rect 9221 96389 9299 96435
rect 9345 96389 9423 96435
rect 9469 96389 9547 96435
rect 9593 96389 9671 96435
rect 9717 96389 9795 96435
rect 9841 96389 9919 96435
rect 9965 96389 10043 96435
rect 10089 96389 10167 96435
rect 10213 96389 10291 96435
rect 10337 96389 10415 96435
rect 10461 96389 10539 96435
rect 10585 96389 10663 96435
rect 10709 96389 10787 96435
rect 10833 96389 10911 96435
rect 10957 96389 11035 96435
rect 11081 96389 11159 96435
rect 11205 96389 11283 96435
rect 11329 96389 11407 96435
rect 11453 96389 11531 96435
rect 11577 96389 11655 96435
rect 11701 96389 11779 96435
rect 11825 96389 11903 96435
rect 11949 96389 12027 96435
rect 12073 96389 12151 96435
rect 12197 96389 12275 96435
rect 12321 96389 12399 96435
rect 12445 96389 12523 96435
rect 12569 96389 12647 96435
rect 12693 96389 12771 96435
rect 12817 96389 12895 96435
rect 12941 96389 13019 96435
rect 13065 96389 13143 96435
rect 13189 96389 13267 96435
rect 13313 96389 13391 96435
rect 13437 96389 13515 96435
rect 13561 96389 13639 96435
rect 13685 96389 13763 96435
rect 13809 96389 13887 96435
rect 13933 96389 14011 96435
rect 14057 96389 14135 96435
rect 14181 96389 14259 96435
rect 14305 96389 14383 96435
rect 14429 96389 14507 96435
rect 14553 96389 14631 96435
rect 14677 96389 14755 96435
rect 14801 96389 14879 96435
rect 14925 96389 15003 96435
rect 15049 96389 15127 96435
rect 15173 96389 15251 96435
rect 15297 96389 15375 96435
rect 15421 96389 15499 96435
rect 15545 96389 15623 96435
rect 15669 96389 15747 96435
rect 15793 96389 15871 96435
rect 15917 96389 15995 96435
rect 16041 96389 16119 96435
rect 16165 96389 16243 96435
rect 16289 96389 16367 96435
rect 16413 96389 16491 96435
rect 16537 96389 16615 96435
rect 16661 96389 16739 96435
rect 16785 96389 16863 96435
rect 16909 96389 16987 96435
rect 17033 96389 17111 96435
rect 17157 96389 17235 96435
rect 17281 96389 17359 96435
rect 17405 96389 17483 96435
rect 17529 96389 17607 96435
rect 17653 96389 17731 96435
rect 17777 96389 17855 96435
rect 17901 96389 17979 96435
rect 18025 96389 18103 96435
rect 18149 96389 18227 96435
rect 18273 96389 18351 96435
rect 18397 96389 18475 96435
rect 18521 96389 18599 96435
rect 18645 96389 18723 96435
rect 18769 96389 18847 96435
rect 18893 96389 18971 96435
rect 19017 96389 19095 96435
rect 19141 96389 19219 96435
rect 19265 96389 19343 96435
rect 19389 96389 19467 96435
rect 19513 96389 19591 96435
rect 19637 96389 19715 96435
rect 19761 96389 19839 96435
rect 19885 96389 19963 96435
rect 20009 96389 20087 96435
rect 20133 96389 20211 96435
rect 20257 96389 20335 96435
rect 20381 96389 20459 96435
rect 20505 96389 20583 96435
rect 20629 96389 20707 96435
rect 20753 96389 20831 96435
rect 20877 96389 20955 96435
rect 21001 96389 21079 96435
rect 21125 96389 21203 96435
rect 21249 96389 21327 96435
rect 21373 96389 21451 96435
rect 21497 96389 21575 96435
rect 21621 96389 21699 96435
rect 21745 96389 21823 96435
rect 21869 96389 21947 96435
rect 21993 96389 22071 96435
rect 22117 96389 22195 96435
rect 22241 96389 22319 96435
rect 22365 96389 22443 96435
rect 22489 96389 22567 96435
rect 22613 96389 22691 96435
rect 22737 96389 22815 96435
rect 22861 96389 22939 96435
rect 22985 96389 23063 96435
rect 23109 96389 23187 96435
rect 23233 96389 23311 96435
rect 23357 96389 23435 96435
rect 23481 96389 23559 96435
rect 23605 96389 23683 96435
rect 23729 96389 23807 96435
rect 23853 96389 23931 96435
rect 23977 96389 24055 96435
rect 24101 96389 24179 96435
rect 24225 96389 24303 96435
rect 24349 96389 24427 96435
rect 24473 96389 24551 96435
rect 24597 96389 24675 96435
rect 24721 96389 24799 96435
rect 24845 96389 24923 96435
rect 24969 96389 25047 96435
rect 25093 96389 25171 96435
rect 25217 96389 25295 96435
rect 25341 96389 25419 96435
rect 25465 96389 25543 96435
rect 25589 96389 25667 96435
rect 25713 96389 25791 96435
rect 25837 96389 25915 96435
rect 25961 96389 26039 96435
rect 26085 96389 26163 96435
rect 26209 96389 26287 96435
rect 26333 96389 26411 96435
rect 26457 96389 26535 96435
rect 26581 96389 26659 96435
rect 26705 96389 26783 96435
rect 26829 96389 26907 96435
rect 26953 96389 27031 96435
rect 27077 96389 27155 96435
rect 27201 96389 27279 96435
rect 27325 96389 27403 96435
rect 27449 96389 27527 96435
rect 27573 96389 27651 96435
rect 27697 96389 27775 96435
rect 27821 96389 27899 96435
rect 27945 96389 28023 96435
rect 28069 96389 28147 96435
rect 28193 96389 28271 96435
rect 28317 96389 28395 96435
rect 28441 96389 28519 96435
rect 28565 96389 28643 96435
rect 28689 96389 28767 96435
rect 28813 96389 28891 96435
rect 28937 96389 29015 96435
rect 29061 96389 29139 96435
rect 29185 96389 29263 96435
rect 29309 96389 29387 96435
rect 29433 96389 29511 96435
rect 29557 96389 29635 96435
rect 29681 96389 29759 96435
rect 29805 96389 29883 96435
rect 29929 96389 30007 96435
rect 30053 96389 30131 96435
rect 30177 96389 30255 96435
rect 30301 96389 30379 96435
rect 30425 96389 30503 96435
rect 30549 96389 30627 96435
rect 30673 96389 30751 96435
rect 30797 96389 30875 96435
rect 30921 96389 30999 96435
rect 31045 96389 31123 96435
rect 31169 96389 31247 96435
rect 31293 96389 31371 96435
rect 31417 96389 31495 96435
rect 31541 96389 31619 96435
rect 31665 96389 31743 96435
rect 31789 96389 31867 96435
rect 31913 96389 31991 96435
rect 32037 96389 32115 96435
rect 32161 96389 32239 96435
rect 32285 96389 32363 96435
rect 32409 96389 32487 96435
rect 32533 96389 32611 96435
rect 32657 96389 32735 96435
rect 32781 96389 32859 96435
rect 32905 96389 32983 96435
rect 33029 96389 33107 96435
rect 33153 96389 33231 96435
rect 33277 96389 33355 96435
rect 33401 96389 33479 96435
rect 33525 96389 33603 96435
rect 33649 96389 33727 96435
rect 33773 96389 33851 96435
rect 33897 96389 33975 96435
rect 34021 96389 34099 96435
rect 34145 96389 34223 96435
rect 34269 96389 34347 96435
rect 34393 96389 34471 96435
rect 34517 96389 34595 96435
rect 34641 96389 34719 96435
rect 34765 96389 34843 96435
rect 34889 96389 34967 96435
rect 35013 96389 35091 96435
rect 35137 96389 35215 96435
rect 35261 96389 35339 96435
rect 35385 96389 35463 96435
rect 35509 96389 35587 96435
rect 35633 96389 35711 96435
rect 35757 96389 35835 96435
rect 35881 96389 35959 96435
rect 36005 96389 36083 96435
rect 36129 96389 36207 96435
rect 36253 96389 36331 96435
rect 36377 96389 36455 96435
rect 36501 96389 36579 96435
rect 36625 96389 36703 96435
rect 36749 96389 36827 96435
rect 36873 96389 36951 96435
rect 36997 96389 37075 96435
rect 37121 96389 37199 96435
rect 37245 96389 37323 96435
rect 37369 96389 37447 96435
rect 37493 96389 37571 96435
rect 37617 96389 37695 96435
rect 37741 96389 37819 96435
rect 37865 96389 37943 96435
rect 37989 96389 38067 96435
rect 38113 96389 38191 96435
rect 38237 96389 38315 96435
rect 38361 96389 38439 96435
rect 38485 96389 38563 96435
rect 38609 96389 38687 96435
rect 38733 96389 38811 96435
rect 38857 96389 38935 96435
rect 38981 96389 39059 96435
rect 39105 96389 39183 96435
rect 39229 96389 39307 96435
rect 39353 96389 39431 96435
rect 39477 96389 39555 96435
rect 39601 96389 39679 96435
rect 39725 96389 39803 96435
rect 39849 96389 39927 96435
rect 39973 96389 40051 96435
rect 40097 96389 40175 96435
rect 40221 96389 40299 96435
rect 40345 96389 40423 96435
rect 40469 96389 40547 96435
rect 40593 96389 40671 96435
rect 40717 96389 40795 96435
rect 40841 96389 40919 96435
rect 40965 96389 41043 96435
rect 41089 96389 41167 96435
rect 41213 96389 41291 96435
rect 41337 96389 41415 96435
rect 41461 96389 41539 96435
rect 41585 96389 41663 96435
rect 41709 96389 41787 96435
rect 41833 96389 41911 96435
rect 41957 96389 42035 96435
rect 42081 96389 42159 96435
rect 42205 96389 42283 96435
rect 42329 96389 42407 96435
rect 42453 96389 42531 96435
rect 42577 96389 42655 96435
rect 42701 96389 42779 96435
rect 42825 96389 42903 96435
rect 42949 96389 43027 96435
rect 43073 96389 43151 96435
rect 43197 96389 43275 96435
rect 43321 96389 43399 96435
rect 43445 96389 43523 96435
rect 43569 96389 43647 96435
rect 43693 96389 43771 96435
rect 43817 96389 43895 96435
rect 43941 96389 44019 96435
rect 44065 96389 44143 96435
rect 44189 96389 44267 96435
rect 44313 96389 44391 96435
rect 44437 96389 44515 96435
rect 44561 96389 44639 96435
rect 44685 96389 44763 96435
rect 44809 96389 44887 96435
rect 44933 96389 45011 96435
rect 45057 96389 45135 96435
rect 45181 96389 45259 96435
rect 45305 96389 45383 96435
rect 45429 96389 45507 96435
rect 45553 96389 45631 96435
rect 45677 96389 45755 96435
rect 45801 96389 45879 96435
rect 45925 96389 46003 96435
rect 46049 96389 46127 96435
rect 46173 96389 46251 96435
rect 46297 96389 46375 96435
rect 46421 96389 46499 96435
rect 46545 96389 46623 96435
rect 46669 96389 46747 96435
rect 46793 96389 46871 96435
rect 46917 96389 46995 96435
rect 47041 96389 47119 96435
rect 47165 96389 47243 96435
rect 47289 96389 47367 96435
rect 47413 96389 47491 96435
rect 47537 96389 47615 96435
rect 47661 96389 47739 96435
rect 47785 96389 47863 96435
rect 47909 96389 47987 96435
rect 48033 96389 48111 96435
rect 48157 96389 48235 96435
rect 48281 96389 48359 96435
rect 48405 96389 48483 96435
rect 48529 96389 48607 96435
rect 48653 96389 48731 96435
rect 48777 96389 48855 96435
rect 48901 96389 48979 96435
rect 49025 96389 49103 96435
rect 49149 96389 49227 96435
rect 49273 96389 49351 96435
rect 49397 96389 49475 96435
rect 49521 96389 49599 96435
rect 49645 96389 49723 96435
rect 49769 96389 49847 96435
rect 49893 96389 49971 96435
rect 50017 96389 50095 96435
rect 50141 96389 50219 96435
rect 50265 96389 50343 96435
rect 50389 96389 50467 96435
rect 50513 96389 50591 96435
rect 50637 96389 50715 96435
rect 50761 96389 50839 96435
rect 50885 96389 50963 96435
rect 51009 96389 51087 96435
rect 51133 96389 51211 96435
rect 51257 96389 51335 96435
rect 51381 96389 51459 96435
rect 51505 96389 51583 96435
rect 51629 96389 51707 96435
rect 51753 96389 51831 96435
rect 51877 96389 51955 96435
rect 52001 96389 52079 96435
rect 52125 96389 52203 96435
rect 52249 96389 52327 96435
rect 52373 96389 52451 96435
rect 52497 96389 52575 96435
rect 52621 96389 52699 96435
rect 52745 96389 52823 96435
rect 52869 96389 52947 96435
rect 52993 96389 53071 96435
rect 53117 96389 53195 96435
rect 53241 96389 53319 96435
rect 53365 96389 53443 96435
rect 53489 96389 53567 96435
rect 53613 96389 53691 96435
rect 53737 96389 53815 96435
rect 53861 96389 53939 96435
rect 53985 96389 54063 96435
rect 54109 96389 54187 96435
rect 54233 96389 54311 96435
rect 54357 96389 54435 96435
rect 54481 96389 54559 96435
rect 54605 96389 54683 96435
rect 54729 96389 54807 96435
rect 54853 96389 54931 96435
rect 54977 96389 55055 96435
rect 55101 96389 55179 96435
rect 55225 96389 55303 96435
rect 55349 96389 55427 96435
rect 55473 96389 55551 96435
rect 55597 96389 55675 96435
rect 55721 96389 55799 96435
rect 55845 96389 55923 96435
rect 55969 96389 56047 96435
rect 56093 96389 56171 96435
rect 56217 96389 56295 96435
rect 56341 96389 56419 96435
rect 56465 96389 56543 96435
rect 56589 96389 56667 96435
rect 56713 96389 56791 96435
rect 56837 96389 56915 96435
rect 56961 96389 57039 96435
rect 57085 96389 57163 96435
rect 57209 96389 57287 96435
rect 57333 96389 57411 96435
rect 57457 96389 57535 96435
rect 57581 96389 57659 96435
rect 57705 96389 57783 96435
rect 57829 96389 57907 96435
rect 57953 96389 58031 96435
rect 58077 96389 58155 96435
rect 58201 96389 58279 96435
rect 58325 96389 58403 96435
rect 58449 96389 58527 96435
rect 58573 96389 58651 96435
rect 58697 96389 58775 96435
rect 58821 96389 58899 96435
rect 58945 96389 59023 96435
rect 59069 96389 59147 96435
rect 59193 96389 59271 96435
rect 59317 96389 59395 96435
rect 59441 96389 59519 96435
rect 59565 96389 59643 96435
rect 59689 96389 59767 96435
rect 59813 96389 59891 96435
rect 59937 96389 60015 96435
rect 60061 96389 60139 96435
rect 60185 96389 60263 96435
rect 60309 96389 60387 96435
rect 60433 96389 60511 96435
rect 60557 96389 60635 96435
rect 60681 96389 60759 96435
rect 60805 96389 60883 96435
rect 60929 96389 61007 96435
rect 61053 96389 61131 96435
rect 61177 96389 61255 96435
rect 61301 96389 61379 96435
rect 61425 96389 61503 96435
rect 61549 96389 61627 96435
rect 61673 96389 61751 96435
rect 61797 96389 61875 96435
rect 61921 96389 61999 96435
rect 62045 96389 62123 96435
rect 62169 96389 62247 96435
rect 62293 96389 62371 96435
rect 62417 96389 62495 96435
rect 62541 96389 62619 96435
rect 62665 96389 62743 96435
rect 62789 96389 62867 96435
rect 62913 96389 62991 96435
rect 63037 96389 63115 96435
rect 63161 96389 63239 96435
rect 63285 96389 63363 96435
rect 63409 96389 63487 96435
rect 63533 96389 63611 96435
rect 63657 96389 63735 96435
rect 63781 96389 63859 96435
rect 63905 96389 63983 96435
rect 64029 96389 64107 96435
rect 64153 96389 64231 96435
rect 64277 96389 64355 96435
rect 64401 96389 64479 96435
rect 64525 96389 64603 96435
rect 64649 96389 64727 96435
rect 64773 96389 64851 96435
rect 64897 96389 64975 96435
rect 65021 96389 65099 96435
rect 65145 96389 65223 96435
rect 65269 96389 65347 96435
rect 65393 96389 65471 96435
rect 65517 96389 65595 96435
rect 65641 96389 65719 96435
rect 65765 96389 65843 96435
rect 65889 96389 65967 96435
rect 66013 96389 66091 96435
rect 66137 96389 66215 96435
rect 66261 96389 66339 96435
rect 66385 96389 66463 96435
rect 66509 96389 66587 96435
rect 66633 96389 66711 96435
rect 66757 96389 66835 96435
rect 66881 96389 66959 96435
rect 67005 96389 67083 96435
rect 67129 96389 67207 96435
rect 67253 96389 67331 96435
rect 67377 96389 67455 96435
rect 67501 96389 67579 96435
rect 67625 96389 67703 96435
rect 67749 96389 67827 96435
rect 67873 96389 67951 96435
rect 67997 96389 68075 96435
rect 68121 96389 68199 96435
rect 68245 96389 68323 96435
rect 68369 96389 68447 96435
rect 68493 96389 68571 96435
rect 68617 96389 68695 96435
rect 68741 96389 68819 96435
rect 68865 96389 68943 96435
rect 68989 96389 69067 96435
rect 69113 96389 69191 96435
rect 69237 96389 69315 96435
rect 69361 96389 69439 96435
rect 69485 96389 69563 96435
rect 69609 96389 69687 96435
rect 69733 96389 69811 96435
rect 69857 96389 69935 96435
rect 69981 96389 70059 96435
rect 70105 96389 70183 96435
rect 70229 96389 70307 96435
rect 70353 96389 70431 96435
rect 70477 96389 70555 96435
rect 70601 96389 70679 96435
rect 70725 96389 70803 96435
rect 70849 96389 70927 96435
rect 70973 96389 71051 96435
rect 71097 96389 71175 96435
rect 71221 96389 71299 96435
rect 71345 96389 71423 96435
rect 71469 96389 71547 96435
rect 71593 96389 71671 96435
rect 71717 96389 71795 96435
rect 71841 96389 71919 96435
rect 71965 96389 72043 96435
rect 72089 96389 72167 96435
rect 72213 96389 72291 96435
rect 72337 96389 72415 96435
rect 72461 96389 72539 96435
rect 72585 96389 72663 96435
rect 72709 96389 72787 96435
rect 72833 96389 72911 96435
rect 72957 96389 73035 96435
rect 73081 96389 73159 96435
rect 73205 96389 73283 96435
rect 73329 96389 73407 96435
rect 73453 96389 73531 96435
rect 73577 96389 73655 96435
rect 73701 96389 73779 96435
rect 73825 96389 73903 96435
rect 73949 96389 74027 96435
rect 74073 96389 74151 96435
rect 74197 96389 74275 96435
rect 74321 96389 74399 96435
rect 74445 96389 74523 96435
rect 74569 96389 74647 96435
rect 74693 96389 74771 96435
rect 74817 96389 74895 96435
rect 74941 96389 75019 96435
rect 75065 96389 75143 96435
rect 75189 96389 75267 96435
rect 75313 96389 75391 96435
rect 75437 96389 75515 96435
rect 75561 96389 75639 96435
rect 75685 96389 75763 96435
rect 75809 96389 75887 96435
rect 75933 96389 76011 96435
rect 76057 96389 76135 96435
rect 76181 96389 76259 96435
rect 76305 96389 76383 96435
rect 76429 96389 76507 96435
rect 76553 96389 76631 96435
rect 76677 96389 76755 96435
rect 76801 96389 76879 96435
rect 76925 96389 77003 96435
rect 77049 96389 77127 96435
rect 77173 96389 77251 96435
rect 77297 96389 77375 96435
rect 77421 96389 77499 96435
rect 77545 96389 77623 96435
rect 77669 96389 77747 96435
rect 77793 96389 77871 96435
rect 77917 96389 77995 96435
rect 78041 96389 78119 96435
rect 78165 96389 78243 96435
rect 78289 96389 78367 96435
rect 78413 96389 78491 96435
rect 78537 96389 78615 96435
rect 78661 96389 78739 96435
rect 78785 96389 78863 96435
rect 78909 96389 78987 96435
rect 79033 96389 79111 96435
rect 79157 96389 79235 96435
rect 79281 96389 79359 96435
rect 79405 96389 79483 96435
rect 79529 96389 79607 96435
rect 79653 96389 79731 96435
rect 79777 96389 79855 96435
rect 79901 96389 79979 96435
rect 80025 96389 80103 96435
rect 80149 96389 80227 96435
rect 80273 96389 80351 96435
rect 80397 96389 80475 96435
rect 80521 96389 80599 96435
rect 80645 96389 80723 96435
rect 80769 96389 80847 96435
rect 80893 96389 80971 96435
rect 81017 96389 81095 96435
rect 81141 96389 81219 96435
rect 81265 96389 81343 96435
rect 81389 96389 81467 96435
rect 81513 96389 81591 96435
rect 81637 96389 81715 96435
rect 81761 96389 81839 96435
rect 81885 96389 81963 96435
rect 82009 96389 82087 96435
rect 82133 96389 82211 96435
rect 82257 96389 82335 96435
rect 82381 96389 82459 96435
rect 82505 96389 82583 96435
rect 82629 96389 82707 96435
rect 82753 96389 82831 96435
rect 82877 96389 82955 96435
rect 83001 96389 83079 96435
rect 83125 96389 83203 96435
rect 83249 96389 83327 96435
rect 83373 96389 83451 96435
rect 83497 96389 83575 96435
rect 83621 96389 83699 96435
rect 83745 96389 83823 96435
rect 83869 96389 83947 96435
rect 83993 96389 84071 96435
rect 84117 96389 84195 96435
rect 84241 96389 84319 96435
rect 84365 96389 84443 96435
rect 84489 96389 84567 96435
rect 84613 96389 84691 96435
rect 84737 96389 84815 96435
rect 84861 96389 84939 96435
rect 84985 96389 85063 96435
rect 85109 96389 85187 96435
rect 85233 96389 85311 96435
rect 85357 96389 85435 96435
rect 85481 96389 85559 96435
rect 85605 96389 85683 96435
rect 85729 96389 85807 96435
rect 85853 96389 85931 96435
rect 85977 96389 86090 96435
rect 282 96311 86090 96389
rect 282 96265 371 96311
rect 417 96265 495 96311
rect 541 96265 619 96311
rect 665 96265 743 96311
rect 789 96265 867 96311
rect 913 96265 991 96311
rect 1037 96265 1115 96311
rect 1161 96265 1239 96311
rect 1285 96265 1363 96311
rect 1409 96265 1487 96311
rect 1533 96265 1611 96311
rect 1657 96265 1735 96311
rect 1781 96265 1859 96311
rect 1905 96265 1983 96311
rect 2029 96265 2107 96311
rect 2153 96265 2231 96311
rect 2277 96265 2355 96311
rect 2401 96265 2479 96311
rect 2525 96265 2603 96311
rect 2649 96265 2727 96311
rect 2773 96265 2851 96311
rect 2897 96265 2975 96311
rect 3021 96265 3099 96311
rect 3145 96265 3223 96311
rect 3269 96265 3347 96311
rect 3393 96265 3471 96311
rect 3517 96265 3595 96311
rect 3641 96265 3719 96311
rect 3765 96265 3843 96311
rect 3889 96265 3967 96311
rect 4013 96265 4091 96311
rect 4137 96265 4215 96311
rect 4261 96265 4339 96311
rect 4385 96265 4463 96311
rect 4509 96265 4587 96311
rect 4633 96265 4711 96311
rect 4757 96265 4835 96311
rect 4881 96265 4959 96311
rect 5005 96265 5083 96311
rect 5129 96265 5207 96311
rect 5253 96265 5331 96311
rect 5377 96265 5455 96311
rect 5501 96265 5579 96311
rect 5625 96265 5703 96311
rect 5749 96265 5827 96311
rect 5873 96265 5951 96311
rect 5997 96265 6075 96311
rect 6121 96265 6199 96311
rect 6245 96265 6323 96311
rect 6369 96265 6447 96311
rect 6493 96265 6571 96311
rect 6617 96265 6695 96311
rect 6741 96265 6819 96311
rect 6865 96265 6943 96311
rect 6989 96265 7067 96311
rect 7113 96265 7191 96311
rect 7237 96265 7315 96311
rect 7361 96265 7439 96311
rect 7485 96265 7563 96311
rect 7609 96265 7687 96311
rect 7733 96265 7811 96311
rect 7857 96265 7935 96311
rect 7981 96265 8059 96311
rect 8105 96265 8183 96311
rect 8229 96265 8307 96311
rect 8353 96265 8431 96311
rect 8477 96265 8555 96311
rect 8601 96265 8679 96311
rect 8725 96265 8803 96311
rect 8849 96265 8927 96311
rect 8973 96265 9051 96311
rect 9097 96265 9175 96311
rect 9221 96265 9299 96311
rect 9345 96265 9423 96311
rect 9469 96265 9547 96311
rect 9593 96265 9671 96311
rect 9717 96265 9795 96311
rect 9841 96265 9919 96311
rect 9965 96265 10043 96311
rect 10089 96265 10167 96311
rect 10213 96265 10291 96311
rect 10337 96265 10415 96311
rect 10461 96265 10539 96311
rect 10585 96265 10663 96311
rect 10709 96265 10787 96311
rect 10833 96265 10911 96311
rect 10957 96265 11035 96311
rect 11081 96265 11159 96311
rect 11205 96265 11283 96311
rect 11329 96265 11407 96311
rect 11453 96265 11531 96311
rect 11577 96265 11655 96311
rect 11701 96265 11779 96311
rect 11825 96265 11903 96311
rect 11949 96265 12027 96311
rect 12073 96265 12151 96311
rect 12197 96265 12275 96311
rect 12321 96265 12399 96311
rect 12445 96265 12523 96311
rect 12569 96265 12647 96311
rect 12693 96265 12771 96311
rect 12817 96265 12895 96311
rect 12941 96265 13019 96311
rect 13065 96265 13143 96311
rect 13189 96265 13267 96311
rect 13313 96265 13391 96311
rect 13437 96265 13515 96311
rect 13561 96265 13639 96311
rect 13685 96265 13763 96311
rect 13809 96265 13887 96311
rect 13933 96265 14011 96311
rect 14057 96265 14135 96311
rect 14181 96265 14259 96311
rect 14305 96265 14383 96311
rect 14429 96265 14507 96311
rect 14553 96265 14631 96311
rect 14677 96265 14755 96311
rect 14801 96265 14879 96311
rect 14925 96265 15003 96311
rect 15049 96265 15127 96311
rect 15173 96265 15251 96311
rect 15297 96265 15375 96311
rect 15421 96265 15499 96311
rect 15545 96265 15623 96311
rect 15669 96265 15747 96311
rect 15793 96265 15871 96311
rect 15917 96265 15995 96311
rect 16041 96265 16119 96311
rect 16165 96265 16243 96311
rect 16289 96265 16367 96311
rect 16413 96265 16491 96311
rect 16537 96265 16615 96311
rect 16661 96265 16739 96311
rect 16785 96265 16863 96311
rect 16909 96265 16987 96311
rect 17033 96265 17111 96311
rect 17157 96265 17235 96311
rect 17281 96265 17359 96311
rect 17405 96265 17483 96311
rect 17529 96265 17607 96311
rect 17653 96265 17731 96311
rect 17777 96265 17855 96311
rect 17901 96265 17979 96311
rect 18025 96265 18103 96311
rect 18149 96265 18227 96311
rect 18273 96265 18351 96311
rect 18397 96265 18475 96311
rect 18521 96265 18599 96311
rect 18645 96265 18723 96311
rect 18769 96265 18847 96311
rect 18893 96265 18971 96311
rect 19017 96265 19095 96311
rect 19141 96265 19219 96311
rect 19265 96265 19343 96311
rect 19389 96265 19467 96311
rect 19513 96265 19591 96311
rect 19637 96265 19715 96311
rect 19761 96265 19839 96311
rect 19885 96265 19963 96311
rect 20009 96265 20087 96311
rect 20133 96265 20211 96311
rect 20257 96265 20335 96311
rect 20381 96265 20459 96311
rect 20505 96265 20583 96311
rect 20629 96265 20707 96311
rect 20753 96265 20831 96311
rect 20877 96265 20955 96311
rect 21001 96265 21079 96311
rect 21125 96265 21203 96311
rect 21249 96265 21327 96311
rect 21373 96265 21451 96311
rect 21497 96265 21575 96311
rect 21621 96265 21699 96311
rect 21745 96265 21823 96311
rect 21869 96265 21947 96311
rect 21993 96265 22071 96311
rect 22117 96265 22195 96311
rect 22241 96265 22319 96311
rect 22365 96265 22443 96311
rect 22489 96265 22567 96311
rect 22613 96265 22691 96311
rect 22737 96265 22815 96311
rect 22861 96265 22939 96311
rect 22985 96265 23063 96311
rect 23109 96265 23187 96311
rect 23233 96265 23311 96311
rect 23357 96265 23435 96311
rect 23481 96265 23559 96311
rect 23605 96265 23683 96311
rect 23729 96265 23807 96311
rect 23853 96265 23931 96311
rect 23977 96265 24055 96311
rect 24101 96265 24179 96311
rect 24225 96265 24303 96311
rect 24349 96265 24427 96311
rect 24473 96265 24551 96311
rect 24597 96265 24675 96311
rect 24721 96265 24799 96311
rect 24845 96265 24923 96311
rect 24969 96265 25047 96311
rect 25093 96265 25171 96311
rect 25217 96265 25295 96311
rect 25341 96265 25419 96311
rect 25465 96265 25543 96311
rect 25589 96265 25667 96311
rect 25713 96265 25791 96311
rect 25837 96265 25915 96311
rect 25961 96265 26039 96311
rect 26085 96265 26163 96311
rect 26209 96265 26287 96311
rect 26333 96265 26411 96311
rect 26457 96265 26535 96311
rect 26581 96265 26659 96311
rect 26705 96265 26783 96311
rect 26829 96265 26907 96311
rect 26953 96265 27031 96311
rect 27077 96265 27155 96311
rect 27201 96265 27279 96311
rect 27325 96265 27403 96311
rect 27449 96265 27527 96311
rect 27573 96265 27651 96311
rect 27697 96265 27775 96311
rect 27821 96265 27899 96311
rect 27945 96265 28023 96311
rect 28069 96265 28147 96311
rect 28193 96265 28271 96311
rect 28317 96265 28395 96311
rect 28441 96265 28519 96311
rect 28565 96265 28643 96311
rect 28689 96265 28767 96311
rect 28813 96265 28891 96311
rect 28937 96265 29015 96311
rect 29061 96265 29139 96311
rect 29185 96265 29263 96311
rect 29309 96265 29387 96311
rect 29433 96265 29511 96311
rect 29557 96265 29635 96311
rect 29681 96265 29759 96311
rect 29805 96265 29883 96311
rect 29929 96265 30007 96311
rect 30053 96265 30131 96311
rect 30177 96265 30255 96311
rect 30301 96265 30379 96311
rect 30425 96265 30503 96311
rect 30549 96265 30627 96311
rect 30673 96265 30751 96311
rect 30797 96265 30875 96311
rect 30921 96265 30999 96311
rect 31045 96265 31123 96311
rect 31169 96265 31247 96311
rect 31293 96265 31371 96311
rect 31417 96265 31495 96311
rect 31541 96265 31619 96311
rect 31665 96265 31743 96311
rect 31789 96265 31867 96311
rect 31913 96265 31991 96311
rect 32037 96265 32115 96311
rect 32161 96265 32239 96311
rect 32285 96265 32363 96311
rect 32409 96265 32487 96311
rect 32533 96265 32611 96311
rect 32657 96265 32735 96311
rect 32781 96265 32859 96311
rect 32905 96265 32983 96311
rect 33029 96265 33107 96311
rect 33153 96265 33231 96311
rect 33277 96265 33355 96311
rect 33401 96265 33479 96311
rect 33525 96265 33603 96311
rect 33649 96265 33727 96311
rect 33773 96265 33851 96311
rect 33897 96265 33975 96311
rect 34021 96265 34099 96311
rect 34145 96265 34223 96311
rect 34269 96265 34347 96311
rect 34393 96265 34471 96311
rect 34517 96265 34595 96311
rect 34641 96265 34719 96311
rect 34765 96265 34843 96311
rect 34889 96265 34967 96311
rect 35013 96265 35091 96311
rect 35137 96265 35215 96311
rect 35261 96265 35339 96311
rect 35385 96265 35463 96311
rect 35509 96265 35587 96311
rect 35633 96265 35711 96311
rect 35757 96265 35835 96311
rect 35881 96265 35959 96311
rect 36005 96265 36083 96311
rect 36129 96265 36207 96311
rect 36253 96265 36331 96311
rect 36377 96265 36455 96311
rect 36501 96265 36579 96311
rect 36625 96265 36703 96311
rect 36749 96265 36827 96311
rect 36873 96265 36951 96311
rect 36997 96265 37075 96311
rect 37121 96265 37199 96311
rect 37245 96265 37323 96311
rect 37369 96265 37447 96311
rect 37493 96265 37571 96311
rect 37617 96265 37695 96311
rect 37741 96265 37819 96311
rect 37865 96265 37943 96311
rect 37989 96265 38067 96311
rect 38113 96265 38191 96311
rect 38237 96265 38315 96311
rect 38361 96265 38439 96311
rect 38485 96265 38563 96311
rect 38609 96265 38687 96311
rect 38733 96265 38811 96311
rect 38857 96265 38935 96311
rect 38981 96265 39059 96311
rect 39105 96265 39183 96311
rect 39229 96265 39307 96311
rect 39353 96265 39431 96311
rect 39477 96265 39555 96311
rect 39601 96265 39679 96311
rect 39725 96265 39803 96311
rect 39849 96265 39927 96311
rect 39973 96265 40051 96311
rect 40097 96265 40175 96311
rect 40221 96265 40299 96311
rect 40345 96265 40423 96311
rect 40469 96265 40547 96311
rect 40593 96265 40671 96311
rect 40717 96265 40795 96311
rect 40841 96265 40919 96311
rect 40965 96265 41043 96311
rect 41089 96265 41167 96311
rect 41213 96265 41291 96311
rect 41337 96265 41415 96311
rect 41461 96265 41539 96311
rect 41585 96265 41663 96311
rect 41709 96265 41787 96311
rect 41833 96265 41911 96311
rect 41957 96265 42035 96311
rect 42081 96265 42159 96311
rect 42205 96265 42283 96311
rect 42329 96265 42407 96311
rect 42453 96265 42531 96311
rect 42577 96265 42655 96311
rect 42701 96265 42779 96311
rect 42825 96265 42903 96311
rect 42949 96265 43027 96311
rect 43073 96265 43151 96311
rect 43197 96265 43275 96311
rect 43321 96265 43399 96311
rect 43445 96265 43523 96311
rect 43569 96265 43647 96311
rect 43693 96265 43771 96311
rect 43817 96265 43895 96311
rect 43941 96265 44019 96311
rect 44065 96265 44143 96311
rect 44189 96265 44267 96311
rect 44313 96265 44391 96311
rect 44437 96265 44515 96311
rect 44561 96265 44639 96311
rect 44685 96265 44763 96311
rect 44809 96265 44887 96311
rect 44933 96265 45011 96311
rect 45057 96265 45135 96311
rect 45181 96265 45259 96311
rect 45305 96265 45383 96311
rect 45429 96265 45507 96311
rect 45553 96265 45631 96311
rect 45677 96265 45755 96311
rect 45801 96265 45879 96311
rect 45925 96265 46003 96311
rect 46049 96265 46127 96311
rect 46173 96265 46251 96311
rect 46297 96265 46375 96311
rect 46421 96265 46499 96311
rect 46545 96265 46623 96311
rect 46669 96265 46747 96311
rect 46793 96265 46871 96311
rect 46917 96265 46995 96311
rect 47041 96265 47119 96311
rect 47165 96265 47243 96311
rect 47289 96265 47367 96311
rect 47413 96265 47491 96311
rect 47537 96265 47615 96311
rect 47661 96265 47739 96311
rect 47785 96265 47863 96311
rect 47909 96265 47987 96311
rect 48033 96265 48111 96311
rect 48157 96265 48235 96311
rect 48281 96265 48359 96311
rect 48405 96265 48483 96311
rect 48529 96265 48607 96311
rect 48653 96265 48731 96311
rect 48777 96265 48855 96311
rect 48901 96265 48979 96311
rect 49025 96265 49103 96311
rect 49149 96265 49227 96311
rect 49273 96265 49351 96311
rect 49397 96265 49475 96311
rect 49521 96265 49599 96311
rect 49645 96265 49723 96311
rect 49769 96265 49847 96311
rect 49893 96265 49971 96311
rect 50017 96265 50095 96311
rect 50141 96265 50219 96311
rect 50265 96265 50343 96311
rect 50389 96265 50467 96311
rect 50513 96265 50591 96311
rect 50637 96265 50715 96311
rect 50761 96265 50839 96311
rect 50885 96265 50963 96311
rect 51009 96265 51087 96311
rect 51133 96265 51211 96311
rect 51257 96265 51335 96311
rect 51381 96265 51459 96311
rect 51505 96265 51583 96311
rect 51629 96265 51707 96311
rect 51753 96265 51831 96311
rect 51877 96265 51955 96311
rect 52001 96265 52079 96311
rect 52125 96265 52203 96311
rect 52249 96265 52327 96311
rect 52373 96265 52451 96311
rect 52497 96265 52575 96311
rect 52621 96265 52699 96311
rect 52745 96265 52823 96311
rect 52869 96265 52947 96311
rect 52993 96265 53071 96311
rect 53117 96265 53195 96311
rect 53241 96265 53319 96311
rect 53365 96265 53443 96311
rect 53489 96265 53567 96311
rect 53613 96265 53691 96311
rect 53737 96265 53815 96311
rect 53861 96265 53939 96311
rect 53985 96265 54063 96311
rect 54109 96265 54187 96311
rect 54233 96265 54311 96311
rect 54357 96265 54435 96311
rect 54481 96265 54559 96311
rect 54605 96265 54683 96311
rect 54729 96265 54807 96311
rect 54853 96265 54931 96311
rect 54977 96265 55055 96311
rect 55101 96265 55179 96311
rect 55225 96265 55303 96311
rect 55349 96265 55427 96311
rect 55473 96265 55551 96311
rect 55597 96265 55675 96311
rect 55721 96265 55799 96311
rect 55845 96265 55923 96311
rect 55969 96265 56047 96311
rect 56093 96265 56171 96311
rect 56217 96265 56295 96311
rect 56341 96265 56419 96311
rect 56465 96265 56543 96311
rect 56589 96265 56667 96311
rect 56713 96265 56791 96311
rect 56837 96265 56915 96311
rect 56961 96265 57039 96311
rect 57085 96265 57163 96311
rect 57209 96265 57287 96311
rect 57333 96265 57411 96311
rect 57457 96265 57535 96311
rect 57581 96265 57659 96311
rect 57705 96265 57783 96311
rect 57829 96265 57907 96311
rect 57953 96265 58031 96311
rect 58077 96265 58155 96311
rect 58201 96265 58279 96311
rect 58325 96265 58403 96311
rect 58449 96265 58527 96311
rect 58573 96265 58651 96311
rect 58697 96265 58775 96311
rect 58821 96265 58899 96311
rect 58945 96265 59023 96311
rect 59069 96265 59147 96311
rect 59193 96265 59271 96311
rect 59317 96265 59395 96311
rect 59441 96265 59519 96311
rect 59565 96265 59643 96311
rect 59689 96265 59767 96311
rect 59813 96265 59891 96311
rect 59937 96265 60015 96311
rect 60061 96265 60139 96311
rect 60185 96265 60263 96311
rect 60309 96265 60387 96311
rect 60433 96265 60511 96311
rect 60557 96265 60635 96311
rect 60681 96265 60759 96311
rect 60805 96265 60883 96311
rect 60929 96265 61007 96311
rect 61053 96265 61131 96311
rect 61177 96265 61255 96311
rect 61301 96265 61379 96311
rect 61425 96265 61503 96311
rect 61549 96265 61627 96311
rect 61673 96265 61751 96311
rect 61797 96265 61875 96311
rect 61921 96265 61999 96311
rect 62045 96265 62123 96311
rect 62169 96265 62247 96311
rect 62293 96265 62371 96311
rect 62417 96265 62495 96311
rect 62541 96265 62619 96311
rect 62665 96265 62743 96311
rect 62789 96265 62867 96311
rect 62913 96265 62991 96311
rect 63037 96265 63115 96311
rect 63161 96265 63239 96311
rect 63285 96265 63363 96311
rect 63409 96265 63487 96311
rect 63533 96265 63611 96311
rect 63657 96265 63735 96311
rect 63781 96265 63859 96311
rect 63905 96265 63983 96311
rect 64029 96265 64107 96311
rect 64153 96265 64231 96311
rect 64277 96265 64355 96311
rect 64401 96265 64479 96311
rect 64525 96265 64603 96311
rect 64649 96265 64727 96311
rect 64773 96265 64851 96311
rect 64897 96265 64975 96311
rect 65021 96265 65099 96311
rect 65145 96265 65223 96311
rect 65269 96265 65347 96311
rect 65393 96265 65471 96311
rect 65517 96265 65595 96311
rect 65641 96265 65719 96311
rect 65765 96265 65843 96311
rect 65889 96265 65967 96311
rect 66013 96265 66091 96311
rect 66137 96265 66215 96311
rect 66261 96265 66339 96311
rect 66385 96265 66463 96311
rect 66509 96265 66587 96311
rect 66633 96265 66711 96311
rect 66757 96265 66835 96311
rect 66881 96265 66959 96311
rect 67005 96265 67083 96311
rect 67129 96265 67207 96311
rect 67253 96265 67331 96311
rect 67377 96265 67455 96311
rect 67501 96265 67579 96311
rect 67625 96265 67703 96311
rect 67749 96265 67827 96311
rect 67873 96265 67951 96311
rect 67997 96265 68075 96311
rect 68121 96265 68199 96311
rect 68245 96265 68323 96311
rect 68369 96265 68447 96311
rect 68493 96265 68571 96311
rect 68617 96265 68695 96311
rect 68741 96265 68819 96311
rect 68865 96265 68943 96311
rect 68989 96265 69067 96311
rect 69113 96265 69191 96311
rect 69237 96265 69315 96311
rect 69361 96265 69439 96311
rect 69485 96265 69563 96311
rect 69609 96265 69687 96311
rect 69733 96265 69811 96311
rect 69857 96265 69935 96311
rect 69981 96265 70059 96311
rect 70105 96265 70183 96311
rect 70229 96265 70307 96311
rect 70353 96265 70431 96311
rect 70477 96265 70555 96311
rect 70601 96265 70679 96311
rect 70725 96265 70803 96311
rect 70849 96265 70927 96311
rect 70973 96265 71051 96311
rect 71097 96265 71175 96311
rect 71221 96265 71299 96311
rect 71345 96265 71423 96311
rect 71469 96265 71547 96311
rect 71593 96265 71671 96311
rect 71717 96265 71795 96311
rect 71841 96265 71919 96311
rect 71965 96265 72043 96311
rect 72089 96265 72167 96311
rect 72213 96265 72291 96311
rect 72337 96265 72415 96311
rect 72461 96265 72539 96311
rect 72585 96265 72663 96311
rect 72709 96265 72787 96311
rect 72833 96265 72911 96311
rect 72957 96265 73035 96311
rect 73081 96265 73159 96311
rect 73205 96265 73283 96311
rect 73329 96265 73407 96311
rect 73453 96265 73531 96311
rect 73577 96265 73655 96311
rect 73701 96265 73779 96311
rect 73825 96265 73903 96311
rect 73949 96265 74027 96311
rect 74073 96265 74151 96311
rect 74197 96265 74275 96311
rect 74321 96265 74399 96311
rect 74445 96265 74523 96311
rect 74569 96265 74647 96311
rect 74693 96265 74771 96311
rect 74817 96265 74895 96311
rect 74941 96265 75019 96311
rect 75065 96265 75143 96311
rect 75189 96265 75267 96311
rect 75313 96265 75391 96311
rect 75437 96265 75515 96311
rect 75561 96265 75639 96311
rect 75685 96265 75763 96311
rect 75809 96265 75887 96311
rect 75933 96265 76011 96311
rect 76057 96265 76135 96311
rect 76181 96265 76259 96311
rect 76305 96265 76383 96311
rect 76429 96265 76507 96311
rect 76553 96265 76631 96311
rect 76677 96265 76755 96311
rect 76801 96265 76879 96311
rect 76925 96265 77003 96311
rect 77049 96265 77127 96311
rect 77173 96265 77251 96311
rect 77297 96265 77375 96311
rect 77421 96265 77499 96311
rect 77545 96265 77623 96311
rect 77669 96265 77747 96311
rect 77793 96265 77871 96311
rect 77917 96265 77995 96311
rect 78041 96265 78119 96311
rect 78165 96265 78243 96311
rect 78289 96265 78367 96311
rect 78413 96265 78491 96311
rect 78537 96265 78615 96311
rect 78661 96265 78739 96311
rect 78785 96265 78863 96311
rect 78909 96265 78987 96311
rect 79033 96265 79111 96311
rect 79157 96265 79235 96311
rect 79281 96265 79359 96311
rect 79405 96265 79483 96311
rect 79529 96265 79607 96311
rect 79653 96265 79731 96311
rect 79777 96265 79855 96311
rect 79901 96265 79979 96311
rect 80025 96265 80103 96311
rect 80149 96265 80227 96311
rect 80273 96265 80351 96311
rect 80397 96265 80475 96311
rect 80521 96265 80599 96311
rect 80645 96265 80723 96311
rect 80769 96265 80847 96311
rect 80893 96265 80971 96311
rect 81017 96265 81095 96311
rect 81141 96265 81219 96311
rect 81265 96265 81343 96311
rect 81389 96265 81467 96311
rect 81513 96265 81591 96311
rect 81637 96265 81715 96311
rect 81761 96265 81839 96311
rect 81885 96265 81963 96311
rect 82009 96265 82087 96311
rect 82133 96265 82211 96311
rect 82257 96265 82335 96311
rect 82381 96265 82459 96311
rect 82505 96265 82583 96311
rect 82629 96265 82707 96311
rect 82753 96265 82831 96311
rect 82877 96265 82955 96311
rect 83001 96265 83079 96311
rect 83125 96265 83203 96311
rect 83249 96265 83327 96311
rect 83373 96265 83451 96311
rect 83497 96265 83575 96311
rect 83621 96265 83699 96311
rect 83745 96265 83823 96311
rect 83869 96265 83947 96311
rect 83993 96265 84071 96311
rect 84117 96265 84195 96311
rect 84241 96265 84319 96311
rect 84365 96265 84443 96311
rect 84489 96265 84567 96311
rect 84613 96265 84691 96311
rect 84737 96265 84815 96311
rect 84861 96265 84939 96311
rect 84985 96265 85063 96311
rect 85109 96265 85187 96311
rect 85233 96265 85311 96311
rect 85357 96265 85435 96311
rect 85481 96265 85559 96311
rect 85605 96265 85683 96311
rect 85729 96265 85807 96311
rect 85853 96265 85931 96311
rect 85977 96265 86090 96311
rect 282 96163 86090 96265
rect 282 1117 371 96163
rect 717 95694 27398 96163
rect 717 1282 1282 95694
rect 25312 94773 26039 95694
rect 25312 94721 25388 94773
rect 25440 94721 25512 94773
rect 25564 94721 25636 94773
rect 25688 94721 25760 94773
rect 25812 94721 25884 94773
rect 25936 94721 26039 94773
rect 25312 94649 26039 94721
rect 25312 94597 25388 94649
rect 25440 94597 25512 94649
rect 25564 94597 25636 94649
rect 25688 94597 25760 94649
rect 25812 94597 25884 94649
rect 25936 94597 26039 94649
rect 25312 94525 26039 94597
rect 25312 94473 25388 94525
rect 25440 94473 25512 94525
rect 25564 94473 25636 94525
rect 25688 94473 25760 94525
rect 25812 94473 25884 94525
rect 25936 94473 26039 94525
rect 25312 94454 26039 94473
rect 25376 34990 25948 35002
rect 25376 34938 25388 34990
rect 25440 34938 25512 34990
rect 25564 34938 25636 34990
rect 25688 34938 25760 34990
rect 25812 34938 25884 34990
rect 25936 34938 25948 34990
rect 25376 34866 25948 34938
rect 25376 34814 25388 34866
rect 25440 34814 25512 34866
rect 25564 34814 25636 34866
rect 25688 34814 25760 34866
rect 25812 34814 25884 34866
rect 25936 34814 25948 34866
rect 25376 34742 25948 34814
rect 25376 34690 25388 34742
rect 25440 34690 25512 34742
rect 25564 34690 25636 34742
rect 25688 34690 25760 34742
rect 25812 34690 25884 34742
rect 25936 34690 25948 34742
rect 25376 34618 25948 34690
rect 27387 34631 27398 95694
rect 27744 96142 57306 96163
rect 27744 94653 27822 96142
rect 28668 95694 56382 96142
rect 28668 94653 29197 95694
rect 34227 94671 35013 95694
rect 40062 94671 40590 95694
rect 43738 94671 44564 95694
rect 27744 94601 27790 94653
rect 28686 94601 28845 94653
rect 28897 94601 29056 94653
rect 29108 94601 29197 94653
rect 27744 92853 27822 94601
rect 28668 92853 29197 94601
rect 50098 94485 50913 95694
rect 55927 94653 56382 95694
rect 57228 94653 57306 96142
rect 57652 95694 85733 96163
rect 55927 94601 56015 94653
rect 56067 94601 56226 94653
rect 56278 94601 56382 94653
rect 57228 94601 57281 94653
rect 27744 92801 27790 92853
rect 28686 92801 28845 92853
rect 28897 92801 29056 92853
rect 29108 92801 29197 92853
rect 27744 91053 27822 92801
rect 28668 91053 29197 92801
rect 27744 91001 27790 91053
rect 28686 91001 28845 91053
rect 28897 91001 29056 91053
rect 29108 91001 29197 91053
rect 27744 89253 27822 91001
rect 28668 89253 29197 91001
rect 27744 89201 27790 89253
rect 28686 89201 28845 89253
rect 28897 89201 29056 89253
rect 29108 89201 29197 89253
rect 27744 87453 27822 89201
rect 28668 87453 29197 89201
rect 27744 87401 27790 87453
rect 28686 87401 28845 87453
rect 28897 87401 29056 87453
rect 29108 87401 29197 87453
rect 27744 85653 27822 87401
rect 28668 85653 29197 87401
rect 27744 85601 27790 85653
rect 28686 85601 28845 85653
rect 28897 85601 29056 85653
rect 29108 85601 29197 85653
rect 27744 83853 27822 85601
rect 28668 83853 29197 85601
rect 27744 83801 27790 83853
rect 28686 83801 28845 83853
rect 28897 83801 29056 83853
rect 29108 83801 29197 83853
rect 27744 82053 27822 83801
rect 28668 82053 29197 83801
rect 27744 82001 27790 82053
rect 28686 82001 28845 82053
rect 28897 82001 29056 82053
rect 29108 82001 29197 82053
rect 27744 80253 27822 82001
rect 28668 80253 29197 82001
rect 27744 80201 27790 80253
rect 28686 80201 28845 80253
rect 28897 80201 29056 80253
rect 29108 80201 29197 80253
rect 27744 78453 27822 80201
rect 28668 78453 29197 80201
rect 27744 78401 27790 78453
rect 28686 78401 28845 78453
rect 28897 78401 29056 78453
rect 29108 78401 29197 78453
rect 27744 76653 27822 78401
rect 28668 76653 29197 78401
rect 27744 76601 27790 76653
rect 28686 76601 28845 76653
rect 28897 76601 29056 76653
rect 29108 76601 29197 76653
rect 27744 74853 27822 76601
rect 28668 74853 29197 76601
rect 27744 74801 27790 74853
rect 28686 74801 28845 74853
rect 28897 74801 29056 74853
rect 29108 74801 29197 74853
rect 27744 73053 27822 74801
rect 28668 73053 29197 74801
rect 27744 73001 27790 73053
rect 28686 73001 28845 73053
rect 28897 73001 29056 73053
rect 29108 73001 29197 73053
rect 27744 71253 27822 73001
rect 28668 71253 29197 73001
rect 27744 71201 27790 71253
rect 28686 71201 28845 71253
rect 28897 71201 29056 71253
rect 29108 71201 29197 71253
rect 27744 69453 27822 71201
rect 28668 69453 29197 71201
rect 27744 69401 27790 69453
rect 28686 69401 28845 69453
rect 28897 69401 29056 69453
rect 29108 69401 29197 69453
rect 27744 67653 27822 69401
rect 28668 67653 29197 69401
rect 27744 67601 27790 67653
rect 28686 67601 28845 67653
rect 28897 67601 29056 67653
rect 29108 67601 29197 67653
rect 27744 65853 27822 67601
rect 28668 65853 29197 67601
rect 27744 65801 27790 65853
rect 28686 65801 28845 65853
rect 28897 65801 29056 65853
rect 29108 65801 29197 65853
rect 27744 64053 27822 65801
rect 28668 64053 29197 65801
rect 27744 64001 27790 64053
rect 28686 64001 28845 64053
rect 28897 64001 29056 64053
rect 29108 64001 29197 64053
rect 27744 62253 27822 64001
rect 28668 62253 29197 64001
rect 27744 62201 27790 62253
rect 28686 62201 28845 62253
rect 28897 62201 29056 62253
rect 29108 62201 29197 62253
rect 27744 60453 27822 62201
rect 28668 60453 29197 62201
rect 27744 60401 27790 60453
rect 28686 60401 28845 60453
rect 28897 60401 29056 60453
rect 29108 60401 29197 60453
rect 27744 58653 27822 60401
rect 28668 58653 29197 60401
rect 27744 58601 27790 58653
rect 28686 58601 28845 58653
rect 28897 58601 29056 58653
rect 29108 58601 29197 58653
rect 27744 56853 27822 58601
rect 28668 56853 29197 58601
rect 27744 56801 27790 56853
rect 28686 56801 28845 56853
rect 28897 56801 29056 56853
rect 29108 56801 29197 56853
rect 27744 55053 27822 56801
rect 28668 55053 29197 56801
rect 27744 55001 27790 55053
rect 28686 55001 28845 55053
rect 28897 55001 29056 55053
rect 29108 55001 29197 55053
rect 27744 53253 27822 55001
rect 28668 53253 29197 55001
rect 27744 53201 27790 53253
rect 28686 53201 28845 53253
rect 28897 53201 29056 53253
rect 29108 53201 29197 53253
rect 27744 51453 27822 53201
rect 28668 51453 29197 53201
rect 27744 51401 27790 51453
rect 28686 51401 28845 51453
rect 28897 51401 29056 51453
rect 29108 51401 29197 51453
rect 27744 49653 27822 51401
rect 28668 49653 29197 51401
rect 27744 49601 27790 49653
rect 28686 49601 28845 49653
rect 28897 49601 29056 49653
rect 29108 49601 29197 49653
rect 27744 47853 27822 49601
rect 28668 47853 29197 49601
rect 27744 47801 27790 47853
rect 28686 47801 28845 47853
rect 28897 47801 29056 47853
rect 29108 47801 29197 47853
rect 27744 46053 27822 47801
rect 28668 46053 29197 47801
rect 27744 46001 27790 46053
rect 28686 46001 28845 46053
rect 28897 46001 29056 46053
rect 29108 46001 29197 46053
rect 27744 44253 27822 46001
rect 28668 44253 29197 46001
rect 27744 44201 27790 44253
rect 28686 44201 28845 44253
rect 28897 44201 29056 44253
rect 29108 44201 29197 44253
rect 27744 42453 27822 44201
rect 28668 42453 29197 44201
rect 27744 42401 27790 42453
rect 28686 42401 28845 42453
rect 28897 42401 29056 42453
rect 29108 42401 29197 42453
rect 27744 40653 27822 42401
rect 28668 40653 29197 42401
rect 27744 40601 27790 40653
rect 28686 40601 28845 40653
rect 28897 40601 29056 40653
rect 29108 40601 29197 40653
rect 27744 38853 27822 40601
rect 28668 38853 29197 40601
rect 27744 38801 27790 38853
rect 28686 38801 28845 38853
rect 28897 38801 29056 38853
rect 29108 38801 29197 38853
rect 27744 37053 27822 38801
rect 28668 37053 29197 38801
rect 27744 37001 27790 37053
rect 28686 37001 28845 37053
rect 28897 37001 29056 37053
rect 29108 37001 29197 37053
rect 27744 35996 27822 37001
rect 28668 35996 29197 37001
rect 27744 35985 29197 35996
rect 55927 92853 56382 94601
rect 57228 92853 57306 94601
rect 55927 92801 56015 92853
rect 56067 92801 56226 92853
rect 56278 92801 56382 92853
rect 57228 92801 57281 92853
rect 55927 91053 56382 92801
rect 57228 91053 57306 92801
rect 55927 91001 56015 91053
rect 56067 91001 56226 91053
rect 56278 91001 56382 91053
rect 57228 91001 57281 91053
rect 55927 89253 56382 91001
rect 57228 89253 57306 91001
rect 55927 89201 56015 89253
rect 56067 89201 56226 89253
rect 56278 89201 56382 89253
rect 57228 89201 57281 89253
rect 55927 87453 56382 89201
rect 57228 87453 57306 89201
rect 55927 87401 56015 87453
rect 56067 87401 56226 87453
rect 56278 87401 56382 87453
rect 57228 87401 57281 87453
rect 55927 85653 56382 87401
rect 57228 85653 57306 87401
rect 55927 85601 56015 85653
rect 56067 85601 56226 85653
rect 56278 85601 56382 85653
rect 57228 85601 57281 85653
rect 55927 83853 56382 85601
rect 57228 83853 57306 85601
rect 55927 83801 56015 83853
rect 56067 83801 56226 83853
rect 56278 83801 56382 83853
rect 57228 83801 57281 83853
rect 55927 82053 56382 83801
rect 57228 82053 57306 83801
rect 55927 82001 56015 82053
rect 56067 82001 56226 82053
rect 56278 82001 56382 82053
rect 57228 82001 57281 82053
rect 55927 80253 56382 82001
rect 57228 80253 57306 82001
rect 55927 80201 56015 80253
rect 56067 80201 56226 80253
rect 56278 80201 56382 80253
rect 57228 80201 57281 80253
rect 55927 78453 56382 80201
rect 57228 78453 57306 80201
rect 55927 78401 56015 78453
rect 56067 78401 56226 78453
rect 56278 78401 56382 78453
rect 57228 78401 57281 78453
rect 55927 76653 56382 78401
rect 57228 76653 57306 78401
rect 55927 76601 56015 76653
rect 56067 76601 56226 76653
rect 56278 76601 56382 76653
rect 57228 76601 57281 76653
rect 55927 74853 56382 76601
rect 57228 74853 57306 76601
rect 55927 74801 56015 74853
rect 56067 74801 56226 74853
rect 56278 74801 56382 74853
rect 57228 74801 57281 74853
rect 55927 73053 56382 74801
rect 57228 73053 57306 74801
rect 55927 73001 56015 73053
rect 56067 73001 56226 73053
rect 56278 73001 56382 73053
rect 57228 73001 57281 73053
rect 55927 71253 56382 73001
rect 57228 71253 57306 73001
rect 55927 71201 56015 71253
rect 56067 71201 56226 71253
rect 56278 71201 56382 71253
rect 57228 71201 57281 71253
rect 55927 69453 56382 71201
rect 57228 69453 57306 71201
rect 55927 69401 56015 69453
rect 56067 69401 56226 69453
rect 56278 69401 56382 69453
rect 57228 69401 57281 69453
rect 55927 67653 56382 69401
rect 57228 67653 57306 69401
rect 55927 67601 56015 67653
rect 56067 67601 56226 67653
rect 56278 67601 56382 67653
rect 57228 67601 57281 67653
rect 55927 65853 56382 67601
rect 57228 65853 57306 67601
rect 55927 65801 56015 65853
rect 56067 65801 56226 65853
rect 56278 65801 56382 65853
rect 57228 65801 57281 65853
rect 55927 64053 56382 65801
rect 57228 64053 57306 65801
rect 55927 64001 56015 64053
rect 56067 64001 56226 64053
rect 56278 64001 56382 64053
rect 57228 64001 57281 64053
rect 55927 62253 56382 64001
rect 57228 62253 57306 64001
rect 55927 62201 56015 62253
rect 56067 62201 56226 62253
rect 56278 62201 56382 62253
rect 57228 62201 57281 62253
rect 55927 60453 56382 62201
rect 57228 60453 57306 62201
rect 55927 60401 56015 60453
rect 56067 60401 56226 60453
rect 56278 60401 56382 60453
rect 57228 60401 57281 60453
rect 55927 58653 56382 60401
rect 57228 58653 57306 60401
rect 55927 58601 56015 58653
rect 56067 58601 56226 58653
rect 56278 58601 56382 58653
rect 57228 58601 57281 58653
rect 55927 56853 56382 58601
rect 57228 56853 57306 58601
rect 55927 56801 56015 56853
rect 56067 56801 56226 56853
rect 56278 56801 56382 56853
rect 57228 56801 57281 56853
rect 55927 55053 56382 56801
rect 57228 55053 57306 56801
rect 55927 55001 56015 55053
rect 56067 55001 56226 55053
rect 56278 55001 56382 55053
rect 57228 55001 57281 55053
rect 55927 53253 56382 55001
rect 57228 53253 57306 55001
rect 55927 53201 56015 53253
rect 56067 53201 56226 53253
rect 56278 53201 56382 53253
rect 57228 53201 57281 53253
rect 55927 51453 56382 53201
rect 57228 51453 57306 53201
rect 55927 51401 56015 51453
rect 56067 51401 56226 51453
rect 56278 51401 56382 51453
rect 57228 51401 57281 51453
rect 55927 49653 56382 51401
rect 57228 49653 57306 51401
rect 55927 49601 56015 49653
rect 56067 49601 56226 49653
rect 56278 49601 56382 49653
rect 57228 49601 57281 49653
rect 55927 47853 56382 49601
rect 57228 47853 57306 49601
rect 55927 47801 56015 47853
rect 56067 47801 56226 47853
rect 56278 47801 56382 47853
rect 57228 47801 57281 47853
rect 55927 46053 56382 47801
rect 57228 46053 57306 47801
rect 55927 46001 56015 46053
rect 56067 46001 56226 46053
rect 56278 46001 56382 46053
rect 57228 46001 57281 46053
rect 55927 44253 56382 46001
rect 57228 44253 57306 46001
rect 55927 44201 56015 44253
rect 56067 44201 56226 44253
rect 56278 44201 56382 44253
rect 57228 44201 57281 44253
rect 55927 42453 56382 44201
rect 57228 42453 57306 44201
rect 55927 42401 56015 42453
rect 56067 42401 56226 42453
rect 56278 42401 56382 42453
rect 57228 42401 57281 42453
rect 55927 40653 56382 42401
rect 57228 40653 57306 42401
rect 55927 40601 56015 40653
rect 56067 40601 56226 40653
rect 56278 40601 56382 40653
rect 57228 40601 57281 40653
rect 55927 38853 56382 40601
rect 57228 38853 57306 40601
rect 55927 38801 56015 38853
rect 56067 38801 56226 38853
rect 56278 38801 56382 38853
rect 57228 38801 57281 38853
rect 55927 37053 56382 38801
rect 57228 37053 57306 38801
rect 55927 37001 56015 37053
rect 56067 37001 56226 37053
rect 56278 37001 56382 37053
rect 57228 37001 57281 37053
rect 55927 35996 56382 37001
rect 57228 35996 57306 37001
rect 55927 35985 57306 35996
rect 27744 34990 27828 35985
rect 27749 34938 27828 34990
rect 27744 34866 27828 34938
rect 27749 34814 27828 34866
rect 27744 34742 27828 34814
rect 27749 34690 27828 34742
rect 25376 34566 25388 34618
rect 25440 34566 25512 34618
rect 25564 34566 25636 34618
rect 25688 34566 25760 34618
rect 25812 34566 25884 34618
rect 25936 34566 25948 34618
rect 25376 34554 25948 34566
rect 27386 34163 27398 34631
rect 27744 34631 27828 34690
rect 57295 34631 57306 35985
rect 27744 34620 57306 34631
rect 27744 34618 27822 34620
rect 27749 34566 27822 34618
rect 26772 33432 27214 33519
rect 26772 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27214 33432
rect 26772 33215 27214 33380
rect 26772 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27214 33215
rect 26772 32997 27214 33163
rect 26772 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27214 32997
rect 26772 32779 27214 32945
rect 26772 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27214 32779
rect 26772 32562 27214 32727
rect 26772 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27214 32562
rect 26772 32344 27214 32510
rect 26772 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27214 32344
rect 26772 32127 27214 32292
rect 26772 32075 26861 32127
rect 26913 32075 27073 32127
rect 27125 32075 27214 32127
rect 26772 31909 27214 32075
rect 26772 31857 26861 31909
rect 26913 31857 27073 31909
rect 27125 31857 27214 31909
rect 26772 31691 27214 31857
rect 26772 31639 26861 31691
rect 26913 31639 27073 31691
rect 27125 31639 27214 31691
rect 26772 31474 27214 31639
rect 26772 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27214 31474
rect 26772 31256 27214 31422
rect 26772 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27214 31256
rect 26772 31038 27214 31204
rect 26772 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27214 31038
rect 26772 30821 27214 30986
rect 26772 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27214 30821
rect 26772 30603 27214 30769
rect 26772 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27214 30603
rect 26772 30386 27214 30551
rect 26772 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27214 30386
rect 26772 30168 27214 30334
rect 26772 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27214 30168
rect 26772 29950 27214 30116
rect 26772 29898 26861 29950
rect 26913 29898 27073 29950
rect 27125 29898 27214 29950
rect 26772 29733 27214 29898
rect 26772 29681 26861 29733
rect 26913 29681 27073 29733
rect 27125 29681 27214 29733
rect 26772 29515 27214 29681
rect 26772 29463 26861 29515
rect 26913 29463 27073 29515
rect 27125 29463 27214 29515
rect 26772 29297 27214 29463
rect 26772 29245 26861 29297
rect 26913 29245 27073 29297
rect 27125 29245 27214 29297
rect 26772 29080 27214 29245
rect 26772 29028 26861 29080
rect 26913 29028 27073 29080
rect 27125 29028 27214 29080
rect 26772 28862 27214 29028
rect 26772 28810 26861 28862
rect 26913 28810 27073 28862
rect 27125 28810 27214 28862
rect 26772 28644 27214 28810
rect 26772 28592 26861 28644
rect 26913 28592 27073 28644
rect 27125 28592 27214 28644
rect 26772 28427 27214 28592
rect 26772 28375 26861 28427
rect 26913 28375 27073 28427
rect 27125 28375 27214 28427
rect 26772 28209 27214 28375
rect 26772 28157 26861 28209
rect 26913 28157 27073 28209
rect 27125 28157 27214 28209
rect 26772 27992 27214 28157
rect 26772 27940 26861 27992
rect 26913 27940 27073 27992
rect 27125 27940 27214 27992
rect 26772 27774 27214 27940
rect 26772 27722 26861 27774
rect 26913 27722 27073 27774
rect 27125 27722 27214 27774
rect 26772 27556 27214 27722
rect 26772 27504 26861 27556
rect 26913 27504 27073 27556
rect 27125 27504 27214 27556
rect 26772 27339 27214 27504
rect 26772 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27214 27339
rect 26772 27121 27214 27287
rect 26772 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27214 27121
rect 26772 26903 27214 27069
rect 26772 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27214 26903
rect 26772 26686 27214 26851
rect 26772 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27214 26686
rect 26772 26468 27214 26634
rect 26772 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27214 26468
rect 26772 26250 27214 26416
rect 26772 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27214 26250
rect 26772 26033 27214 26198
rect 26772 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27214 26033
rect 26772 25815 27214 25981
rect 26772 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27214 25815
rect 26772 25598 27214 25763
rect 26772 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27214 25598
rect 26772 25380 27214 25546
rect 26772 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27214 25380
rect 26772 25162 27214 25328
rect 26772 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27214 25162
rect 26772 24945 27214 25110
rect 26772 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27214 24945
rect 26772 24727 27214 24893
rect 26772 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27214 24727
rect 26772 24509 27214 24675
rect 26772 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27214 24509
rect 26772 24292 27214 24457
rect 26772 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27214 24292
rect 26772 24074 27214 24240
rect 26772 24022 26861 24074
rect 26913 24022 27073 24074
rect 27125 24022 27214 24074
rect 26772 23857 27214 24022
rect 26772 23805 26861 23857
rect 26913 23805 27073 23857
rect 27125 23805 27214 23857
rect 26772 23639 27214 23805
rect 26772 23587 26861 23639
rect 26913 23587 27073 23639
rect 27125 23587 27214 23639
rect 26772 23421 27214 23587
rect 26772 23369 26861 23421
rect 26913 23369 27073 23421
rect 27125 23369 27214 23421
rect 26772 23204 27214 23369
rect 26772 23152 26861 23204
rect 26913 23152 27073 23204
rect 27125 23152 27214 23204
rect 26772 22986 27214 23152
rect 26772 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27214 22986
rect 26772 22768 27214 22934
rect 26772 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27214 22768
rect 26772 22551 27214 22716
rect 26772 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27214 22551
rect 26772 22333 27214 22499
rect 26772 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27214 22333
rect 26772 22115 27214 22281
rect 26772 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27214 22115
rect 26772 21898 27214 22063
rect 26772 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27214 21898
rect 26772 21680 27214 21846
rect 26772 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27214 21680
rect 26772 21463 27214 21628
rect 26772 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27214 21463
rect 26772 21245 27214 21411
rect 26772 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27214 21245
rect 26772 21027 27214 21193
rect 26772 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27214 21027
rect 26772 20810 27214 20975
rect 26772 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27214 20810
rect 26772 20592 27214 20758
rect 26772 20540 26861 20592
rect 26913 20540 27073 20592
rect 27125 20540 27214 20592
rect 26772 20374 27214 20540
rect 26772 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27214 20374
rect 26772 20157 27214 20322
rect 26772 20105 26861 20157
rect 26913 20105 27073 20157
rect 27125 20105 27214 20157
rect 26772 19939 27214 20105
rect 26772 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27214 19939
rect 26772 19722 27214 19887
rect 26772 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27214 19722
rect 26772 19504 27214 19670
rect 26772 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27214 19504
rect 26772 19286 27214 19452
rect 26772 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27214 19286
rect 26772 19068 27214 19234
rect 26772 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27214 19068
rect 26772 18851 27214 19016
rect 26772 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27214 18851
rect 26772 18633 27214 18799
rect 26772 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27214 18633
rect 26772 18416 27214 18581
rect 26772 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27214 18416
rect 26772 18198 27214 18364
rect 26772 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27214 18198
rect 26772 17980 27214 18146
rect 26772 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27214 17980
rect 26772 17763 27214 17928
rect 26772 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27214 17763
rect 26772 17545 27214 17711
rect 26772 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27214 17545
rect 26772 17327 27214 17493
rect 26772 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27214 17327
rect 26772 17110 27214 17275
rect 26772 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27214 17110
rect 26772 16892 27214 17058
rect 26772 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27214 16892
rect 26772 16675 27214 16840
rect 26772 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27214 16675
rect 26772 16457 27214 16623
rect 26772 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27214 16457
rect 26772 16239 27214 16405
rect 26772 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27214 16239
rect 26772 16022 27214 16187
rect 26772 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27214 16022
rect 26772 15804 27214 15970
rect 26772 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27214 15804
rect 26772 15586 27214 15752
rect 26772 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27214 15586
rect 26772 15369 27214 15534
rect 26772 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27214 15369
rect 26772 15151 27214 15317
rect 26772 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27214 15151
rect 26772 14933 27214 15099
rect 26772 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27214 14933
rect 26772 14716 27214 14881
rect 26772 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27214 14716
rect 26772 14498 27214 14664
rect 26772 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27214 14498
rect 26772 14281 27214 14446
rect 26772 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27214 14281
rect 26772 14063 27214 14229
rect 26772 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27214 14063
rect 26772 13845 27214 14011
rect 26772 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27214 13845
rect 26772 13628 27214 13793
rect 26772 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27214 13628
rect 26772 13410 27214 13576
rect 26772 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27214 13410
rect 26772 13192 27214 13358
rect 26772 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27214 13192
rect 26772 12975 27214 13140
rect 26772 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27214 12975
rect 26772 12757 27214 12923
rect 26772 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27214 12757
rect 26772 12540 27214 12705
rect 26772 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27214 12540
rect 26772 12322 27214 12488
rect 26772 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27214 12322
rect 26772 12104 27214 12270
rect 26772 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27214 12104
rect 26772 11887 27214 12052
rect 26772 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27214 11887
rect 26772 11669 27214 11835
rect 26772 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27214 11669
rect 26772 11451 27214 11617
rect 26772 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27214 11451
rect 26772 11234 27214 11399
rect 26772 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27214 11234
rect 26772 11016 27214 11182
rect 26772 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27214 11016
rect 26772 10798 27214 10964
rect 26772 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27214 10798
rect 26772 10581 27214 10746
rect 26772 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27214 10581
rect 26772 10363 27214 10529
rect 26772 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27214 10363
rect 26772 10146 27214 10311
rect 26772 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27214 10146
rect 26772 9928 27214 10094
rect 26772 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27214 9928
rect 26772 9710 27214 9876
rect 26772 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27214 9710
rect 26772 9493 27214 9658
rect 26772 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27214 9493
rect 26772 9275 27214 9441
rect 26772 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27214 9275
rect 26772 9057 27214 9223
rect 26772 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27214 9057
rect 26772 8840 27214 9005
rect 26772 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27214 8840
rect 26772 8622 27214 8788
rect 26772 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27214 8622
rect 26772 8404 27214 8570
rect 26772 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27214 8404
rect 26772 8187 27214 8352
rect 26772 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27214 8187
rect 26772 7969 27214 8135
rect 26772 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27214 7969
rect 26772 7752 27214 7917
rect 26772 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27214 7752
rect 26772 7534 27214 7700
rect 26772 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27214 7534
rect 26772 7316 27214 7482
rect 26772 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27214 7316
rect 26772 7099 27214 7264
rect 26772 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27214 7099
rect 26772 6881 27214 7047
rect 26772 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27214 6881
rect 26772 6663 27214 6829
rect 26772 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27214 6663
rect 26772 6446 27214 6611
rect 26772 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27214 6446
rect 26772 6228 27214 6394
rect 26772 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27214 6228
rect 26772 6011 27214 6176
rect 26772 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27214 6011
rect 26772 5793 27214 5959
rect 26772 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27214 5793
rect 26772 5575 27214 5741
rect 26772 5523 26861 5575
rect 26913 5523 27073 5575
rect 27125 5523 27214 5575
rect 26772 5358 27214 5523
rect 26772 5306 26861 5358
rect 26913 5306 27073 5358
rect 27125 5306 27214 5358
rect 26772 4587 27214 5306
rect 26772 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27214 4587
rect 26772 4370 27214 4535
rect 26772 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27214 4370
rect 26772 4152 27214 4318
rect 26772 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27214 4152
rect 26772 3934 27214 4100
rect 26772 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27214 3934
rect 26772 3717 27214 3882
rect 26772 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27214 3717
rect 26772 1777 27214 3665
rect 2562 1689 2742 1701
rect 2562 1637 2574 1689
rect 2730 1637 2742 1689
rect 2562 1625 2742 1637
rect 12627 1689 12807 1701
rect 12627 1637 12639 1689
rect 12795 1637 12807 1689
rect 12627 1625 12807 1637
rect 13077 1689 13257 1701
rect 13077 1637 13089 1689
rect 13245 1637 13257 1689
rect 13077 1625 13257 1637
rect 23427 1689 23607 1701
rect 23427 1637 23439 1689
rect 23595 1637 23607 1689
rect 23427 1625 23607 1637
rect 27387 1282 27398 34163
rect 27744 34174 27822 34566
rect 57168 34174 57306 34620
rect 27744 34163 57306 34174
rect 717 1117 27398 1282
rect 27744 1925 27828 34163
rect 49896 6349 50076 6361
rect 49896 6347 49908 6349
rect 49728 6301 49908 6347
rect 49896 6297 49908 6301
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 51642 5199 51822 5211
rect 51642 5196 51654 5199
rect 49963 5150 51654 5196
rect 51642 5147 51654 5150
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 28628 3906 40180 3917
rect 28628 3860 28639 3906
rect 28685 3860 28755 3906
rect 28801 3860 28871 3906
rect 28917 3860 28987 3906
rect 29033 3860 29103 3906
rect 29149 3860 29219 3906
rect 29265 3860 29335 3906
rect 29381 3860 29451 3906
rect 29497 3860 29567 3906
rect 29613 3860 29683 3906
rect 29729 3860 29799 3906
rect 29845 3860 29915 3906
rect 29961 3860 30031 3906
rect 30077 3860 30147 3906
rect 30193 3860 30263 3906
rect 30309 3860 30379 3906
rect 30425 3860 30495 3906
rect 30541 3860 30611 3906
rect 30657 3860 30727 3906
rect 30773 3860 30843 3906
rect 30889 3860 30959 3906
rect 31005 3860 31075 3906
rect 31121 3860 31191 3906
rect 31237 3860 31307 3906
rect 31353 3860 31423 3906
rect 31469 3860 31539 3906
rect 31585 3860 31655 3906
rect 31701 3860 31771 3906
rect 31817 3860 31887 3906
rect 31933 3860 32003 3906
rect 32049 3860 32119 3906
rect 32165 3860 32235 3906
rect 32281 3860 32351 3906
rect 32397 3860 32467 3906
rect 32513 3860 32583 3906
rect 32629 3860 32699 3906
rect 32745 3860 32815 3906
rect 32861 3860 32931 3906
rect 32977 3860 33047 3906
rect 33093 3860 33163 3906
rect 33209 3860 33279 3906
rect 33325 3860 33395 3906
rect 33441 3860 33511 3906
rect 33557 3860 33627 3906
rect 33673 3860 33743 3906
rect 33789 3860 33859 3906
rect 33905 3860 33975 3906
rect 34021 3860 34091 3906
rect 34137 3860 34207 3906
rect 34253 3860 34323 3906
rect 34369 3860 34439 3906
rect 34485 3860 34555 3906
rect 34601 3860 34671 3906
rect 34717 3860 34787 3906
rect 34833 3860 34903 3906
rect 34949 3860 35019 3906
rect 35065 3860 35135 3906
rect 35181 3860 35251 3906
rect 35297 3860 35367 3906
rect 35413 3860 35483 3906
rect 35529 3860 35599 3906
rect 35645 3860 35715 3906
rect 35761 3860 35831 3906
rect 35877 3860 35947 3906
rect 35993 3860 36063 3906
rect 36109 3860 36179 3906
rect 36225 3860 36295 3906
rect 36341 3860 36411 3906
rect 36457 3860 36527 3906
rect 36573 3860 36643 3906
rect 36689 3860 36759 3906
rect 36805 3860 36875 3906
rect 36921 3860 36991 3906
rect 37037 3860 37107 3906
rect 37153 3860 37223 3906
rect 37269 3860 37339 3906
rect 37385 3860 37455 3906
rect 37501 3860 37571 3906
rect 37617 3860 37687 3906
rect 37733 3860 37803 3906
rect 37849 3860 37919 3906
rect 37965 3860 38035 3906
rect 38081 3860 38151 3906
rect 38197 3860 38267 3906
rect 38313 3860 38383 3906
rect 38429 3860 38499 3906
rect 38545 3860 38615 3906
rect 38661 3860 38731 3906
rect 38777 3860 38847 3906
rect 38893 3860 38963 3906
rect 39009 3860 39079 3906
rect 39125 3860 39195 3906
rect 39241 3860 39311 3906
rect 39357 3860 39427 3906
rect 39473 3860 39543 3906
rect 39589 3860 39659 3906
rect 39705 3860 39775 3906
rect 39821 3860 39891 3906
rect 39937 3860 40007 3906
rect 40053 3860 40123 3906
rect 40169 3860 40180 3906
rect 28628 3790 40180 3860
rect 28628 3744 28639 3790
rect 28685 3744 28755 3790
rect 28801 3744 28871 3790
rect 28917 3744 28987 3790
rect 29033 3744 29103 3790
rect 29149 3744 29219 3790
rect 29265 3744 29335 3790
rect 29381 3744 29451 3790
rect 29497 3744 29567 3790
rect 29613 3744 29683 3790
rect 29729 3744 29799 3790
rect 29845 3744 29915 3790
rect 29961 3744 30031 3790
rect 30077 3744 30147 3790
rect 30193 3744 30263 3790
rect 30309 3744 30379 3790
rect 30425 3744 30495 3790
rect 30541 3744 30611 3790
rect 30657 3744 30727 3790
rect 30773 3744 30843 3790
rect 30889 3744 30959 3790
rect 31005 3744 31075 3790
rect 31121 3744 31191 3790
rect 31237 3744 31307 3790
rect 31353 3744 31423 3790
rect 31469 3744 31539 3790
rect 31585 3744 31655 3790
rect 31701 3744 31771 3790
rect 31817 3744 31887 3790
rect 31933 3744 32003 3790
rect 32049 3744 32119 3790
rect 32165 3744 32235 3790
rect 32281 3744 32351 3790
rect 32397 3744 32467 3790
rect 32513 3744 32583 3790
rect 32629 3744 32699 3790
rect 32745 3744 32815 3790
rect 32861 3744 32931 3790
rect 32977 3744 33047 3790
rect 33093 3744 33163 3790
rect 33209 3744 33279 3790
rect 33325 3744 33395 3790
rect 33441 3744 33511 3790
rect 33557 3744 33627 3790
rect 33673 3744 33743 3790
rect 33789 3744 33859 3790
rect 33905 3744 33975 3790
rect 34021 3744 34091 3790
rect 34137 3744 34207 3790
rect 34253 3744 34323 3790
rect 34369 3744 34439 3790
rect 34485 3744 34555 3790
rect 34601 3744 34671 3790
rect 34717 3744 34787 3790
rect 34833 3744 34903 3790
rect 34949 3744 35019 3790
rect 35065 3744 35135 3790
rect 35181 3744 35251 3790
rect 35297 3744 35367 3790
rect 35413 3744 35483 3790
rect 35529 3744 35599 3790
rect 35645 3744 35715 3790
rect 35761 3744 35831 3790
rect 35877 3744 35947 3790
rect 35993 3744 36063 3790
rect 36109 3744 36179 3790
rect 36225 3744 36295 3790
rect 36341 3744 36411 3790
rect 36457 3744 36527 3790
rect 36573 3744 36643 3790
rect 36689 3744 36759 3790
rect 36805 3744 36875 3790
rect 36921 3744 36991 3790
rect 37037 3744 37107 3790
rect 37153 3744 37223 3790
rect 37269 3744 37339 3790
rect 37385 3744 37455 3790
rect 37501 3744 37571 3790
rect 37617 3744 37687 3790
rect 37733 3744 37803 3790
rect 37849 3744 37919 3790
rect 37965 3744 38035 3790
rect 38081 3744 38151 3790
rect 38197 3744 38267 3790
rect 38313 3744 38383 3790
rect 38429 3744 38499 3790
rect 38545 3744 38615 3790
rect 38661 3744 38731 3790
rect 38777 3744 38847 3790
rect 38893 3744 38963 3790
rect 39009 3744 39079 3790
rect 39125 3744 39195 3790
rect 39241 3744 39311 3790
rect 39357 3744 39427 3790
rect 39473 3744 39543 3790
rect 39589 3744 39659 3790
rect 39705 3744 39775 3790
rect 39821 3744 39891 3790
rect 39937 3744 40007 3790
rect 40053 3744 40123 3790
rect 40169 3744 40180 3790
rect 28628 3674 40180 3744
rect 28628 3628 28639 3674
rect 28685 3628 28755 3674
rect 28801 3628 28871 3674
rect 28917 3628 28987 3674
rect 29033 3628 29103 3674
rect 29149 3628 29219 3674
rect 29265 3628 29335 3674
rect 29381 3628 29451 3674
rect 29497 3628 29567 3674
rect 29613 3628 29683 3674
rect 29729 3628 29799 3674
rect 29845 3628 29915 3674
rect 29961 3628 30031 3674
rect 30077 3628 30147 3674
rect 30193 3628 30263 3674
rect 30309 3628 30379 3674
rect 30425 3628 30495 3674
rect 30541 3628 30611 3674
rect 30657 3628 30727 3674
rect 30773 3628 30843 3674
rect 30889 3628 30959 3674
rect 31005 3628 31075 3674
rect 31121 3628 31191 3674
rect 31237 3628 31307 3674
rect 31353 3628 31423 3674
rect 31469 3628 31539 3674
rect 31585 3628 31655 3674
rect 31701 3628 31771 3674
rect 31817 3628 31887 3674
rect 31933 3628 32003 3674
rect 32049 3628 32119 3674
rect 32165 3628 32235 3674
rect 32281 3628 32351 3674
rect 32397 3628 32467 3674
rect 32513 3628 32583 3674
rect 32629 3628 32699 3674
rect 32745 3628 32815 3674
rect 32861 3628 32931 3674
rect 32977 3628 33047 3674
rect 33093 3628 33163 3674
rect 33209 3628 33279 3674
rect 33325 3628 33395 3674
rect 33441 3628 33511 3674
rect 33557 3628 33627 3674
rect 33673 3628 33743 3674
rect 33789 3628 33859 3674
rect 33905 3628 33975 3674
rect 34021 3628 34091 3674
rect 34137 3628 34207 3674
rect 34253 3628 34323 3674
rect 34369 3628 34439 3674
rect 34485 3628 34555 3674
rect 34601 3628 34671 3674
rect 34717 3628 34787 3674
rect 34833 3628 34903 3674
rect 34949 3628 35019 3674
rect 35065 3628 35135 3674
rect 35181 3628 35251 3674
rect 35297 3628 35367 3674
rect 35413 3628 35483 3674
rect 35529 3628 35599 3674
rect 35645 3628 35715 3674
rect 35761 3628 35831 3674
rect 35877 3628 35947 3674
rect 35993 3628 36063 3674
rect 36109 3628 36179 3674
rect 36225 3628 36295 3674
rect 36341 3628 36411 3674
rect 36457 3628 36527 3674
rect 36573 3628 36643 3674
rect 36689 3628 36759 3674
rect 36805 3628 36875 3674
rect 36921 3628 36991 3674
rect 37037 3628 37107 3674
rect 37153 3628 37223 3674
rect 37269 3628 37339 3674
rect 37385 3628 37455 3674
rect 37501 3628 37571 3674
rect 37617 3628 37687 3674
rect 37733 3628 37803 3674
rect 37849 3628 37919 3674
rect 37965 3628 38035 3674
rect 38081 3628 38151 3674
rect 38197 3628 38267 3674
rect 38313 3628 38383 3674
rect 38429 3628 38499 3674
rect 38545 3628 38615 3674
rect 38661 3628 38731 3674
rect 38777 3628 38847 3674
rect 38893 3628 38963 3674
rect 39009 3628 39079 3674
rect 39125 3628 39195 3674
rect 39241 3628 39311 3674
rect 39357 3628 39427 3674
rect 39473 3628 39543 3674
rect 39589 3628 39659 3674
rect 39705 3628 39775 3674
rect 39821 3628 39891 3674
rect 39937 3628 40007 3674
rect 40053 3628 40123 3674
rect 40169 3628 40180 3674
rect 28628 3558 40180 3628
rect 28628 3512 28639 3558
rect 28685 3512 28755 3558
rect 28801 3512 28871 3558
rect 28917 3512 28987 3558
rect 29033 3512 29103 3558
rect 29149 3512 29219 3558
rect 29265 3512 29335 3558
rect 29381 3512 29451 3558
rect 29497 3512 29567 3558
rect 29613 3512 29683 3558
rect 29729 3512 29799 3558
rect 29845 3512 29915 3558
rect 29961 3512 30031 3558
rect 30077 3512 30147 3558
rect 30193 3512 30263 3558
rect 30309 3512 30379 3558
rect 30425 3512 30495 3558
rect 30541 3512 30611 3558
rect 30657 3512 30727 3558
rect 30773 3512 30843 3558
rect 30889 3512 30959 3558
rect 31005 3512 31075 3558
rect 31121 3512 31191 3558
rect 31237 3512 31307 3558
rect 31353 3512 31423 3558
rect 31469 3512 31539 3558
rect 31585 3512 31655 3558
rect 31701 3512 31771 3558
rect 31817 3512 31887 3558
rect 31933 3512 32003 3558
rect 32049 3512 32119 3558
rect 32165 3512 32235 3558
rect 32281 3512 32351 3558
rect 32397 3512 32467 3558
rect 32513 3512 32583 3558
rect 32629 3512 32699 3558
rect 32745 3512 32815 3558
rect 32861 3512 32931 3558
rect 32977 3512 33047 3558
rect 33093 3512 33163 3558
rect 33209 3512 33279 3558
rect 33325 3512 33395 3558
rect 33441 3512 33511 3558
rect 33557 3512 33627 3558
rect 33673 3512 33743 3558
rect 33789 3512 33859 3558
rect 33905 3512 33975 3558
rect 34021 3512 34091 3558
rect 34137 3512 34207 3558
rect 34253 3512 34323 3558
rect 34369 3512 34439 3558
rect 34485 3512 34555 3558
rect 34601 3512 34671 3558
rect 34717 3512 34787 3558
rect 34833 3512 34903 3558
rect 34949 3512 35019 3558
rect 35065 3512 35135 3558
rect 35181 3512 35251 3558
rect 35297 3512 35367 3558
rect 35413 3512 35483 3558
rect 35529 3512 35599 3558
rect 35645 3512 35715 3558
rect 35761 3512 35831 3558
rect 35877 3512 35947 3558
rect 35993 3512 36063 3558
rect 36109 3512 36179 3558
rect 36225 3512 36295 3558
rect 36341 3512 36411 3558
rect 36457 3512 36527 3558
rect 36573 3512 36643 3558
rect 36689 3512 36759 3558
rect 36805 3512 36875 3558
rect 36921 3512 36991 3558
rect 37037 3512 37107 3558
rect 37153 3512 37223 3558
rect 37269 3512 37339 3558
rect 37385 3512 37455 3558
rect 37501 3512 37571 3558
rect 37617 3512 37687 3558
rect 37733 3512 37803 3558
rect 37849 3512 37919 3558
rect 37965 3512 38035 3558
rect 38081 3512 38151 3558
rect 38197 3512 38267 3558
rect 38313 3512 38383 3558
rect 38429 3512 38499 3558
rect 38545 3512 38615 3558
rect 38661 3512 38731 3558
rect 38777 3512 38847 3558
rect 38893 3512 38963 3558
rect 39009 3512 39079 3558
rect 39125 3512 39195 3558
rect 39241 3512 39311 3558
rect 39357 3512 39427 3558
rect 39473 3512 39543 3558
rect 39589 3512 39659 3558
rect 39705 3512 39775 3558
rect 39821 3512 39891 3558
rect 39937 3512 40007 3558
rect 40053 3512 40123 3558
rect 40169 3512 40180 3558
rect 28628 3442 40180 3512
rect 28628 3396 28639 3442
rect 28685 3396 28755 3442
rect 28801 3396 28871 3442
rect 28917 3396 28987 3442
rect 29033 3396 29103 3442
rect 29149 3396 29219 3442
rect 29265 3396 29335 3442
rect 29381 3396 29451 3442
rect 29497 3396 29567 3442
rect 29613 3396 29683 3442
rect 29729 3396 29799 3442
rect 29845 3396 29915 3442
rect 29961 3396 30031 3442
rect 30077 3396 30147 3442
rect 30193 3396 30263 3442
rect 30309 3396 30379 3442
rect 30425 3396 30495 3442
rect 30541 3396 30611 3442
rect 30657 3396 30727 3442
rect 30773 3396 30843 3442
rect 30889 3396 30959 3442
rect 31005 3396 31075 3442
rect 31121 3396 31191 3442
rect 31237 3396 31307 3442
rect 31353 3396 31423 3442
rect 31469 3396 31539 3442
rect 31585 3396 31655 3442
rect 31701 3396 31771 3442
rect 31817 3396 31887 3442
rect 31933 3396 32003 3442
rect 32049 3396 32119 3442
rect 32165 3396 32235 3442
rect 32281 3396 32351 3442
rect 32397 3396 32467 3442
rect 32513 3396 32583 3442
rect 32629 3396 32699 3442
rect 32745 3396 32815 3442
rect 32861 3396 32931 3442
rect 32977 3396 33047 3442
rect 33093 3396 33163 3442
rect 33209 3396 33279 3442
rect 33325 3396 33395 3442
rect 33441 3396 33511 3442
rect 33557 3396 33627 3442
rect 33673 3396 33743 3442
rect 33789 3396 33859 3442
rect 33905 3396 33975 3442
rect 34021 3396 34091 3442
rect 34137 3396 34207 3442
rect 34253 3396 34323 3442
rect 34369 3396 34439 3442
rect 34485 3396 34555 3442
rect 34601 3396 34671 3442
rect 34717 3396 34787 3442
rect 34833 3396 34903 3442
rect 34949 3396 35019 3442
rect 35065 3396 35135 3442
rect 35181 3396 35251 3442
rect 35297 3396 35367 3442
rect 35413 3396 35483 3442
rect 35529 3396 35599 3442
rect 35645 3396 35715 3442
rect 35761 3396 35831 3442
rect 35877 3396 35947 3442
rect 35993 3396 36063 3442
rect 36109 3396 36179 3442
rect 36225 3396 36295 3442
rect 36341 3396 36411 3442
rect 36457 3396 36527 3442
rect 36573 3396 36643 3442
rect 36689 3396 36759 3442
rect 36805 3396 36875 3442
rect 36921 3396 36991 3442
rect 37037 3396 37107 3442
rect 37153 3396 37223 3442
rect 37269 3396 37339 3442
rect 37385 3396 37455 3442
rect 37501 3396 37571 3442
rect 37617 3396 37687 3442
rect 37733 3396 37803 3442
rect 37849 3396 37919 3442
rect 37965 3396 38035 3442
rect 38081 3396 38151 3442
rect 38197 3396 38267 3442
rect 38313 3396 38383 3442
rect 38429 3396 38499 3442
rect 38545 3396 38615 3442
rect 38661 3396 38731 3442
rect 38777 3396 38847 3442
rect 38893 3396 38963 3442
rect 39009 3396 39079 3442
rect 39125 3396 39195 3442
rect 39241 3396 39311 3442
rect 39357 3396 39427 3442
rect 39473 3396 39543 3442
rect 39589 3396 39659 3442
rect 39705 3396 39775 3442
rect 39821 3396 39891 3442
rect 39937 3396 40007 3442
rect 40053 3396 40123 3442
rect 40169 3396 40180 3442
rect 28628 3326 40180 3396
rect 28628 3280 28639 3326
rect 28685 3280 28755 3326
rect 28801 3280 28871 3326
rect 28917 3280 28987 3326
rect 29033 3280 29103 3326
rect 29149 3280 29219 3326
rect 29265 3280 29335 3326
rect 29381 3280 29451 3326
rect 29497 3280 29567 3326
rect 29613 3280 29683 3326
rect 29729 3280 29799 3326
rect 29845 3280 29915 3326
rect 29961 3280 30031 3326
rect 30077 3280 30147 3326
rect 30193 3280 30263 3326
rect 30309 3280 30379 3326
rect 30425 3280 30495 3326
rect 30541 3280 30611 3326
rect 30657 3280 30727 3326
rect 30773 3280 30843 3326
rect 30889 3280 30959 3326
rect 31005 3280 31075 3326
rect 31121 3280 31191 3326
rect 31237 3280 31307 3326
rect 31353 3280 31423 3326
rect 31469 3280 31539 3326
rect 31585 3280 31655 3326
rect 31701 3280 31771 3326
rect 31817 3280 31887 3326
rect 31933 3280 32003 3326
rect 32049 3280 32119 3326
rect 32165 3280 32235 3326
rect 32281 3280 32351 3326
rect 32397 3280 32467 3326
rect 32513 3280 32583 3326
rect 32629 3280 32699 3326
rect 32745 3280 32815 3326
rect 32861 3280 32931 3326
rect 32977 3280 33047 3326
rect 33093 3280 33163 3326
rect 33209 3280 33279 3326
rect 33325 3280 33395 3326
rect 33441 3280 33511 3326
rect 33557 3280 33627 3326
rect 33673 3280 33743 3326
rect 33789 3280 33859 3326
rect 33905 3280 33975 3326
rect 34021 3280 34091 3326
rect 34137 3280 34207 3326
rect 34253 3280 34323 3326
rect 34369 3280 34439 3326
rect 34485 3280 34555 3326
rect 34601 3280 34671 3326
rect 34717 3280 34787 3326
rect 34833 3280 34903 3326
rect 34949 3280 35019 3326
rect 35065 3280 35135 3326
rect 35181 3280 35251 3326
rect 35297 3280 35367 3326
rect 35413 3280 35483 3326
rect 35529 3280 35599 3326
rect 35645 3280 35715 3326
rect 35761 3280 35831 3326
rect 35877 3280 35947 3326
rect 35993 3280 36063 3326
rect 36109 3280 36179 3326
rect 36225 3280 36295 3326
rect 36341 3280 36411 3326
rect 36457 3280 36527 3326
rect 36573 3280 36643 3326
rect 36689 3280 36759 3326
rect 36805 3280 36875 3326
rect 36921 3280 36991 3326
rect 37037 3280 37107 3326
rect 37153 3280 37223 3326
rect 37269 3280 37339 3326
rect 37385 3280 37455 3326
rect 37501 3280 37571 3326
rect 37617 3280 37687 3326
rect 37733 3280 37803 3326
rect 37849 3280 37919 3326
rect 37965 3280 38035 3326
rect 38081 3280 38151 3326
rect 38197 3280 38267 3326
rect 38313 3280 38383 3326
rect 38429 3280 38499 3326
rect 38545 3280 38615 3326
rect 38661 3280 38731 3326
rect 38777 3280 38847 3326
rect 38893 3280 38963 3326
rect 39009 3280 39079 3326
rect 39125 3280 39195 3326
rect 39241 3280 39311 3326
rect 39357 3280 39427 3326
rect 39473 3280 39543 3326
rect 39589 3280 39659 3326
rect 39705 3280 39775 3326
rect 39821 3280 39891 3326
rect 39937 3280 40007 3326
rect 40053 3280 40123 3326
rect 40169 3280 40180 3326
rect 50834 3906 56586 3917
rect 50834 3860 50845 3906
rect 50891 3860 50961 3906
rect 51007 3860 51077 3906
rect 51123 3860 51193 3906
rect 51239 3860 51309 3906
rect 51355 3860 51425 3906
rect 51471 3860 51541 3906
rect 51587 3860 51657 3906
rect 51703 3860 51773 3906
rect 51819 3860 51889 3906
rect 51935 3860 52005 3906
rect 52051 3860 52121 3906
rect 52167 3860 52237 3906
rect 52283 3860 52353 3906
rect 52399 3860 52469 3906
rect 52515 3860 52585 3906
rect 52631 3860 52701 3906
rect 52747 3860 52817 3906
rect 52863 3860 52933 3906
rect 52979 3860 53049 3906
rect 53095 3860 53165 3906
rect 53211 3860 53281 3906
rect 53327 3860 53397 3906
rect 53443 3860 53513 3906
rect 53559 3860 53629 3906
rect 53675 3860 53745 3906
rect 53791 3860 53861 3906
rect 53907 3860 53977 3906
rect 54023 3860 54093 3906
rect 54139 3860 54209 3906
rect 54255 3860 54325 3906
rect 54371 3860 54441 3906
rect 54487 3860 54557 3906
rect 54603 3860 54673 3906
rect 54719 3860 54789 3906
rect 54835 3860 54905 3906
rect 54951 3860 55021 3906
rect 55067 3860 55137 3906
rect 55183 3860 55253 3906
rect 55299 3860 55369 3906
rect 55415 3860 55485 3906
rect 55531 3860 55601 3906
rect 55647 3860 55717 3906
rect 55763 3860 55833 3906
rect 55879 3860 55949 3906
rect 55995 3860 56065 3906
rect 56111 3860 56181 3906
rect 56227 3860 56297 3906
rect 56343 3860 56413 3906
rect 56459 3860 56529 3906
rect 56575 3860 56586 3906
rect 50834 3790 56586 3860
rect 50834 3744 50845 3790
rect 50891 3744 50961 3790
rect 51007 3744 51077 3790
rect 51123 3744 51193 3790
rect 51239 3744 51309 3790
rect 51355 3744 51425 3790
rect 51471 3744 51541 3790
rect 51587 3744 51657 3790
rect 51703 3744 51773 3790
rect 51819 3744 51889 3790
rect 51935 3744 52005 3790
rect 52051 3744 52121 3790
rect 52167 3744 52237 3790
rect 52283 3744 52353 3790
rect 52399 3744 52469 3790
rect 52515 3744 52585 3790
rect 52631 3744 52701 3790
rect 52747 3744 52817 3790
rect 52863 3744 52933 3790
rect 52979 3744 53049 3790
rect 53095 3744 53165 3790
rect 53211 3744 53281 3790
rect 53327 3744 53397 3790
rect 53443 3744 53513 3790
rect 53559 3744 53629 3790
rect 53675 3744 53745 3790
rect 53791 3744 53861 3790
rect 53907 3744 53977 3790
rect 54023 3744 54093 3790
rect 54139 3744 54209 3790
rect 54255 3744 54325 3790
rect 54371 3744 54441 3790
rect 54487 3744 54557 3790
rect 54603 3744 54673 3790
rect 54719 3744 54789 3790
rect 54835 3744 54905 3790
rect 54951 3744 55021 3790
rect 55067 3744 55137 3790
rect 55183 3744 55253 3790
rect 55299 3744 55369 3790
rect 55415 3744 55485 3790
rect 55531 3744 55601 3790
rect 55647 3744 55717 3790
rect 55763 3744 55833 3790
rect 55879 3744 55949 3790
rect 55995 3744 56065 3790
rect 56111 3744 56181 3790
rect 56227 3744 56297 3790
rect 56343 3744 56413 3790
rect 56459 3744 56529 3790
rect 56575 3744 56586 3790
rect 50834 3674 56586 3744
rect 50834 3628 50845 3674
rect 50891 3628 50961 3674
rect 51007 3628 51077 3674
rect 51123 3628 51193 3674
rect 51239 3628 51309 3674
rect 51355 3628 51425 3674
rect 51471 3628 51541 3674
rect 51587 3628 51657 3674
rect 51703 3628 51773 3674
rect 51819 3628 51889 3674
rect 51935 3628 52005 3674
rect 52051 3628 52121 3674
rect 52167 3628 52237 3674
rect 52283 3628 52353 3674
rect 52399 3628 52469 3674
rect 52515 3628 52585 3674
rect 52631 3628 52701 3674
rect 52747 3628 52817 3674
rect 52863 3628 52933 3674
rect 52979 3628 53049 3674
rect 53095 3628 53165 3674
rect 53211 3628 53281 3674
rect 53327 3628 53397 3674
rect 53443 3628 53513 3674
rect 53559 3628 53629 3674
rect 53675 3628 53745 3674
rect 53791 3628 53861 3674
rect 53907 3628 53977 3674
rect 54023 3628 54093 3674
rect 54139 3628 54209 3674
rect 54255 3628 54325 3674
rect 54371 3628 54441 3674
rect 54487 3628 54557 3674
rect 54603 3628 54673 3674
rect 54719 3628 54789 3674
rect 54835 3628 54905 3674
rect 54951 3628 55021 3674
rect 55067 3628 55137 3674
rect 55183 3628 55253 3674
rect 55299 3628 55369 3674
rect 55415 3628 55485 3674
rect 55531 3628 55601 3674
rect 55647 3628 55717 3674
rect 55763 3628 55833 3674
rect 55879 3628 55949 3674
rect 55995 3628 56065 3674
rect 56111 3628 56181 3674
rect 56227 3628 56297 3674
rect 56343 3628 56413 3674
rect 56459 3628 56529 3674
rect 56575 3628 56586 3674
rect 50834 3558 56586 3628
rect 50834 3512 50845 3558
rect 50891 3512 50961 3558
rect 51007 3512 51077 3558
rect 51123 3512 51193 3558
rect 51239 3512 51309 3558
rect 51355 3512 51425 3558
rect 51471 3512 51541 3558
rect 51587 3512 51657 3558
rect 51703 3512 51773 3558
rect 51819 3512 51889 3558
rect 51935 3512 52005 3558
rect 52051 3512 52121 3558
rect 52167 3512 52237 3558
rect 52283 3512 52353 3558
rect 52399 3512 52469 3558
rect 52515 3512 52585 3558
rect 52631 3512 52701 3558
rect 52747 3512 52817 3558
rect 52863 3512 52933 3558
rect 52979 3512 53049 3558
rect 53095 3512 53165 3558
rect 53211 3512 53281 3558
rect 53327 3512 53397 3558
rect 53443 3512 53513 3558
rect 53559 3512 53629 3558
rect 53675 3512 53745 3558
rect 53791 3512 53861 3558
rect 53907 3512 53977 3558
rect 54023 3512 54093 3558
rect 54139 3512 54209 3558
rect 54255 3512 54325 3558
rect 54371 3512 54441 3558
rect 54487 3512 54557 3558
rect 54603 3512 54673 3558
rect 54719 3512 54789 3558
rect 54835 3512 54905 3558
rect 54951 3512 55021 3558
rect 55067 3512 55137 3558
rect 55183 3512 55253 3558
rect 55299 3512 55369 3558
rect 55415 3512 55485 3558
rect 55531 3512 55601 3558
rect 55647 3512 55717 3558
rect 55763 3512 55833 3558
rect 55879 3512 55949 3558
rect 55995 3512 56065 3558
rect 56111 3512 56181 3558
rect 56227 3512 56297 3558
rect 56343 3512 56413 3558
rect 56459 3512 56529 3558
rect 56575 3512 56586 3558
rect 50834 3442 56586 3512
rect 50834 3396 50845 3442
rect 50891 3396 50961 3442
rect 51007 3396 51077 3442
rect 51123 3396 51193 3442
rect 51239 3396 51309 3442
rect 51355 3396 51425 3442
rect 51471 3396 51541 3442
rect 51587 3396 51657 3442
rect 51703 3396 51773 3442
rect 51819 3396 51889 3442
rect 51935 3396 52005 3442
rect 52051 3396 52121 3442
rect 52167 3396 52237 3442
rect 52283 3396 52353 3442
rect 52399 3396 52469 3442
rect 52515 3396 52585 3442
rect 52631 3396 52701 3442
rect 52747 3396 52817 3442
rect 52863 3396 52933 3442
rect 52979 3396 53049 3442
rect 53095 3396 53165 3442
rect 53211 3396 53281 3442
rect 53327 3396 53397 3442
rect 53443 3396 53513 3442
rect 53559 3396 53629 3442
rect 53675 3396 53745 3442
rect 53791 3396 53861 3442
rect 53907 3396 53977 3442
rect 54023 3396 54093 3442
rect 54139 3396 54209 3442
rect 54255 3396 54325 3442
rect 54371 3396 54441 3442
rect 54487 3396 54557 3442
rect 54603 3396 54673 3442
rect 54719 3396 54789 3442
rect 54835 3396 54905 3442
rect 54951 3396 55021 3442
rect 55067 3396 55137 3442
rect 55183 3396 55253 3442
rect 55299 3396 55369 3442
rect 55415 3396 55485 3442
rect 55531 3396 55601 3442
rect 55647 3396 55717 3442
rect 55763 3396 55833 3442
rect 55879 3396 55949 3442
rect 55995 3396 56065 3442
rect 56111 3396 56181 3442
rect 56227 3396 56297 3442
rect 56343 3396 56413 3442
rect 56459 3396 56529 3442
rect 56575 3396 56586 3442
rect 50834 3326 56586 3396
rect 28628 3210 40180 3280
rect 40611 3282 40791 3294
rect 40611 3230 40623 3282
rect 40779 3230 40791 3282
rect 40611 3218 40791 3230
rect 50834 3280 50845 3326
rect 50891 3280 50961 3326
rect 51007 3280 51077 3326
rect 51123 3280 51193 3326
rect 51239 3280 51309 3326
rect 51355 3280 51425 3326
rect 51471 3280 51541 3326
rect 51587 3280 51657 3326
rect 51703 3280 51773 3326
rect 51819 3280 51889 3326
rect 51935 3280 52005 3326
rect 52051 3280 52121 3326
rect 52167 3280 52237 3326
rect 52283 3280 52353 3326
rect 52399 3280 52469 3326
rect 52515 3280 52585 3326
rect 52631 3280 52701 3326
rect 52747 3280 52817 3326
rect 52863 3280 52933 3326
rect 52979 3280 53049 3326
rect 53095 3280 53165 3326
rect 53211 3280 53281 3326
rect 53327 3280 53397 3326
rect 53443 3280 53513 3326
rect 53559 3280 53629 3326
rect 53675 3280 53745 3326
rect 53791 3280 53861 3326
rect 53907 3280 53977 3326
rect 54023 3280 54093 3326
rect 54139 3280 54209 3326
rect 54255 3280 54325 3326
rect 54371 3280 54441 3326
rect 54487 3280 54557 3326
rect 54603 3280 54673 3326
rect 54719 3280 54789 3326
rect 54835 3280 54905 3326
rect 54951 3280 55021 3326
rect 55067 3280 55137 3326
rect 55183 3280 55253 3326
rect 55299 3280 55369 3326
rect 55415 3280 55485 3326
rect 55531 3280 55601 3326
rect 55647 3280 55717 3326
rect 55763 3280 55833 3326
rect 55879 3280 55949 3326
rect 55995 3280 56065 3326
rect 56111 3280 56181 3326
rect 56227 3280 56297 3326
rect 56343 3280 56413 3326
rect 56459 3280 56529 3326
rect 56575 3280 56586 3326
rect 28628 3164 28639 3210
rect 28685 3164 28755 3210
rect 28801 3164 28871 3210
rect 28917 3164 28987 3210
rect 29033 3164 29103 3210
rect 29149 3164 29219 3210
rect 29265 3164 29335 3210
rect 29381 3164 29451 3210
rect 29497 3164 29567 3210
rect 29613 3164 29683 3210
rect 29729 3164 29799 3210
rect 29845 3164 29915 3210
rect 29961 3164 30031 3210
rect 30077 3164 30147 3210
rect 30193 3164 30263 3210
rect 30309 3164 30379 3210
rect 30425 3164 30495 3210
rect 30541 3164 30611 3210
rect 30657 3164 30727 3210
rect 30773 3164 30843 3210
rect 30889 3164 30959 3210
rect 31005 3164 31075 3210
rect 31121 3164 31191 3210
rect 31237 3164 31307 3210
rect 31353 3164 31423 3210
rect 31469 3164 31539 3210
rect 31585 3164 31655 3210
rect 31701 3164 31771 3210
rect 31817 3164 31887 3210
rect 31933 3164 32003 3210
rect 32049 3164 32119 3210
rect 32165 3164 32235 3210
rect 32281 3164 32351 3210
rect 32397 3164 32467 3210
rect 32513 3164 32583 3210
rect 32629 3164 32699 3210
rect 32745 3164 32815 3210
rect 32861 3164 32931 3210
rect 32977 3164 33047 3210
rect 33093 3164 33163 3210
rect 33209 3164 33279 3210
rect 33325 3164 33395 3210
rect 33441 3164 33511 3210
rect 33557 3164 33627 3210
rect 33673 3164 33743 3210
rect 33789 3164 33859 3210
rect 33905 3164 33975 3210
rect 34021 3164 34091 3210
rect 34137 3164 34207 3210
rect 34253 3164 34323 3210
rect 34369 3164 34439 3210
rect 34485 3164 34555 3210
rect 34601 3164 34671 3210
rect 34717 3164 34787 3210
rect 34833 3164 34903 3210
rect 34949 3164 35019 3210
rect 35065 3164 35135 3210
rect 35181 3164 35251 3210
rect 35297 3164 35367 3210
rect 35413 3164 35483 3210
rect 35529 3164 35599 3210
rect 35645 3164 35715 3210
rect 35761 3164 35831 3210
rect 35877 3164 35947 3210
rect 35993 3164 36063 3210
rect 36109 3164 36179 3210
rect 36225 3164 36295 3210
rect 36341 3164 36411 3210
rect 36457 3164 36527 3210
rect 36573 3164 36643 3210
rect 36689 3164 36759 3210
rect 36805 3164 36875 3210
rect 36921 3164 36991 3210
rect 37037 3164 37107 3210
rect 37153 3164 37223 3210
rect 37269 3164 37339 3210
rect 37385 3164 37455 3210
rect 37501 3164 37571 3210
rect 37617 3164 37687 3210
rect 37733 3164 37803 3210
rect 37849 3164 37919 3210
rect 37965 3164 38035 3210
rect 38081 3164 38151 3210
rect 38197 3164 38267 3210
rect 38313 3164 38383 3210
rect 38429 3164 38499 3210
rect 38545 3164 38615 3210
rect 38661 3164 38731 3210
rect 38777 3164 38847 3210
rect 38893 3164 38963 3210
rect 39009 3164 39079 3210
rect 39125 3164 39195 3210
rect 39241 3164 39311 3210
rect 39357 3164 39427 3210
rect 39473 3164 39543 3210
rect 39589 3164 39659 3210
rect 39705 3164 39775 3210
rect 39821 3164 39891 3210
rect 39937 3164 40007 3210
rect 40053 3164 40123 3210
rect 40169 3164 40180 3210
rect 28628 3094 40180 3164
rect 28628 3048 28639 3094
rect 28685 3048 28755 3094
rect 28801 3048 28871 3094
rect 28917 3048 28987 3094
rect 29033 3048 29103 3094
rect 29149 3048 29219 3094
rect 29265 3048 29335 3094
rect 29381 3048 29451 3094
rect 29497 3048 29567 3094
rect 29613 3048 29683 3094
rect 29729 3048 29799 3094
rect 29845 3048 29915 3094
rect 29961 3048 30031 3094
rect 30077 3048 30147 3094
rect 30193 3048 30263 3094
rect 30309 3048 30379 3094
rect 30425 3048 30495 3094
rect 30541 3048 30611 3094
rect 30657 3048 30727 3094
rect 30773 3048 30843 3094
rect 30889 3048 30959 3094
rect 31005 3048 31075 3094
rect 31121 3048 31191 3094
rect 31237 3048 31307 3094
rect 31353 3048 31423 3094
rect 31469 3048 31539 3094
rect 31585 3048 31655 3094
rect 31701 3048 31771 3094
rect 31817 3048 31887 3094
rect 31933 3048 32003 3094
rect 32049 3048 32119 3094
rect 32165 3048 32235 3094
rect 32281 3048 32351 3094
rect 32397 3048 32467 3094
rect 32513 3048 32583 3094
rect 32629 3048 32699 3094
rect 32745 3048 32815 3094
rect 32861 3048 32931 3094
rect 32977 3048 33047 3094
rect 33093 3048 33163 3094
rect 33209 3048 33279 3094
rect 33325 3048 33395 3094
rect 33441 3048 33511 3094
rect 33557 3048 33627 3094
rect 33673 3048 33743 3094
rect 33789 3048 33859 3094
rect 33905 3048 33975 3094
rect 34021 3048 34091 3094
rect 34137 3048 34207 3094
rect 34253 3048 34323 3094
rect 34369 3048 34439 3094
rect 34485 3048 34555 3094
rect 34601 3048 34671 3094
rect 34717 3048 34787 3094
rect 34833 3048 34903 3094
rect 34949 3048 35019 3094
rect 35065 3048 35135 3094
rect 35181 3048 35251 3094
rect 35297 3048 35367 3094
rect 35413 3048 35483 3094
rect 35529 3048 35599 3094
rect 35645 3048 35715 3094
rect 35761 3048 35831 3094
rect 35877 3048 35947 3094
rect 35993 3048 36063 3094
rect 36109 3048 36179 3094
rect 36225 3048 36295 3094
rect 36341 3048 36411 3094
rect 36457 3048 36527 3094
rect 36573 3048 36643 3094
rect 36689 3048 36759 3094
rect 36805 3048 36875 3094
rect 36921 3048 36991 3094
rect 37037 3048 37107 3094
rect 37153 3048 37223 3094
rect 37269 3048 37339 3094
rect 37385 3048 37455 3094
rect 37501 3048 37571 3094
rect 37617 3048 37687 3094
rect 37733 3048 37803 3094
rect 37849 3048 37919 3094
rect 37965 3048 38035 3094
rect 38081 3048 38151 3094
rect 38197 3048 38267 3094
rect 38313 3048 38383 3094
rect 38429 3048 38499 3094
rect 38545 3048 38615 3094
rect 38661 3048 38731 3094
rect 38777 3048 38847 3094
rect 38893 3048 38963 3094
rect 39009 3048 39079 3094
rect 39125 3048 39195 3094
rect 39241 3048 39311 3094
rect 39357 3048 39427 3094
rect 39473 3048 39543 3094
rect 39589 3048 39659 3094
rect 39705 3048 39775 3094
rect 39821 3048 39891 3094
rect 39937 3048 40007 3094
rect 40053 3048 40123 3094
rect 40169 3048 40180 3094
rect 28628 2978 40180 3048
rect 28628 2932 28639 2978
rect 28685 2932 28755 2978
rect 28801 2932 28871 2978
rect 28917 2932 28987 2978
rect 29033 2932 29103 2978
rect 29149 2932 29219 2978
rect 29265 2932 29335 2978
rect 29381 2932 29451 2978
rect 29497 2932 29567 2978
rect 29613 2932 29683 2978
rect 29729 2932 29799 2978
rect 29845 2932 29915 2978
rect 29961 2932 30031 2978
rect 30077 2932 30147 2978
rect 30193 2932 30263 2978
rect 30309 2932 30379 2978
rect 30425 2932 30495 2978
rect 30541 2932 30611 2978
rect 30657 2932 30727 2978
rect 30773 2932 30843 2978
rect 30889 2932 30959 2978
rect 31005 2932 31075 2978
rect 31121 2932 31191 2978
rect 31237 2932 31307 2978
rect 31353 2932 31423 2978
rect 31469 2932 31539 2978
rect 31585 2932 31655 2978
rect 31701 2932 31771 2978
rect 31817 2932 31887 2978
rect 31933 2932 32003 2978
rect 32049 2932 32119 2978
rect 32165 2932 32235 2978
rect 32281 2932 32351 2978
rect 32397 2932 32467 2978
rect 32513 2932 32583 2978
rect 32629 2932 32699 2978
rect 32745 2932 32815 2978
rect 32861 2932 32931 2978
rect 32977 2932 33047 2978
rect 33093 2932 33163 2978
rect 33209 2932 33279 2978
rect 33325 2932 33395 2978
rect 33441 2932 33511 2978
rect 33557 2932 33627 2978
rect 33673 2932 33743 2978
rect 33789 2932 33859 2978
rect 33905 2932 33975 2978
rect 34021 2932 34091 2978
rect 34137 2932 34207 2978
rect 34253 2932 34323 2978
rect 34369 2932 34439 2978
rect 34485 2932 34555 2978
rect 34601 2932 34671 2978
rect 34717 2932 34787 2978
rect 34833 2932 34903 2978
rect 34949 2932 35019 2978
rect 35065 2932 35135 2978
rect 35181 2932 35251 2978
rect 35297 2932 35367 2978
rect 35413 2932 35483 2978
rect 35529 2932 35599 2978
rect 35645 2932 35715 2978
rect 35761 2932 35831 2978
rect 35877 2932 35947 2978
rect 35993 2932 36063 2978
rect 36109 2932 36179 2978
rect 36225 2932 36295 2978
rect 36341 2932 36411 2978
rect 36457 2932 36527 2978
rect 36573 2932 36643 2978
rect 36689 2932 36759 2978
rect 36805 2932 36875 2978
rect 36921 2932 36991 2978
rect 37037 2932 37107 2978
rect 37153 2932 37223 2978
rect 37269 2932 37339 2978
rect 37385 2932 37455 2978
rect 37501 2932 37571 2978
rect 37617 2932 37687 2978
rect 37733 2932 37803 2978
rect 37849 2932 37919 2978
rect 37965 2932 38035 2978
rect 38081 2932 38151 2978
rect 38197 2932 38267 2978
rect 38313 2932 38383 2978
rect 38429 2932 38499 2978
rect 38545 2932 38615 2978
rect 38661 2932 38731 2978
rect 38777 2932 38847 2978
rect 38893 2932 38963 2978
rect 39009 2932 39079 2978
rect 39125 2932 39195 2978
rect 39241 2932 39311 2978
rect 39357 2932 39427 2978
rect 39473 2932 39543 2978
rect 39589 2932 39659 2978
rect 39705 2932 39775 2978
rect 39821 2932 39891 2978
rect 39937 2932 40007 2978
rect 40053 2932 40123 2978
rect 40169 2932 40180 2978
rect 28628 2862 40180 2932
rect 28628 2816 28639 2862
rect 28685 2816 28755 2862
rect 28801 2816 28871 2862
rect 28917 2816 28987 2862
rect 29033 2816 29103 2862
rect 29149 2816 29219 2862
rect 29265 2816 29335 2862
rect 29381 2816 29451 2862
rect 29497 2816 29567 2862
rect 29613 2816 29683 2862
rect 29729 2816 29799 2862
rect 29845 2816 29915 2862
rect 29961 2816 30031 2862
rect 30077 2816 30147 2862
rect 30193 2816 30263 2862
rect 30309 2816 30379 2862
rect 30425 2816 30495 2862
rect 30541 2816 30611 2862
rect 30657 2816 30727 2862
rect 30773 2816 30843 2862
rect 30889 2816 30959 2862
rect 31005 2816 31075 2862
rect 31121 2816 31191 2862
rect 31237 2816 31307 2862
rect 31353 2816 31423 2862
rect 31469 2816 31539 2862
rect 31585 2816 31655 2862
rect 31701 2816 31771 2862
rect 31817 2816 31887 2862
rect 31933 2816 32003 2862
rect 32049 2816 32119 2862
rect 32165 2816 32235 2862
rect 32281 2816 32351 2862
rect 32397 2816 32467 2862
rect 32513 2816 32583 2862
rect 32629 2816 32699 2862
rect 32745 2816 32815 2862
rect 32861 2816 32931 2862
rect 32977 2816 33047 2862
rect 33093 2816 33163 2862
rect 33209 2816 33279 2862
rect 33325 2816 33395 2862
rect 33441 2816 33511 2862
rect 33557 2816 33627 2862
rect 33673 2816 33743 2862
rect 33789 2816 33859 2862
rect 33905 2816 33975 2862
rect 34021 2816 34091 2862
rect 34137 2816 34207 2862
rect 34253 2816 34323 2862
rect 34369 2816 34439 2862
rect 34485 2816 34555 2862
rect 34601 2816 34671 2862
rect 34717 2816 34787 2862
rect 34833 2816 34903 2862
rect 34949 2816 35019 2862
rect 35065 2816 35135 2862
rect 35181 2816 35251 2862
rect 35297 2816 35367 2862
rect 35413 2816 35483 2862
rect 35529 2816 35599 2862
rect 35645 2816 35715 2862
rect 35761 2816 35831 2862
rect 35877 2816 35947 2862
rect 35993 2816 36063 2862
rect 36109 2816 36179 2862
rect 36225 2816 36295 2862
rect 36341 2816 36411 2862
rect 36457 2816 36527 2862
rect 36573 2816 36643 2862
rect 36689 2816 36759 2862
rect 36805 2816 36875 2862
rect 36921 2816 36991 2862
rect 37037 2816 37107 2862
rect 37153 2816 37223 2862
rect 37269 2816 37339 2862
rect 37385 2816 37455 2862
rect 37501 2816 37571 2862
rect 37617 2816 37687 2862
rect 37733 2816 37803 2862
rect 37849 2816 37919 2862
rect 37965 2816 38035 2862
rect 38081 2816 38151 2862
rect 38197 2816 38267 2862
rect 38313 2816 38383 2862
rect 38429 2816 38499 2862
rect 38545 2816 38615 2862
rect 38661 2816 38731 2862
rect 38777 2816 38847 2862
rect 38893 2816 38963 2862
rect 39009 2816 39079 2862
rect 39125 2816 39195 2862
rect 39241 2816 39311 2862
rect 39357 2816 39427 2862
rect 39473 2816 39543 2862
rect 39589 2816 39659 2862
rect 39705 2816 39775 2862
rect 39821 2816 39891 2862
rect 39937 2816 40007 2862
rect 40053 2816 40123 2862
rect 40169 2816 40180 2862
rect 28628 2746 40180 2816
rect 28628 2700 28639 2746
rect 28685 2700 28755 2746
rect 28801 2700 28871 2746
rect 28917 2700 28987 2746
rect 29033 2700 29103 2746
rect 29149 2700 29219 2746
rect 29265 2700 29335 2746
rect 29381 2700 29451 2746
rect 29497 2700 29567 2746
rect 29613 2700 29683 2746
rect 29729 2700 29799 2746
rect 29845 2700 29915 2746
rect 29961 2700 30031 2746
rect 30077 2700 30147 2746
rect 30193 2700 30263 2746
rect 30309 2700 30379 2746
rect 30425 2700 30495 2746
rect 30541 2700 30611 2746
rect 30657 2700 30727 2746
rect 30773 2700 30843 2746
rect 30889 2700 30959 2746
rect 31005 2700 31075 2746
rect 31121 2700 31191 2746
rect 31237 2700 31307 2746
rect 31353 2700 31423 2746
rect 31469 2700 31539 2746
rect 31585 2700 31655 2746
rect 31701 2700 31771 2746
rect 31817 2700 31887 2746
rect 31933 2700 32003 2746
rect 32049 2700 32119 2746
rect 32165 2700 32235 2746
rect 32281 2700 32351 2746
rect 32397 2700 32467 2746
rect 32513 2700 32583 2746
rect 32629 2700 32699 2746
rect 32745 2700 32815 2746
rect 32861 2700 32931 2746
rect 32977 2700 33047 2746
rect 33093 2700 33163 2746
rect 33209 2700 33279 2746
rect 33325 2700 33395 2746
rect 33441 2700 33511 2746
rect 33557 2700 33627 2746
rect 33673 2700 33743 2746
rect 33789 2700 33859 2746
rect 33905 2700 33975 2746
rect 34021 2700 34091 2746
rect 34137 2700 34207 2746
rect 34253 2700 34323 2746
rect 34369 2700 34439 2746
rect 34485 2700 34555 2746
rect 34601 2700 34671 2746
rect 34717 2700 34787 2746
rect 34833 2700 34903 2746
rect 34949 2700 35019 2746
rect 35065 2700 35135 2746
rect 35181 2700 35251 2746
rect 35297 2700 35367 2746
rect 35413 2700 35483 2746
rect 35529 2700 35599 2746
rect 35645 2700 35715 2746
rect 35761 2700 35831 2746
rect 35877 2700 35947 2746
rect 35993 2700 36063 2746
rect 36109 2700 36179 2746
rect 36225 2700 36295 2746
rect 36341 2700 36411 2746
rect 36457 2700 36527 2746
rect 36573 2700 36643 2746
rect 36689 2700 36759 2746
rect 36805 2700 36875 2746
rect 36921 2700 36991 2746
rect 37037 2700 37107 2746
rect 37153 2700 37223 2746
rect 37269 2700 37339 2746
rect 37385 2700 37455 2746
rect 37501 2700 37571 2746
rect 37617 2700 37687 2746
rect 37733 2700 37803 2746
rect 37849 2700 37919 2746
rect 37965 2700 38035 2746
rect 38081 2700 38151 2746
rect 38197 2700 38267 2746
rect 38313 2700 38383 2746
rect 38429 2700 38499 2746
rect 38545 2700 38615 2746
rect 38661 2700 38731 2746
rect 38777 2700 38847 2746
rect 38893 2700 38963 2746
rect 39009 2700 39079 2746
rect 39125 2700 39195 2746
rect 39241 2700 39311 2746
rect 39357 2700 39427 2746
rect 39473 2700 39543 2746
rect 39589 2700 39659 2746
rect 39705 2700 39775 2746
rect 39821 2700 39891 2746
rect 39937 2700 40007 2746
rect 40053 2700 40123 2746
rect 40169 2700 40180 2746
rect 28628 2630 40180 2700
rect 28628 2584 28639 2630
rect 28685 2584 28755 2630
rect 28801 2584 28871 2630
rect 28917 2584 28987 2630
rect 29033 2584 29103 2630
rect 29149 2584 29219 2630
rect 29265 2584 29335 2630
rect 29381 2584 29451 2630
rect 29497 2584 29567 2630
rect 29613 2584 29683 2630
rect 29729 2584 29799 2630
rect 29845 2584 29915 2630
rect 29961 2584 30031 2630
rect 30077 2584 30147 2630
rect 30193 2584 30263 2630
rect 30309 2584 30379 2630
rect 30425 2584 30495 2630
rect 30541 2584 30611 2630
rect 30657 2584 30727 2630
rect 30773 2584 30843 2630
rect 30889 2584 30959 2630
rect 31005 2584 31075 2630
rect 31121 2584 31191 2630
rect 31237 2584 31307 2630
rect 31353 2584 31423 2630
rect 31469 2584 31539 2630
rect 31585 2584 31655 2630
rect 31701 2584 31771 2630
rect 31817 2584 31887 2630
rect 31933 2584 32003 2630
rect 32049 2584 32119 2630
rect 32165 2584 32235 2630
rect 32281 2584 32351 2630
rect 32397 2584 32467 2630
rect 32513 2584 32583 2630
rect 32629 2584 32699 2630
rect 32745 2584 32815 2630
rect 32861 2584 32931 2630
rect 32977 2584 33047 2630
rect 33093 2584 33163 2630
rect 33209 2584 33279 2630
rect 33325 2584 33395 2630
rect 33441 2584 33511 2630
rect 33557 2584 33627 2630
rect 33673 2584 33743 2630
rect 33789 2584 33859 2630
rect 33905 2584 33975 2630
rect 34021 2584 34091 2630
rect 34137 2584 34207 2630
rect 34253 2584 34323 2630
rect 34369 2584 34439 2630
rect 34485 2584 34555 2630
rect 34601 2584 34671 2630
rect 34717 2584 34787 2630
rect 34833 2584 34903 2630
rect 34949 2584 35019 2630
rect 35065 2584 35135 2630
rect 35181 2584 35251 2630
rect 35297 2584 35367 2630
rect 35413 2584 35483 2630
rect 35529 2584 35599 2630
rect 35645 2584 35715 2630
rect 35761 2584 35831 2630
rect 35877 2584 35947 2630
rect 35993 2584 36063 2630
rect 36109 2584 36179 2630
rect 36225 2584 36295 2630
rect 36341 2584 36411 2630
rect 36457 2584 36527 2630
rect 36573 2584 36643 2630
rect 36689 2584 36759 2630
rect 36805 2584 36875 2630
rect 36921 2584 36991 2630
rect 37037 2584 37107 2630
rect 37153 2584 37223 2630
rect 37269 2584 37339 2630
rect 37385 2584 37455 2630
rect 37501 2584 37571 2630
rect 37617 2584 37687 2630
rect 37733 2584 37803 2630
rect 37849 2584 37919 2630
rect 37965 2584 38035 2630
rect 38081 2584 38151 2630
rect 38197 2584 38267 2630
rect 38313 2584 38383 2630
rect 38429 2584 38499 2630
rect 38545 2584 38615 2630
rect 38661 2584 38731 2630
rect 38777 2584 38847 2630
rect 38893 2584 38963 2630
rect 39009 2584 39079 2630
rect 39125 2584 39195 2630
rect 39241 2584 39311 2630
rect 39357 2584 39427 2630
rect 39473 2584 39543 2630
rect 39589 2584 39659 2630
rect 39705 2584 39775 2630
rect 39821 2584 39891 2630
rect 39937 2584 40007 2630
rect 40053 2584 40123 2630
rect 40169 2584 40180 2630
rect 28628 2514 40180 2584
rect 28628 2468 28639 2514
rect 28685 2468 28755 2514
rect 28801 2468 28871 2514
rect 28917 2468 28987 2514
rect 29033 2468 29103 2514
rect 29149 2468 29219 2514
rect 29265 2468 29335 2514
rect 29381 2468 29451 2514
rect 29497 2468 29567 2514
rect 29613 2468 29683 2514
rect 29729 2468 29799 2514
rect 29845 2468 29915 2514
rect 29961 2468 30031 2514
rect 30077 2468 30147 2514
rect 30193 2468 30263 2514
rect 30309 2468 30379 2514
rect 30425 2468 30495 2514
rect 30541 2468 30611 2514
rect 30657 2468 30727 2514
rect 30773 2468 30843 2514
rect 30889 2468 30959 2514
rect 31005 2468 31075 2514
rect 31121 2468 31191 2514
rect 31237 2468 31307 2514
rect 31353 2468 31423 2514
rect 31469 2468 31539 2514
rect 31585 2468 31655 2514
rect 31701 2468 31771 2514
rect 31817 2468 31887 2514
rect 31933 2468 32003 2514
rect 32049 2468 32119 2514
rect 32165 2468 32235 2514
rect 32281 2468 32351 2514
rect 32397 2468 32467 2514
rect 32513 2468 32583 2514
rect 32629 2468 32699 2514
rect 32745 2468 32815 2514
rect 32861 2468 32931 2514
rect 32977 2468 33047 2514
rect 33093 2468 33163 2514
rect 33209 2468 33279 2514
rect 33325 2468 33395 2514
rect 33441 2468 33511 2514
rect 33557 2468 33627 2514
rect 33673 2468 33743 2514
rect 33789 2468 33859 2514
rect 33905 2468 33975 2514
rect 34021 2468 34091 2514
rect 34137 2468 34207 2514
rect 34253 2468 34323 2514
rect 34369 2468 34439 2514
rect 34485 2468 34555 2514
rect 34601 2468 34671 2514
rect 34717 2468 34787 2514
rect 34833 2468 34903 2514
rect 34949 2468 35019 2514
rect 35065 2468 35135 2514
rect 35181 2468 35251 2514
rect 35297 2468 35367 2514
rect 35413 2468 35483 2514
rect 35529 2468 35599 2514
rect 35645 2468 35715 2514
rect 35761 2468 35831 2514
rect 35877 2468 35947 2514
rect 35993 2468 36063 2514
rect 36109 2468 36179 2514
rect 36225 2468 36295 2514
rect 36341 2468 36411 2514
rect 36457 2468 36527 2514
rect 36573 2468 36643 2514
rect 36689 2468 36759 2514
rect 36805 2468 36875 2514
rect 36921 2468 36991 2514
rect 37037 2468 37107 2514
rect 37153 2468 37223 2514
rect 37269 2468 37339 2514
rect 37385 2468 37455 2514
rect 37501 2468 37571 2514
rect 37617 2468 37687 2514
rect 37733 2468 37803 2514
rect 37849 2468 37919 2514
rect 37965 2468 38035 2514
rect 38081 2468 38151 2514
rect 38197 2468 38267 2514
rect 38313 2468 38383 2514
rect 38429 2468 38499 2514
rect 38545 2468 38615 2514
rect 38661 2468 38731 2514
rect 38777 2468 38847 2514
rect 38893 2468 38963 2514
rect 39009 2468 39079 2514
rect 39125 2468 39195 2514
rect 39241 2468 39311 2514
rect 39357 2468 39427 2514
rect 39473 2468 39543 2514
rect 39589 2468 39659 2514
rect 39705 2468 39775 2514
rect 39821 2468 39891 2514
rect 39937 2468 40007 2514
rect 40053 2468 40123 2514
rect 40169 2468 40180 2514
rect 28628 2398 40180 2468
rect 28628 2352 28639 2398
rect 28685 2352 28755 2398
rect 28801 2352 28871 2398
rect 28917 2352 28987 2398
rect 29033 2352 29103 2398
rect 29149 2352 29219 2398
rect 29265 2352 29335 2398
rect 29381 2352 29451 2398
rect 29497 2352 29567 2398
rect 29613 2352 29683 2398
rect 29729 2352 29799 2398
rect 29845 2352 29915 2398
rect 29961 2352 30031 2398
rect 30077 2352 30147 2398
rect 30193 2352 30263 2398
rect 30309 2352 30379 2398
rect 30425 2352 30495 2398
rect 30541 2352 30611 2398
rect 30657 2352 30727 2398
rect 30773 2352 30843 2398
rect 30889 2352 30959 2398
rect 31005 2352 31075 2398
rect 31121 2352 31191 2398
rect 31237 2352 31307 2398
rect 31353 2352 31423 2398
rect 31469 2352 31539 2398
rect 31585 2352 31655 2398
rect 31701 2352 31771 2398
rect 31817 2352 31887 2398
rect 31933 2352 32003 2398
rect 32049 2352 32119 2398
rect 32165 2352 32235 2398
rect 32281 2352 32351 2398
rect 32397 2352 32467 2398
rect 32513 2352 32583 2398
rect 32629 2352 32699 2398
rect 32745 2352 32815 2398
rect 32861 2352 32931 2398
rect 32977 2352 33047 2398
rect 33093 2352 33163 2398
rect 33209 2352 33279 2398
rect 33325 2352 33395 2398
rect 33441 2352 33511 2398
rect 33557 2352 33627 2398
rect 33673 2352 33743 2398
rect 33789 2352 33859 2398
rect 33905 2352 33975 2398
rect 34021 2352 34091 2398
rect 34137 2352 34207 2398
rect 34253 2352 34323 2398
rect 34369 2352 34439 2398
rect 34485 2352 34555 2398
rect 34601 2352 34671 2398
rect 34717 2352 34787 2398
rect 34833 2352 34903 2398
rect 34949 2352 35019 2398
rect 35065 2352 35135 2398
rect 35181 2352 35251 2398
rect 35297 2352 35367 2398
rect 35413 2352 35483 2398
rect 35529 2352 35599 2398
rect 35645 2352 35715 2398
rect 35761 2352 35831 2398
rect 35877 2352 35947 2398
rect 35993 2352 36063 2398
rect 36109 2352 36179 2398
rect 36225 2352 36295 2398
rect 36341 2352 36411 2398
rect 36457 2352 36527 2398
rect 36573 2352 36643 2398
rect 36689 2352 36759 2398
rect 36805 2352 36875 2398
rect 36921 2352 36991 2398
rect 37037 2352 37107 2398
rect 37153 2352 37223 2398
rect 37269 2352 37339 2398
rect 37385 2352 37455 2398
rect 37501 2352 37571 2398
rect 37617 2352 37687 2398
rect 37733 2352 37803 2398
rect 37849 2352 37919 2398
rect 37965 2352 38035 2398
rect 38081 2352 38151 2398
rect 38197 2352 38267 2398
rect 38313 2352 38383 2398
rect 38429 2352 38499 2398
rect 38545 2352 38615 2398
rect 38661 2352 38731 2398
rect 38777 2352 38847 2398
rect 38893 2352 38963 2398
rect 39009 2352 39079 2398
rect 39125 2352 39195 2398
rect 39241 2352 39311 2398
rect 39357 2352 39427 2398
rect 39473 2352 39543 2398
rect 39589 2352 39659 2398
rect 39705 2352 39775 2398
rect 39821 2352 39891 2398
rect 39937 2352 40007 2398
rect 40053 2352 40123 2398
rect 40169 2352 40180 2398
rect 28628 2282 40180 2352
rect 28628 2236 28639 2282
rect 28685 2236 28755 2282
rect 28801 2236 28871 2282
rect 28917 2236 28987 2282
rect 29033 2236 29103 2282
rect 29149 2236 29219 2282
rect 29265 2236 29335 2282
rect 29381 2236 29451 2282
rect 29497 2236 29567 2282
rect 29613 2236 29683 2282
rect 29729 2236 29799 2282
rect 29845 2236 29915 2282
rect 29961 2236 30031 2282
rect 30077 2236 30147 2282
rect 30193 2236 30263 2282
rect 30309 2236 30379 2282
rect 30425 2236 30495 2282
rect 30541 2236 30611 2282
rect 30657 2236 30727 2282
rect 30773 2236 30843 2282
rect 30889 2236 30959 2282
rect 31005 2236 31075 2282
rect 31121 2236 31191 2282
rect 31237 2236 31307 2282
rect 31353 2236 31423 2282
rect 31469 2236 31539 2282
rect 31585 2236 31655 2282
rect 31701 2236 31771 2282
rect 31817 2236 31887 2282
rect 31933 2236 32003 2282
rect 32049 2236 32119 2282
rect 32165 2236 32235 2282
rect 32281 2236 32351 2282
rect 32397 2236 32467 2282
rect 32513 2236 32583 2282
rect 32629 2236 32699 2282
rect 32745 2236 32815 2282
rect 32861 2236 32931 2282
rect 32977 2236 33047 2282
rect 33093 2236 33163 2282
rect 33209 2236 33279 2282
rect 33325 2236 33395 2282
rect 33441 2236 33511 2282
rect 33557 2236 33627 2282
rect 33673 2236 33743 2282
rect 33789 2236 33859 2282
rect 33905 2236 33975 2282
rect 34021 2236 34091 2282
rect 34137 2236 34207 2282
rect 34253 2236 34323 2282
rect 34369 2236 34439 2282
rect 34485 2236 34555 2282
rect 34601 2236 34671 2282
rect 34717 2236 34787 2282
rect 34833 2236 34903 2282
rect 34949 2236 35019 2282
rect 35065 2236 35135 2282
rect 35181 2236 35251 2282
rect 35297 2236 35367 2282
rect 35413 2236 35483 2282
rect 35529 2236 35599 2282
rect 35645 2236 35715 2282
rect 35761 2236 35831 2282
rect 35877 2236 35947 2282
rect 35993 2236 36063 2282
rect 36109 2236 36179 2282
rect 36225 2236 36295 2282
rect 36341 2236 36411 2282
rect 36457 2236 36527 2282
rect 36573 2236 36643 2282
rect 36689 2236 36759 2282
rect 36805 2236 36875 2282
rect 36921 2236 36991 2282
rect 37037 2236 37107 2282
rect 37153 2236 37223 2282
rect 37269 2236 37339 2282
rect 37385 2236 37455 2282
rect 37501 2236 37571 2282
rect 37617 2236 37687 2282
rect 37733 2236 37803 2282
rect 37849 2236 37919 2282
rect 37965 2236 38035 2282
rect 38081 2236 38151 2282
rect 38197 2236 38267 2282
rect 38313 2236 38383 2282
rect 38429 2236 38499 2282
rect 38545 2236 38615 2282
rect 38661 2236 38731 2282
rect 38777 2236 38847 2282
rect 38893 2236 38963 2282
rect 39009 2236 39079 2282
rect 39125 2236 39195 2282
rect 39241 2236 39311 2282
rect 39357 2236 39427 2282
rect 39473 2236 39543 2282
rect 39589 2236 39659 2282
rect 39705 2236 39775 2282
rect 39821 2236 39891 2282
rect 39937 2236 40007 2282
rect 40053 2236 40123 2282
rect 40169 2236 40180 2282
rect 28628 2166 40180 2236
rect 28628 2120 28639 2166
rect 28685 2120 28755 2166
rect 28801 2120 28871 2166
rect 28917 2120 28987 2166
rect 29033 2120 29103 2166
rect 29149 2120 29219 2166
rect 29265 2120 29335 2166
rect 29381 2120 29451 2166
rect 29497 2120 29567 2166
rect 29613 2120 29683 2166
rect 29729 2120 29799 2166
rect 29845 2120 29915 2166
rect 29961 2120 30031 2166
rect 30077 2120 30147 2166
rect 30193 2120 30263 2166
rect 30309 2120 30379 2166
rect 30425 2120 30495 2166
rect 30541 2120 30611 2166
rect 30657 2120 30727 2166
rect 30773 2120 30843 2166
rect 30889 2120 30959 2166
rect 31005 2120 31075 2166
rect 31121 2120 31191 2166
rect 31237 2120 31307 2166
rect 31353 2120 31423 2166
rect 31469 2120 31539 2166
rect 31585 2120 31655 2166
rect 31701 2120 31771 2166
rect 31817 2120 31887 2166
rect 31933 2120 32003 2166
rect 32049 2120 32119 2166
rect 32165 2120 32235 2166
rect 32281 2120 32351 2166
rect 32397 2120 32467 2166
rect 32513 2120 32583 2166
rect 32629 2120 32699 2166
rect 32745 2120 32815 2166
rect 32861 2120 32931 2166
rect 32977 2120 33047 2166
rect 33093 2120 33163 2166
rect 33209 2120 33279 2166
rect 33325 2120 33395 2166
rect 33441 2120 33511 2166
rect 33557 2120 33627 2166
rect 33673 2120 33743 2166
rect 33789 2120 33859 2166
rect 33905 2120 33975 2166
rect 34021 2120 34091 2166
rect 34137 2120 34207 2166
rect 34253 2120 34323 2166
rect 34369 2120 34439 2166
rect 34485 2120 34555 2166
rect 34601 2120 34671 2166
rect 34717 2120 34787 2166
rect 34833 2120 34903 2166
rect 34949 2120 35019 2166
rect 35065 2120 35135 2166
rect 35181 2120 35251 2166
rect 35297 2120 35367 2166
rect 35413 2120 35483 2166
rect 35529 2120 35599 2166
rect 35645 2120 35715 2166
rect 35761 2120 35831 2166
rect 35877 2120 35947 2166
rect 35993 2120 36063 2166
rect 36109 2120 36179 2166
rect 36225 2120 36295 2166
rect 36341 2120 36411 2166
rect 36457 2120 36527 2166
rect 36573 2120 36643 2166
rect 36689 2120 36759 2166
rect 36805 2120 36875 2166
rect 36921 2120 36991 2166
rect 37037 2120 37107 2166
rect 37153 2120 37223 2166
rect 37269 2120 37339 2166
rect 37385 2120 37455 2166
rect 37501 2120 37571 2166
rect 37617 2120 37687 2166
rect 37733 2120 37803 2166
rect 37849 2120 37919 2166
rect 37965 2120 38035 2166
rect 38081 2120 38151 2166
rect 38197 2120 38267 2166
rect 38313 2120 38383 2166
rect 38429 2120 38499 2166
rect 38545 2120 38615 2166
rect 38661 2120 38731 2166
rect 38777 2120 38847 2166
rect 38893 2120 38963 2166
rect 39009 2120 39079 2166
rect 39125 2120 39195 2166
rect 39241 2120 39311 2166
rect 39357 2120 39427 2166
rect 39473 2120 39543 2166
rect 39589 2120 39659 2166
rect 39705 2120 39775 2166
rect 39821 2120 39891 2166
rect 39937 2120 40007 2166
rect 40053 2120 40123 2166
rect 40169 2120 40180 2166
rect 28628 2050 40180 2120
rect 28628 2004 28639 2050
rect 28685 2004 28755 2050
rect 28801 2004 28871 2050
rect 28917 2004 28987 2050
rect 29033 2004 29103 2050
rect 29149 2004 29219 2050
rect 29265 2004 29335 2050
rect 29381 2004 29451 2050
rect 29497 2004 29567 2050
rect 29613 2004 29683 2050
rect 29729 2004 29799 2050
rect 29845 2004 29915 2050
rect 29961 2004 30031 2050
rect 30077 2004 30147 2050
rect 30193 2004 30263 2050
rect 30309 2004 30379 2050
rect 30425 2004 30495 2050
rect 30541 2004 30611 2050
rect 30657 2004 30727 2050
rect 30773 2004 30843 2050
rect 30889 2004 30959 2050
rect 31005 2004 31075 2050
rect 31121 2004 31191 2050
rect 31237 2004 31307 2050
rect 31353 2004 31423 2050
rect 31469 2004 31539 2050
rect 31585 2004 31655 2050
rect 31701 2004 31771 2050
rect 31817 2004 31887 2050
rect 31933 2004 32003 2050
rect 32049 2004 32119 2050
rect 32165 2004 32235 2050
rect 32281 2004 32351 2050
rect 32397 2004 32467 2050
rect 32513 2004 32583 2050
rect 32629 2004 32699 2050
rect 32745 2004 32815 2050
rect 32861 2004 32931 2050
rect 32977 2004 33047 2050
rect 33093 2004 33163 2050
rect 33209 2004 33279 2050
rect 33325 2004 33395 2050
rect 33441 2004 33511 2050
rect 33557 2004 33627 2050
rect 33673 2004 33743 2050
rect 33789 2004 33859 2050
rect 33905 2004 33975 2050
rect 34021 2004 34091 2050
rect 34137 2004 34207 2050
rect 34253 2004 34323 2050
rect 34369 2004 34439 2050
rect 34485 2004 34555 2050
rect 34601 2004 34671 2050
rect 34717 2004 34787 2050
rect 34833 2004 34903 2050
rect 34949 2004 35019 2050
rect 35065 2004 35135 2050
rect 35181 2004 35251 2050
rect 35297 2004 35367 2050
rect 35413 2004 35483 2050
rect 35529 2004 35599 2050
rect 35645 2004 35715 2050
rect 35761 2004 35831 2050
rect 35877 2004 35947 2050
rect 35993 2004 36063 2050
rect 36109 2004 36179 2050
rect 36225 2004 36295 2050
rect 36341 2004 36411 2050
rect 36457 2004 36527 2050
rect 36573 2004 36643 2050
rect 36689 2004 36759 2050
rect 36805 2004 36875 2050
rect 36921 2004 36991 2050
rect 37037 2004 37107 2050
rect 37153 2004 37223 2050
rect 37269 2004 37339 2050
rect 37385 2004 37455 2050
rect 37501 2004 37571 2050
rect 37617 2004 37687 2050
rect 37733 2004 37803 2050
rect 37849 2004 37919 2050
rect 37965 2004 38035 2050
rect 38081 2004 38151 2050
rect 38197 2004 38267 2050
rect 38313 2004 38383 2050
rect 38429 2004 38499 2050
rect 38545 2004 38615 2050
rect 38661 2004 38731 2050
rect 38777 2004 38847 2050
rect 38893 2004 38963 2050
rect 39009 2004 39079 2050
rect 39125 2004 39195 2050
rect 39241 2004 39311 2050
rect 39357 2004 39427 2050
rect 39473 2004 39543 2050
rect 39589 2004 39659 2050
rect 39705 2004 39775 2050
rect 39821 2004 39891 2050
rect 39937 2004 40007 2050
rect 40053 2004 40123 2050
rect 40169 2004 40180 2050
rect 28628 1934 40180 2004
rect 28628 1925 28639 1934
rect 27744 1888 28639 1925
rect 28685 1888 28755 1934
rect 28801 1888 28871 1934
rect 28917 1888 28987 1934
rect 29033 1888 29103 1934
rect 29149 1888 29219 1934
rect 29265 1888 29335 1934
rect 29381 1888 29451 1934
rect 29497 1888 29567 1934
rect 29613 1888 29683 1934
rect 29729 1888 29799 1934
rect 29845 1888 29915 1934
rect 29961 1888 30031 1934
rect 30077 1888 30147 1934
rect 30193 1888 30263 1934
rect 30309 1888 30379 1934
rect 30425 1888 30495 1934
rect 30541 1888 30611 1934
rect 30657 1888 30727 1934
rect 30773 1888 30843 1934
rect 30889 1888 30959 1934
rect 31005 1888 31075 1934
rect 31121 1888 31191 1934
rect 31237 1888 31307 1934
rect 31353 1888 31423 1934
rect 31469 1888 31539 1934
rect 31585 1888 31655 1934
rect 31701 1888 31771 1934
rect 31817 1888 31887 1934
rect 31933 1888 32003 1934
rect 32049 1888 32119 1934
rect 32165 1888 32235 1934
rect 32281 1888 32351 1934
rect 32397 1888 32467 1934
rect 32513 1888 32583 1934
rect 32629 1888 32699 1934
rect 32745 1888 32815 1934
rect 32861 1888 32931 1934
rect 32977 1888 33047 1934
rect 33093 1888 33163 1934
rect 33209 1888 33279 1934
rect 33325 1888 33395 1934
rect 33441 1888 33511 1934
rect 33557 1888 33627 1934
rect 33673 1888 33743 1934
rect 33789 1888 33859 1934
rect 33905 1888 33975 1934
rect 34021 1888 34091 1934
rect 34137 1888 34207 1934
rect 34253 1888 34323 1934
rect 34369 1888 34439 1934
rect 34485 1888 34555 1934
rect 34601 1888 34671 1934
rect 34717 1888 34787 1934
rect 34833 1888 34903 1934
rect 34949 1888 35019 1934
rect 35065 1888 35135 1934
rect 35181 1888 35251 1934
rect 35297 1888 35367 1934
rect 35413 1888 35483 1934
rect 35529 1888 35599 1934
rect 35645 1888 35715 1934
rect 35761 1888 35831 1934
rect 35877 1888 35947 1934
rect 35993 1888 36063 1934
rect 36109 1888 36179 1934
rect 36225 1888 36295 1934
rect 36341 1888 36411 1934
rect 36457 1888 36527 1934
rect 36573 1888 36643 1934
rect 36689 1888 36759 1934
rect 36805 1888 36875 1934
rect 36921 1888 36991 1934
rect 37037 1888 37107 1934
rect 37153 1888 37223 1934
rect 37269 1888 37339 1934
rect 37385 1888 37455 1934
rect 37501 1888 37571 1934
rect 37617 1888 37687 1934
rect 37733 1888 37803 1934
rect 37849 1888 37919 1934
rect 37965 1888 38035 1934
rect 38081 1888 38151 1934
rect 38197 1888 38267 1934
rect 38313 1888 38383 1934
rect 38429 1888 38499 1934
rect 38545 1888 38615 1934
rect 38661 1888 38731 1934
rect 38777 1888 38847 1934
rect 38893 1888 38963 1934
rect 39009 1888 39079 1934
rect 39125 1888 39195 1934
rect 39241 1888 39311 1934
rect 39357 1888 39427 1934
rect 39473 1888 39543 1934
rect 39589 1888 39659 1934
rect 39705 1888 39775 1934
rect 39821 1888 39891 1934
rect 39937 1888 40007 1934
rect 40053 1888 40123 1934
rect 40169 1925 40180 1934
rect 50834 3210 56586 3280
rect 50834 3164 50845 3210
rect 50891 3164 50961 3210
rect 51007 3164 51077 3210
rect 51123 3164 51193 3210
rect 51239 3164 51309 3210
rect 51355 3164 51425 3210
rect 51471 3164 51541 3210
rect 51587 3164 51657 3210
rect 51703 3164 51773 3210
rect 51819 3164 51889 3210
rect 51935 3164 52005 3210
rect 52051 3164 52121 3210
rect 52167 3164 52237 3210
rect 52283 3164 52353 3210
rect 52399 3164 52469 3210
rect 52515 3164 52585 3210
rect 52631 3164 52701 3210
rect 52747 3164 52817 3210
rect 52863 3164 52933 3210
rect 52979 3164 53049 3210
rect 53095 3164 53165 3210
rect 53211 3164 53281 3210
rect 53327 3164 53397 3210
rect 53443 3164 53513 3210
rect 53559 3164 53629 3210
rect 53675 3164 53745 3210
rect 53791 3164 53861 3210
rect 53907 3164 53977 3210
rect 54023 3164 54093 3210
rect 54139 3164 54209 3210
rect 54255 3164 54325 3210
rect 54371 3164 54441 3210
rect 54487 3164 54557 3210
rect 54603 3164 54673 3210
rect 54719 3164 54789 3210
rect 54835 3164 54905 3210
rect 54951 3164 55021 3210
rect 55067 3164 55137 3210
rect 55183 3164 55253 3210
rect 55299 3164 55369 3210
rect 55415 3164 55485 3210
rect 55531 3164 55601 3210
rect 55647 3164 55717 3210
rect 55763 3164 55833 3210
rect 55879 3164 55949 3210
rect 55995 3164 56065 3210
rect 56111 3164 56181 3210
rect 56227 3164 56297 3210
rect 56343 3164 56413 3210
rect 56459 3164 56529 3210
rect 56575 3164 56586 3210
rect 50834 3094 56586 3164
rect 50834 3048 50845 3094
rect 50891 3048 50961 3094
rect 51007 3048 51077 3094
rect 51123 3048 51193 3094
rect 51239 3048 51309 3094
rect 51355 3048 51425 3094
rect 51471 3048 51541 3094
rect 51587 3048 51657 3094
rect 51703 3048 51773 3094
rect 51819 3048 51889 3094
rect 51935 3048 52005 3094
rect 52051 3048 52121 3094
rect 52167 3048 52237 3094
rect 52283 3048 52353 3094
rect 52399 3048 52469 3094
rect 52515 3048 52585 3094
rect 52631 3048 52701 3094
rect 52747 3048 52817 3094
rect 52863 3048 52933 3094
rect 52979 3048 53049 3094
rect 53095 3048 53165 3094
rect 53211 3048 53281 3094
rect 53327 3048 53397 3094
rect 53443 3048 53513 3094
rect 53559 3048 53629 3094
rect 53675 3048 53745 3094
rect 53791 3048 53861 3094
rect 53907 3048 53977 3094
rect 54023 3048 54093 3094
rect 54139 3048 54209 3094
rect 54255 3048 54325 3094
rect 54371 3048 54441 3094
rect 54487 3048 54557 3094
rect 54603 3048 54673 3094
rect 54719 3048 54789 3094
rect 54835 3048 54905 3094
rect 54951 3048 55021 3094
rect 55067 3048 55137 3094
rect 55183 3048 55253 3094
rect 55299 3048 55369 3094
rect 55415 3048 55485 3094
rect 55531 3048 55601 3094
rect 55647 3048 55717 3094
rect 55763 3048 55833 3094
rect 55879 3048 55949 3094
rect 55995 3048 56065 3094
rect 56111 3048 56181 3094
rect 56227 3048 56297 3094
rect 56343 3048 56413 3094
rect 56459 3048 56529 3094
rect 56575 3048 56586 3094
rect 50834 2978 56586 3048
rect 50834 2932 50845 2978
rect 50891 2932 50961 2978
rect 51007 2932 51077 2978
rect 51123 2932 51193 2978
rect 51239 2932 51309 2978
rect 51355 2932 51425 2978
rect 51471 2932 51541 2978
rect 51587 2932 51657 2978
rect 51703 2932 51773 2978
rect 51819 2932 51889 2978
rect 51935 2932 52005 2978
rect 52051 2932 52121 2978
rect 52167 2932 52237 2978
rect 52283 2932 52353 2978
rect 52399 2932 52469 2978
rect 52515 2932 52585 2978
rect 52631 2932 52701 2978
rect 52747 2932 52817 2978
rect 52863 2932 52933 2978
rect 52979 2932 53049 2978
rect 53095 2932 53165 2978
rect 53211 2932 53281 2978
rect 53327 2932 53397 2978
rect 53443 2932 53513 2978
rect 53559 2932 53629 2978
rect 53675 2932 53745 2978
rect 53791 2932 53861 2978
rect 53907 2932 53977 2978
rect 54023 2932 54093 2978
rect 54139 2932 54209 2978
rect 54255 2932 54325 2978
rect 54371 2932 54441 2978
rect 54487 2932 54557 2978
rect 54603 2932 54673 2978
rect 54719 2932 54789 2978
rect 54835 2932 54905 2978
rect 54951 2932 55021 2978
rect 55067 2932 55137 2978
rect 55183 2932 55253 2978
rect 55299 2932 55369 2978
rect 55415 2932 55485 2978
rect 55531 2932 55601 2978
rect 55647 2932 55717 2978
rect 55763 2932 55833 2978
rect 55879 2932 55949 2978
rect 55995 2932 56065 2978
rect 56111 2932 56181 2978
rect 56227 2932 56297 2978
rect 56343 2932 56413 2978
rect 56459 2932 56529 2978
rect 56575 2932 56586 2978
rect 50834 2862 56586 2932
rect 50834 2816 50845 2862
rect 50891 2816 50961 2862
rect 51007 2816 51077 2862
rect 51123 2816 51193 2862
rect 51239 2816 51309 2862
rect 51355 2816 51425 2862
rect 51471 2816 51541 2862
rect 51587 2816 51657 2862
rect 51703 2816 51773 2862
rect 51819 2816 51889 2862
rect 51935 2816 52005 2862
rect 52051 2816 52121 2862
rect 52167 2816 52237 2862
rect 52283 2816 52353 2862
rect 52399 2816 52469 2862
rect 52515 2816 52585 2862
rect 52631 2816 52701 2862
rect 52747 2816 52817 2862
rect 52863 2816 52933 2862
rect 52979 2816 53049 2862
rect 53095 2816 53165 2862
rect 53211 2816 53281 2862
rect 53327 2816 53397 2862
rect 53443 2816 53513 2862
rect 53559 2816 53629 2862
rect 53675 2816 53745 2862
rect 53791 2816 53861 2862
rect 53907 2816 53977 2862
rect 54023 2816 54093 2862
rect 54139 2816 54209 2862
rect 54255 2816 54325 2862
rect 54371 2816 54441 2862
rect 54487 2816 54557 2862
rect 54603 2816 54673 2862
rect 54719 2816 54789 2862
rect 54835 2816 54905 2862
rect 54951 2816 55021 2862
rect 55067 2816 55137 2862
rect 55183 2816 55253 2862
rect 55299 2816 55369 2862
rect 55415 2816 55485 2862
rect 55531 2816 55601 2862
rect 55647 2816 55717 2862
rect 55763 2816 55833 2862
rect 55879 2816 55949 2862
rect 55995 2816 56065 2862
rect 56111 2816 56181 2862
rect 56227 2816 56297 2862
rect 56343 2816 56413 2862
rect 56459 2816 56529 2862
rect 56575 2816 56586 2862
rect 50834 2746 56586 2816
rect 50834 2700 50845 2746
rect 50891 2700 50961 2746
rect 51007 2700 51077 2746
rect 51123 2700 51193 2746
rect 51239 2700 51309 2746
rect 51355 2700 51425 2746
rect 51471 2700 51541 2746
rect 51587 2700 51657 2746
rect 51703 2700 51773 2746
rect 51819 2700 51889 2746
rect 51935 2700 52005 2746
rect 52051 2700 52121 2746
rect 52167 2700 52237 2746
rect 52283 2700 52353 2746
rect 52399 2700 52469 2746
rect 52515 2700 52585 2746
rect 52631 2700 52701 2746
rect 52747 2700 52817 2746
rect 52863 2700 52933 2746
rect 52979 2700 53049 2746
rect 53095 2700 53165 2746
rect 53211 2700 53281 2746
rect 53327 2700 53397 2746
rect 53443 2700 53513 2746
rect 53559 2700 53629 2746
rect 53675 2700 53745 2746
rect 53791 2700 53861 2746
rect 53907 2700 53977 2746
rect 54023 2700 54093 2746
rect 54139 2700 54209 2746
rect 54255 2700 54325 2746
rect 54371 2700 54441 2746
rect 54487 2700 54557 2746
rect 54603 2700 54673 2746
rect 54719 2700 54789 2746
rect 54835 2700 54905 2746
rect 54951 2700 55021 2746
rect 55067 2700 55137 2746
rect 55183 2700 55253 2746
rect 55299 2700 55369 2746
rect 55415 2700 55485 2746
rect 55531 2700 55601 2746
rect 55647 2700 55717 2746
rect 55763 2700 55833 2746
rect 55879 2700 55949 2746
rect 55995 2700 56065 2746
rect 56111 2700 56181 2746
rect 56227 2700 56297 2746
rect 56343 2700 56413 2746
rect 56459 2700 56529 2746
rect 56575 2700 56586 2746
rect 50834 2630 56586 2700
rect 50834 2584 50845 2630
rect 50891 2584 50961 2630
rect 51007 2584 51077 2630
rect 51123 2584 51193 2630
rect 51239 2584 51309 2630
rect 51355 2584 51425 2630
rect 51471 2584 51541 2630
rect 51587 2584 51657 2630
rect 51703 2584 51773 2630
rect 51819 2584 51889 2630
rect 51935 2584 52005 2630
rect 52051 2584 52121 2630
rect 52167 2584 52237 2630
rect 52283 2584 52353 2630
rect 52399 2584 52469 2630
rect 52515 2584 52585 2630
rect 52631 2584 52701 2630
rect 52747 2584 52817 2630
rect 52863 2584 52933 2630
rect 52979 2584 53049 2630
rect 53095 2584 53165 2630
rect 53211 2584 53281 2630
rect 53327 2584 53397 2630
rect 53443 2584 53513 2630
rect 53559 2584 53629 2630
rect 53675 2584 53745 2630
rect 53791 2584 53861 2630
rect 53907 2584 53977 2630
rect 54023 2584 54093 2630
rect 54139 2584 54209 2630
rect 54255 2584 54325 2630
rect 54371 2584 54441 2630
rect 54487 2584 54557 2630
rect 54603 2584 54673 2630
rect 54719 2584 54789 2630
rect 54835 2584 54905 2630
rect 54951 2584 55021 2630
rect 55067 2584 55137 2630
rect 55183 2584 55253 2630
rect 55299 2584 55369 2630
rect 55415 2584 55485 2630
rect 55531 2584 55601 2630
rect 55647 2584 55717 2630
rect 55763 2584 55833 2630
rect 55879 2584 55949 2630
rect 55995 2584 56065 2630
rect 56111 2584 56181 2630
rect 56227 2584 56297 2630
rect 56343 2584 56413 2630
rect 56459 2584 56529 2630
rect 56575 2584 56586 2630
rect 50834 2514 56586 2584
rect 50834 2468 50845 2514
rect 50891 2468 50961 2514
rect 51007 2468 51077 2514
rect 51123 2468 51193 2514
rect 51239 2468 51309 2514
rect 51355 2468 51425 2514
rect 51471 2468 51541 2514
rect 51587 2468 51657 2514
rect 51703 2468 51773 2514
rect 51819 2468 51889 2514
rect 51935 2468 52005 2514
rect 52051 2468 52121 2514
rect 52167 2468 52237 2514
rect 52283 2468 52353 2514
rect 52399 2468 52469 2514
rect 52515 2468 52585 2514
rect 52631 2468 52701 2514
rect 52747 2468 52817 2514
rect 52863 2468 52933 2514
rect 52979 2468 53049 2514
rect 53095 2468 53165 2514
rect 53211 2468 53281 2514
rect 53327 2468 53397 2514
rect 53443 2468 53513 2514
rect 53559 2468 53629 2514
rect 53675 2468 53745 2514
rect 53791 2468 53861 2514
rect 53907 2468 53977 2514
rect 54023 2468 54093 2514
rect 54139 2468 54209 2514
rect 54255 2468 54325 2514
rect 54371 2468 54441 2514
rect 54487 2468 54557 2514
rect 54603 2468 54673 2514
rect 54719 2468 54789 2514
rect 54835 2468 54905 2514
rect 54951 2468 55021 2514
rect 55067 2468 55137 2514
rect 55183 2468 55253 2514
rect 55299 2468 55369 2514
rect 55415 2468 55485 2514
rect 55531 2468 55601 2514
rect 55647 2468 55717 2514
rect 55763 2468 55833 2514
rect 55879 2468 55949 2514
rect 55995 2468 56065 2514
rect 56111 2468 56181 2514
rect 56227 2468 56297 2514
rect 56343 2468 56413 2514
rect 56459 2468 56529 2514
rect 56575 2468 56586 2514
rect 50834 2398 56586 2468
rect 50834 2352 50845 2398
rect 50891 2352 50961 2398
rect 51007 2352 51077 2398
rect 51123 2352 51193 2398
rect 51239 2352 51309 2398
rect 51355 2352 51425 2398
rect 51471 2352 51541 2398
rect 51587 2352 51657 2398
rect 51703 2352 51773 2398
rect 51819 2352 51889 2398
rect 51935 2352 52005 2398
rect 52051 2352 52121 2398
rect 52167 2352 52237 2398
rect 52283 2352 52353 2398
rect 52399 2352 52469 2398
rect 52515 2352 52585 2398
rect 52631 2352 52701 2398
rect 52747 2352 52817 2398
rect 52863 2352 52933 2398
rect 52979 2352 53049 2398
rect 53095 2352 53165 2398
rect 53211 2352 53281 2398
rect 53327 2352 53397 2398
rect 53443 2352 53513 2398
rect 53559 2352 53629 2398
rect 53675 2352 53745 2398
rect 53791 2352 53861 2398
rect 53907 2352 53977 2398
rect 54023 2352 54093 2398
rect 54139 2352 54209 2398
rect 54255 2352 54325 2398
rect 54371 2352 54441 2398
rect 54487 2352 54557 2398
rect 54603 2352 54673 2398
rect 54719 2352 54789 2398
rect 54835 2352 54905 2398
rect 54951 2352 55021 2398
rect 55067 2352 55137 2398
rect 55183 2352 55253 2398
rect 55299 2352 55369 2398
rect 55415 2352 55485 2398
rect 55531 2352 55601 2398
rect 55647 2352 55717 2398
rect 55763 2352 55833 2398
rect 55879 2352 55949 2398
rect 55995 2352 56065 2398
rect 56111 2352 56181 2398
rect 56227 2352 56297 2398
rect 56343 2352 56413 2398
rect 56459 2352 56529 2398
rect 56575 2352 56586 2398
rect 50834 2282 56586 2352
rect 50834 2236 50845 2282
rect 50891 2236 50961 2282
rect 51007 2236 51077 2282
rect 51123 2236 51193 2282
rect 51239 2236 51309 2282
rect 51355 2236 51425 2282
rect 51471 2236 51541 2282
rect 51587 2236 51657 2282
rect 51703 2236 51773 2282
rect 51819 2236 51889 2282
rect 51935 2236 52005 2282
rect 52051 2236 52121 2282
rect 52167 2236 52237 2282
rect 52283 2236 52353 2282
rect 52399 2236 52469 2282
rect 52515 2236 52585 2282
rect 52631 2236 52701 2282
rect 52747 2236 52817 2282
rect 52863 2236 52933 2282
rect 52979 2236 53049 2282
rect 53095 2236 53165 2282
rect 53211 2236 53281 2282
rect 53327 2236 53397 2282
rect 53443 2236 53513 2282
rect 53559 2236 53629 2282
rect 53675 2236 53745 2282
rect 53791 2236 53861 2282
rect 53907 2236 53977 2282
rect 54023 2236 54093 2282
rect 54139 2236 54209 2282
rect 54255 2236 54325 2282
rect 54371 2236 54441 2282
rect 54487 2236 54557 2282
rect 54603 2236 54673 2282
rect 54719 2236 54789 2282
rect 54835 2236 54905 2282
rect 54951 2236 55021 2282
rect 55067 2236 55137 2282
rect 55183 2236 55253 2282
rect 55299 2236 55369 2282
rect 55415 2236 55485 2282
rect 55531 2236 55601 2282
rect 55647 2236 55717 2282
rect 55763 2236 55833 2282
rect 55879 2236 55949 2282
rect 55995 2236 56065 2282
rect 56111 2236 56181 2282
rect 56227 2236 56297 2282
rect 56343 2236 56413 2282
rect 56459 2236 56529 2282
rect 56575 2236 56586 2282
rect 50834 2166 56586 2236
rect 50834 2120 50845 2166
rect 50891 2120 50961 2166
rect 51007 2120 51077 2166
rect 51123 2120 51193 2166
rect 51239 2120 51309 2166
rect 51355 2120 51425 2166
rect 51471 2120 51541 2166
rect 51587 2120 51657 2166
rect 51703 2120 51773 2166
rect 51819 2120 51889 2166
rect 51935 2120 52005 2166
rect 52051 2120 52121 2166
rect 52167 2120 52237 2166
rect 52283 2120 52353 2166
rect 52399 2120 52469 2166
rect 52515 2120 52585 2166
rect 52631 2120 52701 2166
rect 52747 2120 52817 2166
rect 52863 2120 52933 2166
rect 52979 2120 53049 2166
rect 53095 2120 53165 2166
rect 53211 2120 53281 2166
rect 53327 2120 53397 2166
rect 53443 2120 53513 2166
rect 53559 2120 53629 2166
rect 53675 2120 53745 2166
rect 53791 2120 53861 2166
rect 53907 2120 53977 2166
rect 54023 2120 54093 2166
rect 54139 2120 54209 2166
rect 54255 2120 54325 2166
rect 54371 2120 54441 2166
rect 54487 2120 54557 2166
rect 54603 2120 54673 2166
rect 54719 2120 54789 2166
rect 54835 2120 54905 2166
rect 54951 2120 55021 2166
rect 55067 2120 55137 2166
rect 55183 2120 55253 2166
rect 55299 2120 55369 2166
rect 55415 2120 55485 2166
rect 55531 2120 55601 2166
rect 55647 2120 55717 2166
rect 55763 2120 55833 2166
rect 55879 2120 55949 2166
rect 55995 2120 56065 2166
rect 56111 2120 56181 2166
rect 56227 2120 56297 2166
rect 56343 2120 56413 2166
rect 56459 2120 56529 2166
rect 56575 2120 56586 2166
rect 50834 2050 56586 2120
rect 50834 2004 50845 2050
rect 50891 2004 50961 2050
rect 51007 2004 51077 2050
rect 51123 2004 51193 2050
rect 51239 2004 51309 2050
rect 51355 2004 51425 2050
rect 51471 2004 51541 2050
rect 51587 2004 51657 2050
rect 51703 2004 51773 2050
rect 51819 2004 51889 2050
rect 51935 2004 52005 2050
rect 52051 2004 52121 2050
rect 52167 2004 52237 2050
rect 52283 2004 52353 2050
rect 52399 2004 52469 2050
rect 52515 2004 52585 2050
rect 52631 2004 52701 2050
rect 52747 2004 52817 2050
rect 52863 2004 52933 2050
rect 52979 2004 53049 2050
rect 53095 2004 53165 2050
rect 53211 2004 53281 2050
rect 53327 2004 53397 2050
rect 53443 2004 53513 2050
rect 53559 2004 53629 2050
rect 53675 2004 53745 2050
rect 53791 2004 53861 2050
rect 53907 2004 53977 2050
rect 54023 2004 54093 2050
rect 54139 2004 54209 2050
rect 54255 2004 54325 2050
rect 54371 2004 54441 2050
rect 54487 2004 54557 2050
rect 54603 2004 54673 2050
rect 54719 2004 54789 2050
rect 54835 2004 54905 2050
rect 54951 2004 55021 2050
rect 55067 2004 55137 2050
rect 55183 2004 55253 2050
rect 55299 2004 55369 2050
rect 55415 2004 55485 2050
rect 55531 2004 55601 2050
rect 55647 2004 55717 2050
rect 55763 2004 55833 2050
rect 55879 2004 55949 2050
rect 55995 2004 56065 2050
rect 56111 2004 56181 2050
rect 56227 2004 56297 2050
rect 56343 2004 56413 2050
rect 56459 2004 56529 2050
rect 56575 2004 56586 2050
rect 50834 1934 56586 2004
rect 50834 1925 50845 1934
rect 40169 1888 50845 1925
rect 50891 1888 50961 1934
rect 51007 1888 51077 1934
rect 51123 1888 51193 1934
rect 51239 1888 51309 1934
rect 51355 1888 51425 1934
rect 51471 1888 51541 1934
rect 51587 1888 51657 1934
rect 51703 1888 51773 1934
rect 51819 1888 51889 1934
rect 51935 1888 52005 1934
rect 52051 1888 52121 1934
rect 52167 1888 52237 1934
rect 52283 1888 52353 1934
rect 52399 1888 52469 1934
rect 52515 1888 52585 1934
rect 52631 1888 52701 1934
rect 52747 1888 52817 1934
rect 52863 1888 52933 1934
rect 52979 1888 53049 1934
rect 53095 1888 53165 1934
rect 53211 1888 53281 1934
rect 53327 1888 53397 1934
rect 53443 1888 53513 1934
rect 53559 1888 53629 1934
rect 53675 1888 53745 1934
rect 53791 1888 53861 1934
rect 53907 1888 53977 1934
rect 54023 1888 54093 1934
rect 54139 1888 54209 1934
rect 54255 1888 54325 1934
rect 54371 1888 54441 1934
rect 54487 1888 54557 1934
rect 54603 1888 54673 1934
rect 54719 1888 54789 1934
rect 54835 1888 54905 1934
rect 54951 1888 55021 1934
rect 55067 1888 55137 1934
rect 55183 1888 55253 1934
rect 55299 1888 55369 1934
rect 55415 1888 55485 1934
rect 55531 1888 55601 1934
rect 55647 1888 55717 1934
rect 55763 1888 55833 1934
rect 55879 1888 55949 1934
rect 55995 1888 56065 1934
rect 56111 1888 56181 1934
rect 56227 1888 56297 1934
rect 56343 1888 56413 1934
rect 56459 1888 56529 1934
rect 56575 1925 56586 1934
rect 57295 1925 57306 34163
rect 56575 1888 57306 1925
rect 27744 1818 57306 1888
rect 27744 1772 28639 1818
rect 28685 1772 28755 1818
rect 28801 1772 28871 1818
rect 28917 1772 28987 1818
rect 29033 1772 29103 1818
rect 29149 1772 29219 1818
rect 29265 1772 29335 1818
rect 29381 1772 29451 1818
rect 29497 1772 29567 1818
rect 29613 1772 29683 1818
rect 29729 1772 29799 1818
rect 29845 1772 29915 1818
rect 29961 1772 30031 1818
rect 30077 1772 30147 1818
rect 30193 1772 30263 1818
rect 30309 1772 30379 1818
rect 30425 1772 30495 1818
rect 30541 1772 30611 1818
rect 30657 1772 30727 1818
rect 30773 1772 30843 1818
rect 30889 1772 30959 1818
rect 31005 1772 31075 1818
rect 31121 1772 31191 1818
rect 31237 1772 31307 1818
rect 31353 1772 31423 1818
rect 31469 1772 31539 1818
rect 31585 1772 31655 1818
rect 31701 1772 31771 1818
rect 31817 1772 31887 1818
rect 31933 1772 32003 1818
rect 32049 1772 32119 1818
rect 32165 1772 32235 1818
rect 32281 1772 32351 1818
rect 32397 1772 32467 1818
rect 32513 1772 32583 1818
rect 32629 1772 32699 1818
rect 32745 1772 32815 1818
rect 32861 1772 32931 1818
rect 32977 1772 33047 1818
rect 33093 1772 33163 1818
rect 33209 1772 33279 1818
rect 33325 1772 33395 1818
rect 33441 1772 33511 1818
rect 33557 1772 33627 1818
rect 33673 1772 33743 1818
rect 33789 1772 33859 1818
rect 33905 1772 33975 1818
rect 34021 1772 34091 1818
rect 34137 1772 34207 1818
rect 34253 1772 34323 1818
rect 34369 1772 34439 1818
rect 34485 1772 34555 1818
rect 34601 1772 34671 1818
rect 34717 1772 34787 1818
rect 34833 1772 34903 1818
rect 34949 1772 35019 1818
rect 35065 1772 35135 1818
rect 35181 1772 35251 1818
rect 35297 1772 35367 1818
rect 35413 1772 35483 1818
rect 35529 1772 35599 1818
rect 35645 1772 35715 1818
rect 35761 1772 35831 1818
rect 35877 1772 35947 1818
rect 35993 1772 36063 1818
rect 36109 1772 36179 1818
rect 36225 1772 36295 1818
rect 36341 1772 36411 1818
rect 36457 1772 36527 1818
rect 36573 1772 36643 1818
rect 36689 1772 36759 1818
rect 36805 1772 36875 1818
rect 36921 1772 36991 1818
rect 37037 1772 37107 1818
rect 37153 1772 37223 1818
rect 37269 1772 37339 1818
rect 37385 1772 37455 1818
rect 37501 1772 37571 1818
rect 37617 1772 37687 1818
rect 37733 1772 37803 1818
rect 37849 1772 37919 1818
rect 37965 1772 38035 1818
rect 38081 1772 38151 1818
rect 38197 1772 38267 1818
rect 38313 1772 38383 1818
rect 38429 1772 38499 1818
rect 38545 1772 38615 1818
rect 38661 1772 38731 1818
rect 38777 1772 38847 1818
rect 38893 1772 38963 1818
rect 39009 1772 39079 1818
rect 39125 1772 39195 1818
rect 39241 1772 39311 1818
rect 39357 1772 39427 1818
rect 39473 1772 39543 1818
rect 39589 1772 39659 1818
rect 39705 1772 39775 1818
rect 39821 1772 39891 1818
rect 39937 1772 40007 1818
rect 40053 1772 40123 1818
rect 40169 1772 50845 1818
rect 50891 1772 50961 1818
rect 51007 1772 51077 1818
rect 51123 1772 51193 1818
rect 51239 1772 51309 1818
rect 51355 1772 51425 1818
rect 51471 1772 51541 1818
rect 51587 1772 51657 1818
rect 51703 1772 51773 1818
rect 51819 1772 51889 1818
rect 51935 1772 52005 1818
rect 52051 1772 52121 1818
rect 52167 1772 52237 1818
rect 52283 1772 52353 1818
rect 52399 1772 52469 1818
rect 52515 1772 52585 1818
rect 52631 1772 52701 1818
rect 52747 1772 52817 1818
rect 52863 1772 52933 1818
rect 52979 1772 53049 1818
rect 53095 1772 53165 1818
rect 53211 1772 53281 1818
rect 53327 1772 53397 1818
rect 53443 1772 53513 1818
rect 53559 1772 53629 1818
rect 53675 1772 53745 1818
rect 53791 1772 53861 1818
rect 53907 1772 53977 1818
rect 54023 1772 54093 1818
rect 54139 1772 54209 1818
rect 54255 1772 54325 1818
rect 54371 1772 54441 1818
rect 54487 1772 54557 1818
rect 54603 1772 54673 1818
rect 54719 1772 54789 1818
rect 54835 1772 54905 1818
rect 54951 1772 55021 1818
rect 55067 1772 55137 1818
rect 55183 1772 55253 1818
rect 55299 1772 55369 1818
rect 55415 1772 55485 1818
rect 55531 1772 55601 1818
rect 55647 1772 55717 1818
rect 55763 1772 55833 1818
rect 55879 1772 55949 1818
rect 55995 1772 56065 1818
rect 56111 1772 56181 1818
rect 56227 1772 56297 1818
rect 56343 1772 56413 1818
rect 56459 1772 56529 1818
rect 56575 1772 57306 1818
rect 27744 1702 57306 1772
rect 27744 1656 28639 1702
rect 28685 1656 28755 1702
rect 28801 1656 28871 1702
rect 28917 1656 28987 1702
rect 29033 1656 29103 1702
rect 29149 1656 29219 1702
rect 29265 1656 29335 1702
rect 29381 1656 29451 1702
rect 29497 1656 29567 1702
rect 29613 1656 29683 1702
rect 29729 1656 29799 1702
rect 29845 1656 29915 1702
rect 29961 1656 30031 1702
rect 30077 1656 30147 1702
rect 30193 1656 30263 1702
rect 30309 1656 30379 1702
rect 30425 1656 30495 1702
rect 30541 1656 30611 1702
rect 30657 1656 30727 1702
rect 30773 1656 30843 1702
rect 30889 1656 30959 1702
rect 31005 1656 31075 1702
rect 31121 1656 31191 1702
rect 31237 1656 31307 1702
rect 31353 1656 31423 1702
rect 31469 1656 31539 1702
rect 31585 1656 31655 1702
rect 31701 1656 31771 1702
rect 31817 1656 31887 1702
rect 31933 1656 32003 1702
rect 32049 1656 32119 1702
rect 32165 1656 32235 1702
rect 32281 1656 32351 1702
rect 32397 1656 32467 1702
rect 32513 1656 32583 1702
rect 32629 1656 32699 1702
rect 32745 1656 32815 1702
rect 32861 1656 32931 1702
rect 32977 1656 33047 1702
rect 33093 1656 33163 1702
rect 33209 1656 33279 1702
rect 33325 1656 33395 1702
rect 33441 1656 33511 1702
rect 33557 1656 33627 1702
rect 33673 1656 33743 1702
rect 33789 1656 33859 1702
rect 33905 1656 33975 1702
rect 34021 1656 34091 1702
rect 34137 1656 34207 1702
rect 34253 1656 34323 1702
rect 34369 1656 34439 1702
rect 34485 1656 34555 1702
rect 34601 1656 34671 1702
rect 34717 1656 34787 1702
rect 34833 1656 34903 1702
rect 34949 1656 35019 1702
rect 35065 1656 35135 1702
rect 35181 1656 35251 1702
rect 35297 1656 35367 1702
rect 35413 1656 35483 1702
rect 35529 1656 35599 1702
rect 35645 1656 35715 1702
rect 35761 1656 35831 1702
rect 35877 1656 35947 1702
rect 35993 1656 36063 1702
rect 36109 1656 36179 1702
rect 36225 1656 36295 1702
rect 36341 1656 36411 1702
rect 36457 1656 36527 1702
rect 36573 1656 36643 1702
rect 36689 1656 36759 1702
rect 36805 1656 36875 1702
rect 36921 1656 36991 1702
rect 37037 1656 37107 1702
rect 37153 1656 37223 1702
rect 37269 1656 37339 1702
rect 37385 1656 37455 1702
rect 37501 1656 37571 1702
rect 37617 1656 37687 1702
rect 37733 1656 37803 1702
rect 37849 1656 37919 1702
rect 37965 1656 38035 1702
rect 38081 1656 38151 1702
rect 38197 1656 38267 1702
rect 38313 1656 38383 1702
rect 38429 1656 38499 1702
rect 38545 1656 38615 1702
rect 38661 1656 38731 1702
rect 38777 1656 38847 1702
rect 38893 1656 38963 1702
rect 39009 1656 39079 1702
rect 39125 1656 39195 1702
rect 39241 1656 39311 1702
rect 39357 1656 39427 1702
rect 39473 1656 39543 1702
rect 39589 1656 39659 1702
rect 39705 1656 39775 1702
rect 39821 1656 39891 1702
rect 39937 1656 40007 1702
rect 40053 1656 40123 1702
rect 40169 1656 50845 1702
rect 50891 1656 50961 1702
rect 51007 1656 51077 1702
rect 51123 1656 51193 1702
rect 51239 1656 51309 1702
rect 51355 1656 51425 1702
rect 51471 1656 51541 1702
rect 51587 1656 51657 1702
rect 51703 1656 51773 1702
rect 51819 1656 51889 1702
rect 51935 1656 52005 1702
rect 52051 1656 52121 1702
rect 52167 1656 52237 1702
rect 52283 1656 52353 1702
rect 52399 1656 52469 1702
rect 52515 1656 52585 1702
rect 52631 1656 52701 1702
rect 52747 1656 52817 1702
rect 52863 1656 52933 1702
rect 52979 1656 53049 1702
rect 53095 1656 53165 1702
rect 53211 1656 53281 1702
rect 53327 1656 53397 1702
rect 53443 1656 53513 1702
rect 53559 1656 53629 1702
rect 53675 1656 53745 1702
rect 53791 1656 53861 1702
rect 53907 1656 53977 1702
rect 54023 1656 54093 1702
rect 54139 1656 54209 1702
rect 54255 1656 54325 1702
rect 54371 1656 54441 1702
rect 54487 1656 54557 1702
rect 54603 1656 54673 1702
rect 54719 1656 54789 1702
rect 54835 1656 54905 1702
rect 54951 1656 55021 1702
rect 55067 1656 55137 1702
rect 55183 1656 55253 1702
rect 55299 1656 55369 1702
rect 55415 1656 55485 1702
rect 55531 1656 55601 1702
rect 55647 1656 55717 1702
rect 55763 1656 55833 1702
rect 55879 1656 55949 1702
rect 55995 1656 56065 1702
rect 56111 1656 56181 1702
rect 56227 1656 56297 1702
rect 56343 1656 56413 1702
rect 56459 1656 56529 1702
rect 56575 1656 57306 1702
rect 27744 1117 57306 1656
rect 57652 3584 57736 95694
rect 58791 94773 59518 95694
rect 58791 94721 58867 94773
rect 58919 94721 58991 94773
rect 59043 94721 59115 94773
rect 59167 94721 59239 94773
rect 59291 94721 59363 94773
rect 59415 94721 59518 94773
rect 58791 94649 59518 94721
rect 58791 94597 58867 94649
rect 58919 94597 58991 94649
rect 59043 94597 59115 94649
rect 59167 94597 59239 94649
rect 59291 94597 59363 94649
rect 59415 94597 59518 94649
rect 58791 94525 59518 94597
rect 58791 94473 58867 94525
rect 58919 94473 58991 94525
rect 59043 94473 59115 94525
rect 59167 94473 59239 94525
rect 59291 94473 59363 94525
rect 59415 94473 59518 94525
rect 58791 94454 59518 94473
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 85090 35484 85733 95694
rect 84242 35364 85733 35484
rect 60563 35326 60639 35338
rect 57909 33432 58351 33519
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33215 58351 33380
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 32997 58351 33163
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32779 58351 32945
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32562 58351 32727
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32344 58351 32510
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32075 57998 32127
rect 58050 32075 58210 32127
rect 58262 32075 58351 32127
rect 57909 31909 58351 32075
rect 83398 32048 83834 32122
rect 57909 31857 57998 31909
rect 58050 31857 58210 31909
rect 58262 31857 58351 31909
rect 57909 31691 58351 31857
rect 57909 31639 57998 31691
rect 58050 31639 58210 31691
rect 58262 31639 58351 31691
rect 57909 31474 58351 31639
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29950 58351 30116
rect 57909 29898 57998 29950
rect 58050 29898 58210 29950
rect 58262 29898 58351 29950
rect 57909 29733 58351 29898
rect 57909 29681 57998 29733
rect 58050 29681 58210 29733
rect 58262 29681 58351 29733
rect 57909 29515 58351 29681
rect 57909 29463 57998 29515
rect 58050 29463 58210 29515
rect 58262 29463 58351 29515
rect 57909 29297 58351 29463
rect 57909 29245 57998 29297
rect 58050 29245 58210 29297
rect 58262 29245 58351 29297
rect 57909 29080 58351 29245
rect 57909 29028 57998 29080
rect 58050 29028 58210 29080
rect 58262 29028 58351 29080
rect 57909 28862 58351 29028
rect 57909 28810 57998 28862
rect 58050 28810 58210 28862
rect 58262 28810 58351 28862
rect 57909 28644 58351 28810
rect 57909 28592 57998 28644
rect 58050 28592 58210 28644
rect 58262 28592 58351 28644
rect 57909 28427 58351 28592
rect 57909 28375 57998 28427
rect 58050 28375 58210 28427
rect 58262 28375 58351 28427
rect 57909 28209 58351 28375
rect 57909 28157 57998 28209
rect 58050 28157 58210 28209
rect 58262 28157 58351 28209
rect 57909 27992 58351 28157
rect 57909 27940 57998 27992
rect 58050 27940 58210 27992
rect 58262 27940 58351 27992
rect 57909 27774 58351 27940
rect 57909 27722 57998 27774
rect 58050 27722 58210 27774
rect 58262 27722 58351 27774
rect 57909 27556 58351 27722
rect 57909 27504 57998 27556
rect 58050 27504 58210 27556
rect 58262 27504 58351 27556
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24074 58351 24240
rect 57909 24022 57998 24074
rect 58050 24022 58210 24074
rect 58262 24022 58351 24074
rect 57909 23857 58351 24022
rect 57909 23805 57998 23857
rect 58050 23805 58210 23857
rect 58262 23805 58351 23857
rect 57909 23639 58351 23805
rect 57909 23587 57998 23639
rect 58050 23587 58210 23639
rect 58262 23587 58351 23639
rect 57909 23421 58351 23587
rect 57909 23369 57998 23421
rect 58050 23369 58210 23421
rect 58262 23369 58351 23421
rect 57909 23204 58351 23369
rect 57909 23152 57998 23204
rect 58050 23152 58210 23204
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20540 58210 20592
rect 58262 20540 58351 20592
rect 57909 20374 58351 20540
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20157 58351 20322
rect 57909 20105 57998 20157
rect 58050 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 19939 58351 20105
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13628 58351 13793
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13410 58351 13576
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13192 58351 13358
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 12975 58351 13140
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12757 58351 12923
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12540 58351 12705
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12322 58351 12488
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12104 58351 12270
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 11887 58351 12052
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11669 58351 11835
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9275 58351 9441
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9057 58351 9223
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8840 58351 9005
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8622 58351 8788
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8404 58351 8570
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8187 58351 8352
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5523 57998 5575
rect 58050 5523 58210 5575
rect 58262 5523 58351 5575
rect 57909 5358 58351 5523
rect 57909 5306 57998 5358
rect 58050 5306 58210 5358
rect 58262 5306 58351 5358
rect 57909 4587 58351 5306
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4370 58351 4535
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4152 58351 4318
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57652 1282 57737 3584
rect 57909 1777 58351 3665
rect 62138 1689 62318 1701
rect 62138 1637 62150 1689
rect 62306 1637 62318 1689
rect 62138 1625 62318 1637
rect 72203 1689 72383 1701
rect 72203 1637 72215 1689
rect 72371 1637 72383 1689
rect 72203 1625 72383 1637
rect 72653 1689 72833 1701
rect 72653 1637 72665 1689
rect 72821 1637 72833 1689
rect 72653 1625 72833 1637
rect 82718 1689 82898 1701
rect 82718 1637 82730 1689
rect 82886 1637 82898 1689
rect 82718 1625 82898 1637
rect 85090 1282 85733 35364
rect 57652 1117 85733 1282
rect 86079 1117 86090 96163
rect 282 1015 86090 1117
rect 282 969 371 1015
rect 417 969 495 1015
rect 541 969 619 1015
rect 665 969 743 1015
rect 789 969 867 1015
rect 913 969 991 1015
rect 1037 969 1115 1015
rect 1161 969 1239 1015
rect 1285 969 1363 1015
rect 1409 969 1487 1015
rect 1533 969 1611 1015
rect 1657 969 1735 1015
rect 1781 969 1859 1015
rect 1905 969 1983 1015
rect 2029 969 2107 1015
rect 2153 969 2231 1015
rect 2277 969 2355 1015
rect 2401 969 2479 1015
rect 2525 969 2603 1015
rect 2649 969 2727 1015
rect 2773 969 2851 1015
rect 2897 969 2975 1015
rect 3021 969 3099 1015
rect 3145 969 3223 1015
rect 3269 969 3347 1015
rect 3393 969 3471 1015
rect 3517 969 3595 1015
rect 3641 969 3719 1015
rect 3765 969 3843 1015
rect 3889 969 3967 1015
rect 4013 969 4091 1015
rect 4137 969 4215 1015
rect 4261 969 4339 1015
rect 4385 969 4463 1015
rect 4509 969 4587 1015
rect 4633 969 4711 1015
rect 4757 969 4835 1015
rect 4881 969 4959 1015
rect 5005 969 5083 1015
rect 5129 969 5207 1015
rect 5253 969 5331 1015
rect 5377 969 5455 1015
rect 5501 969 5579 1015
rect 5625 969 5703 1015
rect 5749 969 5827 1015
rect 5873 969 5951 1015
rect 5997 969 6075 1015
rect 6121 969 6199 1015
rect 6245 969 6323 1015
rect 6369 969 6447 1015
rect 6493 969 6571 1015
rect 6617 969 6695 1015
rect 6741 969 6819 1015
rect 6865 969 6943 1015
rect 6989 969 7067 1015
rect 7113 969 7191 1015
rect 7237 969 7315 1015
rect 7361 969 7439 1015
rect 7485 969 7563 1015
rect 7609 969 7687 1015
rect 7733 969 7811 1015
rect 7857 969 7935 1015
rect 7981 969 8059 1015
rect 8105 969 8183 1015
rect 8229 969 8307 1015
rect 8353 969 8431 1015
rect 8477 969 8555 1015
rect 8601 969 8679 1015
rect 8725 969 8803 1015
rect 8849 969 8927 1015
rect 8973 969 9051 1015
rect 9097 969 9175 1015
rect 9221 969 9299 1015
rect 9345 969 9423 1015
rect 9469 969 9547 1015
rect 9593 969 9671 1015
rect 9717 969 9795 1015
rect 9841 969 9919 1015
rect 9965 969 10043 1015
rect 10089 969 10167 1015
rect 10213 969 10291 1015
rect 10337 969 10415 1015
rect 10461 969 10539 1015
rect 10585 969 10663 1015
rect 10709 969 10787 1015
rect 10833 969 10911 1015
rect 10957 969 11035 1015
rect 11081 969 11159 1015
rect 11205 969 11283 1015
rect 11329 969 11407 1015
rect 11453 969 11531 1015
rect 11577 969 11655 1015
rect 11701 969 11779 1015
rect 11825 969 11903 1015
rect 11949 969 12027 1015
rect 12073 969 12151 1015
rect 12197 969 12275 1015
rect 12321 969 12399 1015
rect 12445 969 12523 1015
rect 12569 969 12647 1015
rect 12693 969 12771 1015
rect 12817 969 12895 1015
rect 12941 969 13019 1015
rect 13065 969 13143 1015
rect 13189 969 13267 1015
rect 13313 969 13391 1015
rect 13437 969 13515 1015
rect 13561 969 13639 1015
rect 13685 969 13763 1015
rect 13809 969 13887 1015
rect 13933 969 14011 1015
rect 14057 969 14135 1015
rect 14181 969 14259 1015
rect 14305 969 14383 1015
rect 14429 969 14507 1015
rect 14553 969 14631 1015
rect 14677 969 14755 1015
rect 14801 969 14879 1015
rect 14925 969 15003 1015
rect 15049 969 15127 1015
rect 15173 969 15251 1015
rect 15297 969 15375 1015
rect 15421 969 15499 1015
rect 15545 969 15623 1015
rect 15669 969 15747 1015
rect 15793 969 15871 1015
rect 15917 969 15995 1015
rect 16041 969 16119 1015
rect 16165 969 16243 1015
rect 16289 969 16367 1015
rect 16413 969 16491 1015
rect 16537 969 16615 1015
rect 16661 969 16739 1015
rect 16785 969 16863 1015
rect 16909 969 16987 1015
rect 17033 969 17111 1015
rect 17157 969 17235 1015
rect 17281 969 17359 1015
rect 17405 969 17483 1015
rect 17529 969 17607 1015
rect 17653 969 17731 1015
rect 17777 969 17855 1015
rect 17901 969 17979 1015
rect 18025 969 18103 1015
rect 18149 969 18227 1015
rect 18273 969 18351 1015
rect 18397 969 18475 1015
rect 18521 969 18599 1015
rect 18645 969 18723 1015
rect 18769 969 18847 1015
rect 18893 969 18971 1015
rect 19017 969 19095 1015
rect 19141 969 19219 1015
rect 19265 969 19343 1015
rect 19389 969 19467 1015
rect 19513 969 19591 1015
rect 19637 969 19715 1015
rect 19761 969 19839 1015
rect 19885 969 19963 1015
rect 20009 969 20087 1015
rect 20133 969 20211 1015
rect 20257 969 20335 1015
rect 20381 969 20459 1015
rect 20505 969 20583 1015
rect 20629 969 20707 1015
rect 20753 969 20831 1015
rect 20877 969 20955 1015
rect 21001 969 21079 1015
rect 21125 969 21203 1015
rect 21249 969 21327 1015
rect 21373 969 21451 1015
rect 21497 969 21575 1015
rect 21621 969 21699 1015
rect 21745 969 21823 1015
rect 21869 969 21947 1015
rect 21993 969 22071 1015
rect 22117 969 22195 1015
rect 22241 969 22319 1015
rect 22365 969 22443 1015
rect 22489 969 22567 1015
rect 22613 969 22691 1015
rect 22737 969 22815 1015
rect 22861 969 22939 1015
rect 22985 969 23063 1015
rect 23109 969 23187 1015
rect 23233 969 23311 1015
rect 23357 969 23435 1015
rect 23481 969 23559 1015
rect 23605 969 23683 1015
rect 23729 969 23807 1015
rect 23853 969 23931 1015
rect 23977 969 24055 1015
rect 24101 969 24179 1015
rect 24225 969 24303 1015
rect 24349 969 24427 1015
rect 24473 969 24551 1015
rect 24597 969 24675 1015
rect 24721 969 24799 1015
rect 24845 969 24923 1015
rect 24969 969 25047 1015
rect 25093 969 25171 1015
rect 25217 969 25295 1015
rect 25341 969 25419 1015
rect 25465 969 25543 1015
rect 25589 969 25667 1015
rect 25713 969 25791 1015
rect 25837 969 25915 1015
rect 25961 969 26039 1015
rect 26085 969 26163 1015
rect 26209 969 26287 1015
rect 26333 969 26411 1015
rect 26457 969 26535 1015
rect 26581 969 26659 1015
rect 26705 969 26783 1015
rect 26829 969 26907 1015
rect 26953 969 27031 1015
rect 27077 969 27155 1015
rect 27201 969 27279 1015
rect 27325 969 27403 1015
rect 27449 969 27527 1015
rect 27573 969 27651 1015
rect 27697 969 27775 1015
rect 27821 969 27899 1015
rect 27945 969 28023 1015
rect 28069 969 28147 1015
rect 28193 969 28271 1015
rect 28317 969 28395 1015
rect 28441 969 28519 1015
rect 28565 969 28643 1015
rect 28689 969 28767 1015
rect 28813 969 28891 1015
rect 28937 969 29015 1015
rect 29061 969 29139 1015
rect 29185 969 29263 1015
rect 29309 969 29387 1015
rect 29433 969 29511 1015
rect 29557 969 29635 1015
rect 29681 969 29759 1015
rect 29805 969 29883 1015
rect 29929 969 30007 1015
rect 30053 969 30131 1015
rect 30177 969 30255 1015
rect 30301 969 30379 1015
rect 30425 969 30503 1015
rect 30549 969 30627 1015
rect 30673 969 30751 1015
rect 30797 969 30875 1015
rect 30921 969 30999 1015
rect 31045 969 31123 1015
rect 31169 969 31247 1015
rect 31293 969 31371 1015
rect 31417 969 31495 1015
rect 31541 969 31619 1015
rect 31665 969 31743 1015
rect 31789 969 31867 1015
rect 31913 969 31991 1015
rect 32037 969 32115 1015
rect 32161 969 32239 1015
rect 32285 969 32363 1015
rect 32409 969 32487 1015
rect 32533 969 32611 1015
rect 32657 969 32735 1015
rect 32781 969 32859 1015
rect 32905 969 32983 1015
rect 33029 969 33107 1015
rect 33153 969 33231 1015
rect 33277 969 33355 1015
rect 33401 969 33479 1015
rect 33525 969 33603 1015
rect 33649 969 33727 1015
rect 33773 969 33851 1015
rect 33897 969 33975 1015
rect 34021 969 34099 1015
rect 34145 969 34223 1015
rect 34269 969 34347 1015
rect 34393 969 34471 1015
rect 34517 969 34595 1015
rect 34641 969 34719 1015
rect 34765 969 34843 1015
rect 34889 969 34967 1015
rect 35013 969 35091 1015
rect 35137 969 35215 1015
rect 35261 969 35339 1015
rect 35385 969 35463 1015
rect 35509 969 35587 1015
rect 35633 969 35711 1015
rect 35757 969 35835 1015
rect 35881 969 35959 1015
rect 36005 969 36083 1015
rect 36129 969 36207 1015
rect 36253 969 36331 1015
rect 36377 969 36455 1015
rect 36501 969 36579 1015
rect 36625 969 36703 1015
rect 36749 969 36827 1015
rect 36873 969 36951 1015
rect 36997 969 37075 1015
rect 37121 969 37199 1015
rect 37245 969 37323 1015
rect 37369 969 37447 1015
rect 37493 969 37571 1015
rect 37617 969 37695 1015
rect 37741 969 37819 1015
rect 37865 969 37943 1015
rect 37989 969 38067 1015
rect 38113 969 38191 1015
rect 38237 969 38315 1015
rect 38361 969 38439 1015
rect 38485 969 38563 1015
rect 38609 969 38687 1015
rect 38733 969 38811 1015
rect 38857 969 38935 1015
rect 38981 969 39059 1015
rect 39105 969 39183 1015
rect 39229 969 39307 1015
rect 39353 969 39431 1015
rect 39477 969 39555 1015
rect 39601 969 39679 1015
rect 39725 969 39803 1015
rect 39849 969 39927 1015
rect 39973 969 40051 1015
rect 40097 969 40175 1015
rect 40221 969 40299 1015
rect 40345 969 40423 1015
rect 40469 969 40547 1015
rect 40593 969 40671 1015
rect 40717 969 40795 1015
rect 40841 969 40919 1015
rect 40965 969 41043 1015
rect 41089 969 41167 1015
rect 41213 969 41291 1015
rect 41337 969 41415 1015
rect 41461 969 41539 1015
rect 41585 969 41663 1015
rect 41709 969 41787 1015
rect 41833 969 41911 1015
rect 41957 969 42035 1015
rect 42081 969 42159 1015
rect 42205 969 42283 1015
rect 42329 969 42407 1015
rect 42453 969 42531 1015
rect 42577 969 42655 1015
rect 42701 969 42779 1015
rect 42825 969 42903 1015
rect 42949 969 43027 1015
rect 43073 969 43151 1015
rect 43197 969 43275 1015
rect 43321 969 43399 1015
rect 43445 969 43523 1015
rect 43569 969 43647 1015
rect 43693 969 43771 1015
rect 43817 969 43895 1015
rect 43941 969 44019 1015
rect 44065 969 44143 1015
rect 44189 969 44267 1015
rect 44313 969 44391 1015
rect 44437 969 44515 1015
rect 44561 969 44639 1015
rect 44685 969 44763 1015
rect 44809 969 44887 1015
rect 44933 969 45011 1015
rect 45057 969 45135 1015
rect 45181 969 45259 1015
rect 45305 969 45383 1015
rect 45429 969 45507 1015
rect 45553 969 45631 1015
rect 45677 969 45755 1015
rect 45801 969 45879 1015
rect 45925 969 46003 1015
rect 46049 969 46127 1015
rect 46173 969 46251 1015
rect 46297 969 46375 1015
rect 46421 969 46499 1015
rect 46545 969 46623 1015
rect 46669 969 46747 1015
rect 46793 969 46871 1015
rect 46917 969 46995 1015
rect 47041 969 47119 1015
rect 47165 969 47243 1015
rect 47289 969 47367 1015
rect 47413 969 47491 1015
rect 47537 969 47615 1015
rect 47661 969 47739 1015
rect 47785 969 47863 1015
rect 47909 969 47987 1015
rect 48033 969 48111 1015
rect 48157 969 48235 1015
rect 48281 969 48359 1015
rect 48405 969 48483 1015
rect 48529 969 48607 1015
rect 48653 969 48731 1015
rect 48777 969 48855 1015
rect 48901 969 48979 1015
rect 49025 969 49103 1015
rect 49149 969 49227 1015
rect 49273 969 49351 1015
rect 49397 969 49475 1015
rect 49521 969 49599 1015
rect 49645 969 49723 1015
rect 49769 969 49847 1015
rect 49893 969 49971 1015
rect 50017 969 50095 1015
rect 50141 969 50219 1015
rect 50265 969 50343 1015
rect 50389 969 50467 1015
rect 50513 969 50591 1015
rect 50637 969 50715 1015
rect 50761 969 50839 1015
rect 50885 969 50963 1015
rect 51009 969 51087 1015
rect 51133 969 51211 1015
rect 51257 969 51335 1015
rect 51381 969 51459 1015
rect 51505 969 51583 1015
rect 51629 969 51707 1015
rect 51753 969 51831 1015
rect 51877 969 51955 1015
rect 52001 969 52079 1015
rect 52125 969 52203 1015
rect 52249 969 52327 1015
rect 52373 969 52451 1015
rect 52497 969 52575 1015
rect 52621 969 52699 1015
rect 52745 969 52823 1015
rect 52869 969 52947 1015
rect 52993 969 53071 1015
rect 53117 969 53195 1015
rect 53241 969 53319 1015
rect 53365 969 53443 1015
rect 53489 969 53567 1015
rect 53613 969 53691 1015
rect 53737 969 53815 1015
rect 53861 969 53939 1015
rect 53985 969 54063 1015
rect 54109 969 54187 1015
rect 54233 969 54311 1015
rect 54357 969 54435 1015
rect 54481 969 54559 1015
rect 54605 969 54683 1015
rect 54729 969 54807 1015
rect 54853 969 54931 1015
rect 54977 969 55055 1015
rect 55101 969 55179 1015
rect 55225 969 55303 1015
rect 55349 969 55427 1015
rect 55473 969 55551 1015
rect 55597 969 55675 1015
rect 55721 969 55799 1015
rect 55845 969 55923 1015
rect 55969 969 56047 1015
rect 56093 969 56171 1015
rect 56217 969 56295 1015
rect 56341 969 56419 1015
rect 56465 969 56543 1015
rect 56589 969 56667 1015
rect 56713 969 56791 1015
rect 56837 969 56915 1015
rect 56961 969 57039 1015
rect 57085 969 57163 1015
rect 57209 969 57287 1015
rect 57333 969 57411 1015
rect 57457 969 57535 1015
rect 57581 969 57659 1015
rect 57705 969 57783 1015
rect 57829 969 57907 1015
rect 57953 969 58031 1015
rect 58077 969 58155 1015
rect 58201 969 58279 1015
rect 58325 969 58403 1015
rect 58449 969 58527 1015
rect 58573 969 58651 1015
rect 58697 969 58775 1015
rect 58821 969 58899 1015
rect 58945 969 59023 1015
rect 59069 969 59147 1015
rect 59193 969 59271 1015
rect 59317 969 59395 1015
rect 59441 969 59519 1015
rect 59565 969 59643 1015
rect 59689 969 59767 1015
rect 59813 969 59891 1015
rect 59937 969 60015 1015
rect 60061 969 60139 1015
rect 60185 969 60263 1015
rect 60309 969 60387 1015
rect 60433 969 60511 1015
rect 60557 969 60635 1015
rect 60681 969 60759 1015
rect 60805 969 60883 1015
rect 60929 969 61007 1015
rect 61053 969 61131 1015
rect 61177 969 61255 1015
rect 61301 969 61379 1015
rect 61425 969 61503 1015
rect 61549 969 61627 1015
rect 61673 969 61751 1015
rect 61797 969 61875 1015
rect 61921 969 61999 1015
rect 62045 969 62123 1015
rect 62169 969 62247 1015
rect 62293 969 62371 1015
rect 62417 969 62495 1015
rect 62541 969 62619 1015
rect 62665 969 62743 1015
rect 62789 969 62867 1015
rect 62913 969 62991 1015
rect 63037 969 63115 1015
rect 63161 969 63239 1015
rect 63285 969 63363 1015
rect 63409 969 63487 1015
rect 63533 969 63611 1015
rect 63657 969 63735 1015
rect 63781 969 63859 1015
rect 63905 969 63983 1015
rect 64029 969 64107 1015
rect 64153 969 64231 1015
rect 64277 969 64355 1015
rect 64401 969 64479 1015
rect 64525 969 64603 1015
rect 64649 969 64727 1015
rect 64773 969 64851 1015
rect 64897 969 64975 1015
rect 65021 969 65099 1015
rect 65145 969 65223 1015
rect 65269 969 65347 1015
rect 65393 969 65471 1015
rect 65517 969 65595 1015
rect 65641 969 65719 1015
rect 65765 969 65843 1015
rect 65889 969 65967 1015
rect 66013 969 66091 1015
rect 66137 969 66215 1015
rect 66261 969 66339 1015
rect 66385 969 66463 1015
rect 66509 969 66587 1015
rect 66633 969 66711 1015
rect 66757 969 66835 1015
rect 66881 969 66959 1015
rect 67005 969 67083 1015
rect 67129 969 67207 1015
rect 67253 969 67331 1015
rect 67377 969 67455 1015
rect 67501 969 67579 1015
rect 67625 969 67703 1015
rect 67749 969 67827 1015
rect 67873 969 67951 1015
rect 67997 969 68075 1015
rect 68121 969 68199 1015
rect 68245 969 68323 1015
rect 68369 969 68447 1015
rect 68493 969 68571 1015
rect 68617 969 68695 1015
rect 68741 969 68819 1015
rect 68865 969 68943 1015
rect 68989 969 69067 1015
rect 69113 969 69191 1015
rect 69237 969 69315 1015
rect 69361 969 69439 1015
rect 69485 969 69563 1015
rect 69609 969 69687 1015
rect 69733 969 69811 1015
rect 69857 969 69935 1015
rect 69981 969 70059 1015
rect 70105 969 70183 1015
rect 70229 969 70307 1015
rect 70353 969 70431 1015
rect 70477 969 70555 1015
rect 70601 969 70679 1015
rect 70725 969 70803 1015
rect 70849 969 70927 1015
rect 70973 969 71051 1015
rect 71097 969 71175 1015
rect 71221 969 71299 1015
rect 71345 969 71423 1015
rect 71469 969 71547 1015
rect 71593 969 71671 1015
rect 71717 969 71795 1015
rect 71841 969 71919 1015
rect 71965 969 72043 1015
rect 72089 969 72167 1015
rect 72213 969 72291 1015
rect 72337 969 72415 1015
rect 72461 969 72539 1015
rect 72585 969 72663 1015
rect 72709 969 72787 1015
rect 72833 969 72911 1015
rect 72957 969 73035 1015
rect 73081 969 73159 1015
rect 73205 969 73283 1015
rect 73329 969 73407 1015
rect 73453 969 73531 1015
rect 73577 969 73655 1015
rect 73701 969 73779 1015
rect 73825 969 73903 1015
rect 73949 969 74027 1015
rect 74073 969 74151 1015
rect 74197 969 74275 1015
rect 74321 969 74399 1015
rect 74445 969 74523 1015
rect 74569 969 74647 1015
rect 74693 969 74771 1015
rect 74817 969 74895 1015
rect 74941 969 75019 1015
rect 75065 969 75143 1015
rect 75189 969 75267 1015
rect 75313 969 75391 1015
rect 75437 969 75515 1015
rect 75561 969 75639 1015
rect 75685 969 75763 1015
rect 75809 969 75887 1015
rect 75933 969 76011 1015
rect 76057 969 76135 1015
rect 76181 969 76259 1015
rect 76305 969 76383 1015
rect 76429 969 76507 1015
rect 76553 969 76631 1015
rect 76677 969 76755 1015
rect 76801 969 76879 1015
rect 76925 969 77003 1015
rect 77049 969 77127 1015
rect 77173 969 77251 1015
rect 77297 969 77375 1015
rect 77421 969 77499 1015
rect 77545 969 77623 1015
rect 77669 969 77747 1015
rect 77793 969 77871 1015
rect 77917 969 77995 1015
rect 78041 969 78119 1015
rect 78165 969 78243 1015
rect 78289 969 78367 1015
rect 78413 969 78491 1015
rect 78537 969 78615 1015
rect 78661 969 78739 1015
rect 78785 969 78863 1015
rect 78909 969 78987 1015
rect 79033 969 79111 1015
rect 79157 969 79235 1015
rect 79281 969 79359 1015
rect 79405 969 79483 1015
rect 79529 969 79607 1015
rect 79653 969 79731 1015
rect 79777 969 79855 1015
rect 79901 969 79979 1015
rect 80025 969 80103 1015
rect 80149 969 80227 1015
rect 80273 969 80351 1015
rect 80397 969 80475 1015
rect 80521 969 80599 1015
rect 80645 969 80723 1015
rect 80769 969 80847 1015
rect 80893 969 80971 1015
rect 81017 969 81095 1015
rect 81141 969 81219 1015
rect 81265 969 81343 1015
rect 81389 969 81467 1015
rect 81513 969 81591 1015
rect 81637 969 81715 1015
rect 81761 969 81839 1015
rect 81885 969 81963 1015
rect 82009 969 82087 1015
rect 82133 969 82211 1015
rect 82257 969 82335 1015
rect 82381 969 82459 1015
rect 82505 969 82583 1015
rect 82629 969 82707 1015
rect 82753 969 82831 1015
rect 82877 969 82955 1015
rect 83001 969 83079 1015
rect 83125 969 83203 1015
rect 83249 969 83327 1015
rect 83373 969 83451 1015
rect 83497 969 83575 1015
rect 83621 969 83699 1015
rect 83745 969 83823 1015
rect 83869 969 83947 1015
rect 83993 969 84071 1015
rect 84117 969 84195 1015
rect 84241 969 84319 1015
rect 84365 969 84443 1015
rect 84489 969 84567 1015
rect 84613 969 84691 1015
rect 84737 969 84815 1015
rect 84861 969 84939 1015
rect 84985 969 85063 1015
rect 85109 969 85187 1015
rect 85233 969 85311 1015
rect 85357 969 85435 1015
rect 85481 969 85559 1015
rect 85605 969 85683 1015
rect 85729 969 85807 1015
rect 85853 969 85931 1015
rect 85977 969 86090 1015
rect 282 891 86090 969
rect 282 845 371 891
rect 417 845 495 891
rect 541 845 619 891
rect 665 845 743 891
rect 789 845 867 891
rect 913 845 991 891
rect 1037 845 1115 891
rect 1161 845 1239 891
rect 1285 845 1363 891
rect 1409 845 1487 891
rect 1533 845 1611 891
rect 1657 845 1735 891
rect 1781 845 1859 891
rect 1905 845 1983 891
rect 2029 845 2107 891
rect 2153 845 2231 891
rect 2277 845 2355 891
rect 2401 845 2479 891
rect 2525 845 2603 891
rect 2649 845 2727 891
rect 2773 845 2851 891
rect 2897 845 2975 891
rect 3021 845 3099 891
rect 3145 845 3223 891
rect 3269 845 3347 891
rect 3393 845 3471 891
rect 3517 845 3595 891
rect 3641 845 3719 891
rect 3765 845 3843 891
rect 3889 845 3967 891
rect 4013 845 4091 891
rect 4137 845 4215 891
rect 4261 845 4339 891
rect 4385 845 4463 891
rect 4509 845 4587 891
rect 4633 845 4711 891
rect 4757 845 4835 891
rect 4881 845 4959 891
rect 5005 845 5083 891
rect 5129 845 5207 891
rect 5253 845 5331 891
rect 5377 845 5455 891
rect 5501 845 5579 891
rect 5625 845 5703 891
rect 5749 845 5827 891
rect 5873 845 5951 891
rect 5997 845 6075 891
rect 6121 845 6199 891
rect 6245 845 6323 891
rect 6369 845 6447 891
rect 6493 845 6571 891
rect 6617 845 6695 891
rect 6741 845 6819 891
rect 6865 845 6943 891
rect 6989 845 7067 891
rect 7113 845 7191 891
rect 7237 845 7315 891
rect 7361 845 7439 891
rect 7485 845 7563 891
rect 7609 845 7687 891
rect 7733 845 7811 891
rect 7857 845 7935 891
rect 7981 845 8059 891
rect 8105 845 8183 891
rect 8229 845 8307 891
rect 8353 845 8431 891
rect 8477 845 8555 891
rect 8601 845 8679 891
rect 8725 845 8803 891
rect 8849 845 8927 891
rect 8973 845 9051 891
rect 9097 845 9175 891
rect 9221 845 9299 891
rect 9345 845 9423 891
rect 9469 845 9547 891
rect 9593 845 9671 891
rect 9717 845 9795 891
rect 9841 845 9919 891
rect 9965 845 10043 891
rect 10089 845 10167 891
rect 10213 845 10291 891
rect 10337 845 10415 891
rect 10461 845 10539 891
rect 10585 845 10663 891
rect 10709 845 10787 891
rect 10833 845 10911 891
rect 10957 845 11035 891
rect 11081 845 11159 891
rect 11205 845 11283 891
rect 11329 845 11407 891
rect 11453 845 11531 891
rect 11577 845 11655 891
rect 11701 845 11779 891
rect 11825 845 11903 891
rect 11949 845 12027 891
rect 12073 845 12151 891
rect 12197 845 12275 891
rect 12321 845 12399 891
rect 12445 845 12523 891
rect 12569 845 12647 891
rect 12693 845 12771 891
rect 12817 845 12895 891
rect 12941 845 13019 891
rect 13065 845 13143 891
rect 13189 845 13267 891
rect 13313 845 13391 891
rect 13437 845 13515 891
rect 13561 845 13639 891
rect 13685 845 13763 891
rect 13809 845 13887 891
rect 13933 845 14011 891
rect 14057 845 14135 891
rect 14181 845 14259 891
rect 14305 845 14383 891
rect 14429 845 14507 891
rect 14553 845 14631 891
rect 14677 845 14755 891
rect 14801 845 14879 891
rect 14925 845 15003 891
rect 15049 845 15127 891
rect 15173 845 15251 891
rect 15297 845 15375 891
rect 15421 845 15499 891
rect 15545 845 15623 891
rect 15669 845 15747 891
rect 15793 845 15871 891
rect 15917 845 15995 891
rect 16041 845 16119 891
rect 16165 845 16243 891
rect 16289 845 16367 891
rect 16413 845 16491 891
rect 16537 845 16615 891
rect 16661 845 16739 891
rect 16785 845 16863 891
rect 16909 845 16987 891
rect 17033 845 17111 891
rect 17157 845 17235 891
rect 17281 845 17359 891
rect 17405 845 17483 891
rect 17529 845 17607 891
rect 17653 845 17731 891
rect 17777 845 17855 891
rect 17901 845 17979 891
rect 18025 845 18103 891
rect 18149 845 18227 891
rect 18273 845 18351 891
rect 18397 845 18475 891
rect 18521 845 18599 891
rect 18645 845 18723 891
rect 18769 845 18847 891
rect 18893 845 18971 891
rect 19017 845 19095 891
rect 19141 845 19219 891
rect 19265 845 19343 891
rect 19389 845 19467 891
rect 19513 845 19591 891
rect 19637 845 19715 891
rect 19761 845 19839 891
rect 19885 845 19963 891
rect 20009 845 20087 891
rect 20133 845 20211 891
rect 20257 845 20335 891
rect 20381 845 20459 891
rect 20505 845 20583 891
rect 20629 845 20707 891
rect 20753 845 20831 891
rect 20877 845 20955 891
rect 21001 845 21079 891
rect 21125 845 21203 891
rect 21249 845 21327 891
rect 21373 845 21451 891
rect 21497 845 21575 891
rect 21621 845 21699 891
rect 21745 845 21823 891
rect 21869 845 21947 891
rect 21993 845 22071 891
rect 22117 845 22195 891
rect 22241 845 22319 891
rect 22365 845 22443 891
rect 22489 845 22567 891
rect 22613 845 22691 891
rect 22737 845 22815 891
rect 22861 845 22939 891
rect 22985 845 23063 891
rect 23109 845 23187 891
rect 23233 845 23311 891
rect 23357 845 23435 891
rect 23481 845 23559 891
rect 23605 845 23683 891
rect 23729 845 23807 891
rect 23853 845 23931 891
rect 23977 845 24055 891
rect 24101 845 24179 891
rect 24225 845 24303 891
rect 24349 845 24427 891
rect 24473 845 24551 891
rect 24597 845 24675 891
rect 24721 845 24799 891
rect 24845 845 24923 891
rect 24969 845 25047 891
rect 25093 845 25171 891
rect 25217 845 25295 891
rect 25341 845 25419 891
rect 25465 845 25543 891
rect 25589 845 25667 891
rect 25713 845 25791 891
rect 25837 845 25915 891
rect 25961 845 26039 891
rect 26085 845 26163 891
rect 26209 845 26287 891
rect 26333 845 26411 891
rect 26457 845 26535 891
rect 26581 845 26659 891
rect 26705 845 26783 891
rect 26829 845 26907 891
rect 26953 845 27031 891
rect 27077 845 27155 891
rect 27201 845 27279 891
rect 27325 845 27403 891
rect 27449 845 27527 891
rect 27573 845 27651 891
rect 27697 845 27775 891
rect 27821 845 27899 891
rect 27945 845 28023 891
rect 28069 845 28147 891
rect 28193 845 28271 891
rect 28317 845 28395 891
rect 28441 845 28519 891
rect 28565 845 28643 891
rect 28689 845 28767 891
rect 28813 845 28891 891
rect 28937 845 29015 891
rect 29061 845 29139 891
rect 29185 845 29263 891
rect 29309 845 29387 891
rect 29433 845 29511 891
rect 29557 845 29635 891
rect 29681 845 29759 891
rect 29805 845 29883 891
rect 29929 845 30007 891
rect 30053 845 30131 891
rect 30177 845 30255 891
rect 30301 845 30379 891
rect 30425 845 30503 891
rect 30549 845 30627 891
rect 30673 845 30751 891
rect 30797 845 30875 891
rect 30921 845 30999 891
rect 31045 845 31123 891
rect 31169 845 31247 891
rect 31293 845 31371 891
rect 31417 845 31495 891
rect 31541 845 31619 891
rect 31665 845 31743 891
rect 31789 845 31867 891
rect 31913 845 31991 891
rect 32037 845 32115 891
rect 32161 845 32239 891
rect 32285 845 32363 891
rect 32409 845 32487 891
rect 32533 845 32611 891
rect 32657 845 32735 891
rect 32781 845 32859 891
rect 32905 845 32983 891
rect 33029 845 33107 891
rect 33153 845 33231 891
rect 33277 845 33355 891
rect 33401 845 33479 891
rect 33525 845 33603 891
rect 33649 845 33727 891
rect 33773 845 33851 891
rect 33897 845 33975 891
rect 34021 845 34099 891
rect 34145 845 34223 891
rect 34269 845 34347 891
rect 34393 845 34471 891
rect 34517 845 34595 891
rect 34641 845 34719 891
rect 34765 845 34843 891
rect 34889 845 34967 891
rect 35013 845 35091 891
rect 35137 845 35215 891
rect 35261 845 35339 891
rect 35385 845 35463 891
rect 35509 845 35587 891
rect 35633 845 35711 891
rect 35757 845 35835 891
rect 35881 845 35959 891
rect 36005 845 36083 891
rect 36129 845 36207 891
rect 36253 845 36331 891
rect 36377 845 36455 891
rect 36501 845 36579 891
rect 36625 845 36703 891
rect 36749 845 36827 891
rect 36873 845 36951 891
rect 36997 845 37075 891
rect 37121 845 37199 891
rect 37245 845 37323 891
rect 37369 845 37447 891
rect 37493 845 37571 891
rect 37617 845 37695 891
rect 37741 845 37819 891
rect 37865 845 37943 891
rect 37989 845 38067 891
rect 38113 845 38191 891
rect 38237 845 38315 891
rect 38361 845 38439 891
rect 38485 845 38563 891
rect 38609 845 38687 891
rect 38733 845 38811 891
rect 38857 845 38935 891
rect 38981 845 39059 891
rect 39105 845 39183 891
rect 39229 845 39307 891
rect 39353 845 39431 891
rect 39477 845 39555 891
rect 39601 845 39679 891
rect 39725 845 39803 891
rect 39849 845 39927 891
rect 39973 845 40051 891
rect 40097 845 40175 891
rect 40221 845 40299 891
rect 40345 845 40423 891
rect 40469 845 40547 891
rect 40593 845 40671 891
rect 40717 845 40795 891
rect 40841 845 40919 891
rect 40965 845 41043 891
rect 41089 845 41167 891
rect 41213 845 41291 891
rect 41337 845 41415 891
rect 41461 845 41539 891
rect 41585 845 41663 891
rect 41709 845 41787 891
rect 41833 845 41911 891
rect 41957 845 42035 891
rect 42081 845 42159 891
rect 42205 845 42283 891
rect 42329 845 42407 891
rect 42453 845 42531 891
rect 42577 845 42655 891
rect 42701 845 42779 891
rect 42825 845 42903 891
rect 42949 845 43027 891
rect 43073 845 43151 891
rect 43197 845 43275 891
rect 43321 845 43399 891
rect 43445 845 43523 891
rect 43569 845 43647 891
rect 43693 845 43771 891
rect 43817 845 43895 891
rect 43941 845 44019 891
rect 44065 845 44143 891
rect 44189 845 44267 891
rect 44313 845 44391 891
rect 44437 845 44515 891
rect 44561 845 44639 891
rect 44685 845 44763 891
rect 44809 845 44887 891
rect 44933 845 45011 891
rect 45057 845 45135 891
rect 45181 845 45259 891
rect 45305 845 45383 891
rect 45429 845 45507 891
rect 45553 845 45631 891
rect 45677 845 45755 891
rect 45801 845 45879 891
rect 45925 845 46003 891
rect 46049 845 46127 891
rect 46173 845 46251 891
rect 46297 845 46375 891
rect 46421 845 46499 891
rect 46545 845 46623 891
rect 46669 845 46747 891
rect 46793 845 46871 891
rect 46917 845 46995 891
rect 47041 845 47119 891
rect 47165 845 47243 891
rect 47289 845 47367 891
rect 47413 845 47491 891
rect 47537 845 47615 891
rect 47661 845 47739 891
rect 47785 845 47863 891
rect 47909 845 47987 891
rect 48033 845 48111 891
rect 48157 845 48235 891
rect 48281 845 48359 891
rect 48405 845 48483 891
rect 48529 845 48607 891
rect 48653 845 48731 891
rect 48777 845 48855 891
rect 48901 845 48979 891
rect 49025 845 49103 891
rect 49149 845 49227 891
rect 49273 845 49351 891
rect 49397 845 49475 891
rect 49521 845 49599 891
rect 49645 845 49723 891
rect 49769 845 49847 891
rect 49893 845 49971 891
rect 50017 845 50095 891
rect 50141 845 50219 891
rect 50265 845 50343 891
rect 50389 845 50467 891
rect 50513 845 50591 891
rect 50637 845 50715 891
rect 50761 845 50839 891
rect 50885 845 50963 891
rect 51009 845 51087 891
rect 51133 845 51211 891
rect 51257 845 51335 891
rect 51381 845 51459 891
rect 51505 845 51583 891
rect 51629 845 51707 891
rect 51753 845 51831 891
rect 51877 845 51955 891
rect 52001 845 52079 891
rect 52125 845 52203 891
rect 52249 845 52327 891
rect 52373 845 52451 891
rect 52497 845 52575 891
rect 52621 845 52699 891
rect 52745 845 52823 891
rect 52869 845 52947 891
rect 52993 845 53071 891
rect 53117 845 53195 891
rect 53241 845 53319 891
rect 53365 845 53443 891
rect 53489 845 53567 891
rect 53613 845 53691 891
rect 53737 845 53815 891
rect 53861 845 53939 891
rect 53985 845 54063 891
rect 54109 845 54187 891
rect 54233 845 54311 891
rect 54357 845 54435 891
rect 54481 845 54559 891
rect 54605 845 54683 891
rect 54729 845 54807 891
rect 54853 845 54931 891
rect 54977 845 55055 891
rect 55101 845 55179 891
rect 55225 845 55303 891
rect 55349 845 55427 891
rect 55473 845 55551 891
rect 55597 845 55675 891
rect 55721 845 55799 891
rect 55845 845 55923 891
rect 55969 845 56047 891
rect 56093 845 56171 891
rect 56217 845 56295 891
rect 56341 845 56419 891
rect 56465 845 56543 891
rect 56589 845 56667 891
rect 56713 845 56791 891
rect 56837 845 56915 891
rect 56961 845 57039 891
rect 57085 845 57163 891
rect 57209 845 57287 891
rect 57333 845 57411 891
rect 57457 845 57535 891
rect 57581 845 57659 891
rect 57705 845 57783 891
rect 57829 845 57907 891
rect 57953 845 58031 891
rect 58077 845 58155 891
rect 58201 845 58279 891
rect 58325 845 58403 891
rect 58449 845 58527 891
rect 58573 845 58651 891
rect 58697 845 58775 891
rect 58821 845 58899 891
rect 58945 845 59023 891
rect 59069 845 59147 891
rect 59193 845 59271 891
rect 59317 845 59395 891
rect 59441 845 59519 891
rect 59565 845 59643 891
rect 59689 845 59767 891
rect 59813 845 59891 891
rect 59937 845 60015 891
rect 60061 845 60139 891
rect 60185 845 60263 891
rect 60309 845 60387 891
rect 60433 845 60511 891
rect 60557 845 60635 891
rect 60681 845 60759 891
rect 60805 845 60883 891
rect 60929 845 61007 891
rect 61053 845 61131 891
rect 61177 845 61255 891
rect 61301 845 61379 891
rect 61425 845 61503 891
rect 61549 845 61627 891
rect 61673 845 61751 891
rect 61797 845 61875 891
rect 61921 845 61999 891
rect 62045 845 62123 891
rect 62169 845 62247 891
rect 62293 845 62371 891
rect 62417 845 62495 891
rect 62541 845 62619 891
rect 62665 845 62743 891
rect 62789 845 62867 891
rect 62913 845 62991 891
rect 63037 845 63115 891
rect 63161 845 63239 891
rect 63285 845 63363 891
rect 63409 845 63487 891
rect 63533 845 63611 891
rect 63657 845 63735 891
rect 63781 845 63859 891
rect 63905 845 63983 891
rect 64029 845 64107 891
rect 64153 845 64231 891
rect 64277 845 64355 891
rect 64401 845 64479 891
rect 64525 845 64603 891
rect 64649 845 64727 891
rect 64773 845 64851 891
rect 64897 845 64975 891
rect 65021 845 65099 891
rect 65145 845 65223 891
rect 65269 845 65347 891
rect 65393 845 65471 891
rect 65517 845 65595 891
rect 65641 845 65719 891
rect 65765 845 65843 891
rect 65889 845 65967 891
rect 66013 845 66091 891
rect 66137 845 66215 891
rect 66261 845 66339 891
rect 66385 845 66463 891
rect 66509 845 66587 891
rect 66633 845 66711 891
rect 66757 845 66835 891
rect 66881 845 66959 891
rect 67005 845 67083 891
rect 67129 845 67207 891
rect 67253 845 67331 891
rect 67377 845 67455 891
rect 67501 845 67579 891
rect 67625 845 67703 891
rect 67749 845 67827 891
rect 67873 845 67951 891
rect 67997 845 68075 891
rect 68121 845 68199 891
rect 68245 845 68323 891
rect 68369 845 68447 891
rect 68493 845 68571 891
rect 68617 845 68695 891
rect 68741 845 68819 891
rect 68865 845 68943 891
rect 68989 845 69067 891
rect 69113 845 69191 891
rect 69237 845 69315 891
rect 69361 845 69439 891
rect 69485 845 69563 891
rect 69609 845 69687 891
rect 69733 845 69811 891
rect 69857 845 69935 891
rect 69981 845 70059 891
rect 70105 845 70183 891
rect 70229 845 70307 891
rect 70353 845 70431 891
rect 70477 845 70555 891
rect 70601 845 70679 891
rect 70725 845 70803 891
rect 70849 845 70927 891
rect 70973 845 71051 891
rect 71097 845 71175 891
rect 71221 845 71299 891
rect 71345 845 71423 891
rect 71469 845 71547 891
rect 71593 845 71671 891
rect 71717 845 71795 891
rect 71841 845 71919 891
rect 71965 845 72043 891
rect 72089 845 72167 891
rect 72213 845 72291 891
rect 72337 845 72415 891
rect 72461 845 72539 891
rect 72585 845 72663 891
rect 72709 845 72787 891
rect 72833 845 72911 891
rect 72957 845 73035 891
rect 73081 845 73159 891
rect 73205 845 73283 891
rect 73329 845 73407 891
rect 73453 845 73531 891
rect 73577 845 73655 891
rect 73701 845 73779 891
rect 73825 845 73903 891
rect 73949 845 74027 891
rect 74073 845 74151 891
rect 74197 845 74275 891
rect 74321 845 74399 891
rect 74445 845 74523 891
rect 74569 845 74647 891
rect 74693 845 74771 891
rect 74817 845 74895 891
rect 74941 845 75019 891
rect 75065 845 75143 891
rect 75189 845 75267 891
rect 75313 845 75391 891
rect 75437 845 75515 891
rect 75561 845 75639 891
rect 75685 845 75763 891
rect 75809 845 75887 891
rect 75933 845 76011 891
rect 76057 845 76135 891
rect 76181 845 76259 891
rect 76305 845 76383 891
rect 76429 845 76507 891
rect 76553 845 76631 891
rect 76677 845 76755 891
rect 76801 845 76879 891
rect 76925 845 77003 891
rect 77049 845 77127 891
rect 77173 845 77251 891
rect 77297 845 77375 891
rect 77421 845 77499 891
rect 77545 845 77623 891
rect 77669 845 77747 891
rect 77793 845 77871 891
rect 77917 845 77995 891
rect 78041 845 78119 891
rect 78165 845 78243 891
rect 78289 845 78367 891
rect 78413 845 78491 891
rect 78537 845 78615 891
rect 78661 845 78739 891
rect 78785 845 78863 891
rect 78909 845 78987 891
rect 79033 845 79111 891
rect 79157 845 79235 891
rect 79281 845 79359 891
rect 79405 845 79483 891
rect 79529 845 79607 891
rect 79653 845 79731 891
rect 79777 845 79855 891
rect 79901 845 79979 891
rect 80025 845 80103 891
rect 80149 845 80227 891
rect 80273 845 80351 891
rect 80397 845 80475 891
rect 80521 845 80599 891
rect 80645 845 80723 891
rect 80769 845 80847 891
rect 80893 845 80971 891
rect 81017 845 81095 891
rect 81141 845 81219 891
rect 81265 845 81343 891
rect 81389 845 81467 891
rect 81513 845 81591 891
rect 81637 845 81715 891
rect 81761 845 81839 891
rect 81885 845 81963 891
rect 82009 845 82087 891
rect 82133 845 82211 891
rect 82257 845 82335 891
rect 82381 845 82459 891
rect 82505 845 82583 891
rect 82629 845 82707 891
rect 82753 845 82831 891
rect 82877 845 82955 891
rect 83001 845 83079 891
rect 83125 845 83203 891
rect 83249 845 83327 891
rect 83373 845 83451 891
rect 83497 845 83575 891
rect 83621 845 83699 891
rect 83745 845 83823 891
rect 83869 845 83947 891
rect 83993 845 84071 891
rect 84117 845 84195 891
rect 84241 845 84319 891
rect 84365 845 84443 891
rect 84489 845 84567 891
rect 84613 845 84691 891
rect 84737 845 84815 891
rect 84861 845 84939 891
rect 84985 845 85063 891
rect 85109 845 85187 891
rect 85233 845 85311 891
rect 85357 845 85435 891
rect 85481 845 85559 891
rect 85605 845 85683 891
rect 85729 845 85807 891
rect 85853 845 85931 891
rect 85977 845 86090 891
rect 282 767 86090 845
rect 282 721 371 767
rect 417 721 495 767
rect 541 721 619 767
rect 665 721 743 767
rect 789 721 867 767
rect 913 721 991 767
rect 1037 721 1115 767
rect 1161 721 1239 767
rect 1285 721 1363 767
rect 1409 721 1487 767
rect 1533 721 1611 767
rect 1657 721 1735 767
rect 1781 721 1859 767
rect 1905 721 1983 767
rect 2029 721 2107 767
rect 2153 721 2231 767
rect 2277 721 2355 767
rect 2401 721 2479 767
rect 2525 721 2603 767
rect 2649 721 2727 767
rect 2773 721 2851 767
rect 2897 721 2975 767
rect 3021 721 3099 767
rect 3145 721 3223 767
rect 3269 721 3347 767
rect 3393 721 3471 767
rect 3517 721 3595 767
rect 3641 721 3719 767
rect 3765 721 3843 767
rect 3889 721 3967 767
rect 4013 721 4091 767
rect 4137 721 4215 767
rect 4261 721 4339 767
rect 4385 721 4463 767
rect 4509 721 4587 767
rect 4633 721 4711 767
rect 4757 721 4835 767
rect 4881 721 4959 767
rect 5005 721 5083 767
rect 5129 721 5207 767
rect 5253 721 5331 767
rect 5377 721 5455 767
rect 5501 721 5579 767
rect 5625 721 5703 767
rect 5749 721 5827 767
rect 5873 721 5951 767
rect 5997 721 6075 767
rect 6121 721 6199 767
rect 6245 721 6323 767
rect 6369 721 6447 767
rect 6493 721 6571 767
rect 6617 721 6695 767
rect 6741 721 6819 767
rect 6865 721 6943 767
rect 6989 721 7067 767
rect 7113 721 7191 767
rect 7237 721 7315 767
rect 7361 721 7439 767
rect 7485 721 7563 767
rect 7609 721 7687 767
rect 7733 721 7811 767
rect 7857 721 7935 767
rect 7981 721 8059 767
rect 8105 721 8183 767
rect 8229 721 8307 767
rect 8353 721 8431 767
rect 8477 721 8555 767
rect 8601 721 8679 767
rect 8725 721 8803 767
rect 8849 721 8927 767
rect 8973 721 9051 767
rect 9097 721 9175 767
rect 9221 721 9299 767
rect 9345 721 9423 767
rect 9469 721 9547 767
rect 9593 721 9671 767
rect 9717 721 9795 767
rect 9841 721 9919 767
rect 9965 721 10043 767
rect 10089 721 10167 767
rect 10213 721 10291 767
rect 10337 721 10415 767
rect 10461 721 10539 767
rect 10585 721 10663 767
rect 10709 721 10787 767
rect 10833 721 10911 767
rect 10957 721 11035 767
rect 11081 721 11159 767
rect 11205 721 11283 767
rect 11329 721 11407 767
rect 11453 721 11531 767
rect 11577 721 11655 767
rect 11701 721 11779 767
rect 11825 721 11903 767
rect 11949 721 12027 767
rect 12073 721 12151 767
rect 12197 721 12275 767
rect 12321 721 12399 767
rect 12445 721 12523 767
rect 12569 721 12647 767
rect 12693 721 12771 767
rect 12817 721 12895 767
rect 12941 721 13019 767
rect 13065 721 13143 767
rect 13189 721 13267 767
rect 13313 721 13391 767
rect 13437 721 13515 767
rect 13561 721 13639 767
rect 13685 721 13763 767
rect 13809 721 13887 767
rect 13933 721 14011 767
rect 14057 721 14135 767
rect 14181 721 14259 767
rect 14305 721 14383 767
rect 14429 721 14507 767
rect 14553 721 14631 767
rect 14677 721 14755 767
rect 14801 721 14879 767
rect 14925 721 15003 767
rect 15049 721 15127 767
rect 15173 721 15251 767
rect 15297 721 15375 767
rect 15421 721 15499 767
rect 15545 721 15623 767
rect 15669 721 15747 767
rect 15793 721 15871 767
rect 15917 721 15995 767
rect 16041 721 16119 767
rect 16165 721 16243 767
rect 16289 721 16367 767
rect 16413 721 16491 767
rect 16537 721 16615 767
rect 16661 721 16739 767
rect 16785 721 16863 767
rect 16909 721 16987 767
rect 17033 721 17111 767
rect 17157 721 17235 767
rect 17281 721 17359 767
rect 17405 721 17483 767
rect 17529 721 17607 767
rect 17653 721 17731 767
rect 17777 721 17855 767
rect 17901 721 17979 767
rect 18025 721 18103 767
rect 18149 721 18227 767
rect 18273 721 18351 767
rect 18397 721 18475 767
rect 18521 721 18599 767
rect 18645 721 18723 767
rect 18769 721 18847 767
rect 18893 721 18971 767
rect 19017 721 19095 767
rect 19141 721 19219 767
rect 19265 721 19343 767
rect 19389 721 19467 767
rect 19513 721 19591 767
rect 19637 721 19715 767
rect 19761 721 19839 767
rect 19885 721 19963 767
rect 20009 721 20087 767
rect 20133 721 20211 767
rect 20257 721 20335 767
rect 20381 721 20459 767
rect 20505 721 20583 767
rect 20629 721 20707 767
rect 20753 721 20831 767
rect 20877 721 20955 767
rect 21001 721 21079 767
rect 21125 721 21203 767
rect 21249 721 21327 767
rect 21373 721 21451 767
rect 21497 721 21575 767
rect 21621 721 21699 767
rect 21745 721 21823 767
rect 21869 721 21947 767
rect 21993 721 22071 767
rect 22117 721 22195 767
rect 22241 721 22319 767
rect 22365 721 22443 767
rect 22489 721 22567 767
rect 22613 721 22691 767
rect 22737 721 22815 767
rect 22861 721 22939 767
rect 22985 721 23063 767
rect 23109 721 23187 767
rect 23233 721 23311 767
rect 23357 721 23435 767
rect 23481 721 23559 767
rect 23605 721 23683 767
rect 23729 721 23807 767
rect 23853 721 23931 767
rect 23977 721 24055 767
rect 24101 721 24179 767
rect 24225 721 24303 767
rect 24349 721 24427 767
rect 24473 721 24551 767
rect 24597 721 24675 767
rect 24721 721 24799 767
rect 24845 721 24923 767
rect 24969 721 25047 767
rect 25093 721 25171 767
rect 25217 721 25295 767
rect 25341 721 25419 767
rect 25465 721 25543 767
rect 25589 721 25667 767
rect 25713 721 25791 767
rect 25837 721 25915 767
rect 25961 721 26039 767
rect 26085 721 26163 767
rect 26209 721 26287 767
rect 26333 721 26411 767
rect 26457 721 26535 767
rect 26581 721 26659 767
rect 26705 721 26783 767
rect 26829 721 26907 767
rect 26953 721 27031 767
rect 27077 721 27155 767
rect 27201 721 27279 767
rect 27325 721 27403 767
rect 27449 721 27527 767
rect 27573 721 27651 767
rect 27697 721 27775 767
rect 27821 721 27899 767
rect 27945 721 28023 767
rect 28069 721 28147 767
rect 28193 721 28271 767
rect 28317 721 28395 767
rect 28441 721 28519 767
rect 28565 721 28643 767
rect 28689 721 28767 767
rect 28813 721 28891 767
rect 28937 721 29015 767
rect 29061 721 29139 767
rect 29185 721 29263 767
rect 29309 721 29387 767
rect 29433 721 29511 767
rect 29557 721 29635 767
rect 29681 721 29759 767
rect 29805 721 29883 767
rect 29929 721 30007 767
rect 30053 721 30131 767
rect 30177 721 30255 767
rect 30301 721 30379 767
rect 30425 721 30503 767
rect 30549 721 30627 767
rect 30673 721 30751 767
rect 30797 721 30875 767
rect 30921 721 30999 767
rect 31045 721 31123 767
rect 31169 721 31247 767
rect 31293 721 31371 767
rect 31417 721 31495 767
rect 31541 721 31619 767
rect 31665 721 31743 767
rect 31789 721 31867 767
rect 31913 721 31991 767
rect 32037 721 32115 767
rect 32161 721 32239 767
rect 32285 721 32363 767
rect 32409 721 32487 767
rect 32533 721 32611 767
rect 32657 721 32735 767
rect 32781 721 32859 767
rect 32905 721 32983 767
rect 33029 721 33107 767
rect 33153 721 33231 767
rect 33277 721 33355 767
rect 33401 721 33479 767
rect 33525 721 33603 767
rect 33649 721 33727 767
rect 33773 721 33851 767
rect 33897 721 33975 767
rect 34021 721 34099 767
rect 34145 721 34223 767
rect 34269 721 34347 767
rect 34393 721 34471 767
rect 34517 721 34595 767
rect 34641 721 34719 767
rect 34765 721 34843 767
rect 34889 721 34967 767
rect 35013 721 35091 767
rect 35137 721 35215 767
rect 35261 721 35339 767
rect 35385 721 35463 767
rect 35509 721 35587 767
rect 35633 721 35711 767
rect 35757 721 35835 767
rect 35881 721 35959 767
rect 36005 721 36083 767
rect 36129 721 36207 767
rect 36253 721 36331 767
rect 36377 721 36455 767
rect 36501 721 36579 767
rect 36625 721 36703 767
rect 36749 721 36827 767
rect 36873 721 36951 767
rect 36997 721 37075 767
rect 37121 721 37199 767
rect 37245 721 37323 767
rect 37369 721 37447 767
rect 37493 721 37571 767
rect 37617 721 37695 767
rect 37741 721 37819 767
rect 37865 721 37943 767
rect 37989 721 38067 767
rect 38113 721 38191 767
rect 38237 721 38315 767
rect 38361 721 38439 767
rect 38485 721 38563 767
rect 38609 721 38687 767
rect 38733 721 38811 767
rect 38857 721 38935 767
rect 38981 721 39059 767
rect 39105 721 39183 767
rect 39229 721 39307 767
rect 39353 721 39431 767
rect 39477 721 39555 767
rect 39601 721 39679 767
rect 39725 721 39803 767
rect 39849 721 39927 767
rect 39973 721 40051 767
rect 40097 721 40175 767
rect 40221 721 40299 767
rect 40345 721 40423 767
rect 40469 721 40547 767
rect 40593 721 40671 767
rect 40717 721 40795 767
rect 40841 721 40919 767
rect 40965 721 41043 767
rect 41089 721 41167 767
rect 41213 721 41291 767
rect 41337 721 41415 767
rect 41461 721 41539 767
rect 41585 721 41663 767
rect 41709 721 41787 767
rect 41833 721 41911 767
rect 41957 721 42035 767
rect 42081 721 42159 767
rect 42205 721 42283 767
rect 42329 721 42407 767
rect 42453 721 42531 767
rect 42577 721 42655 767
rect 42701 721 42779 767
rect 42825 721 42903 767
rect 42949 721 43027 767
rect 43073 721 43151 767
rect 43197 721 43275 767
rect 43321 721 43399 767
rect 43445 721 43523 767
rect 43569 721 43647 767
rect 43693 721 43771 767
rect 43817 721 43895 767
rect 43941 721 44019 767
rect 44065 721 44143 767
rect 44189 721 44267 767
rect 44313 721 44391 767
rect 44437 721 44515 767
rect 44561 721 44639 767
rect 44685 721 44763 767
rect 44809 721 44887 767
rect 44933 721 45011 767
rect 45057 721 45135 767
rect 45181 721 45259 767
rect 45305 721 45383 767
rect 45429 721 45507 767
rect 45553 721 45631 767
rect 45677 721 45755 767
rect 45801 721 45879 767
rect 45925 721 46003 767
rect 46049 721 46127 767
rect 46173 721 46251 767
rect 46297 721 46375 767
rect 46421 721 46499 767
rect 46545 721 46623 767
rect 46669 721 46747 767
rect 46793 721 46871 767
rect 46917 721 46995 767
rect 47041 721 47119 767
rect 47165 721 47243 767
rect 47289 721 47367 767
rect 47413 721 47491 767
rect 47537 721 47615 767
rect 47661 721 47739 767
rect 47785 721 47863 767
rect 47909 721 47987 767
rect 48033 721 48111 767
rect 48157 721 48235 767
rect 48281 721 48359 767
rect 48405 721 48483 767
rect 48529 721 48607 767
rect 48653 721 48731 767
rect 48777 721 48855 767
rect 48901 721 48979 767
rect 49025 721 49103 767
rect 49149 721 49227 767
rect 49273 721 49351 767
rect 49397 721 49475 767
rect 49521 721 49599 767
rect 49645 721 49723 767
rect 49769 721 49847 767
rect 49893 721 49971 767
rect 50017 721 50095 767
rect 50141 721 50219 767
rect 50265 721 50343 767
rect 50389 721 50467 767
rect 50513 721 50591 767
rect 50637 721 50715 767
rect 50761 721 50839 767
rect 50885 721 50963 767
rect 51009 721 51087 767
rect 51133 721 51211 767
rect 51257 721 51335 767
rect 51381 721 51459 767
rect 51505 721 51583 767
rect 51629 721 51707 767
rect 51753 721 51831 767
rect 51877 721 51955 767
rect 52001 721 52079 767
rect 52125 721 52203 767
rect 52249 721 52327 767
rect 52373 721 52451 767
rect 52497 721 52575 767
rect 52621 721 52699 767
rect 52745 721 52823 767
rect 52869 721 52947 767
rect 52993 721 53071 767
rect 53117 721 53195 767
rect 53241 721 53319 767
rect 53365 721 53443 767
rect 53489 721 53567 767
rect 53613 721 53691 767
rect 53737 721 53815 767
rect 53861 721 53939 767
rect 53985 721 54063 767
rect 54109 721 54187 767
rect 54233 721 54311 767
rect 54357 721 54435 767
rect 54481 721 54559 767
rect 54605 721 54683 767
rect 54729 721 54807 767
rect 54853 721 54931 767
rect 54977 721 55055 767
rect 55101 721 55179 767
rect 55225 721 55303 767
rect 55349 721 55427 767
rect 55473 721 55551 767
rect 55597 721 55675 767
rect 55721 721 55799 767
rect 55845 721 55923 767
rect 55969 721 56047 767
rect 56093 721 56171 767
rect 56217 721 56295 767
rect 56341 721 56419 767
rect 56465 721 56543 767
rect 56589 721 56667 767
rect 56713 721 56791 767
rect 56837 721 56915 767
rect 56961 721 57039 767
rect 57085 721 57163 767
rect 57209 721 57287 767
rect 57333 721 57411 767
rect 57457 721 57535 767
rect 57581 721 57659 767
rect 57705 721 57783 767
rect 57829 721 57907 767
rect 57953 721 58031 767
rect 58077 721 58155 767
rect 58201 721 58279 767
rect 58325 721 58403 767
rect 58449 721 58527 767
rect 58573 721 58651 767
rect 58697 721 58775 767
rect 58821 721 58899 767
rect 58945 721 59023 767
rect 59069 721 59147 767
rect 59193 721 59271 767
rect 59317 721 59395 767
rect 59441 721 59519 767
rect 59565 721 59643 767
rect 59689 721 59767 767
rect 59813 721 59891 767
rect 59937 721 60015 767
rect 60061 721 60139 767
rect 60185 721 60263 767
rect 60309 721 60387 767
rect 60433 721 60511 767
rect 60557 721 60635 767
rect 60681 721 60759 767
rect 60805 721 60883 767
rect 60929 721 61007 767
rect 61053 721 61131 767
rect 61177 721 61255 767
rect 61301 721 61379 767
rect 61425 721 61503 767
rect 61549 721 61627 767
rect 61673 721 61751 767
rect 61797 721 61875 767
rect 61921 721 61999 767
rect 62045 721 62123 767
rect 62169 721 62247 767
rect 62293 721 62371 767
rect 62417 721 62495 767
rect 62541 721 62619 767
rect 62665 721 62743 767
rect 62789 721 62867 767
rect 62913 721 62991 767
rect 63037 721 63115 767
rect 63161 721 63239 767
rect 63285 721 63363 767
rect 63409 721 63487 767
rect 63533 721 63611 767
rect 63657 721 63735 767
rect 63781 721 63859 767
rect 63905 721 63983 767
rect 64029 721 64107 767
rect 64153 721 64231 767
rect 64277 721 64355 767
rect 64401 721 64479 767
rect 64525 721 64603 767
rect 64649 721 64727 767
rect 64773 721 64851 767
rect 64897 721 64975 767
rect 65021 721 65099 767
rect 65145 721 65223 767
rect 65269 721 65347 767
rect 65393 721 65471 767
rect 65517 721 65595 767
rect 65641 721 65719 767
rect 65765 721 65843 767
rect 65889 721 65967 767
rect 66013 721 66091 767
rect 66137 721 66215 767
rect 66261 721 66339 767
rect 66385 721 66463 767
rect 66509 721 66587 767
rect 66633 721 66711 767
rect 66757 721 66835 767
rect 66881 721 66959 767
rect 67005 721 67083 767
rect 67129 721 67207 767
rect 67253 721 67331 767
rect 67377 721 67455 767
rect 67501 721 67579 767
rect 67625 721 67703 767
rect 67749 721 67827 767
rect 67873 721 67951 767
rect 67997 721 68075 767
rect 68121 721 68199 767
rect 68245 721 68323 767
rect 68369 721 68447 767
rect 68493 721 68571 767
rect 68617 721 68695 767
rect 68741 721 68819 767
rect 68865 721 68943 767
rect 68989 721 69067 767
rect 69113 721 69191 767
rect 69237 721 69315 767
rect 69361 721 69439 767
rect 69485 721 69563 767
rect 69609 721 69687 767
rect 69733 721 69811 767
rect 69857 721 69935 767
rect 69981 721 70059 767
rect 70105 721 70183 767
rect 70229 721 70307 767
rect 70353 721 70431 767
rect 70477 721 70555 767
rect 70601 721 70679 767
rect 70725 721 70803 767
rect 70849 721 70927 767
rect 70973 721 71051 767
rect 71097 721 71175 767
rect 71221 721 71299 767
rect 71345 721 71423 767
rect 71469 721 71547 767
rect 71593 721 71671 767
rect 71717 721 71795 767
rect 71841 721 71919 767
rect 71965 721 72043 767
rect 72089 721 72167 767
rect 72213 721 72291 767
rect 72337 721 72415 767
rect 72461 721 72539 767
rect 72585 721 72663 767
rect 72709 721 72787 767
rect 72833 721 72911 767
rect 72957 721 73035 767
rect 73081 721 73159 767
rect 73205 721 73283 767
rect 73329 721 73407 767
rect 73453 721 73531 767
rect 73577 721 73655 767
rect 73701 721 73779 767
rect 73825 721 73903 767
rect 73949 721 74027 767
rect 74073 721 74151 767
rect 74197 721 74275 767
rect 74321 721 74399 767
rect 74445 721 74523 767
rect 74569 721 74647 767
rect 74693 721 74771 767
rect 74817 721 74895 767
rect 74941 721 75019 767
rect 75065 721 75143 767
rect 75189 721 75267 767
rect 75313 721 75391 767
rect 75437 721 75515 767
rect 75561 721 75639 767
rect 75685 721 75763 767
rect 75809 721 75887 767
rect 75933 721 76011 767
rect 76057 721 76135 767
rect 76181 721 76259 767
rect 76305 721 76383 767
rect 76429 721 76507 767
rect 76553 721 76631 767
rect 76677 721 76755 767
rect 76801 721 76879 767
rect 76925 721 77003 767
rect 77049 721 77127 767
rect 77173 721 77251 767
rect 77297 721 77375 767
rect 77421 721 77499 767
rect 77545 721 77623 767
rect 77669 721 77747 767
rect 77793 721 77871 767
rect 77917 721 77995 767
rect 78041 721 78119 767
rect 78165 721 78243 767
rect 78289 721 78367 767
rect 78413 721 78491 767
rect 78537 721 78615 767
rect 78661 721 78739 767
rect 78785 721 78863 767
rect 78909 721 78987 767
rect 79033 721 79111 767
rect 79157 721 79235 767
rect 79281 721 79359 767
rect 79405 721 79483 767
rect 79529 721 79607 767
rect 79653 721 79731 767
rect 79777 721 79855 767
rect 79901 721 79979 767
rect 80025 721 80103 767
rect 80149 721 80227 767
rect 80273 721 80351 767
rect 80397 721 80475 767
rect 80521 721 80599 767
rect 80645 721 80723 767
rect 80769 721 80847 767
rect 80893 721 80971 767
rect 81017 721 81095 767
rect 81141 721 81219 767
rect 81265 721 81343 767
rect 81389 721 81467 767
rect 81513 721 81591 767
rect 81637 721 81715 767
rect 81761 721 81839 767
rect 81885 721 81963 767
rect 82009 721 82087 767
rect 82133 721 82211 767
rect 82257 721 82335 767
rect 82381 721 82459 767
rect 82505 721 82583 767
rect 82629 721 82707 767
rect 82753 721 82831 767
rect 82877 721 82955 767
rect 83001 721 83079 767
rect 83125 721 83203 767
rect 83249 721 83327 767
rect 83373 721 83451 767
rect 83497 721 83575 767
rect 83621 721 83699 767
rect 83745 721 83823 767
rect 83869 721 83947 767
rect 83993 721 84071 767
rect 84117 721 84195 767
rect 84241 721 84319 767
rect 84365 721 84443 767
rect 84489 721 84567 767
rect 84613 721 84691 767
rect 84737 721 84815 767
rect 84861 721 84939 767
rect 84985 721 85063 767
rect 85109 721 85187 767
rect 85233 721 85311 767
rect 85357 721 85435 767
rect 85481 721 85559 767
rect 85605 721 85683 767
rect 85729 721 85807 767
rect 85853 721 85931 767
rect 85977 721 86090 767
rect 282 643 86090 721
rect 282 597 371 643
rect 417 597 495 643
rect 541 597 619 643
rect 665 597 743 643
rect 789 597 867 643
rect 913 597 991 643
rect 1037 597 1115 643
rect 1161 597 1239 643
rect 1285 597 1363 643
rect 1409 597 1487 643
rect 1533 597 1611 643
rect 1657 597 1735 643
rect 1781 597 1859 643
rect 1905 597 1983 643
rect 2029 597 2107 643
rect 2153 597 2231 643
rect 2277 597 2355 643
rect 2401 597 2479 643
rect 2525 597 2603 643
rect 2649 597 2727 643
rect 2773 597 2851 643
rect 2897 597 2975 643
rect 3021 597 3099 643
rect 3145 597 3223 643
rect 3269 597 3347 643
rect 3393 597 3471 643
rect 3517 597 3595 643
rect 3641 597 3719 643
rect 3765 597 3843 643
rect 3889 597 3967 643
rect 4013 597 4091 643
rect 4137 597 4215 643
rect 4261 597 4339 643
rect 4385 597 4463 643
rect 4509 597 4587 643
rect 4633 597 4711 643
rect 4757 597 4835 643
rect 4881 597 4959 643
rect 5005 597 5083 643
rect 5129 597 5207 643
rect 5253 597 5331 643
rect 5377 597 5455 643
rect 5501 597 5579 643
rect 5625 597 5703 643
rect 5749 597 5827 643
rect 5873 597 5951 643
rect 5997 597 6075 643
rect 6121 597 6199 643
rect 6245 597 6323 643
rect 6369 597 6447 643
rect 6493 597 6571 643
rect 6617 597 6695 643
rect 6741 597 6819 643
rect 6865 597 6943 643
rect 6989 597 7067 643
rect 7113 597 7191 643
rect 7237 597 7315 643
rect 7361 597 7439 643
rect 7485 597 7563 643
rect 7609 597 7687 643
rect 7733 597 7811 643
rect 7857 597 7935 643
rect 7981 597 8059 643
rect 8105 597 8183 643
rect 8229 597 8307 643
rect 8353 597 8431 643
rect 8477 597 8555 643
rect 8601 597 8679 643
rect 8725 597 8803 643
rect 8849 597 8927 643
rect 8973 597 9051 643
rect 9097 597 9175 643
rect 9221 597 9299 643
rect 9345 597 9423 643
rect 9469 597 9547 643
rect 9593 597 9671 643
rect 9717 597 9795 643
rect 9841 597 9919 643
rect 9965 597 10043 643
rect 10089 597 10167 643
rect 10213 597 10291 643
rect 10337 597 10415 643
rect 10461 597 10539 643
rect 10585 597 10663 643
rect 10709 597 10787 643
rect 10833 597 10911 643
rect 10957 597 11035 643
rect 11081 597 11159 643
rect 11205 597 11283 643
rect 11329 597 11407 643
rect 11453 597 11531 643
rect 11577 597 11655 643
rect 11701 597 11779 643
rect 11825 597 11903 643
rect 11949 597 12027 643
rect 12073 597 12151 643
rect 12197 597 12275 643
rect 12321 597 12399 643
rect 12445 597 12523 643
rect 12569 597 12647 643
rect 12693 597 12771 643
rect 12817 597 12895 643
rect 12941 597 13019 643
rect 13065 597 13143 643
rect 13189 597 13267 643
rect 13313 597 13391 643
rect 13437 597 13515 643
rect 13561 597 13639 643
rect 13685 597 13763 643
rect 13809 597 13887 643
rect 13933 597 14011 643
rect 14057 597 14135 643
rect 14181 597 14259 643
rect 14305 597 14383 643
rect 14429 597 14507 643
rect 14553 597 14631 643
rect 14677 597 14755 643
rect 14801 597 14879 643
rect 14925 597 15003 643
rect 15049 597 15127 643
rect 15173 597 15251 643
rect 15297 597 15375 643
rect 15421 597 15499 643
rect 15545 597 15623 643
rect 15669 597 15747 643
rect 15793 597 15871 643
rect 15917 597 15995 643
rect 16041 597 16119 643
rect 16165 597 16243 643
rect 16289 597 16367 643
rect 16413 597 16491 643
rect 16537 597 16615 643
rect 16661 597 16739 643
rect 16785 597 16863 643
rect 16909 597 16987 643
rect 17033 597 17111 643
rect 17157 597 17235 643
rect 17281 597 17359 643
rect 17405 597 17483 643
rect 17529 597 17607 643
rect 17653 597 17731 643
rect 17777 597 17855 643
rect 17901 597 17979 643
rect 18025 597 18103 643
rect 18149 597 18227 643
rect 18273 597 18351 643
rect 18397 597 18475 643
rect 18521 597 18599 643
rect 18645 597 18723 643
rect 18769 597 18847 643
rect 18893 597 18971 643
rect 19017 597 19095 643
rect 19141 597 19219 643
rect 19265 597 19343 643
rect 19389 597 19467 643
rect 19513 597 19591 643
rect 19637 597 19715 643
rect 19761 597 19839 643
rect 19885 597 19963 643
rect 20009 597 20087 643
rect 20133 597 20211 643
rect 20257 597 20335 643
rect 20381 597 20459 643
rect 20505 597 20583 643
rect 20629 597 20707 643
rect 20753 597 20831 643
rect 20877 597 20955 643
rect 21001 597 21079 643
rect 21125 597 21203 643
rect 21249 597 21327 643
rect 21373 597 21451 643
rect 21497 597 21575 643
rect 21621 597 21699 643
rect 21745 597 21823 643
rect 21869 597 21947 643
rect 21993 597 22071 643
rect 22117 597 22195 643
rect 22241 597 22319 643
rect 22365 597 22443 643
rect 22489 597 22567 643
rect 22613 597 22691 643
rect 22737 597 22815 643
rect 22861 597 22939 643
rect 22985 597 23063 643
rect 23109 597 23187 643
rect 23233 597 23311 643
rect 23357 597 23435 643
rect 23481 597 23559 643
rect 23605 597 23683 643
rect 23729 597 23807 643
rect 23853 597 23931 643
rect 23977 597 24055 643
rect 24101 597 24179 643
rect 24225 597 24303 643
rect 24349 597 24427 643
rect 24473 597 24551 643
rect 24597 597 24675 643
rect 24721 597 24799 643
rect 24845 597 24923 643
rect 24969 597 25047 643
rect 25093 597 25171 643
rect 25217 597 25295 643
rect 25341 597 25419 643
rect 25465 597 25543 643
rect 25589 597 25667 643
rect 25713 597 25791 643
rect 25837 597 25915 643
rect 25961 597 26039 643
rect 26085 597 26163 643
rect 26209 597 26287 643
rect 26333 597 26411 643
rect 26457 597 26535 643
rect 26581 597 26659 643
rect 26705 597 26783 643
rect 26829 597 26907 643
rect 26953 597 27031 643
rect 27077 597 27155 643
rect 27201 597 27279 643
rect 27325 597 27403 643
rect 27449 597 27527 643
rect 27573 597 27651 643
rect 27697 597 27775 643
rect 27821 597 27899 643
rect 27945 597 28023 643
rect 28069 597 28147 643
rect 28193 597 28271 643
rect 28317 597 28395 643
rect 28441 597 28519 643
rect 28565 597 28643 643
rect 28689 597 28767 643
rect 28813 597 28891 643
rect 28937 597 29015 643
rect 29061 597 29139 643
rect 29185 597 29263 643
rect 29309 597 29387 643
rect 29433 597 29511 643
rect 29557 597 29635 643
rect 29681 597 29759 643
rect 29805 597 29883 643
rect 29929 597 30007 643
rect 30053 597 30131 643
rect 30177 597 30255 643
rect 30301 597 30379 643
rect 30425 597 30503 643
rect 30549 597 30627 643
rect 30673 597 30751 643
rect 30797 597 30875 643
rect 30921 597 30999 643
rect 31045 597 31123 643
rect 31169 597 31247 643
rect 31293 597 31371 643
rect 31417 597 31495 643
rect 31541 597 31619 643
rect 31665 597 31743 643
rect 31789 597 31867 643
rect 31913 597 31991 643
rect 32037 597 32115 643
rect 32161 597 32239 643
rect 32285 597 32363 643
rect 32409 597 32487 643
rect 32533 597 32611 643
rect 32657 597 32735 643
rect 32781 597 32859 643
rect 32905 597 32983 643
rect 33029 597 33107 643
rect 33153 597 33231 643
rect 33277 597 33355 643
rect 33401 597 33479 643
rect 33525 597 33603 643
rect 33649 597 33727 643
rect 33773 597 33851 643
rect 33897 597 33975 643
rect 34021 597 34099 643
rect 34145 597 34223 643
rect 34269 597 34347 643
rect 34393 597 34471 643
rect 34517 597 34595 643
rect 34641 597 34719 643
rect 34765 597 34843 643
rect 34889 597 34967 643
rect 35013 597 35091 643
rect 35137 597 35215 643
rect 35261 597 35339 643
rect 35385 597 35463 643
rect 35509 597 35587 643
rect 35633 597 35711 643
rect 35757 597 35835 643
rect 35881 597 35959 643
rect 36005 597 36083 643
rect 36129 597 36207 643
rect 36253 597 36331 643
rect 36377 597 36455 643
rect 36501 597 36579 643
rect 36625 597 36703 643
rect 36749 597 36827 643
rect 36873 597 36951 643
rect 36997 597 37075 643
rect 37121 597 37199 643
rect 37245 597 37323 643
rect 37369 597 37447 643
rect 37493 597 37571 643
rect 37617 597 37695 643
rect 37741 597 37819 643
rect 37865 597 37943 643
rect 37989 597 38067 643
rect 38113 597 38191 643
rect 38237 597 38315 643
rect 38361 597 38439 643
rect 38485 597 38563 643
rect 38609 597 38687 643
rect 38733 597 38811 643
rect 38857 597 38935 643
rect 38981 597 39059 643
rect 39105 597 39183 643
rect 39229 597 39307 643
rect 39353 597 39431 643
rect 39477 597 39555 643
rect 39601 597 39679 643
rect 39725 597 39803 643
rect 39849 597 39927 643
rect 39973 597 40051 643
rect 40097 597 40175 643
rect 40221 597 40299 643
rect 40345 597 40423 643
rect 40469 597 40547 643
rect 40593 597 40671 643
rect 40717 597 40795 643
rect 40841 597 40919 643
rect 40965 597 41043 643
rect 41089 597 41167 643
rect 41213 597 41291 643
rect 41337 597 41415 643
rect 41461 597 41539 643
rect 41585 597 41663 643
rect 41709 597 41787 643
rect 41833 597 41911 643
rect 41957 597 42035 643
rect 42081 597 42159 643
rect 42205 597 42283 643
rect 42329 597 42407 643
rect 42453 597 42531 643
rect 42577 597 42655 643
rect 42701 597 42779 643
rect 42825 597 42903 643
rect 42949 597 43027 643
rect 43073 597 43151 643
rect 43197 597 43275 643
rect 43321 597 43399 643
rect 43445 597 43523 643
rect 43569 597 43647 643
rect 43693 597 43771 643
rect 43817 597 43895 643
rect 43941 597 44019 643
rect 44065 597 44143 643
rect 44189 597 44267 643
rect 44313 597 44391 643
rect 44437 597 44515 643
rect 44561 597 44639 643
rect 44685 597 44763 643
rect 44809 597 44887 643
rect 44933 597 45011 643
rect 45057 597 45135 643
rect 45181 597 45259 643
rect 45305 597 45383 643
rect 45429 597 45507 643
rect 45553 597 45631 643
rect 45677 597 45755 643
rect 45801 597 45879 643
rect 45925 597 46003 643
rect 46049 597 46127 643
rect 46173 597 46251 643
rect 46297 597 46375 643
rect 46421 597 46499 643
rect 46545 597 46623 643
rect 46669 597 46747 643
rect 46793 597 46871 643
rect 46917 597 46995 643
rect 47041 597 47119 643
rect 47165 597 47243 643
rect 47289 597 47367 643
rect 47413 597 47491 643
rect 47537 597 47615 643
rect 47661 597 47739 643
rect 47785 597 47863 643
rect 47909 597 47987 643
rect 48033 597 48111 643
rect 48157 597 48235 643
rect 48281 597 48359 643
rect 48405 597 48483 643
rect 48529 597 48607 643
rect 48653 597 48731 643
rect 48777 597 48855 643
rect 48901 597 48979 643
rect 49025 597 49103 643
rect 49149 597 49227 643
rect 49273 597 49351 643
rect 49397 597 49475 643
rect 49521 597 49599 643
rect 49645 597 49723 643
rect 49769 597 49847 643
rect 49893 597 49971 643
rect 50017 597 50095 643
rect 50141 597 50219 643
rect 50265 597 50343 643
rect 50389 597 50467 643
rect 50513 597 50591 643
rect 50637 597 50715 643
rect 50761 597 50839 643
rect 50885 597 50963 643
rect 51009 597 51087 643
rect 51133 597 51211 643
rect 51257 597 51335 643
rect 51381 597 51459 643
rect 51505 597 51583 643
rect 51629 597 51707 643
rect 51753 597 51831 643
rect 51877 597 51955 643
rect 52001 597 52079 643
rect 52125 597 52203 643
rect 52249 597 52327 643
rect 52373 597 52451 643
rect 52497 597 52575 643
rect 52621 597 52699 643
rect 52745 597 52823 643
rect 52869 597 52947 643
rect 52993 597 53071 643
rect 53117 597 53195 643
rect 53241 597 53319 643
rect 53365 597 53443 643
rect 53489 597 53567 643
rect 53613 597 53691 643
rect 53737 597 53815 643
rect 53861 597 53939 643
rect 53985 597 54063 643
rect 54109 597 54187 643
rect 54233 597 54311 643
rect 54357 597 54435 643
rect 54481 597 54559 643
rect 54605 597 54683 643
rect 54729 597 54807 643
rect 54853 597 54931 643
rect 54977 597 55055 643
rect 55101 597 55179 643
rect 55225 597 55303 643
rect 55349 597 55427 643
rect 55473 597 55551 643
rect 55597 597 55675 643
rect 55721 597 55799 643
rect 55845 597 55923 643
rect 55969 597 56047 643
rect 56093 597 56171 643
rect 56217 597 56295 643
rect 56341 597 56419 643
rect 56465 597 56543 643
rect 56589 597 56667 643
rect 56713 597 56791 643
rect 56837 597 56915 643
rect 56961 597 57039 643
rect 57085 597 57163 643
rect 57209 597 57287 643
rect 57333 597 57411 643
rect 57457 597 57535 643
rect 57581 597 57659 643
rect 57705 597 57783 643
rect 57829 597 57907 643
rect 57953 597 58031 643
rect 58077 597 58155 643
rect 58201 597 58279 643
rect 58325 597 58403 643
rect 58449 597 58527 643
rect 58573 597 58651 643
rect 58697 597 58775 643
rect 58821 597 58899 643
rect 58945 597 59023 643
rect 59069 597 59147 643
rect 59193 597 59271 643
rect 59317 597 59395 643
rect 59441 597 59519 643
rect 59565 597 59643 643
rect 59689 597 59767 643
rect 59813 597 59891 643
rect 59937 597 60015 643
rect 60061 597 60139 643
rect 60185 597 60263 643
rect 60309 597 60387 643
rect 60433 597 60511 643
rect 60557 597 60635 643
rect 60681 597 60759 643
rect 60805 597 60883 643
rect 60929 597 61007 643
rect 61053 597 61131 643
rect 61177 597 61255 643
rect 61301 597 61379 643
rect 61425 597 61503 643
rect 61549 597 61627 643
rect 61673 597 61751 643
rect 61797 597 61875 643
rect 61921 597 61999 643
rect 62045 597 62123 643
rect 62169 597 62247 643
rect 62293 597 62371 643
rect 62417 597 62495 643
rect 62541 597 62619 643
rect 62665 597 62743 643
rect 62789 597 62867 643
rect 62913 597 62991 643
rect 63037 597 63115 643
rect 63161 597 63239 643
rect 63285 597 63363 643
rect 63409 597 63487 643
rect 63533 597 63611 643
rect 63657 597 63735 643
rect 63781 597 63859 643
rect 63905 597 63983 643
rect 64029 597 64107 643
rect 64153 597 64231 643
rect 64277 597 64355 643
rect 64401 597 64479 643
rect 64525 597 64603 643
rect 64649 597 64727 643
rect 64773 597 64851 643
rect 64897 597 64975 643
rect 65021 597 65099 643
rect 65145 597 65223 643
rect 65269 597 65347 643
rect 65393 597 65471 643
rect 65517 597 65595 643
rect 65641 597 65719 643
rect 65765 597 65843 643
rect 65889 597 65967 643
rect 66013 597 66091 643
rect 66137 597 66215 643
rect 66261 597 66339 643
rect 66385 597 66463 643
rect 66509 597 66587 643
rect 66633 597 66711 643
rect 66757 597 66835 643
rect 66881 597 66959 643
rect 67005 597 67083 643
rect 67129 597 67207 643
rect 67253 597 67331 643
rect 67377 597 67455 643
rect 67501 597 67579 643
rect 67625 597 67703 643
rect 67749 597 67827 643
rect 67873 597 67951 643
rect 67997 597 68075 643
rect 68121 597 68199 643
rect 68245 597 68323 643
rect 68369 597 68447 643
rect 68493 597 68571 643
rect 68617 597 68695 643
rect 68741 597 68819 643
rect 68865 597 68943 643
rect 68989 597 69067 643
rect 69113 597 69191 643
rect 69237 597 69315 643
rect 69361 597 69439 643
rect 69485 597 69563 643
rect 69609 597 69687 643
rect 69733 597 69811 643
rect 69857 597 69935 643
rect 69981 597 70059 643
rect 70105 597 70183 643
rect 70229 597 70307 643
rect 70353 597 70431 643
rect 70477 597 70555 643
rect 70601 597 70679 643
rect 70725 597 70803 643
rect 70849 597 70927 643
rect 70973 597 71051 643
rect 71097 597 71175 643
rect 71221 597 71299 643
rect 71345 597 71423 643
rect 71469 597 71547 643
rect 71593 597 71671 643
rect 71717 597 71795 643
rect 71841 597 71919 643
rect 71965 597 72043 643
rect 72089 597 72167 643
rect 72213 597 72291 643
rect 72337 597 72415 643
rect 72461 597 72539 643
rect 72585 597 72663 643
rect 72709 597 72787 643
rect 72833 597 72911 643
rect 72957 597 73035 643
rect 73081 597 73159 643
rect 73205 597 73283 643
rect 73329 597 73407 643
rect 73453 597 73531 643
rect 73577 597 73655 643
rect 73701 597 73779 643
rect 73825 597 73903 643
rect 73949 597 74027 643
rect 74073 597 74151 643
rect 74197 597 74275 643
rect 74321 597 74399 643
rect 74445 597 74523 643
rect 74569 597 74647 643
rect 74693 597 74771 643
rect 74817 597 74895 643
rect 74941 597 75019 643
rect 75065 597 75143 643
rect 75189 597 75267 643
rect 75313 597 75391 643
rect 75437 597 75515 643
rect 75561 597 75639 643
rect 75685 597 75763 643
rect 75809 597 75887 643
rect 75933 597 76011 643
rect 76057 597 76135 643
rect 76181 597 76259 643
rect 76305 597 76383 643
rect 76429 597 76507 643
rect 76553 597 76631 643
rect 76677 597 76755 643
rect 76801 597 76879 643
rect 76925 597 77003 643
rect 77049 597 77127 643
rect 77173 597 77251 643
rect 77297 597 77375 643
rect 77421 597 77499 643
rect 77545 597 77623 643
rect 77669 597 77747 643
rect 77793 597 77871 643
rect 77917 597 77995 643
rect 78041 597 78119 643
rect 78165 597 78243 643
rect 78289 597 78367 643
rect 78413 597 78491 643
rect 78537 597 78615 643
rect 78661 597 78739 643
rect 78785 597 78863 643
rect 78909 597 78987 643
rect 79033 597 79111 643
rect 79157 597 79235 643
rect 79281 597 79359 643
rect 79405 597 79483 643
rect 79529 597 79607 643
rect 79653 597 79731 643
rect 79777 597 79855 643
rect 79901 597 79979 643
rect 80025 597 80103 643
rect 80149 597 80227 643
rect 80273 597 80351 643
rect 80397 597 80475 643
rect 80521 597 80599 643
rect 80645 597 80723 643
rect 80769 597 80847 643
rect 80893 597 80971 643
rect 81017 597 81095 643
rect 81141 597 81219 643
rect 81265 597 81343 643
rect 81389 597 81467 643
rect 81513 597 81591 643
rect 81637 597 81715 643
rect 81761 597 81839 643
rect 81885 597 81963 643
rect 82009 597 82087 643
rect 82133 597 82211 643
rect 82257 597 82335 643
rect 82381 597 82459 643
rect 82505 597 82583 643
rect 82629 597 82707 643
rect 82753 597 82831 643
rect 82877 597 82955 643
rect 83001 597 83079 643
rect 83125 597 83203 643
rect 83249 597 83327 643
rect 83373 597 83451 643
rect 83497 597 83575 643
rect 83621 597 83699 643
rect 83745 597 83823 643
rect 83869 597 83947 643
rect 83993 597 84071 643
rect 84117 597 84195 643
rect 84241 597 84319 643
rect 84365 597 84443 643
rect 84489 597 84567 643
rect 84613 597 84691 643
rect 84737 597 84815 643
rect 84861 597 84939 643
rect 84985 597 85063 643
rect 85109 597 85187 643
rect 85233 597 85311 643
rect 85357 597 85435 643
rect 85481 597 85559 643
rect 85605 597 85683 643
rect 85729 597 85807 643
rect 85853 597 85931 643
rect 85977 597 86090 643
rect 282 282 86090 597
<< via1 >>
rect 25388 94721 25440 94773
rect 25512 94721 25564 94773
rect 25636 94721 25688 94773
rect 25760 94721 25812 94773
rect 25884 94721 25936 94773
rect 25388 94597 25440 94649
rect 25512 94597 25564 94649
rect 25636 94597 25688 94649
rect 25760 94597 25812 94649
rect 25884 94597 25936 94649
rect 25388 94473 25440 94525
rect 25512 94473 25564 94525
rect 25636 94473 25688 94525
rect 25760 94473 25812 94525
rect 25884 94473 25936 94525
rect 25388 34938 25440 34990
rect 25512 34938 25564 34990
rect 25636 34938 25688 34990
rect 25760 34938 25812 34990
rect 25884 34938 25936 34990
rect 25388 34814 25440 34866
rect 25512 34814 25564 34866
rect 25636 34814 25688 34866
rect 25760 34814 25812 34866
rect 25884 34814 25936 34866
rect 25388 34690 25440 34742
rect 25512 34690 25564 34742
rect 25636 34690 25688 34742
rect 25760 34690 25812 34742
rect 25884 34690 25936 34742
rect 27790 94601 27822 94653
rect 27822 94601 27842 94653
rect 28001 94601 28053 94653
rect 28212 94601 28264 94653
rect 28423 94601 28475 94653
rect 28634 94601 28668 94653
rect 28668 94601 28686 94653
rect 28845 94601 28897 94653
rect 29056 94601 29108 94653
rect 56015 94601 56067 94653
rect 56226 94601 56278 94653
rect 56437 94601 56489 94653
rect 56648 94601 56700 94653
rect 56859 94601 56911 94653
rect 57070 94601 57122 94653
rect 57281 94601 57306 94653
rect 57306 94601 57333 94653
rect 27790 92801 27822 92853
rect 27822 92801 27842 92853
rect 28001 92801 28053 92853
rect 28212 92801 28264 92853
rect 28423 92801 28475 92853
rect 28634 92801 28668 92853
rect 28668 92801 28686 92853
rect 28845 92801 28897 92853
rect 29056 92801 29108 92853
rect 27790 91001 27822 91053
rect 27822 91001 27842 91053
rect 28001 91001 28053 91053
rect 28212 91001 28264 91053
rect 28423 91001 28475 91053
rect 28634 91001 28668 91053
rect 28668 91001 28686 91053
rect 28845 91001 28897 91053
rect 29056 91001 29108 91053
rect 27790 89201 27822 89253
rect 27822 89201 27842 89253
rect 28001 89201 28053 89253
rect 28212 89201 28264 89253
rect 28423 89201 28475 89253
rect 28634 89201 28668 89253
rect 28668 89201 28686 89253
rect 28845 89201 28897 89253
rect 29056 89201 29108 89253
rect 27790 87401 27822 87453
rect 27822 87401 27842 87453
rect 28001 87401 28053 87453
rect 28212 87401 28264 87453
rect 28423 87401 28475 87453
rect 28634 87401 28668 87453
rect 28668 87401 28686 87453
rect 28845 87401 28897 87453
rect 29056 87401 29108 87453
rect 27790 85601 27822 85653
rect 27822 85601 27842 85653
rect 28001 85601 28053 85653
rect 28212 85601 28264 85653
rect 28423 85601 28475 85653
rect 28634 85601 28668 85653
rect 28668 85601 28686 85653
rect 28845 85601 28897 85653
rect 29056 85601 29108 85653
rect 27790 83801 27822 83853
rect 27822 83801 27842 83853
rect 28001 83801 28053 83853
rect 28212 83801 28264 83853
rect 28423 83801 28475 83853
rect 28634 83801 28668 83853
rect 28668 83801 28686 83853
rect 28845 83801 28897 83853
rect 29056 83801 29108 83853
rect 27790 82001 27822 82053
rect 27822 82001 27842 82053
rect 28001 82001 28053 82053
rect 28212 82001 28264 82053
rect 28423 82001 28475 82053
rect 28634 82001 28668 82053
rect 28668 82001 28686 82053
rect 28845 82001 28897 82053
rect 29056 82001 29108 82053
rect 27790 80201 27822 80253
rect 27822 80201 27842 80253
rect 28001 80201 28053 80253
rect 28212 80201 28264 80253
rect 28423 80201 28475 80253
rect 28634 80201 28668 80253
rect 28668 80201 28686 80253
rect 28845 80201 28897 80253
rect 29056 80201 29108 80253
rect 27790 78401 27822 78453
rect 27822 78401 27842 78453
rect 28001 78401 28053 78453
rect 28212 78401 28264 78453
rect 28423 78401 28475 78453
rect 28634 78401 28668 78453
rect 28668 78401 28686 78453
rect 28845 78401 28897 78453
rect 29056 78401 29108 78453
rect 27790 76601 27822 76653
rect 27822 76601 27842 76653
rect 28001 76601 28053 76653
rect 28212 76601 28264 76653
rect 28423 76601 28475 76653
rect 28634 76601 28668 76653
rect 28668 76601 28686 76653
rect 28845 76601 28897 76653
rect 29056 76601 29108 76653
rect 27790 74801 27822 74853
rect 27822 74801 27842 74853
rect 28001 74801 28053 74853
rect 28212 74801 28264 74853
rect 28423 74801 28475 74853
rect 28634 74801 28668 74853
rect 28668 74801 28686 74853
rect 28845 74801 28897 74853
rect 29056 74801 29108 74853
rect 27790 73001 27822 73053
rect 27822 73001 27842 73053
rect 28001 73001 28053 73053
rect 28212 73001 28264 73053
rect 28423 73001 28475 73053
rect 28634 73001 28668 73053
rect 28668 73001 28686 73053
rect 28845 73001 28897 73053
rect 29056 73001 29108 73053
rect 27790 71201 27822 71253
rect 27822 71201 27842 71253
rect 28001 71201 28053 71253
rect 28212 71201 28264 71253
rect 28423 71201 28475 71253
rect 28634 71201 28668 71253
rect 28668 71201 28686 71253
rect 28845 71201 28897 71253
rect 29056 71201 29108 71253
rect 27790 69401 27822 69453
rect 27822 69401 27842 69453
rect 28001 69401 28053 69453
rect 28212 69401 28264 69453
rect 28423 69401 28475 69453
rect 28634 69401 28668 69453
rect 28668 69401 28686 69453
rect 28845 69401 28897 69453
rect 29056 69401 29108 69453
rect 27790 67601 27822 67653
rect 27822 67601 27842 67653
rect 28001 67601 28053 67653
rect 28212 67601 28264 67653
rect 28423 67601 28475 67653
rect 28634 67601 28668 67653
rect 28668 67601 28686 67653
rect 28845 67601 28897 67653
rect 29056 67601 29108 67653
rect 27790 65801 27822 65853
rect 27822 65801 27842 65853
rect 28001 65801 28053 65853
rect 28212 65801 28264 65853
rect 28423 65801 28475 65853
rect 28634 65801 28668 65853
rect 28668 65801 28686 65853
rect 28845 65801 28897 65853
rect 29056 65801 29108 65853
rect 27790 64001 27822 64053
rect 27822 64001 27842 64053
rect 28001 64001 28053 64053
rect 28212 64001 28264 64053
rect 28423 64001 28475 64053
rect 28634 64001 28668 64053
rect 28668 64001 28686 64053
rect 28845 64001 28897 64053
rect 29056 64001 29108 64053
rect 27790 62201 27822 62253
rect 27822 62201 27842 62253
rect 28001 62201 28053 62253
rect 28212 62201 28264 62253
rect 28423 62201 28475 62253
rect 28634 62201 28668 62253
rect 28668 62201 28686 62253
rect 28845 62201 28897 62253
rect 29056 62201 29108 62253
rect 27790 60401 27822 60453
rect 27822 60401 27842 60453
rect 28001 60401 28053 60453
rect 28212 60401 28264 60453
rect 28423 60401 28475 60453
rect 28634 60401 28668 60453
rect 28668 60401 28686 60453
rect 28845 60401 28897 60453
rect 29056 60401 29108 60453
rect 27790 58601 27822 58653
rect 27822 58601 27842 58653
rect 28001 58601 28053 58653
rect 28212 58601 28264 58653
rect 28423 58601 28475 58653
rect 28634 58601 28668 58653
rect 28668 58601 28686 58653
rect 28845 58601 28897 58653
rect 29056 58601 29108 58653
rect 27790 56801 27822 56853
rect 27822 56801 27842 56853
rect 28001 56801 28053 56853
rect 28212 56801 28264 56853
rect 28423 56801 28475 56853
rect 28634 56801 28668 56853
rect 28668 56801 28686 56853
rect 28845 56801 28897 56853
rect 29056 56801 29108 56853
rect 27790 55001 27822 55053
rect 27822 55001 27842 55053
rect 28001 55001 28053 55053
rect 28212 55001 28264 55053
rect 28423 55001 28475 55053
rect 28634 55001 28668 55053
rect 28668 55001 28686 55053
rect 28845 55001 28897 55053
rect 29056 55001 29108 55053
rect 27790 53201 27822 53253
rect 27822 53201 27842 53253
rect 28001 53201 28053 53253
rect 28212 53201 28264 53253
rect 28423 53201 28475 53253
rect 28634 53201 28668 53253
rect 28668 53201 28686 53253
rect 28845 53201 28897 53253
rect 29056 53201 29108 53253
rect 27790 51401 27822 51453
rect 27822 51401 27842 51453
rect 28001 51401 28053 51453
rect 28212 51401 28264 51453
rect 28423 51401 28475 51453
rect 28634 51401 28668 51453
rect 28668 51401 28686 51453
rect 28845 51401 28897 51453
rect 29056 51401 29108 51453
rect 27790 49601 27822 49653
rect 27822 49601 27842 49653
rect 28001 49601 28053 49653
rect 28212 49601 28264 49653
rect 28423 49601 28475 49653
rect 28634 49601 28668 49653
rect 28668 49601 28686 49653
rect 28845 49601 28897 49653
rect 29056 49601 29108 49653
rect 27790 47801 27822 47853
rect 27822 47801 27842 47853
rect 28001 47801 28053 47853
rect 28212 47801 28264 47853
rect 28423 47801 28475 47853
rect 28634 47801 28668 47853
rect 28668 47801 28686 47853
rect 28845 47801 28897 47853
rect 29056 47801 29108 47853
rect 27790 46001 27822 46053
rect 27822 46001 27842 46053
rect 28001 46001 28053 46053
rect 28212 46001 28264 46053
rect 28423 46001 28475 46053
rect 28634 46001 28668 46053
rect 28668 46001 28686 46053
rect 28845 46001 28897 46053
rect 29056 46001 29108 46053
rect 27790 44201 27822 44253
rect 27822 44201 27842 44253
rect 28001 44201 28053 44253
rect 28212 44201 28264 44253
rect 28423 44201 28475 44253
rect 28634 44201 28668 44253
rect 28668 44201 28686 44253
rect 28845 44201 28897 44253
rect 29056 44201 29108 44253
rect 27790 42401 27822 42453
rect 27822 42401 27842 42453
rect 28001 42401 28053 42453
rect 28212 42401 28264 42453
rect 28423 42401 28475 42453
rect 28634 42401 28668 42453
rect 28668 42401 28686 42453
rect 28845 42401 28897 42453
rect 29056 42401 29108 42453
rect 27790 40601 27822 40653
rect 27822 40601 27842 40653
rect 28001 40601 28053 40653
rect 28212 40601 28264 40653
rect 28423 40601 28475 40653
rect 28634 40601 28668 40653
rect 28668 40601 28686 40653
rect 28845 40601 28897 40653
rect 29056 40601 29108 40653
rect 27790 38801 27822 38853
rect 27822 38801 27842 38853
rect 28001 38801 28053 38853
rect 28212 38801 28264 38853
rect 28423 38801 28475 38853
rect 28634 38801 28668 38853
rect 28668 38801 28686 38853
rect 28845 38801 28897 38853
rect 29056 38801 29108 38853
rect 27790 37001 27822 37053
rect 27822 37001 27842 37053
rect 28001 37001 28053 37053
rect 28212 37001 28264 37053
rect 28423 37001 28475 37053
rect 28634 37001 28668 37053
rect 28668 37001 28686 37053
rect 28845 37001 28897 37053
rect 29056 37001 29108 37053
rect 56015 92801 56067 92853
rect 56226 92801 56278 92853
rect 56437 92801 56489 92853
rect 56648 92801 56700 92853
rect 56859 92801 56911 92853
rect 57070 92801 57122 92853
rect 57281 92801 57306 92853
rect 57306 92801 57333 92853
rect 56015 91001 56067 91053
rect 56226 91001 56278 91053
rect 56437 91001 56489 91053
rect 56648 91001 56700 91053
rect 56859 91001 56911 91053
rect 57070 91001 57122 91053
rect 57281 91001 57306 91053
rect 57306 91001 57333 91053
rect 56015 89201 56067 89253
rect 56226 89201 56278 89253
rect 56437 89201 56489 89253
rect 56648 89201 56700 89253
rect 56859 89201 56911 89253
rect 57070 89201 57122 89253
rect 57281 89201 57306 89253
rect 57306 89201 57333 89253
rect 56015 87401 56067 87453
rect 56226 87401 56278 87453
rect 56437 87401 56489 87453
rect 56648 87401 56700 87453
rect 56859 87401 56911 87453
rect 57070 87401 57122 87453
rect 57281 87401 57306 87453
rect 57306 87401 57333 87453
rect 56015 85601 56067 85653
rect 56226 85601 56278 85653
rect 56437 85601 56489 85653
rect 56648 85601 56700 85653
rect 56859 85601 56911 85653
rect 57070 85601 57122 85653
rect 57281 85601 57306 85653
rect 57306 85601 57333 85653
rect 56015 83801 56067 83853
rect 56226 83801 56278 83853
rect 56437 83801 56489 83853
rect 56648 83801 56700 83853
rect 56859 83801 56911 83853
rect 57070 83801 57122 83853
rect 57281 83801 57306 83853
rect 57306 83801 57333 83853
rect 56015 82001 56067 82053
rect 56226 82001 56278 82053
rect 56437 82001 56489 82053
rect 56648 82001 56700 82053
rect 56859 82001 56911 82053
rect 57070 82001 57122 82053
rect 57281 82001 57306 82053
rect 57306 82001 57333 82053
rect 56015 80201 56067 80253
rect 56226 80201 56278 80253
rect 56437 80201 56489 80253
rect 56648 80201 56700 80253
rect 56859 80201 56911 80253
rect 57070 80201 57122 80253
rect 57281 80201 57306 80253
rect 57306 80201 57333 80253
rect 56015 78401 56067 78453
rect 56226 78401 56278 78453
rect 56437 78401 56489 78453
rect 56648 78401 56700 78453
rect 56859 78401 56911 78453
rect 57070 78401 57122 78453
rect 57281 78401 57306 78453
rect 57306 78401 57333 78453
rect 56015 76601 56067 76653
rect 56226 76601 56278 76653
rect 56437 76601 56489 76653
rect 56648 76601 56700 76653
rect 56859 76601 56911 76653
rect 57070 76601 57122 76653
rect 57281 76601 57306 76653
rect 57306 76601 57333 76653
rect 56015 74801 56067 74853
rect 56226 74801 56278 74853
rect 56437 74801 56489 74853
rect 56648 74801 56700 74853
rect 56859 74801 56911 74853
rect 57070 74801 57122 74853
rect 57281 74801 57306 74853
rect 57306 74801 57333 74853
rect 56015 73001 56067 73053
rect 56226 73001 56278 73053
rect 56437 73001 56489 73053
rect 56648 73001 56700 73053
rect 56859 73001 56911 73053
rect 57070 73001 57122 73053
rect 57281 73001 57306 73053
rect 57306 73001 57333 73053
rect 56015 71201 56067 71253
rect 56226 71201 56278 71253
rect 56437 71201 56489 71253
rect 56648 71201 56700 71253
rect 56859 71201 56911 71253
rect 57070 71201 57122 71253
rect 57281 71201 57306 71253
rect 57306 71201 57333 71253
rect 56015 69401 56067 69453
rect 56226 69401 56278 69453
rect 56437 69401 56489 69453
rect 56648 69401 56700 69453
rect 56859 69401 56911 69453
rect 57070 69401 57122 69453
rect 57281 69401 57306 69453
rect 57306 69401 57333 69453
rect 56015 67601 56067 67653
rect 56226 67601 56278 67653
rect 56437 67601 56489 67653
rect 56648 67601 56700 67653
rect 56859 67601 56911 67653
rect 57070 67601 57122 67653
rect 57281 67601 57306 67653
rect 57306 67601 57333 67653
rect 56015 65801 56067 65853
rect 56226 65801 56278 65853
rect 56437 65801 56489 65853
rect 56648 65801 56700 65853
rect 56859 65801 56911 65853
rect 57070 65801 57122 65853
rect 57281 65801 57306 65853
rect 57306 65801 57333 65853
rect 56015 64001 56067 64053
rect 56226 64001 56278 64053
rect 56437 64001 56489 64053
rect 56648 64001 56700 64053
rect 56859 64001 56911 64053
rect 57070 64001 57122 64053
rect 57281 64001 57306 64053
rect 57306 64001 57333 64053
rect 56015 62201 56067 62253
rect 56226 62201 56278 62253
rect 56437 62201 56489 62253
rect 56648 62201 56700 62253
rect 56859 62201 56911 62253
rect 57070 62201 57122 62253
rect 57281 62201 57306 62253
rect 57306 62201 57333 62253
rect 56015 60401 56067 60453
rect 56226 60401 56278 60453
rect 56437 60401 56489 60453
rect 56648 60401 56700 60453
rect 56859 60401 56911 60453
rect 57070 60401 57122 60453
rect 57281 60401 57306 60453
rect 57306 60401 57333 60453
rect 56015 58601 56067 58653
rect 56226 58601 56278 58653
rect 56437 58601 56489 58653
rect 56648 58601 56700 58653
rect 56859 58601 56911 58653
rect 57070 58601 57122 58653
rect 57281 58601 57306 58653
rect 57306 58601 57333 58653
rect 56015 56801 56067 56853
rect 56226 56801 56278 56853
rect 56437 56801 56489 56853
rect 56648 56801 56700 56853
rect 56859 56801 56911 56853
rect 57070 56801 57122 56853
rect 57281 56801 57306 56853
rect 57306 56801 57333 56853
rect 56015 55001 56067 55053
rect 56226 55001 56278 55053
rect 56437 55001 56489 55053
rect 56648 55001 56700 55053
rect 56859 55001 56911 55053
rect 57070 55001 57122 55053
rect 57281 55001 57306 55053
rect 57306 55001 57333 55053
rect 56015 53201 56067 53253
rect 56226 53201 56278 53253
rect 56437 53201 56489 53253
rect 56648 53201 56700 53253
rect 56859 53201 56911 53253
rect 57070 53201 57122 53253
rect 57281 53201 57306 53253
rect 57306 53201 57333 53253
rect 56015 51401 56067 51453
rect 56226 51401 56278 51453
rect 56437 51401 56489 51453
rect 56648 51401 56700 51453
rect 56859 51401 56911 51453
rect 57070 51401 57122 51453
rect 57281 51401 57306 51453
rect 57306 51401 57333 51453
rect 56015 49601 56067 49653
rect 56226 49601 56278 49653
rect 56437 49601 56489 49653
rect 56648 49601 56700 49653
rect 56859 49601 56911 49653
rect 57070 49601 57122 49653
rect 57281 49601 57306 49653
rect 57306 49601 57333 49653
rect 56015 47801 56067 47853
rect 56226 47801 56278 47853
rect 56437 47801 56489 47853
rect 56648 47801 56700 47853
rect 56859 47801 56911 47853
rect 57070 47801 57122 47853
rect 57281 47801 57306 47853
rect 57306 47801 57333 47853
rect 56015 46001 56067 46053
rect 56226 46001 56278 46053
rect 56437 46001 56489 46053
rect 56648 46001 56700 46053
rect 56859 46001 56911 46053
rect 57070 46001 57122 46053
rect 57281 46001 57306 46053
rect 57306 46001 57333 46053
rect 56015 44201 56067 44253
rect 56226 44201 56278 44253
rect 56437 44201 56489 44253
rect 56648 44201 56700 44253
rect 56859 44201 56911 44253
rect 57070 44201 57122 44253
rect 57281 44201 57306 44253
rect 57306 44201 57333 44253
rect 56015 42401 56067 42453
rect 56226 42401 56278 42453
rect 56437 42401 56489 42453
rect 56648 42401 56700 42453
rect 56859 42401 56911 42453
rect 57070 42401 57122 42453
rect 57281 42401 57306 42453
rect 57306 42401 57333 42453
rect 56015 40601 56067 40653
rect 56226 40601 56278 40653
rect 56437 40601 56489 40653
rect 56648 40601 56700 40653
rect 56859 40601 56911 40653
rect 57070 40601 57122 40653
rect 57281 40601 57306 40653
rect 57306 40601 57333 40653
rect 56015 38801 56067 38853
rect 56226 38801 56278 38853
rect 56437 38801 56489 38853
rect 56648 38801 56700 38853
rect 56859 38801 56911 38853
rect 57070 38801 57122 38853
rect 57281 38801 57306 38853
rect 57306 38801 57333 38853
rect 56015 37001 56067 37053
rect 56226 37001 56278 37053
rect 56437 37001 56489 37053
rect 56648 37001 56700 37053
rect 56859 37001 56911 37053
rect 57070 37001 57122 37053
rect 57281 37001 57306 37053
rect 57306 37001 57333 37053
rect 27449 34938 27501 34990
rect 27573 34938 27625 34990
rect 27697 34938 27744 34990
rect 27744 34938 27749 34990
rect 27449 34814 27501 34866
rect 27573 34814 27625 34866
rect 27697 34814 27744 34866
rect 27744 34814 27749 34866
rect 27449 34690 27501 34742
rect 27573 34690 27625 34742
rect 27697 34690 27744 34742
rect 27744 34690 27749 34742
rect 25388 34566 25440 34618
rect 25512 34566 25564 34618
rect 25636 34566 25688 34618
rect 25760 34566 25812 34618
rect 25884 34566 25936 34618
rect 27449 34566 27501 34618
rect 27573 34566 27625 34618
rect 27697 34566 27744 34618
rect 27744 34566 27749 34618
rect 26861 33380 26913 33432
rect 27073 33380 27125 33432
rect 26861 33163 26913 33215
rect 27073 33163 27125 33215
rect 26861 32945 26913 32997
rect 27073 32945 27125 32997
rect 26861 32727 26913 32779
rect 27073 32727 27125 32779
rect 26861 32510 26913 32562
rect 27073 32510 27125 32562
rect 26861 32292 26913 32344
rect 27073 32292 27125 32344
rect 26861 32075 26913 32127
rect 27073 32075 27125 32127
rect 26861 31857 26913 31909
rect 27073 31857 27125 31909
rect 26861 31639 26913 31691
rect 27073 31639 27125 31691
rect 26861 31422 26913 31474
rect 27073 31422 27125 31474
rect 26861 31204 26913 31256
rect 27073 31204 27125 31256
rect 26861 30986 26913 31038
rect 27073 30986 27125 31038
rect 26861 30769 26913 30821
rect 27073 30769 27125 30821
rect 26861 30551 26913 30603
rect 27073 30551 27125 30603
rect 26861 30334 26913 30386
rect 27073 30334 27125 30386
rect 26861 30116 26913 30168
rect 27073 30116 27125 30168
rect 26861 29898 26913 29950
rect 27073 29898 27125 29950
rect 26861 29681 26913 29733
rect 27073 29681 27125 29733
rect 26861 29463 26913 29515
rect 27073 29463 27125 29515
rect 26861 29245 26913 29297
rect 27073 29245 27125 29297
rect 26861 29028 26913 29080
rect 27073 29028 27125 29080
rect 26861 28810 26913 28862
rect 27073 28810 27125 28862
rect 26861 28592 26913 28644
rect 27073 28592 27125 28644
rect 26861 28375 26913 28427
rect 27073 28375 27125 28427
rect 26861 28157 26913 28209
rect 27073 28157 27125 28209
rect 26861 27940 26913 27992
rect 27073 27940 27125 27992
rect 26861 27722 26913 27774
rect 27073 27722 27125 27774
rect 26861 27504 26913 27556
rect 27073 27504 27125 27556
rect 26861 27287 26913 27339
rect 27073 27287 27125 27339
rect 26861 27069 26913 27121
rect 27073 27069 27125 27121
rect 26861 26851 26913 26903
rect 27073 26851 27125 26903
rect 26861 26634 26913 26686
rect 27073 26634 27125 26686
rect 26861 26416 26913 26468
rect 27073 26416 27125 26468
rect 26861 26198 26913 26250
rect 27073 26198 27125 26250
rect 26861 25981 26913 26033
rect 27073 25981 27125 26033
rect 26861 25763 26913 25815
rect 27073 25763 27125 25815
rect 26861 25546 26913 25598
rect 27073 25546 27125 25598
rect 26861 25328 26913 25380
rect 27073 25328 27125 25380
rect 26861 25110 26913 25162
rect 27073 25110 27125 25162
rect 26861 24893 26913 24945
rect 27073 24893 27125 24945
rect 26861 24675 26913 24727
rect 27073 24675 27125 24727
rect 26861 24457 26913 24509
rect 27073 24457 27125 24509
rect 26861 24240 26913 24292
rect 27073 24240 27125 24292
rect 26861 24022 26913 24074
rect 27073 24022 27125 24074
rect 26861 23805 26913 23857
rect 27073 23805 27125 23857
rect 26861 23587 26913 23639
rect 27073 23587 27125 23639
rect 26861 23369 26913 23421
rect 27073 23369 27125 23421
rect 26861 23152 26913 23204
rect 27073 23152 27125 23204
rect 26861 22934 26913 22986
rect 27073 22934 27125 22986
rect 26861 22716 26913 22768
rect 27073 22716 27125 22768
rect 26861 22499 26913 22551
rect 27073 22499 27125 22551
rect 26861 22281 26913 22333
rect 27073 22281 27125 22333
rect 26861 22063 26913 22115
rect 27073 22063 27125 22115
rect 26861 21846 26913 21898
rect 27073 21846 27125 21898
rect 26861 21628 26913 21680
rect 27073 21628 27125 21680
rect 26861 21411 26913 21463
rect 27073 21411 27125 21463
rect 26861 21193 26913 21245
rect 27073 21193 27125 21245
rect 26861 20975 26913 21027
rect 27073 20975 27125 21027
rect 26861 20758 26913 20810
rect 27073 20758 27125 20810
rect 26861 20540 26913 20592
rect 27073 20540 27125 20592
rect 26861 20322 26913 20374
rect 27073 20322 27125 20374
rect 26861 20105 26913 20157
rect 27073 20105 27125 20157
rect 26861 19887 26913 19939
rect 27073 19887 27125 19939
rect 26861 19670 26913 19722
rect 27073 19670 27125 19722
rect 26861 19452 26913 19504
rect 27073 19452 27125 19504
rect 26861 19234 26913 19286
rect 27073 19234 27125 19286
rect 26861 19016 26913 19068
rect 27073 19016 27125 19068
rect 26861 18799 26913 18851
rect 27073 18799 27125 18851
rect 26861 18581 26913 18633
rect 27073 18581 27125 18633
rect 26861 18364 26913 18416
rect 27073 18364 27125 18416
rect 26861 18146 26913 18198
rect 27073 18146 27125 18198
rect 26861 17928 26913 17980
rect 27073 17928 27125 17980
rect 26861 17711 26913 17763
rect 27073 17711 27125 17763
rect 26861 17493 26913 17545
rect 27073 17493 27125 17545
rect 26861 17275 26913 17327
rect 27073 17275 27125 17327
rect 26861 17058 26913 17110
rect 27073 17058 27125 17110
rect 26861 16840 26913 16892
rect 27073 16840 27125 16892
rect 26861 16623 26913 16675
rect 27073 16623 27125 16675
rect 26861 16405 26913 16457
rect 27073 16405 27125 16457
rect 26861 16187 26913 16239
rect 27073 16187 27125 16239
rect 26861 15970 26913 16022
rect 27073 15970 27125 16022
rect 26861 15752 26913 15804
rect 27073 15752 27125 15804
rect 26861 15534 26913 15586
rect 27073 15534 27125 15586
rect 26861 15317 26913 15369
rect 27073 15317 27125 15369
rect 26861 15099 26913 15151
rect 27073 15099 27125 15151
rect 26861 14881 26913 14933
rect 27073 14881 27125 14933
rect 26861 14664 26913 14716
rect 27073 14664 27125 14716
rect 26861 14446 26913 14498
rect 27073 14446 27125 14498
rect 26861 14229 26913 14281
rect 27073 14229 27125 14281
rect 26861 14011 26913 14063
rect 27073 14011 27125 14063
rect 26861 13793 26913 13845
rect 27073 13793 27125 13845
rect 26861 13576 26913 13628
rect 27073 13576 27125 13628
rect 26861 13358 26913 13410
rect 27073 13358 27125 13410
rect 26861 13140 26913 13192
rect 27073 13140 27125 13192
rect 26861 12923 26913 12975
rect 27073 12923 27125 12975
rect 26861 12705 26913 12757
rect 27073 12705 27125 12757
rect 26861 12488 26913 12540
rect 27073 12488 27125 12540
rect 26861 12270 26913 12322
rect 27073 12270 27125 12322
rect 26861 12052 26913 12104
rect 27073 12052 27125 12104
rect 26861 11835 26913 11887
rect 27073 11835 27125 11887
rect 26861 11617 26913 11669
rect 27073 11617 27125 11669
rect 26861 11399 26913 11451
rect 27073 11399 27125 11451
rect 26861 11182 26913 11234
rect 27073 11182 27125 11234
rect 26861 10964 26913 11016
rect 27073 10964 27125 11016
rect 26861 10746 26913 10798
rect 27073 10746 27125 10798
rect 26861 10529 26913 10581
rect 27073 10529 27125 10581
rect 26861 10311 26913 10363
rect 27073 10311 27125 10363
rect 26861 10094 26913 10146
rect 27073 10094 27125 10146
rect 26861 9876 26913 9928
rect 27073 9876 27125 9928
rect 26861 9658 26913 9710
rect 27073 9658 27125 9710
rect 26861 9441 26913 9493
rect 27073 9441 27125 9493
rect 26861 9223 26913 9275
rect 27073 9223 27125 9275
rect 26861 9005 26913 9057
rect 27073 9005 27125 9057
rect 26861 8788 26913 8840
rect 27073 8788 27125 8840
rect 26861 8570 26913 8622
rect 27073 8570 27125 8622
rect 26861 8352 26913 8404
rect 27073 8352 27125 8404
rect 26861 8135 26913 8187
rect 27073 8135 27125 8187
rect 26861 7917 26913 7969
rect 27073 7917 27125 7969
rect 26861 7700 26913 7752
rect 27073 7700 27125 7752
rect 26861 7482 26913 7534
rect 27073 7482 27125 7534
rect 26861 7264 26913 7316
rect 27073 7264 27125 7316
rect 26861 7047 26913 7099
rect 27073 7047 27125 7099
rect 26861 6829 26913 6881
rect 27073 6829 27125 6881
rect 26861 6611 26913 6663
rect 27073 6611 27125 6663
rect 26861 6394 26913 6446
rect 27073 6394 27125 6446
rect 26861 6176 26913 6228
rect 27073 6176 27125 6228
rect 26861 5959 26913 6011
rect 27073 5959 27125 6011
rect 26861 5741 26913 5793
rect 27073 5741 27125 5793
rect 26861 5523 26913 5575
rect 27073 5523 27125 5575
rect 26861 5306 26913 5358
rect 27073 5306 27125 5358
rect 26861 4535 26913 4587
rect 27073 4535 27125 4587
rect 26861 4318 26913 4370
rect 27073 4318 27125 4370
rect 26861 4100 26913 4152
rect 27073 4100 27125 4152
rect 26861 3882 26913 3934
rect 27073 3882 27125 3934
rect 26861 3665 26913 3717
rect 27073 3665 27125 3717
rect 2574 1637 2730 1689
rect 12639 1637 12795 1689
rect 13089 1637 13245 1689
rect 23439 1637 23595 1689
rect 27476 33380 27528 33432
rect 27688 33380 27740 33432
rect 27476 33163 27528 33215
rect 27688 33163 27740 33215
rect 27476 32945 27528 32997
rect 27688 32945 27740 32997
rect 27476 32727 27528 32779
rect 27688 32727 27740 32779
rect 27476 32510 27528 32562
rect 27688 32510 27740 32562
rect 27476 32292 27528 32344
rect 27688 32292 27740 32344
rect 27476 32075 27528 32127
rect 27688 32075 27740 32127
rect 27476 31857 27528 31909
rect 27688 31857 27740 31909
rect 27476 31639 27528 31691
rect 27688 31639 27740 31691
rect 27476 31422 27528 31474
rect 27688 31422 27740 31474
rect 27476 31204 27528 31256
rect 27688 31204 27740 31256
rect 27476 30986 27528 31038
rect 27688 30986 27740 31038
rect 27476 30769 27528 30821
rect 27688 30769 27740 30821
rect 27476 30551 27528 30603
rect 27688 30551 27740 30603
rect 27476 30334 27528 30386
rect 27688 30334 27740 30386
rect 27476 30116 27528 30168
rect 27688 30116 27740 30168
rect 27476 29898 27528 29950
rect 27688 29898 27740 29950
rect 27476 29681 27528 29733
rect 27688 29681 27740 29733
rect 27476 29463 27528 29515
rect 27688 29463 27740 29515
rect 27476 29245 27528 29297
rect 27688 29245 27740 29297
rect 27476 29028 27528 29080
rect 27688 29028 27740 29080
rect 27476 28810 27528 28862
rect 27688 28810 27740 28862
rect 27476 28592 27528 28644
rect 27688 28592 27740 28644
rect 27476 28375 27528 28427
rect 27688 28375 27740 28427
rect 27476 28157 27528 28209
rect 27688 28157 27740 28209
rect 27476 27940 27528 27992
rect 27688 27940 27740 27992
rect 27476 27722 27528 27774
rect 27688 27722 27740 27774
rect 27476 27504 27528 27556
rect 27688 27504 27740 27556
rect 27476 27287 27528 27339
rect 27688 27287 27740 27339
rect 27476 27069 27528 27121
rect 27688 27069 27740 27121
rect 27476 26851 27528 26903
rect 27688 26851 27740 26903
rect 27476 26634 27528 26686
rect 27688 26634 27740 26686
rect 27476 26416 27528 26468
rect 27688 26416 27740 26468
rect 27476 26198 27528 26250
rect 27688 26198 27740 26250
rect 27476 25981 27528 26033
rect 27688 25981 27740 26033
rect 27476 25763 27528 25815
rect 27688 25763 27740 25815
rect 27476 25546 27528 25598
rect 27688 25546 27740 25598
rect 27476 25328 27528 25380
rect 27688 25328 27740 25380
rect 27476 25110 27528 25162
rect 27688 25110 27740 25162
rect 27476 24893 27528 24945
rect 27688 24893 27740 24945
rect 27476 24675 27528 24727
rect 27688 24675 27740 24727
rect 27476 24457 27528 24509
rect 27688 24457 27740 24509
rect 27476 24240 27528 24292
rect 27688 24240 27740 24292
rect 27476 24022 27528 24074
rect 27688 24022 27740 24074
rect 27476 23805 27528 23857
rect 27688 23805 27740 23857
rect 27476 23587 27528 23639
rect 27688 23587 27740 23639
rect 27476 23369 27528 23421
rect 27688 23369 27740 23421
rect 27476 23152 27528 23204
rect 27688 23152 27740 23204
rect 27476 22934 27528 22986
rect 27688 22934 27740 22986
rect 27476 22716 27528 22768
rect 27688 22716 27740 22768
rect 27476 22499 27528 22551
rect 27688 22499 27740 22551
rect 27476 22281 27528 22333
rect 27688 22281 27740 22333
rect 27476 22063 27528 22115
rect 27688 22063 27740 22115
rect 27476 21846 27528 21898
rect 27688 21846 27740 21898
rect 27476 21628 27528 21680
rect 27688 21628 27740 21680
rect 27476 21411 27528 21463
rect 27688 21411 27740 21463
rect 27476 21193 27528 21245
rect 27688 21193 27740 21245
rect 27476 20975 27528 21027
rect 27688 20975 27740 21027
rect 27476 20758 27528 20810
rect 27688 20758 27740 20810
rect 27476 20540 27528 20592
rect 27688 20540 27740 20592
rect 27476 20322 27528 20374
rect 27688 20322 27740 20374
rect 27476 20105 27528 20157
rect 27688 20105 27740 20157
rect 27476 19887 27528 19939
rect 27688 19887 27740 19939
rect 27476 19670 27528 19722
rect 27688 19670 27740 19722
rect 27476 19452 27528 19504
rect 27688 19452 27740 19504
rect 27476 19234 27528 19286
rect 27688 19234 27740 19286
rect 27476 19016 27528 19068
rect 27688 19016 27740 19068
rect 27476 18799 27528 18851
rect 27688 18799 27740 18851
rect 27476 18581 27528 18633
rect 27688 18581 27740 18633
rect 27476 18364 27528 18416
rect 27688 18364 27740 18416
rect 27476 18146 27528 18198
rect 27688 18146 27740 18198
rect 27476 17928 27528 17980
rect 27688 17928 27740 17980
rect 27476 17711 27528 17763
rect 27688 17711 27740 17763
rect 27476 17493 27528 17545
rect 27688 17493 27740 17545
rect 27476 17275 27528 17327
rect 27688 17275 27740 17327
rect 27476 17058 27528 17110
rect 27688 17058 27740 17110
rect 27476 16840 27528 16892
rect 27688 16840 27740 16892
rect 27476 16623 27528 16675
rect 27688 16623 27740 16675
rect 27476 16405 27528 16457
rect 27688 16405 27740 16457
rect 27476 16187 27528 16239
rect 27688 16187 27740 16239
rect 27476 15970 27528 16022
rect 27688 15970 27740 16022
rect 27476 15752 27528 15804
rect 27688 15752 27740 15804
rect 27476 15534 27528 15586
rect 27688 15534 27740 15586
rect 27476 15317 27528 15369
rect 27688 15317 27740 15369
rect 27476 15099 27528 15151
rect 27688 15099 27740 15151
rect 27476 14881 27528 14933
rect 27688 14881 27740 14933
rect 27476 14664 27528 14716
rect 27688 14664 27740 14716
rect 27476 14446 27528 14498
rect 27688 14446 27740 14498
rect 27476 14229 27528 14281
rect 27688 14229 27740 14281
rect 27476 14011 27528 14063
rect 27688 14011 27740 14063
rect 27476 13793 27528 13845
rect 27688 13793 27740 13845
rect 27476 13576 27528 13628
rect 27688 13576 27740 13628
rect 27476 13358 27528 13410
rect 27688 13358 27740 13410
rect 27476 13140 27528 13192
rect 27688 13140 27740 13192
rect 27476 12923 27528 12975
rect 27688 12923 27740 12975
rect 27476 12705 27528 12757
rect 27688 12705 27740 12757
rect 27476 12488 27528 12540
rect 27688 12488 27740 12540
rect 27476 12270 27528 12322
rect 27688 12270 27740 12322
rect 27476 12052 27528 12104
rect 27688 12052 27740 12104
rect 27476 11835 27528 11887
rect 27688 11835 27740 11887
rect 27476 11617 27528 11669
rect 27688 11617 27740 11669
rect 27476 11399 27528 11451
rect 27688 11399 27740 11451
rect 27476 11182 27528 11234
rect 27688 11182 27740 11234
rect 27476 10964 27528 11016
rect 27688 10964 27740 11016
rect 27476 10746 27528 10798
rect 27688 10746 27740 10798
rect 27476 10529 27528 10581
rect 27688 10529 27740 10581
rect 27476 10311 27528 10363
rect 27688 10311 27740 10363
rect 27476 10094 27528 10146
rect 27688 10094 27740 10146
rect 27476 9876 27528 9928
rect 27688 9876 27740 9928
rect 27476 9658 27528 9710
rect 27688 9658 27740 9710
rect 27476 9441 27528 9493
rect 27688 9441 27740 9493
rect 27476 9223 27528 9275
rect 27688 9223 27740 9275
rect 27476 9005 27528 9057
rect 27688 9005 27740 9057
rect 27476 8788 27528 8840
rect 27688 8788 27740 8840
rect 27476 8570 27528 8622
rect 27688 8570 27740 8622
rect 27476 8352 27528 8404
rect 27688 8352 27740 8404
rect 27476 8135 27528 8187
rect 27688 8135 27740 8187
rect 27476 7917 27528 7969
rect 27688 7917 27740 7969
rect 27476 7700 27528 7752
rect 27688 7700 27740 7752
rect 27476 7482 27528 7534
rect 27688 7482 27740 7534
rect 27476 7264 27528 7316
rect 27688 7264 27740 7316
rect 27476 7047 27528 7099
rect 27688 7047 27740 7099
rect 27476 6829 27528 6881
rect 27688 6829 27740 6881
rect 27476 6611 27528 6663
rect 27688 6611 27740 6663
rect 27476 6394 27528 6446
rect 27688 6394 27740 6446
rect 27476 6176 27528 6228
rect 27688 6176 27740 6228
rect 27476 5959 27528 6011
rect 27688 5959 27740 6011
rect 27476 5741 27528 5793
rect 27688 5741 27740 5793
rect 27476 5523 27528 5575
rect 27688 5523 27740 5575
rect 27476 5306 27528 5358
rect 27688 5306 27740 5358
rect 27476 4535 27528 4587
rect 27688 4535 27740 4587
rect 27476 4318 27528 4370
rect 27688 4318 27740 4370
rect 27476 4100 27528 4152
rect 27688 4100 27740 4152
rect 27476 3882 27528 3934
rect 27688 3882 27740 3934
rect 27476 3665 27528 3717
rect 27688 3665 27740 3717
rect 49908 6297 50064 6349
rect 51654 5147 51810 5199
rect 40623 3230 40779 3282
rect 57383 33380 57435 33432
rect 57595 33380 57647 33432
rect 57383 33163 57435 33215
rect 57595 33163 57647 33215
rect 57383 32945 57435 32997
rect 57595 32945 57647 32997
rect 57383 32727 57435 32779
rect 57595 32727 57647 32779
rect 57383 32510 57435 32562
rect 57595 32510 57647 32562
rect 57383 32292 57435 32344
rect 57595 32292 57647 32344
rect 57383 32075 57435 32127
rect 57595 32075 57647 32127
rect 57383 31857 57435 31909
rect 57595 31857 57647 31909
rect 57383 31639 57435 31691
rect 57595 31639 57647 31691
rect 57383 31422 57435 31474
rect 57595 31422 57647 31474
rect 57383 31204 57435 31256
rect 57595 31204 57647 31256
rect 57383 30986 57435 31038
rect 57595 30986 57647 31038
rect 57383 30769 57435 30821
rect 57595 30769 57647 30821
rect 57383 30551 57435 30603
rect 57595 30551 57647 30603
rect 57383 30334 57435 30386
rect 57595 30334 57647 30386
rect 57383 30116 57435 30168
rect 57595 30116 57647 30168
rect 57383 29898 57435 29950
rect 57595 29898 57647 29950
rect 57383 29681 57435 29733
rect 57595 29681 57647 29733
rect 57383 29463 57435 29515
rect 57595 29463 57647 29515
rect 57383 29245 57435 29297
rect 57595 29245 57647 29297
rect 57383 29028 57435 29080
rect 57595 29028 57647 29080
rect 57383 28810 57435 28862
rect 57595 28810 57647 28862
rect 57383 28592 57435 28644
rect 57595 28592 57647 28644
rect 57383 28375 57435 28427
rect 57595 28375 57647 28427
rect 57383 28157 57435 28209
rect 57595 28157 57647 28209
rect 57383 27940 57435 27992
rect 57595 27940 57647 27992
rect 57383 27722 57435 27774
rect 57595 27722 57647 27774
rect 57383 27504 57435 27556
rect 57595 27504 57647 27556
rect 57383 27287 57435 27339
rect 57595 27287 57647 27339
rect 57383 27069 57435 27121
rect 57595 27069 57647 27121
rect 57383 26851 57435 26903
rect 57595 26851 57647 26903
rect 57383 26634 57435 26686
rect 57595 26634 57647 26686
rect 57383 26416 57435 26468
rect 57595 26416 57647 26468
rect 57383 26198 57435 26250
rect 57595 26198 57647 26250
rect 57383 25981 57435 26033
rect 57595 25981 57647 26033
rect 57383 25763 57435 25815
rect 57595 25763 57647 25815
rect 57383 25546 57435 25598
rect 57595 25546 57647 25598
rect 57383 25328 57435 25380
rect 57595 25328 57647 25380
rect 57383 25110 57435 25162
rect 57595 25110 57647 25162
rect 57383 24893 57435 24945
rect 57595 24893 57647 24945
rect 57383 24675 57435 24727
rect 57595 24675 57647 24727
rect 57383 24457 57435 24509
rect 57595 24457 57647 24509
rect 57383 24240 57435 24292
rect 57595 24240 57647 24292
rect 57383 24022 57435 24074
rect 57595 24022 57647 24074
rect 57383 23805 57435 23857
rect 57595 23805 57647 23857
rect 57383 23587 57435 23639
rect 57595 23587 57647 23639
rect 57383 23369 57435 23421
rect 57595 23369 57647 23421
rect 57383 23152 57435 23204
rect 57595 23152 57647 23204
rect 57383 22934 57435 22986
rect 57595 22934 57647 22986
rect 57383 22716 57435 22768
rect 57595 22716 57647 22768
rect 57383 22499 57435 22551
rect 57595 22499 57647 22551
rect 57383 22281 57435 22333
rect 57595 22281 57647 22333
rect 57383 22063 57435 22115
rect 57595 22063 57647 22115
rect 57383 21846 57435 21898
rect 57595 21846 57647 21898
rect 57383 21628 57435 21680
rect 57595 21628 57647 21680
rect 57383 21411 57435 21463
rect 57595 21411 57647 21463
rect 57383 21193 57435 21245
rect 57595 21193 57647 21245
rect 57383 20975 57435 21027
rect 57595 20975 57647 21027
rect 57383 20758 57435 20810
rect 57595 20758 57647 20810
rect 57383 20540 57435 20592
rect 57595 20540 57647 20592
rect 57383 20322 57435 20374
rect 57595 20322 57647 20374
rect 57383 20105 57435 20157
rect 57595 20105 57647 20157
rect 57383 19887 57435 19939
rect 57595 19887 57647 19939
rect 57383 19670 57435 19722
rect 57595 19670 57647 19722
rect 57383 19452 57435 19504
rect 57595 19452 57647 19504
rect 57383 19234 57435 19286
rect 57595 19234 57647 19286
rect 57383 19016 57435 19068
rect 57595 19016 57647 19068
rect 57383 18799 57435 18851
rect 57595 18799 57647 18851
rect 57383 18581 57435 18633
rect 57595 18581 57647 18633
rect 57383 18364 57435 18416
rect 57595 18364 57647 18416
rect 57383 18146 57435 18198
rect 57595 18146 57647 18198
rect 57383 17928 57435 17980
rect 57595 17928 57647 17980
rect 57383 17711 57435 17763
rect 57595 17711 57647 17763
rect 57383 17493 57435 17545
rect 57595 17493 57647 17545
rect 57383 17275 57435 17327
rect 57595 17275 57647 17327
rect 57383 17058 57435 17110
rect 57595 17058 57647 17110
rect 57383 16840 57435 16892
rect 57595 16840 57647 16892
rect 57383 16623 57435 16675
rect 57595 16623 57647 16675
rect 57383 16405 57435 16457
rect 57595 16405 57647 16457
rect 57383 16187 57435 16239
rect 57595 16187 57647 16239
rect 57383 15970 57435 16022
rect 57595 15970 57647 16022
rect 57383 15752 57435 15804
rect 57595 15752 57647 15804
rect 57383 15534 57435 15586
rect 57595 15534 57647 15586
rect 57383 15317 57435 15369
rect 57595 15317 57647 15369
rect 57383 15099 57435 15151
rect 57595 15099 57647 15151
rect 57383 14881 57435 14933
rect 57595 14881 57647 14933
rect 57383 14664 57435 14716
rect 57595 14664 57647 14716
rect 57383 14446 57435 14498
rect 57595 14446 57647 14498
rect 57383 14229 57435 14281
rect 57595 14229 57647 14281
rect 57383 14011 57435 14063
rect 57595 14011 57647 14063
rect 57383 13793 57435 13845
rect 57595 13793 57647 13845
rect 57383 13576 57435 13628
rect 57595 13576 57647 13628
rect 57383 13358 57435 13410
rect 57595 13358 57647 13410
rect 57383 13140 57435 13192
rect 57595 13140 57647 13192
rect 57383 12923 57435 12975
rect 57595 12923 57647 12975
rect 57383 12705 57435 12757
rect 57595 12705 57647 12757
rect 57383 12488 57435 12540
rect 57595 12488 57647 12540
rect 57383 12270 57435 12322
rect 57595 12270 57647 12322
rect 57383 12052 57435 12104
rect 57595 12052 57647 12104
rect 57383 11835 57435 11887
rect 57595 11835 57647 11887
rect 57383 11617 57435 11669
rect 57595 11617 57647 11669
rect 57383 11399 57435 11451
rect 57595 11399 57647 11451
rect 57383 11182 57435 11234
rect 57595 11182 57647 11234
rect 57383 10964 57435 11016
rect 57595 10964 57647 11016
rect 57383 10746 57435 10798
rect 57595 10746 57647 10798
rect 57383 10529 57435 10581
rect 57595 10529 57647 10581
rect 57383 10311 57435 10363
rect 57595 10311 57647 10363
rect 57383 10094 57435 10146
rect 57595 10094 57647 10146
rect 57383 9876 57435 9928
rect 57595 9876 57647 9928
rect 57383 9658 57435 9710
rect 57595 9658 57647 9710
rect 57383 9441 57435 9493
rect 57595 9441 57647 9493
rect 57383 9223 57435 9275
rect 57595 9223 57647 9275
rect 57383 9005 57435 9057
rect 57595 9005 57647 9057
rect 57383 8788 57435 8840
rect 57595 8788 57647 8840
rect 57383 8570 57435 8622
rect 57595 8570 57647 8622
rect 57383 8352 57435 8404
rect 57595 8352 57647 8404
rect 57383 8135 57435 8187
rect 57595 8135 57647 8187
rect 57383 7917 57435 7969
rect 57595 7917 57647 7969
rect 57383 7700 57435 7752
rect 57595 7700 57647 7752
rect 57383 7482 57435 7534
rect 57595 7482 57647 7534
rect 57383 7264 57435 7316
rect 57595 7264 57647 7316
rect 57383 7047 57435 7099
rect 57595 7047 57647 7099
rect 57383 6829 57435 6881
rect 57595 6829 57647 6881
rect 57383 6611 57435 6663
rect 57595 6611 57647 6663
rect 57383 6394 57435 6446
rect 57595 6394 57647 6446
rect 57383 6176 57435 6228
rect 57595 6176 57647 6228
rect 57383 5959 57435 6011
rect 57595 5959 57647 6011
rect 57383 5741 57435 5793
rect 57595 5741 57647 5793
rect 57383 5523 57435 5575
rect 57595 5523 57647 5575
rect 57383 5306 57435 5358
rect 57595 5306 57647 5358
rect 57383 4535 57435 4587
rect 57595 4535 57647 4587
rect 57383 4318 57435 4370
rect 57595 4318 57647 4370
rect 57383 4100 57435 4152
rect 57595 4100 57647 4152
rect 57383 3882 57435 3934
rect 57595 3882 57647 3934
rect 57383 3665 57435 3717
rect 57595 3665 57647 3717
rect 58867 94721 58919 94773
rect 58991 94721 59043 94773
rect 59115 94721 59167 94773
rect 59239 94721 59291 94773
rect 59363 94721 59415 94773
rect 58867 94597 58919 94649
rect 58991 94597 59043 94649
rect 59115 94597 59167 94649
rect 59239 94597 59291 94649
rect 59363 94597 59415 94649
rect 58867 94473 58919 94525
rect 58991 94473 59043 94525
rect 59115 94473 59167 94525
rect 59239 94473 59291 94525
rect 59363 94473 59415 94525
rect 60575 35338 60627 35494
rect 57998 33380 58050 33432
rect 58210 33380 58262 33432
rect 57998 33163 58050 33215
rect 58210 33163 58262 33215
rect 57998 32945 58050 32997
rect 58210 32945 58262 32997
rect 57998 32727 58050 32779
rect 58210 32727 58262 32779
rect 57998 32510 58050 32562
rect 58210 32510 58262 32562
rect 57998 32292 58050 32344
rect 58210 32292 58262 32344
rect 57998 32075 58050 32127
rect 58210 32075 58262 32127
rect 57998 31857 58050 31909
rect 58210 31857 58262 31909
rect 57998 31639 58050 31691
rect 58210 31639 58262 31691
rect 57998 31422 58050 31474
rect 58210 31422 58262 31474
rect 57998 31204 58050 31256
rect 58210 31204 58262 31256
rect 57998 30986 58050 31038
rect 58210 30986 58262 31038
rect 57998 30769 58050 30821
rect 58210 30769 58262 30821
rect 57998 30551 58050 30603
rect 58210 30551 58262 30603
rect 57998 30334 58050 30386
rect 58210 30334 58262 30386
rect 57998 30116 58050 30168
rect 58210 30116 58262 30168
rect 57998 29898 58050 29950
rect 58210 29898 58262 29950
rect 57998 29681 58050 29733
rect 58210 29681 58262 29733
rect 57998 29463 58050 29515
rect 58210 29463 58262 29515
rect 57998 29245 58050 29297
rect 58210 29245 58262 29297
rect 57998 29028 58050 29080
rect 58210 29028 58262 29080
rect 57998 28810 58050 28862
rect 58210 28810 58262 28862
rect 57998 28592 58050 28644
rect 58210 28592 58262 28644
rect 57998 28375 58050 28427
rect 58210 28375 58262 28427
rect 57998 28157 58050 28209
rect 58210 28157 58262 28209
rect 57998 27940 58050 27992
rect 58210 27940 58262 27992
rect 57998 27722 58050 27774
rect 58210 27722 58262 27774
rect 57998 27504 58050 27556
rect 58210 27504 58262 27556
rect 57998 27287 58050 27339
rect 58210 27287 58262 27339
rect 57998 27069 58050 27121
rect 58210 27069 58262 27121
rect 57998 26851 58050 26903
rect 58210 26851 58262 26903
rect 57998 26634 58050 26686
rect 58210 26634 58262 26686
rect 57998 26416 58050 26468
rect 58210 26416 58262 26468
rect 57998 26198 58050 26250
rect 58210 26198 58262 26250
rect 57998 25981 58050 26033
rect 58210 25981 58262 26033
rect 57998 25763 58050 25815
rect 58210 25763 58262 25815
rect 57998 25546 58050 25598
rect 58210 25546 58262 25598
rect 57998 25328 58050 25380
rect 58210 25328 58262 25380
rect 57998 25110 58050 25162
rect 58210 25110 58262 25162
rect 57998 24893 58050 24945
rect 58210 24893 58262 24945
rect 57998 24675 58050 24727
rect 58210 24675 58262 24727
rect 57998 24457 58050 24509
rect 58210 24457 58262 24509
rect 57998 24240 58050 24292
rect 58210 24240 58262 24292
rect 57998 24022 58050 24074
rect 58210 24022 58262 24074
rect 57998 23805 58050 23857
rect 58210 23805 58262 23857
rect 57998 23587 58050 23639
rect 58210 23587 58262 23639
rect 57998 23369 58050 23421
rect 58210 23369 58262 23421
rect 57998 23152 58050 23204
rect 58210 23152 58262 23204
rect 57998 22934 58050 22986
rect 58210 22934 58262 22986
rect 57998 22716 58050 22768
rect 58210 22716 58262 22768
rect 57998 22499 58050 22551
rect 58210 22499 58262 22551
rect 57998 22281 58050 22333
rect 58210 22281 58262 22333
rect 57998 22063 58050 22115
rect 58210 22063 58262 22115
rect 57998 21846 58050 21898
rect 58210 21846 58262 21898
rect 57998 21628 58050 21680
rect 58210 21628 58262 21680
rect 57998 21411 58050 21463
rect 58210 21411 58262 21463
rect 57998 21193 58050 21245
rect 58210 21193 58262 21245
rect 57998 20975 58050 21027
rect 58210 20975 58262 21027
rect 57998 20758 58050 20810
rect 58210 20758 58262 20810
rect 57998 20540 58050 20592
rect 58210 20540 58262 20592
rect 57998 20322 58050 20374
rect 58210 20322 58262 20374
rect 57998 20105 58050 20157
rect 58210 20105 58262 20157
rect 57998 19887 58050 19939
rect 58210 19887 58262 19939
rect 57998 19670 58050 19722
rect 58210 19670 58262 19722
rect 57998 19452 58050 19504
rect 58210 19452 58262 19504
rect 57998 19234 58050 19286
rect 58210 19234 58262 19286
rect 57998 19016 58050 19068
rect 58210 19016 58262 19068
rect 57998 18799 58050 18851
rect 58210 18799 58262 18851
rect 57998 18581 58050 18633
rect 58210 18581 58262 18633
rect 57998 18364 58050 18416
rect 58210 18364 58262 18416
rect 57998 18146 58050 18198
rect 58210 18146 58262 18198
rect 57998 17928 58050 17980
rect 58210 17928 58262 17980
rect 57998 17711 58050 17763
rect 58210 17711 58262 17763
rect 57998 17493 58050 17545
rect 58210 17493 58262 17545
rect 57998 17275 58050 17327
rect 58210 17275 58262 17327
rect 57998 17058 58050 17110
rect 58210 17058 58262 17110
rect 57998 16840 58050 16892
rect 58210 16840 58262 16892
rect 57998 16623 58050 16675
rect 58210 16623 58262 16675
rect 57998 16405 58050 16457
rect 58210 16405 58262 16457
rect 57998 16187 58050 16239
rect 58210 16187 58262 16239
rect 57998 15970 58050 16022
rect 58210 15970 58262 16022
rect 57998 15752 58050 15804
rect 58210 15752 58262 15804
rect 57998 15534 58050 15586
rect 58210 15534 58262 15586
rect 57998 15317 58050 15369
rect 58210 15317 58262 15369
rect 57998 15099 58050 15151
rect 58210 15099 58262 15151
rect 57998 14881 58050 14933
rect 58210 14881 58262 14933
rect 57998 14664 58050 14716
rect 58210 14664 58262 14716
rect 57998 14446 58050 14498
rect 58210 14446 58262 14498
rect 57998 14229 58050 14281
rect 58210 14229 58262 14281
rect 57998 14011 58050 14063
rect 58210 14011 58262 14063
rect 57998 13793 58050 13845
rect 58210 13793 58262 13845
rect 57998 13576 58050 13628
rect 58210 13576 58262 13628
rect 57998 13358 58050 13410
rect 58210 13358 58262 13410
rect 57998 13140 58050 13192
rect 58210 13140 58262 13192
rect 57998 12923 58050 12975
rect 58210 12923 58262 12975
rect 57998 12705 58050 12757
rect 58210 12705 58262 12757
rect 57998 12488 58050 12540
rect 58210 12488 58262 12540
rect 57998 12270 58050 12322
rect 58210 12270 58262 12322
rect 57998 12052 58050 12104
rect 58210 12052 58262 12104
rect 57998 11835 58050 11887
rect 58210 11835 58262 11887
rect 57998 11617 58050 11669
rect 58210 11617 58262 11669
rect 57998 11399 58050 11451
rect 58210 11399 58262 11451
rect 57998 11182 58050 11234
rect 58210 11182 58262 11234
rect 57998 10964 58050 11016
rect 58210 10964 58262 11016
rect 57998 10746 58050 10798
rect 58210 10746 58262 10798
rect 57998 10529 58050 10581
rect 58210 10529 58262 10581
rect 57998 10311 58050 10363
rect 58210 10311 58262 10363
rect 57998 10094 58050 10146
rect 58210 10094 58262 10146
rect 57998 9876 58050 9928
rect 58210 9876 58262 9928
rect 57998 9658 58050 9710
rect 58210 9658 58262 9710
rect 57998 9441 58050 9493
rect 58210 9441 58262 9493
rect 57998 9223 58050 9275
rect 58210 9223 58262 9275
rect 57998 9005 58050 9057
rect 58210 9005 58262 9057
rect 57998 8788 58050 8840
rect 58210 8788 58262 8840
rect 57998 8570 58050 8622
rect 58210 8570 58262 8622
rect 57998 8352 58050 8404
rect 58210 8352 58262 8404
rect 57998 8135 58050 8187
rect 58210 8135 58262 8187
rect 57998 7917 58050 7969
rect 58210 7917 58262 7969
rect 57998 7700 58050 7752
rect 58210 7700 58262 7752
rect 57998 7482 58050 7534
rect 58210 7482 58262 7534
rect 57998 7264 58050 7316
rect 58210 7264 58262 7316
rect 57998 7047 58050 7099
rect 58210 7047 58262 7099
rect 57998 6829 58050 6881
rect 58210 6829 58262 6881
rect 57998 6611 58050 6663
rect 58210 6611 58262 6663
rect 57998 6394 58050 6446
rect 58210 6394 58262 6446
rect 57998 6176 58050 6228
rect 58210 6176 58262 6228
rect 57998 5959 58050 6011
rect 58210 5959 58262 6011
rect 57998 5741 58050 5793
rect 58210 5741 58262 5793
rect 57998 5523 58050 5575
rect 58210 5523 58262 5575
rect 57998 5306 58050 5358
rect 58210 5306 58262 5358
rect 57998 4535 58050 4587
rect 58210 4535 58262 4587
rect 57998 4318 58050 4370
rect 58210 4318 58262 4370
rect 57998 4100 58050 4152
rect 58210 4100 58262 4152
rect 57998 3882 58050 3934
rect 58210 3882 58262 3934
rect 57998 3665 58050 3717
rect 58210 3665 58262 3717
rect 62150 1637 62306 1689
rect 72215 1637 72371 1689
rect 72665 1637 72821 1689
rect 82730 1637 82886 1689
<< metal2 >>
rect 282 96368 86090 96694
rect 706 95176 85666 96176
rect 706 282 1706 95176
rect 25313 94775 26039 94803
rect 25313 94719 25386 94775
rect 25442 94719 25510 94775
rect 25566 94719 25634 94775
rect 25690 94719 25758 94775
rect 25814 94719 25882 94775
rect 25938 94719 26039 94775
rect 25313 94651 26039 94719
rect 25313 94595 25386 94651
rect 25442 94595 25510 94651
rect 25566 94595 25634 94651
rect 25690 94595 25758 94651
rect 25814 94595 25882 94651
rect 25938 94595 26039 94651
rect 25313 94527 26039 94595
rect 25313 94471 25386 94527
rect 25442 94471 25510 94527
rect 25566 94471 25634 94527
rect 25690 94471 25758 94527
rect 25814 94471 25882 94527
rect 25938 94471 26039 94527
rect 25313 34992 26039 94471
rect 25313 34936 25386 34992
rect 25442 34936 25510 34992
rect 25566 34936 25634 34992
rect 25690 34936 25758 34992
rect 25814 34936 25882 34992
rect 25938 34936 26039 34992
rect 25313 34868 26039 34936
rect 25313 34812 25386 34868
rect 25442 34812 25510 34868
rect 25566 34812 25634 34868
rect 25690 34812 25758 34868
rect 25814 34812 25882 34868
rect 25938 34812 26039 34868
rect 25313 34744 26039 34812
rect 25313 34688 25386 34744
rect 25442 34688 25510 34744
rect 25566 34688 25634 34744
rect 25690 34688 25758 34744
rect 25814 34688 25882 34744
rect 25938 34688 26039 34744
rect 25313 34620 26039 34688
rect 25313 34564 25386 34620
rect 25442 34564 25510 34620
rect 25566 34564 25634 34620
rect 25690 34564 25758 34620
rect 25814 34564 25882 34620
rect 25938 34564 26039 34620
rect 25313 31248 26039 34564
rect 25313 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31192 26039 31248
rect 25313 31124 26039 31192
rect 25313 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 26039 31124
rect 25313 31000 26039 31068
rect 25313 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30944 26039 31000
rect 25313 30793 26039 30944
rect 25313 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30737 26039 30793
rect 25313 30669 26039 30737
rect 25313 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 26039 30669
rect 25313 30545 26039 30613
rect 25313 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30489 26039 30545
rect 25313 28317 26039 30489
rect 25313 28261 25404 28317
rect 25460 28261 25528 28317
rect 25584 28261 25652 28317
rect 25708 28261 25776 28317
rect 25832 28261 25900 28317
rect 25956 28261 26039 28317
rect 25313 28193 26039 28261
rect 25313 28137 25404 28193
rect 25460 28137 25528 28193
rect 25584 28137 25652 28193
rect 25708 28137 25776 28193
rect 25832 28137 25900 28193
rect 25956 28137 26039 28193
rect 25313 28069 26039 28137
rect 25313 28013 25404 28069
rect 25460 28013 25528 28069
rect 25584 28013 25652 28069
rect 25708 28013 25776 28069
rect 25832 28013 25900 28069
rect 25956 28013 26039 28069
rect 25313 27945 26039 28013
rect 25313 27889 25404 27945
rect 25460 27889 25528 27945
rect 25584 27889 25652 27945
rect 25708 27889 25776 27945
rect 25832 27889 25900 27945
rect 25956 27889 26039 27945
rect 25313 27821 26039 27889
rect 25313 27765 25404 27821
rect 25460 27765 25528 27821
rect 25584 27765 25652 27821
rect 25708 27765 25776 27821
rect 25832 27765 25900 27821
rect 25956 27765 26039 27821
rect 25313 27697 26039 27765
rect 25313 27641 25404 27697
rect 25460 27641 25528 27697
rect 25584 27641 25652 27697
rect 25708 27641 25776 27697
rect 25832 27641 25900 27697
rect 25956 27641 26039 27697
rect 25313 27573 26039 27641
rect 25313 27517 25404 27573
rect 25460 27517 25528 27573
rect 25584 27517 25652 27573
rect 25708 27517 25776 27573
rect 25832 27517 25900 27573
rect 25956 27517 26039 27573
rect 25313 27449 26039 27517
rect 25313 27393 25404 27449
rect 25460 27393 25528 27449
rect 25584 27393 25652 27449
rect 25708 27393 25776 27449
rect 25832 27393 25900 27449
rect 25956 27393 26039 27449
rect 25313 27325 26039 27393
rect 26554 34049 26996 95176
rect 27387 94655 29146 94694
rect 27387 94599 27788 94655
rect 27844 94599 27999 94655
rect 28055 94599 28210 94655
rect 28266 94599 28421 94655
rect 28477 94599 28632 94655
rect 28688 94599 28843 94655
rect 28899 94599 29054 94655
rect 29110 94599 29146 94655
rect 27387 94560 29146 94599
rect 27387 92894 27828 94560
rect 29486 94485 30364 95176
rect 30769 94485 32888 95176
rect 35128 94485 36415 95176
rect 38953 94671 39618 95176
rect 48789 94485 49990 95176
rect 52226 94485 54354 95176
rect 54758 94485 55638 95176
rect 55977 94655 57371 94694
rect 55977 94599 56013 94655
rect 56069 94599 56224 94655
rect 56280 94599 56435 94655
rect 56491 94599 56646 94655
rect 56702 94599 56857 94655
rect 56913 94599 57068 94655
rect 57124 94599 57279 94655
rect 57335 94599 57371 94655
rect 55977 94560 57371 94599
rect 27387 92855 29146 92894
rect 27387 92799 27788 92855
rect 27844 92799 27999 92855
rect 28055 92799 28210 92855
rect 28266 92799 28421 92855
rect 28477 92799 28632 92855
rect 28688 92799 28843 92855
rect 28899 92799 29054 92855
rect 29110 92799 29146 92855
rect 27387 92760 29146 92799
rect 55977 92855 57371 92894
rect 55977 92799 56013 92855
rect 56069 92799 56224 92855
rect 56280 92799 56435 92855
rect 56491 92799 56646 92855
rect 56702 92799 56857 92855
rect 56913 92799 57068 92855
rect 57124 92799 57279 92855
rect 57335 92799 57371 92855
rect 55977 92760 57371 92799
rect 27387 91094 27828 92760
rect 27387 91055 29146 91094
rect 27387 90999 27788 91055
rect 27844 90999 27999 91055
rect 28055 90999 28210 91055
rect 28266 90999 28421 91055
rect 28477 90999 28632 91055
rect 28688 90999 28843 91055
rect 28899 90999 29054 91055
rect 29110 90999 29146 91055
rect 27387 90960 29146 90999
rect 55977 91055 57371 91094
rect 55977 90999 56013 91055
rect 56069 90999 56224 91055
rect 56280 90999 56435 91055
rect 56491 90999 56646 91055
rect 56702 90999 56857 91055
rect 56913 90999 57068 91055
rect 57124 90999 57279 91055
rect 57335 90999 57371 91055
rect 55977 90960 57371 90999
rect 27387 89294 27828 90960
rect 27387 89255 29146 89294
rect 27387 89199 27788 89255
rect 27844 89199 27999 89255
rect 28055 89199 28210 89255
rect 28266 89199 28421 89255
rect 28477 89199 28632 89255
rect 28688 89199 28843 89255
rect 28899 89199 29054 89255
rect 29110 89199 29146 89255
rect 27387 89160 29146 89199
rect 55977 89255 57371 89294
rect 55977 89199 56013 89255
rect 56069 89199 56224 89255
rect 56280 89199 56435 89255
rect 56491 89199 56646 89255
rect 56702 89199 56857 89255
rect 56913 89199 57068 89255
rect 57124 89199 57279 89255
rect 57335 89199 57371 89255
rect 55977 89160 57371 89199
rect 27387 87494 27828 89160
rect 27387 87455 29146 87494
rect 27387 87399 27788 87455
rect 27844 87399 27999 87455
rect 28055 87399 28210 87455
rect 28266 87399 28421 87455
rect 28477 87399 28632 87455
rect 28688 87399 28843 87455
rect 28899 87399 29054 87455
rect 29110 87399 29146 87455
rect 27387 87360 29146 87399
rect 55977 87455 57371 87494
rect 55977 87399 56013 87455
rect 56069 87399 56224 87455
rect 56280 87399 56435 87455
rect 56491 87399 56646 87455
rect 56702 87399 56857 87455
rect 56913 87399 57068 87455
rect 57124 87399 57279 87455
rect 57335 87399 57371 87455
rect 55977 87360 57371 87399
rect 27387 85694 27828 87360
rect 27387 85655 29146 85694
rect 27387 85599 27788 85655
rect 27844 85599 27999 85655
rect 28055 85599 28210 85655
rect 28266 85599 28421 85655
rect 28477 85599 28632 85655
rect 28688 85599 28843 85655
rect 28899 85599 29054 85655
rect 29110 85599 29146 85655
rect 27387 85560 29146 85599
rect 55977 85655 57371 85694
rect 55977 85599 56013 85655
rect 56069 85599 56224 85655
rect 56280 85599 56435 85655
rect 56491 85599 56646 85655
rect 56702 85599 56857 85655
rect 56913 85599 57068 85655
rect 57124 85599 57279 85655
rect 57335 85599 57371 85655
rect 55977 85560 57371 85599
rect 27387 83894 27828 85560
rect 27387 83855 29146 83894
rect 27387 83799 27788 83855
rect 27844 83799 27999 83855
rect 28055 83799 28210 83855
rect 28266 83799 28421 83855
rect 28477 83799 28632 83855
rect 28688 83799 28843 83855
rect 28899 83799 29054 83855
rect 29110 83799 29146 83855
rect 27387 83760 29146 83799
rect 55977 83855 57371 83894
rect 55977 83799 56013 83855
rect 56069 83799 56224 83855
rect 56280 83799 56435 83855
rect 56491 83799 56646 83855
rect 56702 83799 56857 83855
rect 56913 83799 57068 83855
rect 57124 83799 57279 83855
rect 57335 83799 57371 83855
rect 55977 83760 57371 83799
rect 27387 82094 27828 83760
rect 27387 82055 29146 82094
rect 27387 81999 27788 82055
rect 27844 81999 27999 82055
rect 28055 81999 28210 82055
rect 28266 81999 28421 82055
rect 28477 81999 28632 82055
rect 28688 81999 28843 82055
rect 28899 81999 29054 82055
rect 29110 81999 29146 82055
rect 27387 81960 29146 81999
rect 55977 82055 57371 82094
rect 55977 81999 56013 82055
rect 56069 81999 56224 82055
rect 56280 81999 56435 82055
rect 56491 81999 56646 82055
rect 56702 81999 56857 82055
rect 56913 81999 57068 82055
rect 57124 81999 57279 82055
rect 57335 81999 57371 82055
rect 55977 81960 57371 81999
rect 27387 80294 27828 81960
rect 27387 80255 29146 80294
rect 27387 80199 27788 80255
rect 27844 80199 27999 80255
rect 28055 80199 28210 80255
rect 28266 80199 28421 80255
rect 28477 80199 28632 80255
rect 28688 80199 28843 80255
rect 28899 80199 29054 80255
rect 29110 80199 29146 80255
rect 27387 80160 29146 80199
rect 55977 80255 57371 80294
rect 55977 80199 56013 80255
rect 56069 80199 56224 80255
rect 56280 80199 56435 80255
rect 56491 80199 56646 80255
rect 56702 80199 56857 80255
rect 56913 80199 57068 80255
rect 57124 80199 57279 80255
rect 57335 80199 57371 80255
rect 55977 80160 57371 80199
rect 27387 78494 27828 80160
rect 27387 78455 29146 78494
rect 27387 78399 27788 78455
rect 27844 78399 27999 78455
rect 28055 78399 28210 78455
rect 28266 78399 28421 78455
rect 28477 78399 28632 78455
rect 28688 78399 28843 78455
rect 28899 78399 29054 78455
rect 29110 78399 29146 78455
rect 27387 78360 29146 78399
rect 55977 78455 57371 78494
rect 55977 78399 56013 78455
rect 56069 78399 56224 78455
rect 56280 78399 56435 78455
rect 56491 78399 56646 78455
rect 56702 78399 56857 78455
rect 56913 78399 57068 78455
rect 57124 78399 57279 78455
rect 57335 78399 57371 78455
rect 55977 78360 57371 78399
rect 27387 76694 27828 78360
rect 27387 76655 29146 76694
rect 27387 76599 27788 76655
rect 27844 76599 27999 76655
rect 28055 76599 28210 76655
rect 28266 76599 28421 76655
rect 28477 76599 28632 76655
rect 28688 76599 28843 76655
rect 28899 76599 29054 76655
rect 29110 76599 29146 76655
rect 27387 76560 29146 76599
rect 55977 76655 57371 76694
rect 55977 76599 56013 76655
rect 56069 76599 56224 76655
rect 56280 76599 56435 76655
rect 56491 76599 56646 76655
rect 56702 76599 56857 76655
rect 56913 76599 57068 76655
rect 57124 76599 57279 76655
rect 57335 76599 57371 76655
rect 55977 76560 57371 76599
rect 27387 74894 27828 76560
rect 27387 74855 29146 74894
rect 27387 74799 27788 74855
rect 27844 74799 27999 74855
rect 28055 74799 28210 74855
rect 28266 74799 28421 74855
rect 28477 74799 28632 74855
rect 28688 74799 28843 74855
rect 28899 74799 29054 74855
rect 29110 74799 29146 74855
rect 27387 74760 29146 74799
rect 55977 74855 57371 74894
rect 55977 74799 56013 74855
rect 56069 74799 56224 74855
rect 56280 74799 56435 74855
rect 56491 74799 56646 74855
rect 56702 74799 56857 74855
rect 56913 74799 57068 74855
rect 57124 74799 57279 74855
rect 57335 74799 57371 74855
rect 55977 74760 57371 74799
rect 27387 73094 27828 74760
rect 27387 73055 29146 73094
rect 27387 72999 27788 73055
rect 27844 72999 27999 73055
rect 28055 72999 28210 73055
rect 28266 72999 28421 73055
rect 28477 72999 28632 73055
rect 28688 72999 28843 73055
rect 28899 72999 29054 73055
rect 29110 72999 29146 73055
rect 27387 72960 29146 72999
rect 55977 73055 57371 73094
rect 55977 72999 56013 73055
rect 56069 72999 56224 73055
rect 56280 72999 56435 73055
rect 56491 72999 56646 73055
rect 56702 72999 56857 73055
rect 56913 72999 57068 73055
rect 57124 72999 57279 73055
rect 57335 72999 57371 73055
rect 55977 72960 57371 72999
rect 27387 71294 27828 72960
rect 27387 71255 29146 71294
rect 27387 71199 27788 71255
rect 27844 71199 27999 71255
rect 28055 71199 28210 71255
rect 28266 71199 28421 71255
rect 28477 71199 28632 71255
rect 28688 71199 28843 71255
rect 28899 71199 29054 71255
rect 29110 71199 29146 71255
rect 27387 71160 29146 71199
rect 55977 71255 57371 71294
rect 55977 71199 56013 71255
rect 56069 71199 56224 71255
rect 56280 71199 56435 71255
rect 56491 71199 56646 71255
rect 56702 71199 56857 71255
rect 56913 71199 57068 71255
rect 57124 71199 57279 71255
rect 57335 71199 57371 71255
rect 55977 71160 57371 71199
rect 27387 69494 27828 71160
rect 27387 69455 29146 69494
rect 27387 69399 27788 69455
rect 27844 69399 27999 69455
rect 28055 69399 28210 69455
rect 28266 69399 28421 69455
rect 28477 69399 28632 69455
rect 28688 69399 28843 69455
rect 28899 69399 29054 69455
rect 29110 69399 29146 69455
rect 27387 69360 29146 69399
rect 55977 69455 57371 69494
rect 55977 69399 56013 69455
rect 56069 69399 56224 69455
rect 56280 69399 56435 69455
rect 56491 69399 56646 69455
rect 56702 69399 56857 69455
rect 56913 69399 57068 69455
rect 57124 69399 57279 69455
rect 57335 69399 57371 69455
rect 55977 69360 57371 69399
rect 27387 67694 27828 69360
rect 27387 67655 29146 67694
rect 27387 67599 27788 67655
rect 27844 67599 27999 67655
rect 28055 67599 28210 67655
rect 28266 67599 28421 67655
rect 28477 67599 28632 67655
rect 28688 67599 28843 67655
rect 28899 67599 29054 67655
rect 29110 67599 29146 67655
rect 27387 67560 29146 67599
rect 55977 67655 57371 67694
rect 55977 67599 56013 67655
rect 56069 67599 56224 67655
rect 56280 67599 56435 67655
rect 56491 67599 56646 67655
rect 56702 67599 56857 67655
rect 56913 67599 57068 67655
rect 57124 67599 57279 67655
rect 57335 67599 57371 67655
rect 55977 67560 57371 67599
rect 27387 65894 27828 67560
rect 27387 65855 29146 65894
rect 27387 65799 27788 65855
rect 27844 65799 27999 65855
rect 28055 65799 28210 65855
rect 28266 65799 28421 65855
rect 28477 65799 28632 65855
rect 28688 65799 28843 65855
rect 28899 65799 29054 65855
rect 29110 65799 29146 65855
rect 27387 65760 29146 65799
rect 55977 65855 57371 65894
rect 55977 65799 56013 65855
rect 56069 65799 56224 65855
rect 56280 65799 56435 65855
rect 56491 65799 56646 65855
rect 56702 65799 56857 65855
rect 56913 65799 57068 65855
rect 57124 65799 57279 65855
rect 57335 65799 57371 65855
rect 55977 65760 57371 65799
rect 27387 64094 27828 65760
rect 27387 64055 29146 64094
rect 27387 63999 27788 64055
rect 27844 63999 27999 64055
rect 28055 63999 28210 64055
rect 28266 63999 28421 64055
rect 28477 63999 28632 64055
rect 28688 63999 28843 64055
rect 28899 63999 29054 64055
rect 29110 63999 29146 64055
rect 27387 63960 29146 63999
rect 55977 64055 57371 64094
rect 55977 63999 56013 64055
rect 56069 63999 56224 64055
rect 56280 63999 56435 64055
rect 56491 63999 56646 64055
rect 56702 63999 56857 64055
rect 56913 63999 57068 64055
rect 57124 63999 57279 64055
rect 57335 63999 57371 64055
rect 55977 63960 57371 63999
rect 27387 62294 27828 63960
rect 27387 62255 29146 62294
rect 27387 62199 27788 62255
rect 27844 62199 27999 62255
rect 28055 62199 28210 62255
rect 28266 62199 28421 62255
rect 28477 62199 28632 62255
rect 28688 62199 28843 62255
rect 28899 62199 29054 62255
rect 29110 62199 29146 62255
rect 27387 62160 29146 62199
rect 55977 62255 57371 62294
rect 55977 62199 56013 62255
rect 56069 62199 56224 62255
rect 56280 62199 56435 62255
rect 56491 62199 56646 62255
rect 56702 62199 56857 62255
rect 56913 62199 57068 62255
rect 57124 62199 57279 62255
rect 57335 62199 57371 62255
rect 55977 62160 57371 62199
rect 27387 60494 27828 62160
rect 27387 60455 29146 60494
rect 27387 60399 27788 60455
rect 27844 60399 27999 60455
rect 28055 60399 28210 60455
rect 28266 60399 28421 60455
rect 28477 60399 28632 60455
rect 28688 60399 28843 60455
rect 28899 60399 29054 60455
rect 29110 60399 29146 60455
rect 27387 60360 29146 60399
rect 55977 60455 57371 60494
rect 55977 60399 56013 60455
rect 56069 60399 56224 60455
rect 56280 60399 56435 60455
rect 56491 60399 56646 60455
rect 56702 60399 56857 60455
rect 56913 60399 57068 60455
rect 57124 60399 57279 60455
rect 57335 60399 57371 60455
rect 55977 60360 57371 60399
rect 27387 58694 27828 60360
rect 27387 58655 29146 58694
rect 27387 58599 27788 58655
rect 27844 58599 27999 58655
rect 28055 58599 28210 58655
rect 28266 58599 28421 58655
rect 28477 58599 28632 58655
rect 28688 58599 28843 58655
rect 28899 58599 29054 58655
rect 29110 58599 29146 58655
rect 27387 58560 29146 58599
rect 55977 58655 57371 58694
rect 55977 58599 56013 58655
rect 56069 58599 56224 58655
rect 56280 58599 56435 58655
rect 56491 58599 56646 58655
rect 56702 58599 56857 58655
rect 56913 58599 57068 58655
rect 57124 58599 57279 58655
rect 57335 58599 57371 58655
rect 55977 58560 57371 58599
rect 27387 56894 27828 58560
rect 27387 56855 29146 56894
rect 27387 56799 27788 56855
rect 27844 56799 27999 56855
rect 28055 56799 28210 56855
rect 28266 56799 28421 56855
rect 28477 56799 28632 56855
rect 28688 56799 28843 56855
rect 28899 56799 29054 56855
rect 29110 56799 29146 56855
rect 27387 56760 29146 56799
rect 55977 56855 57371 56894
rect 55977 56799 56013 56855
rect 56069 56799 56224 56855
rect 56280 56799 56435 56855
rect 56491 56799 56646 56855
rect 56702 56799 56857 56855
rect 56913 56799 57068 56855
rect 57124 56799 57279 56855
rect 57335 56799 57371 56855
rect 55977 56760 57371 56799
rect 27387 55094 27828 56760
rect 27387 55055 29146 55094
rect 27387 54999 27788 55055
rect 27844 54999 27999 55055
rect 28055 54999 28210 55055
rect 28266 54999 28421 55055
rect 28477 54999 28632 55055
rect 28688 54999 28843 55055
rect 28899 54999 29054 55055
rect 29110 54999 29146 55055
rect 27387 54960 29146 54999
rect 55977 55055 57371 55094
rect 55977 54999 56013 55055
rect 56069 54999 56224 55055
rect 56280 54999 56435 55055
rect 56491 54999 56646 55055
rect 56702 54999 56857 55055
rect 56913 54999 57068 55055
rect 57124 54999 57279 55055
rect 57335 54999 57371 55055
rect 55977 54960 57371 54999
rect 27387 53294 27828 54960
rect 27387 53255 29146 53294
rect 27387 53199 27788 53255
rect 27844 53199 27999 53255
rect 28055 53199 28210 53255
rect 28266 53199 28421 53255
rect 28477 53199 28632 53255
rect 28688 53199 28843 53255
rect 28899 53199 29054 53255
rect 29110 53199 29146 53255
rect 27387 53160 29146 53199
rect 55977 53255 57371 53294
rect 55977 53199 56013 53255
rect 56069 53199 56224 53255
rect 56280 53199 56435 53255
rect 56491 53199 56646 53255
rect 56702 53199 56857 53255
rect 56913 53199 57068 53255
rect 57124 53199 57279 53255
rect 57335 53199 57371 53255
rect 55977 53160 57371 53199
rect 27387 51494 27828 53160
rect 27387 51455 29146 51494
rect 27387 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 29146 51455
rect 27387 51360 29146 51399
rect 55977 51455 57371 51494
rect 55977 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 57371 51455
rect 55977 51360 57371 51399
rect 27387 49694 27828 51360
rect 27387 49655 29146 49694
rect 27387 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 29146 49655
rect 27387 49560 29146 49599
rect 55977 49655 57371 49694
rect 55977 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 57371 49655
rect 55977 49560 57371 49599
rect 27387 47894 27828 49560
rect 27387 47855 29146 47894
rect 27387 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 29146 47855
rect 27387 47760 29146 47799
rect 55977 47855 57371 47894
rect 55977 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 57371 47855
rect 55977 47760 57371 47799
rect 27387 46094 27828 47760
rect 27387 46055 29146 46094
rect 27387 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 29146 46055
rect 27387 45960 29146 45999
rect 55977 46055 57371 46094
rect 55977 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 57371 46055
rect 55977 45960 57371 45999
rect 27387 44294 27828 45960
rect 27387 44255 29146 44294
rect 27387 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 29146 44255
rect 27387 44160 29146 44199
rect 55977 44255 57371 44294
rect 55977 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 57371 44255
rect 55977 44160 57371 44199
rect 27387 42494 27828 44160
rect 27387 42455 29146 42494
rect 27387 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 29146 42455
rect 27387 42360 29146 42399
rect 55977 42455 57371 42494
rect 55977 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 57371 42455
rect 55977 42360 57371 42399
rect 27387 40694 27828 42360
rect 27387 40655 29146 40694
rect 27387 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 29146 40655
rect 27387 40560 29146 40599
rect 55977 40655 57371 40694
rect 55977 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 57371 40655
rect 55977 40560 57371 40599
rect 27387 38894 27828 40560
rect 27387 38855 29146 38894
rect 27387 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 29146 38855
rect 27387 38760 29146 38799
rect 55977 38855 57371 38894
rect 55977 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 57371 38855
rect 55977 38760 57371 38799
rect 27387 37094 27828 38760
rect 27387 37055 29146 37094
rect 27387 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 29146 37055
rect 27387 36960 29146 36999
rect 55977 37055 57371 37094
rect 55977 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 57371 37055
rect 55977 36960 57371 36999
rect 27387 34992 27828 36960
rect 36863 35881 37743 36650
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 36863 35786 37743 35825
rect 41472 35761 41694 36096
rect 38596 35532 41694 35761
rect 38596 35516 38817 35532
rect 27387 34936 27447 34992
rect 27503 34936 27571 34992
rect 27627 34936 27695 34992
rect 27751 34936 27828 34992
rect 27387 34868 27828 34936
rect 27387 34812 27447 34868
rect 27503 34812 27571 34868
rect 27627 34812 27695 34868
rect 27751 34812 27828 34868
rect 27387 34744 27828 34812
rect 27387 34688 27447 34744
rect 27503 34688 27571 34744
rect 27627 34688 27695 34744
rect 27751 34688 27828 34744
rect 27387 34620 27828 34688
rect 27387 34564 27447 34620
rect 27503 34564 27571 34620
rect 27627 34564 27695 34620
rect 27751 34564 27828 34620
rect 26554 34011 27163 34049
rect 26554 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27163 34011
rect 26554 33793 27163 33955
rect 26554 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27163 33793
rect 26554 33576 27163 33737
rect 26554 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27163 33576
rect 26554 33432 27163 33520
rect 26554 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27163 33432
rect 26554 33358 27163 33380
rect 26554 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27163 33358
rect 26554 33215 27163 33302
rect 26554 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27163 33215
rect 26554 33140 27163 33163
rect 26554 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27163 33140
rect 26554 32997 27163 33084
rect 26554 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27163 32997
rect 26554 32922 27163 32945
rect 26554 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27163 32922
rect 26554 32779 27163 32866
rect 26554 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27163 32779
rect 26554 32705 27163 32727
rect 26554 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27163 32705
rect 26554 32562 27163 32649
rect 26554 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27163 32562
rect 26554 32487 27163 32510
rect 26554 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27163 32487
rect 26554 32344 27163 32431
rect 26554 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27163 32344
rect 26554 32127 27163 32292
rect 26554 32088 26861 32127
rect 26913 32088 27073 32127
rect 27125 32088 27163 32127
rect 26554 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 27163 32088
rect 26554 31909 27163 32032
rect 26554 31870 26861 31909
rect 26913 31870 27073 31909
rect 27125 31870 27163 31909
rect 26554 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 27163 31870
rect 26554 31691 27163 31814
rect 26554 31652 26861 31691
rect 26913 31652 27073 31691
rect 27125 31652 27163 31691
rect 26554 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 27163 31652
rect 26554 31474 27163 31596
rect 26554 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27163 31474
rect 26554 31256 27163 31422
rect 26554 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27163 31256
rect 26554 31038 27163 31204
rect 26554 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27163 31038
rect 26554 30821 27163 30986
rect 26554 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27163 30821
rect 26554 30603 27163 30769
rect 26554 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27163 30603
rect 26554 30386 27163 30551
rect 26554 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27163 30386
rect 26554 30168 27163 30334
rect 26554 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27163 30168
rect 26554 29968 27163 30116
rect 26554 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 27163 29968
rect 26554 29898 26861 29912
rect 26913 29898 27073 29912
rect 27125 29898 27163 29912
rect 26554 29750 27163 29898
rect 26554 29694 26859 29750
rect 26915 29694 27071 29750
rect 27127 29694 27163 29750
rect 26554 29681 26861 29694
rect 26913 29681 27073 29694
rect 27125 29681 27163 29694
rect 26554 29533 27163 29681
rect 26554 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 27163 29533
rect 26554 29463 26861 29477
rect 26913 29463 27073 29477
rect 27125 29463 27163 29477
rect 26554 29315 27163 29463
rect 26554 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 27163 29315
rect 26554 29245 26861 29259
rect 26913 29245 27073 29259
rect 27125 29245 27163 29259
rect 26554 29098 27163 29245
rect 26554 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 27163 29098
rect 26554 29028 26861 29042
rect 26913 29028 27073 29042
rect 27125 29028 27163 29042
rect 26554 28880 27163 29028
rect 26554 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 27163 28880
rect 26554 28810 26861 28824
rect 26913 28810 27073 28824
rect 27125 28810 27163 28824
rect 26554 28662 27163 28810
rect 26554 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 27163 28662
rect 26554 28592 26861 28606
rect 26913 28592 27073 28606
rect 27125 28592 27163 28606
rect 26554 28444 27163 28592
rect 26554 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 27163 28444
rect 26554 28375 26861 28388
rect 26913 28375 27073 28388
rect 27125 28375 27163 28388
rect 26554 28227 27163 28375
rect 26554 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 27163 28227
rect 26554 28157 26861 28171
rect 26913 28157 27073 28171
rect 27125 28157 27163 28171
rect 26554 28009 27163 28157
rect 26554 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 27163 28009
rect 26554 27940 26861 27953
rect 26913 27940 27073 27953
rect 27125 27940 27163 27953
rect 26554 27792 27163 27940
rect 26554 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 27163 27792
rect 26554 27722 26861 27736
rect 26913 27722 27073 27736
rect 27125 27722 27163 27736
rect 26554 27574 27163 27722
rect 26554 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 27163 27574
rect 26554 27504 26861 27518
rect 26913 27504 27073 27518
rect 27125 27504 27163 27518
rect 26554 27382 27163 27504
rect 25313 27269 25404 27325
rect 25460 27269 25528 27325
rect 25584 27269 25652 27325
rect 25708 27269 25776 27325
rect 25832 27269 25900 27325
rect 25956 27269 26039 27325
rect 25313 27201 26039 27269
rect 25313 27145 25404 27201
rect 25460 27145 25528 27201
rect 25584 27145 25652 27201
rect 25708 27145 25776 27201
rect 25832 27145 25900 27201
rect 25956 27145 26039 27201
rect 25313 27077 26039 27145
rect 25313 27021 25404 27077
rect 25460 27021 25528 27077
rect 25584 27021 25652 27077
rect 25708 27021 25776 27077
rect 25832 27021 25900 27077
rect 25956 27021 26039 27077
rect 25313 26953 26039 27021
rect 25313 26897 25404 26953
rect 25460 26897 25528 26953
rect 25584 26897 25652 26953
rect 25708 26897 25776 26953
rect 25832 26897 25900 26953
rect 25956 26897 26039 26953
rect 25313 26829 26039 26897
rect 25313 26773 25404 26829
rect 25460 26773 25528 26829
rect 25584 26773 25652 26829
rect 25708 26773 25776 26829
rect 25832 26773 25900 26829
rect 25956 26773 26039 26829
rect 25313 26705 26039 26773
rect 25313 26649 25404 26705
rect 25460 26649 25528 26705
rect 25584 26649 25652 26705
rect 25708 26649 25776 26705
rect 25832 26649 25900 26705
rect 25956 26649 26039 26705
rect 25313 26581 26039 26649
rect 25313 26525 25404 26581
rect 25460 26525 25528 26581
rect 25584 26525 25652 26581
rect 25708 26525 25776 26581
rect 25832 26525 25900 26581
rect 25956 26525 26039 26581
rect 25313 26433 26039 26525
rect 26823 27339 27163 27382
rect 26823 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27163 27339
rect 26823 27121 27163 27287
rect 26823 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27163 27121
rect 26823 26903 27163 27069
rect 26823 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27163 26903
rect 26823 26686 27163 26851
rect 26823 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27163 26686
rect 26823 26468 27163 26634
rect 26823 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27163 26468
rect 26435 26286 26643 26321
rect 26435 26126 26450 26286
rect 26610 26126 26643 26286
rect 26077 25967 26285 26002
rect 26077 25807 26092 25967
rect 26252 25807 26285 25967
rect 25741 25647 25949 25676
rect 25741 25487 25756 25647
rect 25916 25487 25949 25647
rect 25406 25328 25614 25357
rect 25406 25168 25421 25328
rect 25581 25168 25614 25328
rect 25066 24637 25274 24666
rect 25066 24477 25081 24637
rect 25241 24477 25274 24637
rect 24729 24316 24937 24345
rect 24729 24156 24744 24316
rect 24904 24156 24937 24316
rect 24401 23995 24609 24024
rect 24401 23835 24416 23995
rect 24576 23835 24609 23995
rect 24042 23673 24250 23702
rect 24042 23513 24057 23673
rect 24217 23513 24250 23673
rect 24042 17317 24250 23513
rect 24401 17656 24609 23835
rect 24729 17977 24937 24156
rect 25066 18350 25274 24477
rect 25406 18684 25614 25168
rect 25741 19027 25949 25487
rect 26077 19347 26285 25807
rect 26435 19692 26643 26126
rect 26435 19532 26465 19692
rect 26625 19532 26643 19692
rect 26435 19502 26643 19532
rect 26823 26250 27163 26416
rect 26823 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27163 26250
rect 26823 26033 27163 26198
rect 26823 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27163 26033
rect 26823 25815 27163 25981
rect 26823 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27163 25815
rect 26823 25598 27163 25763
rect 26823 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27163 25598
rect 26823 25380 27163 25546
rect 26823 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27163 25380
rect 26823 25162 27163 25328
rect 26823 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27163 25162
rect 26823 24945 27163 25110
rect 26823 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27163 24945
rect 26823 24727 27163 24893
rect 26823 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27163 24727
rect 26823 24509 27163 24675
rect 26823 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27163 24509
rect 26823 24292 27163 24457
rect 26823 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27163 24292
rect 26823 24075 27163 24240
rect 26823 23187 26858 24075
rect 27122 24074 27163 24075
rect 27125 24022 27163 24074
rect 27122 23857 27163 24022
rect 27125 23805 27163 23857
rect 27122 23639 27163 23805
rect 27125 23587 27163 23639
rect 27122 23421 27163 23587
rect 27125 23369 27163 23421
rect 27122 23204 27163 23369
rect 26823 23152 26861 23187
rect 26913 23152 27073 23187
rect 27125 23152 27163 23204
rect 26823 22986 27163 23152
rect 26823 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27163 22986
rect 26823 22768 27163 22934
rect 26823 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27163 22768
rect 26823 22551 27163 22716
rect 26823 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27163 22551
rect 26823 22333 27163 22499
rect 26823 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27163 22333
rect 26823 22115 27163 22281
rect 26823 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27163 22115
rect 26823 21898 27163 22063
rect 26823 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27163 21898
rect 26823 21680 27163 21846
rect 26823 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27163 21680
rect 26823 21463 27163 21628
rect 26823 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27163 21463
rect 26823 21245 27163 21411
rect 26823 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27163 21245
rect 26823 21027 27163 21193
rect 26823 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27163 21027
rect 26823 20810 27163 20975
rect 26823 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27163 20810
rect 26823 20592 27163 20758
rect 26823 20540 26861 20592
rect 26913 20570 27073 20592
rect 26913 20540 26924 20570
rect 27125 20540 27163 20592
rect 26823 20410 26924 20540
rect 27084 20410 27163 20540
rect 26823 20374 27163 20410
rect 26823 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27163 20374
rect 26823 20226 27163 20322
rect 26823 20157 26924 20226
rect 27084 20157 27163 20226
rect 26823 20105 26861 20157
rect 26913 20105 26924 20157
rect 27125 20105 27163 20157
rect 26823 20066 26924 20105
rect 27084 20066 27163 20105
rect 26823 19939 27163 20066
rect 26823 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27163 19939
rect 26823 19722 27163 19887
rect 26823 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27163 19722
rect 26823 19504 27163 19670
rect 26077 19187 26107 19347
rect 26267 19187 26285 19347
rect 26077 19162 26285 19187
rect 26823 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27163 19504
rect 26823 19286 27163 19452
rect 26823 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27163 19286
rect 25741 18867 25771 19027
rect 25931 18867 25949 19027
rect 25741 18822 25949 18867
rect 26823 19068 27163 19234
rect 26823 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27163 19068
rect 26823 18851 27163 19016
rect 25406 18524 25434 18684
rect 25594 18524 25614 18684
rect 25406 18482 25614 18524
rect 26823 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27163 18851
rect 26823 18633 27163 18799
rect 26823 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27163 18633
rect 25066 18190 25094 18350
rect 25254 18190 25274 18350
rect 25066 18142 25274 18190
rect 26823 18416 27163 18581
rect 26823 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27163 18416
rect 26823 18198 27163 18364
rect 26823 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27163 18198
rect 24729 17817 24757 17977
rect 24917 17817 24937 17977
rect 24729 17803 24937 17817
rect 26823 17980 27163 18146
rect 26823 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27163 17980
rect 24401 17496 24429 17656
rect 24589 17496 24609 17656
rect 24401 17462 24609 17496
rect 26823 17763 27163 17928
rect 26823 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27163 17763
rect 26823 17545 27163 17711
rect 26823 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27163 17545
rect 24042 17157 24069 17317
rect 24229 17157 24250 17317
rect 24042 17122 24250 17157
rect 26823 17327 27163 17493
rect 26823 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27163 17327
rect 26823 17110 27163 17275
rect 26823 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27163 17110
rect 26823 16892 27163 17058
rect 26823 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27163 16892
rect 26823 16675 27163 16840
rect 26823 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27163 16675
rect 26823 16457 27163 16623
rect 26823 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27163 16457
rect 26823 16239 27163 16405
rect 26823 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27163 16239
rect 26823 16022 27163 16187
rect 26823 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27163 16022
rect 26823 15804 27163 15970
rect 26823 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27163 15804
rect 26823 15586 27163 15752
rect 26823 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27163 15586
rect 26823 15369 27163 15534
rect 26823 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27163 15369
rect 26823 15151 27163 15317
rect 26823 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27163 15151
rect 26823 14933 27163 15099
rect 26823 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27163 14933
rect 26823 14716 27163 14881
rect 26823 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27163 14716
rect 26823 14498 27163 14664
rect 26823 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27163 14498
rect 26823 14281 27163 14446
rect 26823 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27163 14281
rect 26823 14119 27163 14229
rect 26823 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27163 14119
rect 26823 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27163 14063
rect 26823 13902 27163 14011
rect 26823 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27163 13902
rect 26823 13845 27163 13846
rect 26823 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27163 13845
rect 26823 13684 27163 13793
rect 26823 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27163 13684
rect 26823 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27163 13628
rect 26823 13467 27163 13576
rect 26823 13411 26859 13467
rect 26915 13411 27071 13467
rect 27127 13411 27163 13467
rect 26823 13410 27163 13411
rect 26823 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27163 13410
rect 26823 13249 27163 13358
rect 26823 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27163 13249
rect 26823 13192 27163 13193
rect 26823 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27163 13192
rect 26823 13031 27163 13140
rect 26823 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27163 13031
rect 26823 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27163 12975
rect 26823 12813 27163 12923
rect 26823 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 27163 12813
rect 26823 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27163 12757
rect 26823 12596 27163 12705
rect 26823 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12540 27163 12596
rect 26823 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27163 12540
rect 26823 12378 27163 12488
rect 26823 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 27163 12378
rect 26823 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27163 12322
rect 26823 12161 27163 12270
rect 26823 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 27163 12161
rect 26823 12104 27163 12105
rect 26823 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27163 12104
rect 26823 11887 27163 12052
rect 26823 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27163 11887
rect 26823 11669 27163 11835
rect 26823 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27163 11669
rect 26823 11451 27163 11617
rect 26823 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27163 11451
rect 26823 11234 27163 11399
rect 26823 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27163 11234
rect 26823 11016 27163 11182
rect 26823 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27163 11016
rect 26823 10798 27163 10964
rect 26823 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27163 10798
rect 26823 10581 27163 10746
rect 26823 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27163 10581
rect 26823 10363 27163 10529
rect 26823 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27163 10363
rect 26823 10146 27163 10311
rect 26823 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27163 10146
rect 26823 9928 27163 10094
rect 26823 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27163 9928
rect 26823 9710 27163 9876
rect 26823 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27163 9710
rect 26823 9493 27163 9658
rect 26823 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27163 9493
rect 26823 9407 27163 9441
rect 26823 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 27163 9407
rect 26823 9275 27163 9351
rect 26823 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27163 9275
rect 26823 9190 27163 9223
rect 26823 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 27163 9190
rect 26823 9057 27163 9134
rect 26823 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27163 9057
rect 26823 8972 27163 9005
rect 26823 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 27163 8972
rect 26823 8840 27163 8916
rect 26823 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27163 8840
rect 26823 8754 27163 8788
rect 26823 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 27163 8754
rect 26823 8622 27163 8698
rect 26823 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27163 8622
rect 26823 8536 27163 8570
rect 26823 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 27163 8536
rect 26823 8404 27163 8480
rect 26823 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27163 8404
rect 26823 8319 27163 8352
rect 26823 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 27163 8319
rect 26823 8187 27163 8263
rect 26823 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27163 8187
rect 26823 7969 27163 8135
rect 26823 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27163 7969
rect 26823 7752 27163 7917
rect 26823 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27163 7752
rect 26823 7534 27163 7700
rect 26823 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27163 7534
rect 26823 7316 27163 7482
rect 26823 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27163 7316
rect 26823 7099 27163 7264
rect 26823 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27163 7099
rect 26823 6881 27163 7047
rect 26823 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27163 6881
rect 26823 6663 27163 6829
rect 26823 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27163 6663
rect 26823 6446 27163 6611
rect 26823 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27163 6446
rect 26823 6228 27163 6394
rect 26823 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27163 6228
rect 26823 6011 27163 6176
rect 26823 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27163 6011
rect 26823 5793 27163 5959
rect 26823 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27163 5793
rect 26823 5575 27163 5741
rect 26823 5539 26861 5575
rect 26913 5539 27073 5575
rect 27125 5539 27163 5575
rect 26823 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27163 5539
rect 26823 5358 27163 5483
rect 26823 5321 26861 5358
rect 26913 5321 27073 5358
rect 27125 5321 27163 5358
rect 26823 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27163 5321
rect 26823 5226 27163 5265
rect 27387 33432 27828 34564
rect 27387 33380 27476 33432
rect 27528 33380 27688 33432
rect 27740 33380 27828 33432
rect 27387 33215 27828 33380
rect 31615 35287 38817 35516
rect 41850 35425 42072 36096
rect 31615 33349 31836 35287
rect 39077 35197 42072 35425
rect 39077 35171 39298 35197
rect 31970 34943 39298 35171
rect 42228 35090 42449 36096
rect 31970 33349 32192 34943
rect 39755 34861 42449 35090
rect 39755 34675 39977 34861
rect 42603 34754 42825 36085
rect 38301 34491 39977 34675
rect 37201 34446 39977 34491
rect 40106 34526 42825 34754
rect 37201 34263 38523 34446
rect 40106 34312 40328 34526
rect 42983 34419 43205 36096
rect 37201 33360 37423 34263
rect 38642 34156 40328 34312
rect 37557 34084 40328 34156
rect 40458 34190 43205 34419
rect 37557 33927 38863 34084
rect 40458 33977 40679 34190
rect 43359 34083 43580 36085
rect 45513 35842 45735 36096
rect 37557 33349 37778 33927
rect 38993 33748 40679 33977
rect 40809 33855 43580 34083
rect 44646 35614 45735 35842
rect 38993 33360 39215 33748
rect 40809 33625 41031 33855
rect 39349 33397 41031 33625
rect 44646 33576 44867 35614
rect 45891 35507 46112 36096
rect 44997 35278 46112 35507
rect 46268 35681 46490 36096
rect 46268 35453 46501 35681
rect 44997 33576 45219 35278
rect 46279 33576 46501 35453
rect 46646 35346 46868 36085
rect 46631 35117 46868 35346
rect 46631 33564 46852 35117
rect 47026 34836 47248 36085
rect 47402 35171 47623 36096
rect 47779 35507 48001 36096
rect 48157 35842 48379 36096
rect 48157 35614 50120 35842
rect 47779 35278 49769 35507
rect 47402 34943 48486 35171
rect 47026 34607 48135 34836
rect 47913 33564 48135 34607
rect 48265 33576 48486 34943
rect 49547 33576 49769 35278
rect 49898 33576 50120 35614
rect 57909 34011 58351 95176
rect 57909 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 58351 34011
rect 57909 33793 58351 33955
rect 57909 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 58351 33793
rect 57909 33576 58351 33737
rect 57909 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 58351 33576
rect 57295 33432 57736 33519
rect 57295 33380 57383 33432
rect 57435 33380 57595 33432
rect 57647 33380 57736 33432
rect 27387 33163 27476 33215
rect 27528 33163 27688 33215
rect 27740 33163 27828 33215
rect 27387 33141 27828 33163
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 27828 33141
rect 27387 32997 27828 33085
rect 27387 32945 27476 32997
rect 27528 32945 27688 32997
rect 27740 32945 27828 32997
rect 27387 32923 27828 32945
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 27828 32923
rect 27387 32779 27828 32867
rect 27387 32727 27476 32779
rect 27528 32727 27688 32779
rect 27740 32727 27828 32779
rect 27387 32705 27828 32727
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 27828 32705
rect 27387 32562 27828 32649
rect 27387 32510 27476 32562
rect 27528 32510 27688 32562
rect 27740 32510 27828 32562
rect 27387 32487 27828 32510
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 27828 32487
rect 27387 32344 27828 32431
rect 27387 32292 27476 32344
rect 27528 32292 27688 32344
rect 27740 32292 27828 32344
rect 27387 32127 27828 32292
rect 27387 32075 27476 32127
rect 27528 32075 27688 32127
rect 27740 32075 27828 32127
rect 27387 31909 27828 32075
rect 27387 31857 27476 31909
rect 27528 31857 27688 31909
rect 27740 31857 27828 31909
rect 27387 31691 27828 31857
rect 27387 31639 27476 31691
rect 27528 31639 27688 31691
rect 27740 31639 27828 31691
rect 27387 31474 27828 31639
rect 27387 31422 27476 31474
rect 27528 31422 27688 31474
rect 27740 31422 27828 31474
rect 27387 31256 27828 31422
rect 27387 31252 27476 31256
rect 27528 31252 27688 31256
rect 27740 31252 27828 31256
rect 27387 31196 27474 31252
rect 27530 31196 27686 31252
rect 27742 31196 27828 31252
rect 27387 31038 27828 31196
rect 27387 31034 27476 31038
rect 27528 31034 27688 31038
rect 27740 31034 27828 31038
rect 27387 30978 27474 31034
rect 27530 30978 27686 31034
rect 27742 30978 27828 31034
rect 27387 30821 27828 30978
rect 27387 30816 27476 30821
rect 27528 30816 27688 30821
rect 27740 30816 27828 30821
rect 27387 30760 27474 30816
rect 27530 30760 27686 30816
rect 27742 30760 27828 30816
rect 27387 30603 27828 30760
rect 27387 30598 27476 30603
rect 27528 30598 27688 30603
rect 27740 30598 27828 30603
rect 27387 30542 27474 30598
rect 27530 30542 27686 30598
rect 27742 30542 27828 30598
rect 27387 30386 27828 30542
rect 27387 30334 27476 30386
rect 27528 30334 27688 30386
rect 27740 30334 27828 30386
rect 27387 30168 27828 30334
rect 27387 30116 27476 30168
rect 27528 30116 27688 30168
rect 27740 30116 27828 30168
rect 27387 29950 27828 30116
rect 27387 29898 27476 29950
rect 27528 29898 27688 29950
rect 27740 29898 27828 29950
rect 27387 29733 27828 29898
rect 27387 29681 27476 29733
rect 27528 29681 27688 29733
rect 27740 29681 27828 29733
rect 27387 29515 27828 29681
rect 27387 29463 27476 29515
rect 27528 29463 27688 29515
rect 27740 29463 27828 29515
rect 27387 29297 27828 29463
rect 27387 29245 27476 29297
rect 27528 29245 27688 29297
rect 27740 29245 27828 29297
rect 27387 29080 27828 29245
rect 27387 29028 27476 29080
rect 27528 29028 27688 29080
rect 27740 29028 27828 29080
rect 27387 28862 27828 29028
rect 27387 28810 27476 28862
rect 27528 28810 27688 28862
rect 27740 28810 27828 28862
rect 27387 28644 27828 28810
rect 27387 28592 27476 28644
rect 27528 28592 27688 28644
rect 27740 28592 27828 28644
rect 27387 28427 27828 28592
rect 27387 28375 27476 28427
rect 27528 28375 27688 28427
rect 27740 28375 27828 28427
rect 27387 28209 27828 28375
rect 27387 28157 27476 28209
rect 27528 28157 27688 28209
rect 27740 28157 27828 28209
rect 27387 27992 27828 28157
rect 27387 27940 27476 27992
rect 27528 27940 27688 27992
rect 27740 27940 27828 27992
rect 27387 27774 27828 27940
rect 27387 27722 27476 27774
rect 27528 27722 27688 27774
rect 27740 27722 27828 27774
rect 27387 27556 27828 27722
rect 27387 27504 27476 27556
rect 27528 27504 27688 27556
rect 27740 27504 27828 27556
rect 27387 27339 27828 27504
rect 27387 27287 27476 27339
rect 27528 27287 27688 27339
rect 27740 27287 27828 27339
rect 27387 27121 27828 27287
rect 27387 27069 27476 27121
rect 27528 27069 27688 27121
rect 27740 27069 27828 27121
rect 27387 26903 27828 27069
rect 27387 26851 27476 26903
rect 27528 26851 27688 26903
rect 27740 26851 27828 26903
rect 27387 26799 27828 26851
rect 27387 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 27387 26686 27828 26743
rect 27387 26634 27476 26686
rect 27528 26634 27688 26686
rect 27740 26634 27828 26686
rect 27387 26581 27828 26634
rect 27387 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 27387 26468 27828 26525
rect 27387 26416 27476 26468
rect 27528 26416 27688 26468
rect 27740 26416 27828 26468
rect 27387 26250 27828 26416
rect 27387 26198 27476 26250
rect 27528 26198 27688 26250
rect 27740 26198 27828 26250
rect 27387 26033 27828 26198
rect 27387 25981 27476 26033
rect 27528 25981 27688 26033
rect 27740 25981 27828 26033
rect 27387 25815 27828 25981
rect 27387 25763 27476 25815
rect 27528 25763 27688 25815
rect 27740 25763 27828 25815
rect 27387 25598 27828 25763
rect 27387 25546 27476 25598
rect 27528 25546 27688 25598
rect 27740 25546 27828 25598
rect 27387 25380 27828 25546
rect 27387 25328 27476 25380
rect 27528 25328 27688 25380
rect 27740 25328 27828 25380
rect 27387 25162 27828 25328
rect 27387 25110 27476 25162
rect 27528 25110 27688 25162
rect 27740 25110 27828 25162
rect 27387 25028 27828 25110
rect 27387 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 27828 25028
rect 27387 24945 27828 24972
rect 27387 24893 27476 24945
rect 27528 24893 27688 24945
rect 27740 24893 27828 24945
rect 27387 24810 27828 24893
rect 27387 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 27828 24810
rect 27387 24727 27828 24754
rect 27387 24675 27476 24727
rect 27528 24675 27688 24727
rect 27740 24675 27828 24727
rect 27387 24509 27828 24675
rect 27387 24457 27476 24509
rect 27528 24457 27688 24509
rect 27740 24457 27828 24509
rect 27387 24292 27828 24457
rect 27387 24240 27476 24292
rect 27528 24240 27688 24292
rect 27740 24240 27828 24292
rect 27387 24074 27828 24240
rect 27387 24022 27476 24074
rect 27528 24022 27688 24074
rect 27740 24022 27828 24074
rect 27387 23857 27828 24022
rect 27387 23805 27476 23857
rect 27528 23805 27688 23857
rect 27740 23805 27828 23857
rect 27387 23639 27828 23805
rect 27387 23587 27476 23639
rect 27528 23587 27688 23639
rect 27740 23587 27828 23639
rect 27387 23421 27828 23587
rect 27387 23369 27476 23421
rect 27528 23369 27688 23421
rect 27740 23369 27828 23421
rect 27387 23204 27828 23369
rect 27387 23152 27476 23204
rect 27528 23152 27688 23204
rect 27740 23152 27828 23204
rect 27387 22986 27828 23152
rect 27387 22936 27476 22986
rect 27528 22936 27688 22986
rect 27387 22048 27475 22936
rect 27740 22934 27828 22986
rect 27739 22768 27828 22934
rect 27740 22716 27828 22768
rect 27739 22551 27828 22716
rect 27740 22499 27828 22551
rect 27739 22333 27828 22499
rect 27740 22281 27828 22333
rect 27739 22115 27828 22281
rect 27740 22063 27828 22115
rect 27739 22048 27828 22063
rect 27387 21898 27828 22048
rect 27387 21846 27476 21898
rect 27528 21846 27688 21898
rect 27740 21846 27828 21898
rect 27387 21680 27828 21846
rect 27387 21628 27476 21680
rect 27528 21628 27688 21680
rect 27740 21628 27828 21680
rect 27387 21463 27828 21628
rect 27387 21411 27476 21463
rect 27528 21411 27688 21463
rect 27740 21411 27828 21463
rect 27387 21245 27828 21411
rect 27387 21193 27476 21245
rect 27528 21193 27688 21245
rect 27740 21193 27828 21245
rect 27387 21027 27828 21193
rect 27387 20975 27476 21027
rect 27528 20975 27688 21027
rect 27740 20975 27828 21027
rect 27387 20810 27828 20975
rect 27387 20758 27476 20810
rect 27528 20758 27688 20810
rect 27740 20758 27828 20810
rect 27387 20592 27828 20758
rect 27387 20540 27476 20592
rect 27528 20540 27688 20592
rect 27740 20540 27828 20592
rect 27387 20374 27828 20540
rect 27387 20322 27476 20374
rect 27528 20322 27688 20374
rect 27740 20322 27828 20374
rect 27387 20157 27828 20322
rect 27387 20105 27476 20157
rect 27528 20105 27688 20157
rect 27740 20105 27828 20157
rect 27387 19939 27828 20105
rect 27387 19887 27476 19939
rect 27528 19887 27688 19939
rect 27740 19887 27828 19939
rect 27387 19722 27828 19887
rect 27387 19670 27476 19722
rect 27528 19670 27688 19722
rect 27740 19670 27828 19722
rect 27387 19504 27828 19670
rect 27387 19452 27476 19504
rect 27528 19452 27688 19504
rect 27740 19452 27828 19504
rect 27387 19286 27828 19452
rect 27387 19234 27476 19286
rect 27528 19234 27688 19286
rect 27740 19234 27828 19286
rect 27387 19068 27828 19234
rect 27387 19016 27476 19068
rect 27528 19016 27688 19068
rect 27740 19016 27828 19068
rect 27387 18851 27828 19016
rect 27387 18799 27476 18851
rect 27528 18799 27688 18851
rect 27740 18799 27828 18851
rect 27387 18633 27828 18799
rect 27387 18581 27476 18633
rect 27528 18581 27688 18633
rect 27740 18581 27828 18633
rect 27387 18416 27828 18581
rect 27387 18364 27476 18416
rect 27528 18364 27688 18416
rect 27740 18364 27828 18416
rect 27387 18198 27828 18364
rect 27387 18146 27476 18198
rect 27528 18146 27688 18198
rect 27740 18146 27828 18198
rect 27387 17980 27828 18146
rect 27387 17928 27476 17980
rect 27528 17928 27688 17980
rect 27740 17928 27828 17980
rect 27387 17763 27828 17928
rect 27387 17711 27476 17763
rect 27528 17711 27688 17763
rect 27740 17711 27828 17763
rect 27387 17545 27828 17711
rect 27387 17493 27476 17545
rect 27528 17493 27688 17545
rect 27740 17493 27828 17545
rect 27387 17327 27828 17493
rect 27387 17275 27476 17327
rect 27528 17275 27688 17327
rect 27740 17275 27828 17327
rect 27387 17110 27828 17275
rect 27387 17058 27476 17110
rect 27528 17058 27688 17110
rect 27740 17058 27828 17110
rect 27387 16892 27828 17058
rect 27387 16840 27476 16892
rect 27528 16840 27688 16892
rect 27740 16840 27828 16892
rect 27387 16675 27828 16840
rect 27387 16623 27476 16675
rect 27528 16623 27688 16675
rect 27740 16623 27828 16675
rect 27387 16470 27828 16623
rect 27387 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 27387 16405 27476 16414
rect 27528 16405 27688 16414
rect 27740 16405 27828 16414
rect 27387 16253 27828 16405
rect 27387 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 27387 16187 27476 16197
rect 27528 16187 27688 16197
rect 27740 16187 27828 16197
rect 27387 16035 27828 16187
rect 27387 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 27387 15970 27476 15979
rect 27528 15970 27688 15979
rect 27740 15970 27828 15979
rect 27387 15818 27828 15970
rect 27387 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 27387 15752 27476 15762
rect 27528 15752 27688 15762
rect 27740 15752 27828 15762
rect 27387 15600 27828 15752
rect 27387 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 27387 15534 27476 15544
rect 27528 15534 27688 15544
rect 27740 15534 27828 15544
rect 27387 15382 27828 15534
rect 27387 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 27387 15317 27476 15326
rect 27528 15317 27688 15326
rect 27740 15317 27828 15326
rect 27387 15164 27828 15317
rect 27387 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 27387 15099 27476 15108
rect 27528 15099 27688 15108
rect 27740 15099 27828 15108
rect 27387 14947 27828 15099
rect 27387 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14891 27828 14947
rect 27387 14881 27476 14891
rect 27528 14881 27688 14891
rect 27740 14881 27828 14891
rect 27387 14729 27828 14881
rect 27387 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 27828 14729
rect 27387 14664 27476 14673
rect 27528 14664 27688 14673
rect 27740 14664 27828 14673
rect 27387 14512 27828 14664
rect 27387 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14456 27828 14512
rect 27387 14446 27476 14456
rect 27528 14446 27688 14456
rect 27740 14446 27828 14456
rect 27387 14281 27828 14446
rect 27387 14231 27476 14281
rect 27528 14231 27688 14281
rect 27740 14231 27828 14281
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 27828 14231
rect 27387 14063 27828 14175
rect 27387 14014 27476 14063
rect 27528 14014 27688 14063
rect 27740 14014 27828 14063
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 27828 14014
rect 27387 13845 27828 13958
rect 27387 13796 27476 13845
rect 27528 13796 27688 13845
rect 27740 13796 27828 13845
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13740 27828 13796
rect 27387 13628 27828 13740
rect 27387 13578 27476 13628
rect 27528 13578 27688 13628
rect 27740 13578 27828 13628
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 27828 13578
rect 27387 13410 27828 13522
rect 27387 13361 27476 13410
rect 27528 13361 27688 13410
rect 27740 13361 27828 13410
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 27828 13361
rect 27387 13192 27828 13305
rect 27387 13140 27476 13192
rect 27528 13140 27688 13192
rect 27740 13140 27828 13192
rect 27387 12975 27828 13140
rect 27387 12923 27476 12975
rect 27528 12923 27688 12975
rect 27740 12923 27828 12975
rect 27387 12757 27828 12923
rect 27387 12705 27476 12757
rect 27528 12705 27688 12757
rect 27740 12705 27828 12757
rect 27387 12540 27828 12705
rect 27387 12488 27476 12540
rect 27528 12488 27688 12540
rect 27740 12488 27828 12540
rect 27387 12322 27828 12488
rect 27387 12270 27476 12322
rect 27528 12270 27688 12322
rect 27740 12270 27828 12322
rect 27387 12104 27828 12270
rect 27387 12052 27476 12104
rect 27528 12052 27688 12104
rect 27740 12052 27828 12104
rect 27387 11887 27828 12052
rect 27387 11835 27476 11887
rect 27528 11835 27688 11887
rect 27740 11835 27828 11887
rect 27387 11669 27828 11835
rect 27387 11617 27476 11669
rect 27528 11617 27688 11669
rect 27740 11617 27828 11669
rect 27387 11451 27828 11617
rect 27387 11406 27476 11451
rect 27528 11406 27688 11451
rect 27740 11406 27828 11451
rect 27387 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 27387 11234 27828 11350
rect 27387 11189 27476 11234
rect 27528 11189 27688 11234
rect 27740 11189 27828 11234
rect 27387 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 27387 11016 27828 11133
rect 27387 10971 27476 11016
rect 27528 10971 27688 11016
rect 27740 10971 27828 11016
rect 27387 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 27387 10798 27828 10915
rect 27387 10753 27476 10798
rect 27528 10753 27688 10798
rect 27740 10753 27828 10798
rect 27387 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 27387 10581 27828 10697
rect 27387 10535 27476 10581
rect 27528 10535 27688 10581
rect 27740 10535 27828 10581
rect 27387 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 27387 10363 27828 10479
rect 27387 10318 27476 10363
rect 27528 10318 27688 10363
rect 27740 10318 27828 10363
rect 27387 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 27387 10146 27828 10262
rect 27387 10094 27476 10146
rect 27528 10094 27688 10146
rect 27740 10094 27828 10146
rect 27387 9928 27828 10094
rect 57295 33215 57736 33380
rect 57295 33163 57383 33215
rect 57435 33163 57595 33215
rect 57647 33163 57736 33215
rect 57295 33141 57736 33163
rect 57295 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 57295 32997 57736 33085
rect 57295 32945 57383 32997
rect 57435 32945 57595 32997
rect 57647 32945 57736 32997
rect 57295 32923 57736 32945
rect 57295 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 57295 32779 57736 32867
rect 57295 32727 57383 32779
rect 57435 32727 57595 32779
rect 57647 32727 57736 32779
rect 57295 32705 57736 32727
rect 57295 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 57295 32562 57736 32649
rect 57295 32510 57383 32562
rect 57435 32510 57595 32562
rect 57647 32510 57736 32562
rect 57295 32487 57736 32510
rect 57295 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 57295 32344 57736 32431
rect 57295 32292 57383 32344
rect 57435 32292 57595 32344
rect 57647 32292 57736 32344
rect 57295 32127 57736 32292
rect 57295 32075 57383 32127
rect 57435 32075 57595 32127
rect 57647 32075 57736 32127
rect 57295 31909 57736 32075
rect 57295 31857 57383 31909
rect 57435 31857 57595 31909
rect 57647 31857 57736 31909
rect 57295 31691 57736 31857
rect 57295 31639 57383 31691
rect 57435 31639 57595 31691
rect 57647 31639 57736 31691
rect 57295 31474 57736 31639
rect 57295 31422 57383 31474
rect 57435 31422 57595 31474
rect 57647 31422 57736 31474
rect 57295 31256 57736 31422
rect 57295 31252 57383 31256
rect 57435 31252 57595 31256
rect 57647 31252 57736 31256
rect 57295 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31196 57736 31252
rect 57295 31038 57736 31196
rect 57295 31034 57383 31038
rect 57435 31034 57595 31038
rect 57647 31034 57736 31038
rect 57295 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30978 57736 31034
rect 57295 30821 57736 30978
rect 57295 30816 57383 30821
rect 57435 30816 57595 30821
rect 57647 30816 57736 30821
rect 57295 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30760 57736 30816
rect 57295 30603 57736 30760
rect 57295 30598 57383 30603
rect 57435 30598 57595 30603
rect 57647 30598 57736 30603
rect 57295 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30542 57736 30598
rect 57295 30386 57736 30542
rect 57295 30334 57383 30386
rect 57435 30334 57595 30386
rect 57647 30334 57736 30386
rect 57295 30168 57736 30334
rect 57295 30116 57383 30168
rect 57435 30116 57595 30168
rect 57647 30116 57736 30168
rect 57295 29950 57736 30116
rect 57295 29898 57383 29950
rect 57435 29898 57595 29950
rect 57647 29898 57736 29950
rect 57295 29733 57736 29898
rect 57295 29681 57383 29733
rect 57435 29681 57595 29733
rect 57647 29681 57736 29733
rect 57295 29515 57736 29681
rect 57295 29463 57383 29515
rect 57435 29463 57595 29515
rect 57647 29463 57736 29515
rect 57295 29297 57736 29463
rect 57295 29245 57383 29297
rect 57435 29245 57595 29297
rect 57647 29245 57736 29297
rect 57295 29080 57736 29245
rect 57295 29028 57383 29080
rect 57435 29028 57595 29080
rect 57647 29028 57736 29080
rect 57295 28862 57736 29028
rect 57295 28810 57383 28862
rect 57435 28810 57595 28862
rect 57647 28810 57736 28862
rect 57295 28644 57736 28810
rect 57295 28592 57383 28644
rect 57435 28592 57595 28644
rect 57647 28592 57736 28644
rect 57295 28427 57736 28592
rect 57295 28375 57383 28427
rect 57435 28375 57595 28427
rect 57647 28375 57736 28427
rect 57295 28209 57736 28375
rect 57295 28157 57383 28209
rect 57435 28157 57595 28209
rect 57647 28157 57736 28209
rect 57295 27992 57736 28157
rect 57295 27940 57383 27992
rect 57435 27940 57595 27992
rect 57647 27940 57736 27992
rect 57295 27774 57736 27940
rect 57295 27722 57383 27774
rect 57435 27722 57595 27774
rect 57647 27722 57736 27774
rect 57295 27556 57736 27722
rect 57295 27504 57383 27556
rect 57435 27504 57595 27556
rect 57647 27504 57736 27556
rect 57295 27339 57736 27504
rect 57295 27287 57383 27339
rect 57435 27287 57595 27339
rect 57647 27287 57736 27339
rect 57295 27121 57736 27287
rect 57295 27069 57383 27121
rect 57435 27069 57595 27121
rect 57647 27069 57736 27121
rect 57295 26903 57736 27069
rect 57295 26851 57383 26903
rect 57435 26851 57595 26903
rect 57647 26851 57736 26903
rect 57295 26799 57736 26851
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 57736 26799
rect 57295 26686 57736 26743
rect 57295 26634 57383 26686
rect 57435 26634 57595 26686
rect 57647 26634 57736 26686
rect 57295 26581 57736 26634
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 57736 26581
rect 57295 26468 57736 26525
rect 57295 26416 57383 26468
rect 57435 26416 57595 26468
rect 57647 26416 57736 26468
rect 57295 26250 57736 26416
rect 57295 26198 57383 26250
rect 57435 26198 57595 26250
rect 57647 26198 57736 26250
rect 57295 26033 57736 26198
rect 57295 25981 57383 26033
rect 57435 25981 57595 26033
rect 57647 25981 57736 26033
rect 57295 25815 57736 25981
rect 57295 25763 57383 25815
rect 57435 25763 57595 25815
rect 57647 25763 57736 25815
rect 57295 25598 57736 25763
rect 57295 25546 57383 25598
rect 57435 25546 57595 25598
rect 57647 25546 57736 25598
rect 57295 25380 57736 25546
rect 57295 25328 57383 25380
rect 57435 25328 57595 25380
rect 57647 25328 57736 25380
rect 57295 25162 57736 25328
rect 57295 25110 57383 25162
rect 57435 25110 57595 25162
rect 57647 25110 57736 25162
rect 57295 24945 57736 25110
rect 57295 24893 57383 24945
rect 57435 24893 57595 24945
rect 57647 24893 57736 24945
rect 57295 24727 57736 24893
rect 57295 24675 57383 24727
rect 57435 24675 57595 24727
rect 57647 24675 57736 24727
rect 57295 24509 57736 24675
rect 57295 24457 57383 24509
rect 57435 24457 57595 24509
rect 57647 24457 57736 24509
rect 57295 24292 57736 24457
rect 57295 24240 57383 24292
rect 57435 24240 57595 24292
rect 57647 24240 57736 24292
rect 57295 24074 57736 24240
rect 57295 24022 57383 24074
rect 57435 24022 57595 24074
rect 57647 24022 57736 24074
rect 57295 23857 57736 24022
rect 57295 23805 57383 23857
rect 57435 23805 57595 23857
rect 57647 23805 57736 23857
rect 57295 23639 57736 23805
rect 57295 23587 57383 23639
rect 57435 23587 57595 23639
rect 57647 23587 57736 23639
rect 57295 23421 57736 23587
rect 57295 23369 57383 23421
rect 57435 23369 57595 23421
rect 57647 23369 57736 23421
rect 57295 23204 57736 23369
rect 57295 23152 57383 23204
rect 57435 23152 57595 23204
rect 57647 23152 57736 23204
rect 57295 22986 57736 23152
rect 57295 22934 57383 22986
rect 57435 22934 57595 22986
rect 57647 22934 57736 22986
rect 57295 22923 57736 22934
rect 57295 22035 57363 22923
rect 57627 22768 57736 22923
rect 57647 22716 57736 22768
rect 57627 22551 57736 22716
rect 57647 22499 57736 22551
rect 57627 22333 57736 22499
rect 57647 22281 57736 22333
rect 57627 22115 57736 22281
rect 57647 22063 57736 22115
rect 57627 22035 57736 22063
rect 57295 21898 57736 22035
rect 57295 21846 57383 21898
rect 57435 21846 57595 21898
rect 57647 21846 57736 21898
rect 57295 21680 57736 21846
rect 57295 21628 57383 21680
rect 57435 21628 57595 21680
rect 57647 21628 57736 21680
rect 57295 21463 57736 21628
rect 57295 21411 57383 21463
rect 57435 21411 57595 21463
rect 57647 21411 57736 21463
rect 57295 21245 57736 21411
rect 57295 21193 57383 21245
rect 57435 21193 57595 21245
rect 57647 21193 57736 21245
rect 57295 21027 57736 21193
rect 57295 20975 57383 21027
rect 57435 20975 57595 21027
rect 57647 20975 57736 21027
rect 57295 20810 57736 20975
rect 57295 20758 57383 20810
rect 57435 20758 57595 20810
rect 57647 20758 57736 20810
rect 57295 20592 57736 20758
rect 57295 20540 57383 20592
rect 57435 20540 57595 20592
rect 57647 20540 57736 20592
rect 57295 20374 57736 20540
rect 57295 20322 57383 20374
rect 57435 20322 57595 20374
rect 57647 20322 57736 20374
rect 57295 20157 57736 20322
rect 57295 20105 57383 20157
rect 57435 20105 57595 20157
rect 57647 20105 57736 20157
rect 57295 19939 57736 20105
rect 57295 19887 57383 19939
rect 57435 19887 57595 19939
rect 57647 19887 57736 19939
rect 57295 19722 57736 19887
rect 57295 19670 57383 19722
rect 57435 19670 57595 19722
rect 57647 19670 57736 19722
rect 57295 19504 57736 19670
rect 57295 19452 57383 19504
rect 57435 19452 57595 19504
rect 57647 19452 57736 19504
rect 57295 19286 57736 19452
rect 57295 19234 57383 19286
rect 57435 19234 57595 19286
rect 57647 19234 57736 19286
rect 57295 19068 57736 19234
rect 57295 19016 57383 19068
rect 57435 19016 57595 19068
rect 57647 19016 57736 19068
rect 57295 18851 57736 19016
rect 57295 18799 57383 18851
rect 57435 18799 57595 18851
rect 57647 18799 57736 18851
rect 57295 18633 57736 18799
rect 57295 18581 57383 18633
rect 57435 18581 57595 18633
rect 57647 18581 57736 18633
rect 57295 18416 57736 18581
rect 57295 18364 57383 18416
rect 57435 18364 57595 18416
rect 57647 18364 57736 18416
rect 57295 18198 57736 18364
rect 57295 18146 57383 18198
rect 57435 18146 57595 18198
rect 57647 18146 57736 18198
rect 57295 17980 57736 18146
rect 57295 17928 57383 17980
rect 57435 17928 57595 17980
rect 57647 17928 57736 17980
rect 57295 17763 57736 17928
rect 57295 17711 57383 17763
rect 57435 17711 57595 17763
rect 57647 17711 57736 17763
rect 57295 17545 57736 17711
rect 57295 17493 57383 17545
rect 57435 17493 57595 17545
rect 57647 17493 57736 17545
rect 57295 17327 57736 17493
rect 57295 17275 57383 17327
rect 57435 17275 57595 17327
rect 57647 17275 57736 17327
rect 57295 17110 57736 17275
rect 57295 17058 57383 17110
rect 57435 17058 57595 17110
rect 57647 17058 57736 17110
rect 57295 16892 57736 17058
rect 57295 16840 57383 16892
rect 57435 16840 57595 16892
rect 57647 16840 57736 16892
rect 57295 16678 57736 16840
rect 57295 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 57736 16678
rect 57295 16461 57736 16622
rect 57295 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 57736 16461
rect 57295 16243 57736 16405
rect 57295 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 57736 16243
rect 57295 16026 57736 16187
rect 57295 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 57736 16026
rect 57295 15808 57736 15970
rect 57295 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 57736 15808
rect 57295 15590 57736 15752
rect 57295 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 57736 15590
rect 57295 15372 57736 15534
rect 57295 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 57736 15372
rect 57295 15155 57736 15316
rect 57295 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 57736 15155
rect 57295 14937 57736 15099
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 57736 14937
rect 57295 14720 57736 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 57736 14720
rect 57295 14498 57736 14664
rect 57295 14446 57383 14498
rect 57435 14446 57595 14498
rect 57647 14446 57736 14498
rect 57295 14281 57736 14446
rect 57295 14229 57383 14281
rect 57435 14229 57595 14281
rect 57647 14229 57736 14281
rect 57295 14063 57736 14229
rect 57295 14011 57383 14063
rect 57435 14011 57595 14063
rect 57647 14011 57736 14063
rect 57295 13845 57736 14011
rect 57295 13793 57383 13845
rect 57435 13793 57595 13845
rect 57647 13793 57736 13845
rect 57295 13628 57736 13793
rect 57295 13576 57383 13628
rect 57435 13576 57595 13628
rect 57647 13576 57736 13628
rect 57295 13410 57736 13576
rect 57295 13358 57383 13410
rect 57435 13358 57595 13410
rect 57647 13358 57736 13410
rect 57295 13192 57736 13358
rect 57295 13140 57383 13192
rect 57435 13140 57595 13192
rect 57647 13140 57736 13192
rect 57295 12975 57736 13140
rect 57295 12923 57383 12975
rect 57435 12923 57595 12975
rect 57647 12923 57736 12975
rect 57295 12757 57736 12923
rect 57295 12705 57383 12757
rect 57435 12705 57595 12757
rect 57647 12705 57736 12757
rect 57295 12540 57736 12705
rect 57295 12488 57383 12540
rect 57435 12488 57595 12540
rect 57647 12488 57736 12540
rect 57295 12322 57736 12488
rect 57295 12270 57383 12322
rect 57435 12270 57595 12322
rect 57647 12270 57736 12322
rect 57295 12104 57736 12270
rect 57295 12052 57383 12104
rect 57435 12052 57595 12104
rect 57647 12052 57736 12104
rect 57295 11887 57736 12052
rect 57295 11835 57383 11887
rect 57435 11835 57595 11887
rect 57647 11835 57736 11887
rect 57295 11669 57736 11835
rect 57295 11617 57383 11669
rect 57435 11617 57595 11669
rect 57647 11617 57736 11669
rect 57295 11451 57736 11617
rect 57295 11406 57383 11451
rect 57435 11406 57595 11451
rect 57647 11406 57736 11451
rect 57295 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 57736 11406
rect 57295 11234 57736 11350
rect 57295 11189 57383 11234
rect 57435 11189 57595 11234
rect 57647 11189 57736 11234
rect 57295 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 57736 11189
rect 57295 11016 57736 11133
rect 57295 10971 57383 11016
rect 57435 10971 57595 11016
rect 57647 10971 57736 11016
rect 57295 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 57736 10971
rect 57295 10798 57736 10915
rect 57295 10753 57383 10798
rect 57435 10753 57595 10798
rect 57647 10753 57736 10798
rect 57295 10697 57381 10753
rect 57437 10697 57593 10753
rect 57649 10697 57736 10753
rect 57295 10581 57736 10697
rect 57295 10535 57383 10581
rect 57435 10535 57595 10581
rect 57647 10535 57736 10581
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 57736 10535
rect 57295 10363 57736 10479
rect 57295 10318 57383 10363
rect 57435 10318 57595 10363
rect 57647 10318 57736 10363
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 57736 10318
rect 57295 10146 57736 10262
rect 57295 10094 57383 10146
rect 57435 10094 57595 10146
rect 57647 10094 57736 10146
rect 27387 9876 27476 9928
rect 27528 9876 27688 9928
rect 27740 9876 27828 9928
rect 27387 9710 27828 9876
rect 51756 9971 51832 9981
rect 51756 9811 51766 9971
rect 51822 9811 51832 9971
rect 51756 9801 51832 9811
rect 57295 9928 57736 10094
rect 57295 9876 57383 9928
rect 57435 9876 57595 9928
rect 57647 9876 57736 9928
rect 27387 9658 27476 9710
rect 27528 9658 27688 9710
rect 27740 9658 27828 9710
rect 27387 9493 27828 9658
rect 27387 9441 27476 9493
rect 27528 9441 27688 9493
rect 27740 9441 27828 9493
rect 27387 9275 27828 9441
rect 27387 9223 27476 9275
rect 27528 9223 27688 9275
rect 27740 9223 27828 9275
rect 27387 9057 27828 9223
rect 27387 9005 27476 9057
rect 27528 9005 27688 9057
rect 27740 9005 27828 9057
rect 27387 8840 27828 9005
rect 49887 8953 50067 8963
rect 49887 8897 49897 8953
rect 50057 8897 50067 8953
rect 49887 8887 50067 8897
rect 27387 8788 27476 8840
rect 27528 8788 27688 8840
rect 27740 8788 27828 8840
rect 27387 8622 27828 8788
rect 27387 8570 27476 8622
rect 27528 8570 27688 8622
rect 27740 8570 27828 8622
rect 27387 8404 27828 8570
rect 27387 8352 27476 8404
rect 27528 8352 27688 8404
rect 27740 8352 27828 8404
rect 27387 8187 27828 8352
rect 27387 8135 27476 8187
rect 27528 8135 27688 8187
rect 27740 8135 27828 8187
rect 27387 7969 27828 8135
rect 27387 7917 27476 7969
rect 27528 7917 27688 7969
rect 27740 7917 27828 7969
rect 27387 7752 27828 7917
rect 27387 7700 27476 7752
rect 27528 7700 27688 7752
rect 27740 7700 27828 7752
rect 27387 7535 27828 7700
rect 27387 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 27387 7317 27828 7479
rect 27387 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 27387 7099 27828 7261
rect 27387 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 27387 6881 27828 7043
rect 27387 6829 27476 6881
rect 27528 6829 27688 6881
rect 27740 6829 27828 6881
rect 27387 6663 27828 6829
rect 27387 6611 27476 6663
rect 27528 6611 27688 6663
rect 27740 6611 27828 6663
rect 27387 6446 27828 6611
rect 27387 6394 27476 6446
rect 27528 6394 27688 6446
rect 27740 6394 27828 6446
rect 27387 6228 27828 6394
rect 28237 6836 28999 6874
rect 28237 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 28999 6836
rect 28237 6618 28999 6780
rect 28237 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 28999 6618
rect 28237 6400 28999 6562
rect 28237 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 28999 6400
rect 49958 6361 50014 8887
rect 28237 6306 28999 6344
rect 49896 6349 50076 6361
rect 49896 6297 49908 6349
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6176 27476 6228
rect 27528 6176 27688 6228
rect 27740 6176 27828 6228
rect 27387 6120 27828 6176
rect 27387 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 27828 6120
rect 27387 6011 27828 6064
rect 27387 5959 27476 6011
rect 27528 5959 27688 6011
rect 27740 5959 27828 6011
rect 27387 5902 27828 5959
rect 27387 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 27828 5902
rect 27387 5793 27828 5846
rect 27387 5741 27476 5793
rect 27528 5741 27688 5793
rect 27740 5741 27828 5793
rect 27387 5575 27828 5741
rect 27387 5523 27476 5575
rect 27528 5523 27688 5575
rect 27740 5523 27828 5575
rect 27387 5358 27828 5523
rect 27387 5306 27476 5358
rect 27528 5306 27688 5358
rect 27740 5306 27828 5358
rect 1864 5024 2509 5135
rect 11727 5073 11783 5140
rect 1864 0 2088 5024
rect 3263 5001 3357 5062
rect 11617 5017 11783 5073
rect 3263 4880 3539 5001
rect 3445 1701 3539 4880
rect 11617 1701 11673 5017
rect 12575 4740 12631 5185
rect 12290 4684 12631 4740
rect 13253 4740 13309 5185
rect 14101 5073 14157 5140
rect 14101 5017 14267 5073
rect 13253 4684 13594 4740
rect 12290 1701 12346 4684
rect 13538 1701 13594 4684
rect 14211 1701 14267 5017
rect 22527 5001 22621 5062
rect 23375 5024 23953 5135
rect 22345 4880 22621 5001
rect 22345 1701 22439 4880
rect 23859 3382 23953 5024
rect 26823 4587 27163 4628
rect 26823 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27163 4587
rect 26823 4528 27163 4535
rect 26823 4472 26859 4528
rect 26915 4472 27071 4528
rect 27127 4472 27163 4528
rect 26823 4370 27163 4472
rect 26823 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27163 4370
rect 26823 4310 27163 4318
rect 26823 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 27163 4310
rect 26823 4152 27163 4254
rect 26823 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27163 4152
rect 26823 3934 27163 4100
rect 26823 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27163 3934
rect 26823 3717 27163 3882
rect 26823 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27163 3717
rect 26823 3624 27163 3665
rect 27387 4587 27828 5306
rect 27387 4535 27476 4587
rect 27528 4535 27688 4587
rect 27740 4535 27828 4587
rect 27387 4370 27828 4535
rect 27387 4318 27476 4370
rect 27528 4318 27688 4370
rect 27740 4318 27828 4370
rect 27387 4152 27828 4318
rect 27387 4100 27476 4152
rect 27528 4100 27688 4152
rect 27740 4100 27828 4152
rect 27387 3934 27828 4100
rect 27387 3882 27476 3934
rect 27528 3882 27688 3934
rect 27740 3882 27828 3934
rect 27387 3837 27828 3882
rect 27387 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 27828 3837
rect 27387 3717 27828 3781
rect 27387 3665 27476 3717
rect 27528 3665 27688 3717
rect 27740 3665 27828 3717
rect 27387 3619 27828 3665
rect 27387 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 27828 3619
rect 27387 3524 27828 3563
rect 28764 3837 28894 3876
rect 28764 3781 28801 3837
rect 28857 3781 28894 3837
rect 28764 3619 28894 3781
rect 28764 3563 28801 3619
rect 28857 3563 28894 3619
rect 28764 3525 28894 3563
rect 2539 1689 2763 1701
rect 2539 1637 2574 1689
rect 2730 1637 2763 1689
rect 2539 0 2763 1637
rect 3380 0 3604 1701
rect 11533 0 11757 1701
rect 12206 0 12430 1701
rect 12604 1689 12828 1701
rect 12604 1637 12639 1689
rect 12795 1637 12828 1689
rect 12604 0 12828 1637
rect 13054 1689 13278 1701
rect 13054 1637 13089 1689
rect 13245 1637 13278 1689
rect 13054 0 13278 1637
rect 13454 0 13678 1701
rect 14127 0 14351 1701
rect 22279 0 22503 1701
rect 23404 1689 23628 1701
rect 23404 1637 23439 1689
rect 23595 1637 23628 1689
rect 23404 0 23628 1637
rect 23795 0 24019 3382
rect 27936 0 28160 3382
rect 29006 2524 29135 3418
rect 29247 3004 29377 3418
rect 29247 2768 29929 3004
rect 29006 0 29230 2524
rect 29705 0 29929 2768
rect 30859 0 31083 6229
rect 32552 0 32776 6229
rect 34243 0 34467 6229
rect 40588 3282 40812 3294
rect 40588 3230 40623 3282
rect 40779 3230 40812 3282
rect 40588 0 40812 3230
rect 43790 3050 43970 3060
rect 43790 2994 43800 3050
rect 43960 2994 43970 3050
rect 43790 2984 43970 2994
rect 50342 0 50566 7278
rect 51766 5211 51822 9801
rect 57295 9710 57736 9876
rect 57295 9658 57383 9710
rect 57435 9658 57595 9710
rect 57647 9658 57736 9710
rect 57295 9493 57736 9658
rect 57295 9441 57383 9493
rect 57435 9441 57595 9493
rect 57647 9441 57736 9493
rect 57295 9275 57736 9441
rect 57295 9223 57383 9275
rect 57435 9223 57595 9275
rect 57647 9223 57736 9275
rect 57295 9057 57736 9223
rect 57295 9005 57383 9057
rect 57435 9005 57595 9057
rect 57647 9005 57736 9057
rect 57295 8843 57736 9005
rect 57295 8787 57381 8843
rect 57437 8787 57593 8843
rect 57649 8787 57736 8843
rect 57295 8625 57736 8787
rect 57295 8569 57381 8625
rect 57437 8569 57593 8625
rect 57649 8569 57736 8625
rect 57295 8408 57736 8569
rect 57295 8352 57381 8408
rect 57437 8352 57593 8408
rect 57649 8352 57736 8408
rect 57295 8190 57736 8352
rect 57295 8134 57381 8190
rect 57437 8134 57593 8190
rect 57649 8134 57736 8190
rect 57295 7972 57736 8134
rect 57295 7916 57381 7972
rect 57437 7916 57593 7972
rect 57649 7916 57736 7972
rect 57295 7755 57736 7916
rect 57295 7699 57381 7755
rect 57437 7699 57593 7755
rect 57649 7699 57736 7755
rect 57295 7537 57736 7699
rect 57295 7481 57381 7537
rect 57437 7481 57593 7537
rect 57649 7481 57736 7537
rect 57295 7319 57736 7481
rect 57295 7263 57381 7319
rect 57437 7263 57593 7319
rect 57649 7263 57736 7319
rect 57295 7102 57736 7263
rect 57295 7046 57381 7102
rect 57437 7046 57593 7102
rect 57649 7046 57736 7102
rect 57295 6881 57736 7046
rect 56124 6836 56886 6874
rect 56124 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 56886 6836
rect 56124 6618 56886 6780
rect 56124 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 56886 6618
rect 56124 6400 56886 6562
rect 56124 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 56886 6400
rect 56124 6306 56886 6344
rect 57295 6829 57383 6881
rect 57435 6829 57595 6881
rect 57647 6829 57736 6881
rect 57295 6663 57736 6829
rect 57295 6611 57383 6663
rect 57435 6611 57595 6663
rect 57647 6611 57736 6663
rect 57295 6446 57736 6611
rect 57295 6394 57383 6446
rect 57435 6394 57595 6446
rect 57647 6394 57736 6446
rect 51642 5199 51822 5211
rect 51642 5147 51654 5199
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 6228 57736 6394
rect 57295 6176 57383 6228
rect 57435 6176 57595 6228
rect 57647 6176 57736 6228
rect 57295 6120 57736 6176
rect 57295 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 57736 6120
rect 57295 6011 57736 6064
rect 57295 5959 57383 6011
rect 57435 5959 57595 6011
rect 57647 5959 57736 6011
rect 57295 5902 57736 5959
rect 57295 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 57736 5902
rect 57295 5793 57736 5846
rect 57295 5741 57383 5793
rect 57435 5741 57595 5793
rect 57647 5741 57736 5793
rect 57295 5575 57736 5741
rect 57295 5523 57383 5575
rect 57435 5523 57595 5575
rect 57647 5523 57736 5575
rect 57295 5358 57736 5523
rect 57295 5306 57383 5358
rect 57435 5306 57595 5358
rect 57647 5306 57736 5358
rect 57295 4587 57736 5306
rect 57295 4535 57383 4587
rect 57435 4535 57595 4587
rect 57647 4535 57736 4587
rect 57295 4370 57736 4535
rect 57295 4318 57383 4370
rect 57435 4318 57595 4370
rect 57647 4318 57736 4370
rect 57295 4152 57736 4318
rect 57295 4100 57383 4152
rect 57435 4100 57595 4152
rect 57647 4100 57736 4152
rect 57295 3934 57736 4100
rect 57295 3882 57383 3934
rect 57435 3882 57595 3934
rect 57647 3882 57736 3934
rect 57295 3837 57736 3882
rect 57295 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 57736 3837
rect 53772 3247 55669 3471
rect 53772 0 53996 3247
rect 55781 3024 55911 3418
rect 54417 2800 55911 3024
rect 54417 0 54641 2800
rect 56023 2540 56152 3418
rect 55164 2316 56152 2540
rect 55164 0 55388 2316
rect 56265 0 56489 3729
rect 57295 3717 57736 3781
rect 57295 3665 57383 3717
rect 57435 3665 57595 3717
rect 57647 3665 57736 3717
rect 57295 3619 57736 3665
rect 57295 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 57736 3619
rect 57295 3524 57736 3563
rect 57909 33432 58351 33520
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33358 58351 33380
rect 57909 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 58351 33358
rect 57909 33215 58351 33302
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 33140 58351 33163
rect 57909 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 58351 33140
rect 57909 32997 58351 33084
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32922 58351 32945
rect 57909 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 58351 32922
rect 57909 32779 58351 32866
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32705 58351 32727
rect 57909 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 58351 32705
rect 57909 32562 58351 32649
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32487 58351 32510
rect 57909 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 58351 32487
rect 57909 32344 58351 32431
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32088 57998 32127
rect 58050 32088 58210 32127
rect 58262 32088 58351 32127
rect 57909 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 57909 31909 58351 32032
rect 57909 31870 57998 31909
rect 58050 31870 58210 31909
rect 58262 31870 58351 31909
rect 57909 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 57909 31691 58351 31814
rect 57909 31652 57998 31691
rect 58050 31652 58210 31691
rect 58262 31652 58351 31691
rect 57909 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 57909 31474 58351 31596
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29968 58351 30116
rect 57909 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 57909 29898 57998 29912
rect 58050 29898 58210 29912
rect 58262 29898 58351 29912
rect 57909 29750 58351 29898
rect 57909 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29694 58351 29750
rect 57909 29681 57998 29694
rect 58050 29681 58210 29694
rect 58262 29681 58351 29694
rect 57909 29533 58351 29681
rect 57909 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 58351 29533
rect 57909 29463 57998 29477
rect 58050 29463 58210 29477
rect 58262 29463 58351 29477
rect 57909 29315 58351 29463
rect 57909 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 57909 29245 57998 29259
rect 58050 29245 58210 29259
rect 58262 29245 58351 29259
rect 57909 29098 58351 29245
rect 57909 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 57909 29028 57998 29042
rect 58050 29028 58210 29042
rect 58262 29028 58351 29042
rect 57909 28880 58351 29028
rect 57909 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 57909 28810 57998 28824
rect 58050 28810 58210 28824
rect 58262 28810 58351 28824
rect 57909 28662 58351 28810
rect 57909 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 57909 28592 57998 28606
rect 58050 28592 58210 28606
rect 58262 28592 58351 28606
rect 57909 28444 58351 28592
rect 57909 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 57909 28375 57998 28388
rect 58050 28375 58210 28388
rect 58262 28375 58351 28388
rect 57909 28227 58351 28375
rect 57909 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 57909 28157 57998 28171
rect 58050 28157 58210 28171
rect 58262 28157 58351 28171
rect 57909 28009 58351 28157
rect 57909 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 57909 27940 57998 27953
rect 58050 27940 58210 27953
rect 58262 27940 58351 27953
rect 57909 27792 58351 27940
rect 57909 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 57909 27722 57998 27736
rect 58050 27722 58210 27736
rect 58262 27722 58351 27736
rect 57909 27574 58351 27722
rect 57909 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 57909 27504 57998 27518
rect 58050 27504 58210 27518
rect 58262 27504 58351 27518
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 58791 94775 59517 94794
rect 58791 94719 58865 94775
rect 58921 94719 58989 94775
rect 59045 94719 59113 94775
rect 59169 94719 59237 94775
rect 59293 94719 59361 94775
rect 59417 94719 59517 94775
rect 58791 94651 59517 94719
rect 58791 94595 58865 94651
rect 58921 94595 58989 94651
rect 59045 94595 59113 94651
rect 59169 94595 59237 94651
rect 59293 94595 59361 94651
rect 59417 94595 59517 94651
rect 58791 94527 59517 94595
rect 58791 94471 58865 94527
rect 58921 94471 58989 94527
rect 59045 94471 59113 94527
rect 59169 94471 59237 94527
rect 59293 94471 59361 94527
rect 59417 94471 59517 94527
rect 58791 34992 59517 94471
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 58791 34936 58816 34992
rect 58872 34936 58940 34992
rect 58996 34936 59064 34992
rect 59120 34936 59188 34992
rect 59244 34936 59312 34992
rect 59368 34936 59436 34992
rect 59492 34936 59517 34992
rect 58791 34868 59517 34936
rect 58791 34812 58816 34868
rect 58872 34812 58940 34868
rect 58996 34812 59064 34868
rect 59120 34812 59188 34868
rect 59244 34812 59312 34868
rect 59368 34812 59436 34868
rect 59492 34812 59517 34868
rect 58791 34744 59517 34812
rect 58791 34688 58816 34744
rect 58872 34688 58940 34744
rect 58996 34688 59064 34744
rect 59120 34688 59188 34744
rect 59244 34688 59312 34744
rect 59368 34688 59436 34744
rect 59492 34688 59517 34744
rect 58791 34620 59517 34688
rect 58791 34564 58816 34620
rect 58872 34564 58940 34620
rect 58996 34564 59064 34620
rect 59120 34564 59188 34620
rect 59244 34564 59312 34620
rect 59368 34564 59436 34620
rect 59492 34564 59517 34620
rect 58791 31298 59517 34564
rect 58791 31242 58873 31298
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59517 31298
rect 58791 31174 59517 31242
rect 58791 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59517 31174
rect 58791 31050 59517 31118
rect 58791 30994 58873 31050
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59517 31050
rect 58791 30853 59517 30994
rect 58791 30797 58873 30853
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59517 30853
rect 58791 30729 59517 30797
rect 58791 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59517 30729
rect 58791 30605 59517 30673
rect 58791 30549 58873 30605
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59517 30605
rect 58791 28295 59517 30549
rect 58791 28239 58859 28295
rect 58915 28239 58983 28295
rect 59039 28239 59107 28295
rect 59163 28239 59231 28295
rect 59287 28239 59355 28295
rect 59411 28239 59517 28295
rect 58791 28171 59517 28239
rect 58791 28115 58859 28171
rect 58915 28115 58983 28171
rect 59039 28115 59107 28171
rect 59163 28115 59231 28171
rect 59287 28115 59355 28171
rect 59411 28115 59517 28171
rect 58791 28047 59517 28115
rect 58791 27991 58859 28047
rect 58915 27991 58983 28047
rect 59039 27991 59107 28047
rect 59163 27991 59231 28047
rect 59287 27991 59355 28047
rect 59411 27991 59517 28047
rect 58791 27923 59517 27991
rect 58791 27867 58859 27923
rect 58915 27867 58983 27923
rect 59039 27867 59107 27923
rect 59163 27867 59231 27923
rect 59287 27867 59355 27923
rect 59411 27867 59517 27923
rect 58791 27799 59517 27867
rect 58791 27743 58859 27799
rect 58915 27743 58983 27799
rect 59039 27743 59107 27799
rect 59163 27743 59231 27799
rect 59287 27743 59355 27799
rect 59411 27743 59517 27799
rect 58791 27675 59517 27743
rect 58791 27619 58859 27675
rect 58915 27619 58983 27675
rect 59039 27619 59107 27675
rect 59163 27619 59231 27675
rect 59287 27619 59355 27675
rect 59411 27619 59517 27675
rect 58791 27551 59517 27619
rect 58791 27495 58859 27551
rect 58915 27495 58983 27551
rect 59039 27495 59107 27551
rect 59163 27495 59231 27551
rect 59287 27495 59355 27551
rect 59411 27495 59517 27551
rect 58791 27427 59517 27495
rect 58791 27371 58859 27427
rect 58915 27371 58983 27427
rect 59039 27371 59107 27427
rect 59163 27371 59231 27427
rect 59287 27371 59355 27427
rect 59411 27371 59517 27427
rect 58791 27303 59517 27371
rect 58791 27247 58859 27303
rect 58915 27247 58983 27303
rect 59039 27247 59107 27303
rect 59163 27247 59231 27303
rect 59287 27247 59355 27303
rect 59411 27247 59517 27303
rect 58791 27179 59517 27247
rect 58791 27123 58859 27179
rect 58915 27123 58983 27179
rect 59039 27123 59107 27179
rect 59163 27123 59231 27179
rect 59287 27123 59355 27179
rect 59411 27123 59517 27179
rect 58791 27055 59517 27123
rect 58791 26999 58859 27055
rect 58915 26999 58983 27055
rect 59039 26999 59107 27055
rect 59163 26999 59231 27055
rect 59287 26999 59355 27055
rect 59411 26999 59517 27055
rect 58791 26931 59517 26999
rect 58791 26875 58859 26931
rect 58915 26875 58983 26931
rect 59039 26875 59107 26931
rect 59163 26875 59231 26931
rect 59287 26875 59355 26931
rect 59411 26875 59517 26931
rect 58791 26807 59517 26875
rect 58791 26751 58859 26807
rect 58915 26751 58983 26807
rect 59039 26751 59107 26807
rect 59163 26751 59231 26807
rect 59287 26751 59355 26807
rect 59411 26751 59517 26807
rect 58791 26683 59517 26751
rect 58791 26627 58859 26683
rect 58915 26627 58983 26683
rect 59039 26627 59107 26683
rect 59163 26627 59231 26683
rect 59287 26627 59355 26683
rect 59411 26627 59517 26683
rect 58791 26559 59517 26627
rect 58791 26503 58859 26559
rect 58915 26503 58983 26559
rect 59039 26503 59107 26559
rect 59163 26503 59231 26559
rect 59287 26503 59355 26559
rect 59411 26503 59517 26559
rect 58791 26433 59517 26503
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24075 58351 24240
rect 57909 23187 57994 24075
rect 58258 24074 58351 24075
rect 58262 24022 58351 24074
rect 58258 23857 58351 24022
rect 58262 23805 58351 23857
rect 58258 23639 58351 23805
rect 58262 23587 58351 23639
rect 58258 23421 58351 23587
rect 58262 23369 58351 23421
rect 58258 23204 58351 23369
rect 57909 23152 57998 23187
rect 58050 23152 58210 23187
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20570 58210 20592
rect 58208 20540 58210 20570
rect 58262 20540 58351 20592
rect 57909 20410 58048 20540
rect 58208 20410 58351 20540
rect 57909 20374 58351 20410
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20226 58351 20322
rect 57909 20157 58048 20226
rect 58208 20157 58351 20226
rect 57909 20105 57998 20157
rect 58208 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 20066 58048 20105
rect 58208 20066 58351 20105
rect 57909 19939 58351 20066
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13790 58351 13793
rect 57909 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 58351 13790
rect 57909 13628 58351 13734
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13573 58351 13576
rect 57909 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 58351 13573
rect 57909 13410 58351 13517
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13355 58351 13358
rect 57909 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58351 13355
rect 57909 13192 58351 13299
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 13138 58351 13140
rect 57909 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58351 13138
rect 57909 12975 58351 13082
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12920 58351 12923
rect 57909 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58351 12920
rect 57909 12757 58351 12864
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12702 58351 12705
rect 57909 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 58351 12702
rect 57909 12540 58351 12646
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12484 58351 12488
rect 57909 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 58351 12484
rect 57909 12322 58351 12428
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12267 58351 12270
rect 57909 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 58351 12267
rect 57909 12104 58351 12211
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 12049 58351 12052
rect 57909 11993 57996 12049
rect 58052 11993 58208 12049
rect 58264 11993 58351 12049
rect 57909 11887 58351 11993
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11832 58351 11835
rect 57909 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 57909 11669 58351 11776
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9407 58351 9441
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 58351 9407
rect 57909 9275 58351 9351
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9190 58351 9223
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 58351 9190
rect 57909 9057 58351 9134
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8972 58351 9005
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 58351 8972
rect 57909 8840 58351 8916
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8754 58351 8788
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 58351 8754
rect 57909 8622 58351 8698
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8536 58351 8570
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 58351 8536
rect 57909 8404 58351 8480
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8319 58351 8352
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 58351 8319
rect 57909 8187 58351 8263
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5539 57998 5575
rect 58050 5539 58210 5575
rect 58262 5539 58351 5575
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 58351 5539
rect 57909 5358 58351 5483
rect 57909 5321 57998 5358
rect 58050 5321 58210 5358
rect 58262 5321 58351 5358
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 58351 5321
rect 57909 4587 58351 5265
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4528 58351 4535
rect 57909 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4472 58351 4528
rect 57909 4370 58351 4472
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4310 58351 4318
rect 57909 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 58351 4310
rect 57909 4152 58351 4254
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57909 3524 58351 3665
rect 61447 5024 62085 5135
rect 71303 5073 71359 5140
rect 61447 0 61671 5024
rect 62839 5001 62933 5062
rect 71193 5017 71359 5073
rect 62839 4880 63115 5001
rect 63021 1701 63115 4880
rect 71193 1701 71249 5017
rect 72151 4740 72207 5185
rect 71866 4684 72207 4740
rect 72829 4740 72885 5185
rect 73677 5073 73733 5140
rect 73677 5017 73843 5073
rect 72829 4684 73170 4740
rect 71866 1701 71922 4684
rect 73114 1701 73170 4684
rect 73787 1701 73843 5017
rect 82103 5001 82197 5062
rect 82951 5024 83596 5135
rect 81921 4880 82197 5001
rect 81921 1701 82015 4880
rect 62115 1689 62339 1701
rect 62115 1637 62150 1689
rect 62306 1637 62339 1689
rect 62115 0 62339 1637
rect 62958 0 63182 1701
rect 71109 0 71333 1701
rect 71782 0 72006 1701
rect 72180 1689 72404 1701
rect 72180 1637 72215 1689
rect 72371 1637 72404 1689
rect 72180 0 72404 1637
rect 72630 1689 72854 1701
rect 72630 1637 72665 1689
rect 72821 1637 72854 1689
rect 72630 0 72854 1637
rect 73030 0 73254 1701
rect 73703 0 73927 1701
rect 81855 0 82079 1701
rect 82695 1689 82919 1701
rect 82695 1637 82730 1689
rect 82886 1637 82919 1689
rect 82695 0 82919 1637
rect 83372 0 83596 5024
rect 84666 282 85666 95176
<< via2 >>
rect 25386 94773 25442 94775
rect 25386 94721 25388 94773
rect 25388 94721 25440 94773
rect 25440 94721 25442 94773
rect 25386 94719 25442 94721
rect 25510 94773 25566 94775
rect 25510 94721 25512 94773
rect 25512 94721 25564 94773
rect 25564 94721 25566 94773
rect 25510 94719 25566 94721
rect 25634 94773 25690 94775
rect 25634 94721 25636 94773
rect 25636 94721 25688 94773
rect 25688 94721 25690 94773
rect 25634 94719 25690 94721
rect 25758 94773 25814 94775
rect 25758 94721 25760 94773
rect 25760 94721 25812 94773
rect 25812 94721 25814 94773
rect 25758 94719 25814 94721
rect 25882 94773 25938 94775
rect 25882 94721 25884 94773
rect 25884 94721 25936 94773
rect 25936 94721 25938 94773
rect 25882 94719 25938 94721
rect 25386 94649 25442 94651
rect 25386 94597 25388 94649
rect 25388 94597 25440 94649
rect 25440 94597 25442 94649
rect 25386 94595 25442 94597
rect 25510 94649 25566 94651
rect 25510 94597 25512 94649
rect 25512 94597 25564 94649
rect 25564 94597 25566 94649
rect 25510 94595 25566 94597
rect 25634 94649 25690 94651
rect 25634 94597 25636 94649
rect 25636 94597 25688 94649
rect 25688 94597 25690 94649
rect 25634 94595 25690 94597
rect 25758 94649 25814 94651
rect 25758 94597 25760 94649
rect 25760 94597 25812 94649
rect 25812 94597 25814 94649
rect 25758 94595 25814 94597
rect 25882 94649 25938 94651
rect 25882 94597 25884 94649
rect 25884 94597 25936 94649
rect 25936 94597 25938 94649
rect 25882 94595 25938 94597
rect 25386 94525 25442 94527
rect 25386 94473 25388 94525
rect 25388 94473 25440 94525
rect 25440 94473 25442 94525
rect 25386 94471 25442 94473
rect 25510 94525 25566 94527
rect 25510 94473 25512 94525
rect 25512 94473 25564 94525
rect 25564 94473 25566 94525
rect 25510 94471 25566 94473
rect 25634 94525 25690 94527
rect 25634 94473 25636 94525
rect 25636 94473 25688 94525
rect 25688 94473 25690 94525
rect 25634 94471 25690 94473
rect 25758 94525 25814 94527
rect 25758 94473 25760 94525
rect 25760 94473 25812 94525
rect 25812 94473 25814 94525
rect 25758 94471 25814 94473
rect 25882 94525 25938 94527
rect 25882 94473 25884 94525
rect 25884 94473 25936 94525
rect 25936 94473 25938 94525
rect 25882 94471 25938 94473
rect 25386 34990 25442 34992
rect 25386 34938 25388 34990
rect 25388 34938 25440 34990
rect 25440 34938 25442 34990
rect 25386 34936 25442 34938
rect 25510 34990 25566 34992
rect 25510 34938 25512 34990
rect 25512 34938 25564 34990
rect 25564 34938 25566 34990
rect 25510 34936 25566 34938
rect 25634 34990 25690 34992
rect 25634 34938 25636 34990
rect 25636 34938 25688 34990
rect 25688 34938 25690 34990
rect 25634 34936 25690 34938
rect 25758 34990 25814 34992
rect 25758 34938 25760 34990
rect 25760 34938 25812 34990
rect 25812 34938 25814 34990
rect 25758 34936 25814 34938
rect 25882 34990 25938 34992
rect 25882 34938 25884 34990
rect 25884 34938 25936 34990
rect 25936 34938 25938 34990
rect 25882 34936 25938 34938
rect 25386 34866 25442 34868
rect 25386 34814 25388 34866
rect 25388 34814 25440 34866
rect 25440 34814 25442 34866
rect 25386 34812 25442 34814
rect 25510 34866 25566 34868
rect 25510 34814 25512 34866
rect 25512 34814 25564 34866
rect 25564 34814 25566 34866
rect 25510 34812 25566 34814
rect 25634 34866 25690 34868
rect 25634 34814 25636 34866
rect 25636 34814 25688 34866
rect 25688 34814 25690 34866
rect 25634 34812 25690 34814
rect 25758 34866 25814 34868
rect 25758 34814 25760 34866
rect 25760 34814 25812 34866
rect 25812 34814 25814 34866
rect 25758 34812 25814 34814
rect 25882 34866 25938 34868
rect 25882 34814 25884 34866
rect 25884 34814 25936 34866
rect 25936 34814 25938 34866
rect 25882 34812 25938 34814
rect 25386 34742 25442 34744
rect 25386 34690 25388 34742
rect 25388 34690 25440 34742
rect 25440 34690 25442 34742
rect 25386 34688 25442 34690
rect 25510 34742 25566 34744
rect 25510 34690 25512 34742
rect 25512 34690 25564 34742
rect 25564 34690 25566 34742
rect 25510 34688 25566 34690
rect 25634 34742 25690 34744
rect 25634 34690 25636 34742
rect 25636 34690 25688 34742
rect 25688 34690 25690 34742
rect 25634 34688 25690 34690
rect 25758 34742 25814 34744
rect 25758 34690 25760 34742
rect 25760 34690 25812 34742
rect 25812 34690 25814 34742
rect 25758 34688 25814 34690
rect 25882 34742 25938 34744
rect 25882 34690 25884 34742
rect 25884 34690 25936 34742
rect 25936 34690 25938 34742
rect 25882 34688 25938 34690
rect 25386 34618 25442 34620
rect 25386 34566 25388 34618
rect 25388 34566 25440 34618
rect 25440 34566 25442 34618
rect 25386 34564 25442 34566
rect 25510 34618 25566 34620
rect 25510 34566 25512 34618
rect 25512 34566 25564 34618
rect 25564 34566 25566 34618
rect 25510 34564 25566 34566
rect 25634 34618 25690 34620
rect 25634 34566 25636 34618
rect 25636 34566 25688 34618
rect 25688 34566 25690 34618
rect 25634 34564 25690 34566
rect 25758 34618 25814 34620
rect 25758 34566 25760 34618
rect 25760 34566 25812 34618
rect 25812 34566 25814 34618
rect 25758 34564 25814 34566
rect 25882 34618 25938 34620
rect 25882 34566 25884 34618
rect 25884 34566 25936 34618
rect 25936 34566 25938 34618
rect 25882 34564 25938 34566
rect 25398 31192 25454 31248
rect 25522 31192 25578 31248
rect 25646 31192 25702 31248
rect 25770 31192 25826 31248
rect 25894 31192 25950 31248
rect 25398 31068 25454 31124
rect 25522 31068 25578 31124
rect 25646 31068 25702 31124
rect 25770 31068 25826 31124
rect 25894 31068 25950 31124
rect 25398 30944 25454 31000
rect 25522 30944 25578 31000
rect 25646 30944 25702 31000
rect 25770 30944 25826 31000
rect 25894 30944 25950 31000
rect 25398 30737 25454 30793
rect 25522 30737 25578 30793
rect 25646 30737 25702 30793
rect 25770 30737 25826 30793
rect 25894 30737 25950 30793
rect 25398 30613 25454 30669
rect 25522 30613 25578 30669
rect 25646 30613 25702 30669
rect 25770 30613 25826 30669
rect 25894 30613 25950 30669
rect 25398 30489 25454 30545
rect 25522 30489 25578 30545
rect 25646 30489 25702 30545
rect 25770 30489 25826 30545
rect 25894 30489 25950 30545
rect 25404 28261 25460 28317
rect 25528 28261 25584 28317
rect 25652 28261 25708 28317
rect 25776 28261 25832 28317
rect 25900 28261 25956 28317
rect 25404 28137 25460 28193
rect 25528 28137 25584 28193
rect 25652 28137 25708 28193
rect 25776 28137 25832 28193
rect 25900 28137 25956 28193
rect 25404 28013 25460 28069
rect 25528 28013 25584 28069
rect 25652 28013 25708 28069
rect 25776 28013 25832 28069
rect 25900 28013 25956 28069
rect 25404 27889 25460 27945
rect 25528 27889 25584 27945
rect 25652 27889 25708 27945
rect 25776 27889 25832 27945
rect 25900 27889 25956 27945
rect 25404 27765 25460 27821
rect 25528 27765 25584 27821
rect 25652 27765 25708 27821
rect 25776 27765 25832 27821
rect 25900 27765 25956 27821
rect 25404 27641 25460 27697
rect 25528 27641 25584 27697
rect 25652 27641 25708 27697
rect 25776 27641 25832 27697
rect 25900 27641 25956 27697
rect 25404 27517 25460 27573
rect 25528 27517 25584 27573
rect 25652 27517 25708 27573
rect 25776 27517 25832 27573
rect 25900 27517 25956 27573
rect 25404 27393 25460 27449
rect 25528 27393 25584 27449
rect 25652 27393 25708 27449
rect 25776 27393 25832 27449
rect 25900 27393 25956 27449
rect 27788 94653 27844 94655
rect 27788 94601 27790 94653
rect 27790 94601 27842 94653
rect 27842 94601 27844 94653
rect 27788 94599 27844 94601
rect 27999 94653 28055 94655
rect 27999 94601 28001 94653
rect 28001 94601 28053 94653
rect 28053 94601 28055 94653
rect 27999 94599 28055 94601
rect 28210 94653 28266 94655
rect 28210 94601 28212 94653
rect 28212 94601 28264 94653
rect 28264 94601 28266 94653
rect 28210 94599 28266 94601
rect 28421 94653 28477 94655
rect 28421 94601 28423 94653
rect 28423 94601 28475 94653
rect 28475 94601 28477 94653
rect 28421 94599 28477 94601
rect 28632 94653 28688 94655
rect 28632 94601 28634 94653
rect 28634 94601 28686 94653
rect 28686 94601 28688 94653
rect 28632 94599 28688 94601
rect 28843 94653 28899 94655
rect 28843 94601 28845 94653
rect 28845 94601 28897 94653
rect 28897 94601 28899 94653
rect 28843 94599 28899 94601
rect 29054 94653 29110 94655
rect 29054 94601 29056 94653
rect 29056 94601 29108 94653
rect 29108 94601 29110 94653
rect 29054 94599 29110 94601
rect 56013 94653 56069 94655
rect 56013 94601 56015 94653
rect 56015 94601 56067 94653
rect 56067 94601 56069 94653
rect 56013 94599 56069 94601
rect 56224 94653 56280 94655
rect 56224 94601 56226 94653
rect 56226 94601 56278 94653
rect 56278 94601 56280 94653
rect 56224 94599 56280 94601
rect 56435 94653 56491 94655
rect 56435 94601 56437 94653
rect 56437 94601 56489 94653
rect 56489 94601 56491 94653
rect 56435 94599 56491 94601
rect 56646 94653 56702 94655
rect 56646 94601 56648 94653
rect 56648 94601 56700 94653
rect 56700 94601 56702 94653
rect 56646 94599 56702 94601
rect 56857 94653 56913 94655
rect 56857 94601 56859 94653
rect 56859 94601 56911 94653
rect 56911 94601 56913 94653
rect 56857 94599 56913 94601
rect 57068 94653 57124 94655
rect 57068 94601 57070 94653
rect 57070 94601 57122 94653
rect 57122 94601 57124 94653
rect 57068 94599 57124 94601
rect 57279 94653 57335 94655
rect 57279 94601 57281 94653
rect 57281 94601 57333 94653
rect 57333 94601 57335 94653
rect 57279 94599 57335 94601
rect 27788 92853 27844 92855
rect 27788 92801 27790 92853
rect 27790 92801 27842 92853
rect 27842 92801 27844 92853
rect 27788 92799 27844 92801
rect 27999 92853 28055 92855
rect 27999 92801 28001 92853
rect 28001 92801 28053 92853
rect 28053 92801 28055 92853
rect 27999 92799 28055 92801
rect 28210 92853 28266 92855
rect 28210 92801 28212 92853
rect 28212 92801 28264 92853
rect 28264 92801 28266 92853
rect 28210 92799 28266 92801
rect 28421 92853 28477 92855
rect 28421 92801 28423 92853
rect 28423 92801 28475 92853
rect 28475 92801 28477 92853
rect 28421 92799 28477 92801
rect 28632 92853 28688 92855
rect 28632 92801 28634 92853
rect 28634 92801 28686 92853
rect 28686 92801 28688 92853
rect 28632 92799 28688 92801
rect 28843 92853 28899 92855
rect 28843 92801 28845 92853
rect 28845 92801 28897 92853
rect 28897 92801 28899 92853
rect 28843 92799 28899 92801
rect 29054 92853 29110 92855
rect 29054 92801 29056 92853
rect 29056 92801 29108 92853
rect 29108 92801 29110 92853
rect 29054 92799 29110 92801
rect 56013 92853 56069 92855
rect 56013 92801 56015 92853
rect 56015 92801 56067 92853
rect 56067 92801 56069 92853
rect 56013 92799 56069 92801
rect 56224 92853 56280 92855
rect 56224 92801 56226 92853
rect 56226 92801 56278 92853
rect 56278 92801 56280 92853
rect 56224 92799 56280 92801
rect 56435 92853 56491 92855
rect 56435 92801 56437 92853
rect 56437 92801 56489 92853
rect 56489 92801 56491 92853
rect 56435 92799 56491 92801
rect 56646 92853 56702 92855
rect 56646 92801 56648 92853
rect 56648 92801 56700 92853
rect 56700 92801 56702 92853
rect 56646 92799 56702 92801
rect 56857 92853 56913 92855
rect 56857 92801 56859 92853
rect 56859 92801 56911 92853
rect 56911 92801 56913 92853
rect 56857 92799 56913 92801
rect 57068 92853 57124 92855
rect 57068 92801 57070 92853
rect 57070 92801 57122 92853
rect 57122 92801 57124 92853
rect 57068 92799 57124 92801
rect 57279 92853 57335 92855
rect 57279 92801 57281 92853
rect 57281 92801 57333 92853
rect 57333 92801 57335 92853
rect 57279 92799 57335 92801
rect 27788 91053 27844 91055
rect 27788 91001 27790 91053
rect 27790 91001 27842 91053
rect 27842 91001 27844 91053
rect 27788 90999 27844 91001
rect 27999 91053 28055 91055
rect 27999 91001 28001 91053
rect 28001 91001 28053 91053
rect 28053 91001 28055 91053
rect 27999 90999 28055 91001
rect 28210 91053 28266 91055
rect 28210 91001 28212 91053
rect 28212 91001 28264 91053
rect 28264 91001 28266 91053
rect 28210 90999 28266 91001
rect 28421 91053 28477 91055
rect 28421 91001 28423 91053
rect 28423 91001 28475 91053
rect 28475 91001 28477 91053
rect 28421 90999 28477 91001
rect 28632 91053 28688 91055
rect 28632 91001 28634 91053
rect 28634 91001 28686 91053
rect 28686 91001 28688 91053
rect 28632 90999 28688 91001
rect 28843 91053 28899 91055
rect 28843 91001 28845 91053
rect 28845 91001 28897 91053
rect 28897 91001 28899 91053
rect 28843 90999 28899 91001
rect 29054 91053 29110 91055
rect 29054 91001 29056 91053
rect 29056 91001 29108 91053
rect 29108 91001 29110 91053
rect 29054 90999 29110 91001
rect 56013 91053 56069 91055
rect 56013 91001 56015 91053
rect 56015 91001 56067 91053
rect 56067 91001 56069 91053
rect 56013 90999 56069 91001
rect 56224 91053 56280 91055
rect 56224 91001 56226 91053
rect 56226 91001 56278 91053
rect 56278 91001 56280 91053
rect 56224 90999 56280 91001
rect 56435 91053 56491 91055
rect 56435 91001 56437 91053
rect 56437 91001 56489 91053
rect 56489 91001 56491 91053
rect 56435 90999 56491 91001
rect 56646 91053 56702 91055
rect 56646 91001 56648 91053
rect 56648 91001 56700 91053
rect 56700 91001 56702 91053
rect 56646 90999 56702 91001
rect 56857 91053 56913 91055
rect 56857 91001 56859 91053
rect 56859 91001 56911 91053
rect 56911 91001 56913 91053
rect 56857 90999 56913 91001
rect 57068 91053 57124 91055
rect 57068 91001 57070 91053
rect 57070 91001 57122 91053
rect 57122 91001 57124 91053
rect 57068 90999 57124 91001
rect 57279 91053 57335 91055
rect 57279 91001 57281 91053
rect 57281 91001 57333 91053
rect 57333 91001 57335 91053
rect 57279 90999 57335 91001
rect 27788 89253 27844 89255
rect 27788 89201 27790 89253
rect 27790 89201 27842 89253
rect 27842 89201 27844 89253
rect 27788 89199 27844 89201
rect 27999 89253 28055 89255
rect 27999 89201 28001 89253
rect 28001 89201 28053 89253
rect 28053 89201 28055 89253
rect 27999 89199 28055 89201
rect 28210 89253 28266 89255
rect 28210 89201 28212 89253
rect 28212 89201 28264 89253
rect 28264 89201 28266 89253
rect 28210 89199 28266 89201
rect 28421 89253 28477 89255
rect 28421 89201 28423 89253
rect 28423 89201 28475 89253
rect 28475 89201 28477 89253
rect 28421 89199 28477 89201
rect 28632 89253 28688 89255
rect 28632 89201 28634 89253
rect 28634 89201 28686 89253
rect 28686 89201 28688 89253
rect 28632 89199 28688 89201
rect 28843 89253 28899 89255
rect 28843 89201 28845 89253
rect 28845 89201 28897 89253
rect 28897 89201 28899 89253
rect 28843 89199 28899 89201
rect 29054 89253 29110 89255
rect 29054 89201 29056 89253
rect 29056 89201 29108 89253
rect 29108 89201 29110 89253
rect 29054 89199 29110 89201
rect 56013 89253 56069 89255
rect 56013 89201 56015 89253
rect 56015 89201 56067 89253
rect 56067 89201 56069 89253
rect 56013 89199 56069 89201
rect 56224 89253 56280 89255
rect 56224 89201 56226 89253
rect 56226 89201 56278 89253
rect 56278 89201 56280 89253
rect 56224 89199 56280 89201
rect 56435 89253 56491 89255
rect 56435 89201 56437 89253
rect 56437 89201 56489 89253
rect 56489 89201 56491 89253
rect 56435 89199 56491 89201
rect 56646 89253 56702 89255
rect 56646 89201 56648 89253
rect 56648 89201 56700 89253
rect 56700 89201 56702 89253
rect 56646 89199 56702 89201
rect 56857 89253 56913 89255
rect 56857 89201 56859 89253
rect 56859 89201 56911 89253
rect 56911 89201 56913 89253
rect 56857 89199 56913 89201
rect 57068 89253 57124 89255
rect 57068 89201 57070 89253
rect 57070 89201 57122 89253
rect 57122 89201 57124 89253
rect 57068 89199 57124 89201
rect 57279 89253 57335 89255
rect 57279 89201 57281 89253
rect 57281 89201 57333 89253
rect 57333 89201 57335 89253
rect 57279 89199 57335 89201
rect 27788 87453 27844 87455
rect 27788 87401 27790 87453
rect 27790 87401 27842 87453
rect 27842 87401 27844 87453
rect 27788 87399 27844 87401
rect 27999 87453 28055 87455
rect 27999 87401 28001 87453
rect 28001 87401 28053 87453
rect 28053 87401 28055 87453
rect 27999 87399 28055 87401
rect 28210 87453 28266 87455
rect 28210 87401 28212 87453
rect 28212 87401 28264 87453
rect 28264 87401 28266 87453
rect 28210 87399 28266 87401
rect 28421 87453 28477 87455
rect 28421 87401 28423 87453
rect 28423 87401 28475 87453
rect 28475 87401 28477 87453
rect 28421 87399 28477 87401
rect 28632 87453 28688 87455
rect 28632 87401 28634 87453
rect 28634 87401 28686 87453
rect 28686 87401 28688 87453
rect 28632 87399 28688 87401
rect 28843 87453 28899 87455
rect 28843 87401 28845 87453
rect 28845 87401 28897 87453
rect 28897 87401 28899 87453
rect 28843 87399 28899 87401
rect 29054 87453 29110 87455
rect 29054 87401 29056 87453
rect 29056 87401 29108 87453
rect 29108 87401 29110 87453
rect 29054 87399 29110 87401
rect 56013 87453 56069 87455
rect 56013 87401 56015 87453
rect 56015 87401 56067 87453
rect 56067 87401 56069 87453
rect 56013 87399 56069 87401
rect 56224 87453 56280 87455
rect 56224 87401 56226 87453
rect 56226 87401 56278 87453
rect 56278 87401 56280 87453
rect 56224 87399 56280 87401
rect 56435 87453 56491 87455
rect 56435 87401 56437 87453
rect 56437 87401 56489 87453
rect 56489 87401 56491 87453
rect 56435 87399 56491 87401
rect 56646 87453 56702 87455
rect 56646 87401 56648 87453
rect 56648 87401 56700 87453
rect 56700 87401 56702 87453
rect 56646 87399 56702 87401
rect 56857 87453 56913 87455
rect 56857 87401 56859 87453
rect 56859 87401 56911 87453
rect 56911 87401 56913 87453
rect 56857 87399 56913 87401
rect 57068 87453 57124 87455
rect 57068 87401 57070 87453
rect 57070 87401 57122 87453
rect 57122 87401 57124 87453
rect 57068 87399 57124 87401
rect 57279 87453 57335 87455
rect 57279 87401 57281 87453
rect 57281 87401 57333 87453
rect 57333 87401 57335 87453
rect 57279 87399 57335 87401
rect 27788 85653 27844 85655
rect 27788 85601 27790 85653
rect 27790 85601 27842 85653
rect 27842 85601 27844 85653
rect 27788 85599 27844 85601
rect 27999 85653 28055 85655
rect 27999 85601 28001 85653
rect 28001 85601 28053 85653
rect 28053 85601 28055 85653
rect 27999 85599 28055 85601
rect 28210 85653 28266 85655
rect 28210 85601 28212 85653
rect 28212 85601 28264 85653
rect 28264 85601 28266 85653
rect 28210 85599 28266 85601
rect 28421 85653 28477 85655
rect 28421 85601 28423 85653
rect 28423 85601 28475 85653
rect 28475 85601 28477 85653
rect 28421 85599 28477 85601
rect 28632 85653 28688 85655
rect 28632 85601 28634 85653
rect 28634 85601 28686 85653
rect 28686 85601 28688 85653
rect 28632 85599 28688 85601
rect 28843 85653 28899 85655
rect 28843 85601 28845 85653
rect 28845 85601 28897 85653
rect 28897 85601 28899 85653
rect 28843 85599 28899 85601
rect 29054 85653 29110 85655
rect 29054 85601 29056 85653
rect 29056 85601 29108 85653
rect 29108 85601 29110 85653
rect 29054 85599 29110 85601
rect 56013 85653 56069 85655
rect 56013 85601 56015 85653
rect 56015 85601 56067 85653
rect 56067 85601 56069 85653
rect 56013 85599 56069 85601
rect 56224 85653 56280 85655
rect 56224 85601 56226 85653
rect 56226 85601 56278 85653
rect 56278 85601 56280 85653
rect 56224 85599 56280 85601
rect 56435 85653 56491 85655
rect 56435 85601 56437 85653
rect 56437 85601 56489 85653
rect 56489 85601 56491 85653
rect 56435 85599 56491 85601
rect 56646 85653 56702 85655
rect 56646 85601 56648 85653
rect 56648 85601 56700 85653
rect 56700 85601 56702 85653
rect 56646 85599 56702 85601
rect 56857 85653 56913 85655
rect 56857 85601 56859 85653
rect 56859 85601 56911 85653
rect 56911 85601 56913 85653
rect 56857 85599 56913 85601
rect 57068 85653 57124 85655
rect 57068 85601 57070 85653
rect 57070 85601 57122 85653
rect 57122 85601 57124 85653
rect 57068 85599 57124 85601
rect 57279 85653 57335 85655
rect 57279 85601 57281 85653
rect 57281 85601 57333 85653
rect 57333 85601 57335 85653
rect 57279 85599 57335 85601
rect 27788 83853 27844 83855
rect 27788 83801 27790 83853
rect 27790 83801 27842 83853
rect 27842 83801 27844 83853
rect 27788 83799 27844 83801
rect 27999 83853 28055 83855
rect 27999 83801 28001 83853
rect 28001 83801 28053 83853
rect 28053 83801 28055 83853
rect 27999 83799 28055 83801
rect 28210 83853 28266 83855
rect 28210 83801 28212 83853
rect 28212 83801 28264 83853
rect 28264 83801 28266 83853
rect 28210 83799 28266 83801
rect 28421 83853 28477 83855
rect 28421 83801 28423 83853
rect 28423 83801 28475 83853
rect 28475 83801 28477 83853
rect 28421 83799 28477 83801
rect 28632 83853 28688 83855
rect 28632 83801 28634 83853
rect 28634 83801 28686 83853
rect 28686 83801 28688 83853
rect 28632 83799 28688 83801
rect 28843 83853 28899 83855
rect 28843 83801 28845 83853
rect 28845 83801 28897 83853
rect 28897 83801 28899 83853
rect 28843 83799 28899 83801
rect 29054 83853 29110 83855
rect 29054 83801 29056 83853
rect 29056 83801 29108 83853
rect 29108 83801 29110 83853
rect 29054 83799 29110 83801
rect 56013 83853 56069 83855
rect 56013 83801 56015 83853
rect 56015 83801 56067 83853
rect 56067 83801 56069 83853
rect 56013 83799 56069 83801
rect 56224 83853 56280 83855
rect 56224 83801 56226 83853
rect 56226 83801 56278 83853
rect 56278 83801 56280 83853
rect 56224 83799 56280 83801
rect 56435 83853 56491 83855
rect 56435 83801 56437 83853
rect 56437 83801 56489 83853
rect 56489 83801 56491 83853
rect 56435 83799 56491 83801
rect 56646 83853 56702 83855
rect 56646 83801 56648 83853
rect 56648 83801 56700 83853
rect 56700 83801 56702 83853
rect 56646 83799 56702 83801
rect 56857 83853 56913 83855
rect 56857 83801 56859 83853
rect 56859 83801 56911 83853
rect 56911 83801 56913 83853
rect 56857 83799 56913 83801
rect 57068 83853 57124 83855
rect 57068 83801 57070 83853
rect 57070 83801 57122 83853
rect 57122 83801 57124 83853
rect 57068 83799 57124 83801
rect 57279 83853 57335 83855
rect 57279 83801 57281 83853
rect 57281 83801 57333 83853
rect 57333 83801 57335 83853
rect 57279 83799 57335 83801
rect 27788 82053 27844 82055
rect 27788 82001 27790 82053
rect 27790 82001 27842 82053
rect 27842 82001 27844 82053
rect 27788 81999 27844 82001
rect 27999 82053 28055 82055
rect 27999 82001 28001 82053
rect 28001 82001 28053 82053
rect 28053 82001 28055 82053
rect 27999 81999 28055 82001
rect 28210 82053 28266 82055
rect 28210 82001 28212 82053
rect 28212 82001 28264 82053
rect 28264 82001 28266 82053
rect 28210 81999 28266 82001
rect 28421 82053 28477 82055
rect 28421 82001 28423 82053
rect 28423 82001 28475 82053
rect 28475 82001 28477 82053
rect 28421 81999 28477 82001
rect 28632 82053 28688 82055
rect 28632 82001 28634 82053
rect 28634 82001 28686 82053
rect 28686 82001 28688 82053
rect 28632 81999 28688 82001
rect 28843 82053 28899 82055
rect 28843 82001 28845 82053
rect 28845 82001 28897 82053
rect 28897 82001 28899 82053
rect 28843 81999 28899 82001
rect 29054 82053 29110 82055
rect 29054 82001 29056 82053
rect 29056 82001 29108 82053
rect 29108 82001 29110 82053
rect 29054 81999 29110 82001
rect 56013 82053 56069 82055
rect 56013 82001 56015 82053
rect 56015 82001 56067 82053
rect 56067 82001 56069 82053
rect 56013 81999 56069 82001
rect 56224 82053 56280 82055
rect 56224 82001 56226 82053
rect 56226 82001 56278 82053
rect 56278 82001 56280 82053
rect 56224 81999 56280 82001
rect 56435 82053 56491 82055
rect 56435 82001 56437 82053
rect 56437 82001 56489 82053
rect 56489 82001 56491 82053
rect 56435 81999 56491 82001
rect 56646 82053 56702 82055
rect 56646 82001 56648 82053
rect 56648 82001 56700 82053
rect 56700 82001 56702 82053
rect 56646 81999 56702 82001
rect 56857 82053 56913 82055
rect 56857 82001 56859 82053
rect 56859 82001 56911 82053
rect 56911 82001 56913 82053
rect 56857 81999 56913 82001
rect 57068 82053 57124 82055
rect 57068 82001 57070 82053
rect 57070 82001 57122 82053
rect 57122 82001 57124 82053
rect 57068 81999 57124 82001
rect 57279 82053 57335 82055
rect 57279 82001 57281 82053
rect 57281 82001 57333 82053
rect 57333 82001 57335 82053
rect 57279 81999 57335 82001
rect 27788 80253 27844 80255
rect 27788 80201 27790 80253
rect 27790 80201 27842 80253
rect 27842 80201 27844 80253
rect 27788 80199 27844 80201
rect 27999 80253 28055 80255
rect 27999 80201 28001 80253
rect 28001 80201 28053 80253
rect 28053 80201 28055 80253
rect 27999 80199 28055 80201
rect 28210 80253 28266 80255
rect 28210 80201 28212 80253
rect 28212 80201 28264 80253
rect 28264 80201 28266 80253
rect 28210 80199 28266 80201
rect 28421 80253 28477 80255
rect 28421 80201 28423 80253
rect 28423 80201 28475 80253
rect 28475 80201 28477 80253
rect 28421 80199 28477 80201
rect 28632 80253 28688 80255
rect 28632 80201 28634 80253
rect 28634 80201 28686 80253
rect 28686 80201 28688 80253
rect 28632 80199 28688 80201
rect 28843 80253 28899 80255
rect 28843 80201 28845 80253
rect 28845 80201 28897 80253
rect 28897 80201 28899 80253
rect 28843 80199 28899 80201
rect 29054 80253 29110 80255
rect 29054 80201 29056 80253
rect 29056 80201 29108 80253
rect 29108 80201 29110 80253
rect 29054 80199 29110 80201
rect 56013 80253 56069 80255
rect 56013 80201 56015 80253
rect 56015 80201 56067 80253
rect 56067 80201 56069 80253
rect 56013 80199 56069 80201
rect 56224 80253 56280 80255
rect 56224 80201 56226 80253
rect 56226 80201 56278 80253
rect 56278 80201 56280 80253
rect 56224 80199 56280 80201
rect 56435 80253 56491 80255
rect 56435 80201 56437 80253
rect 56437 80201 56489 80253
rect 56489 80201 56491 80253
rect 56435 80199 56491 80201
rect 56646 80253 56702 80255
rect 56646 80201 56648 80253
rect 56648 80201 56700 80253
rect 56700 80201 56702 80253
rect 56646 80199 56702 80201
rect 56857 80253 56913 80255
rect 56857 80201 56859 80253
rect 56859 80201 56911 80253
rect 56911 80201 56913 80253
rect 56857 80199 56913 80201
rect 57068 80253 57124 80255
rect 57068 80201 57070 80253
rect 57070 80201 57122 80253
rect 57122 80201 57124 80253
rect 57068 80199 57124 80201
rect 57279 80253 57335 80255
rect 57279 80201 57281 80253
rect 57281 80201 57333 80253
rect 57333 80201 57335 80253
rect 57279 80199 57335 80201
rect 27788 78453 27844 78455
rect 27788 78401 27790 78453
rect 27790 78401 27842 78453
rect 27842 78401 27844 78453
rect 27788 78399 27844 78401
rect 27999 78453 28055 78455
rect 27999 78401 28001 78453
rect 28001 78401 28053 78453
rect 28053 78401 28055 78453
rect 27999 78399 28055 78401
rect 28210 78453 28266 78455
rect 28210 78401 28212 78453
rect 28212 78401 28264 78453
rect 28264 78401 28266 78453
rect 28210 78399 28266 78401
rect 28421 78453 28477 78455
rect 28421 78401 28423 78453
rect 28423 78401 28475 78453
rect 28475 78401 28477 78453
rect 28421 78399 28477 78401
rect 28632 78453 28688 78455
rect 28632 78401 28634 78453
rect 28634 78401 28686 78453
rect 28686 78401 28688 78453
rect 28632 78399 28688 78401
rect 28843 78453 28899 78455
rect 28843 78401 28845 78453
rect 28845 78401 28897 78453
rect 28897 78401 28899 78453
rect 28843 78399 28899 78401
rect 29054 78453 29110 78455
rect 29054 78401 29056 78453
rect 29056 78401 29108 78453
rect 29108 78401 29110 78453
rect 29054 78399 29110 78401
rect 56013 78453 56069 78455
rect 56013 78401 56015 78453
rect 56015 78401 56067 78453
rect 56067 78401 56069 78453
rect 56013 78399 56069 78401
rect 56224 78453 56280 78455
rect 56224 78401 56226 78453
rect 56226 78401 56278 78453
rect 56278 78401 56280 78453
rect 56224 78399 56280 78401
rect 56435 78453 56491 78455
rect 56435 78401 56437 78453
rect 56437 78401 56489 78453
rect 56489 78401 56491 78453
rect 56435 78399 56491 78401
rect 56646 78453 56702 78455
rect 56646 78401 56648 78453
rect 56648 78401 56700 78453
rect 56700 78401 56702 78453
rect 56646 78399 56702 78401
rect 56857 78453 56913 78455
rect 56857 78401 56859 78453
rect 56859 78401 56911 78453
rect 56911 78401 56913 78453
rect 56857 78399 56913 78401
rect 57068 78453 57124 78455
rect 57068 78401 57070 78453
rect 57070 78401 57122 78453
rect 57122 78401 57124 78453
rect 57068 78399 57124 78401
rect 57279 78453 57335 78455
rect 57279 78401 57281 78453
rect 57281 78401 57333 78453
rect 57333 78401 57335 78453
rect 57279 78399 57335 78401
rect 27788 76653 27844 76655
rect 27788 76601 27790 76653
rect 27790 76601 27842 76653
rect 27842 76601 27844 76653
rect 27788 76599 27844 76601
rect 27999 76653 28055 76655
rect 27999 76601 28001 76653
rect 28001 76601 28053 76653
rect 28053 76601 28055 76653
rect 27999 76599 28055 76601
rect 28210 76653 28266 76655
rect 28210 76601 28212 76653
rect 28212 76601 28264 76653
rect 28264 76601 28266 76653
rect 28210 76599 28266 76601
rect 28421 76653 28477 76655
rect 28421 76601 28423 76653
rect 28423 76601 28475 76653
rect 28475 76601 28477 76653
rect 28421 76599 28477 76601
rect 28632 76653 28688 76655
rect 28632 76601 28634 76653
rect 28634 76601 28686 76653
rect 28686 76601 28688 76653
rect 28632 76599 28688 76601
rect 28843 76653 28899 76655
rect 28843 76601 28845 76653
rect 28845 76601 28897 76653
rect 28897 76601 28899 76653
rect 28843 76599 28899 76601
rect 29054 76653 29110 76655
rect 29054 76601 29056 76653
rect 29056 76601 29108 76653
rect 29108 76601 29110 76653
rect 29054 76599 29110 76601
rect 56013 76653 56069 76655
rect 56013 76601 56015 76653
rect 56015 76601 56067 76653
rect 56067 76601 56069 76653
rect 56013 76599 56069 76601
rect 56224 76653 56280 76655
rect 56224 76601 56226 76653
rect 56226 76601 56278 76653
rect 56278 76601 56280 76653
rect 56224 76599 56280 76601
rect 56435 76653 56491 76655
rect 56435 76601 56437 76653
rect 56437 76601 56489 76653
rect 56489 76601 56491 76653
rect 56435 76599 56491 76601
rect 56646 76653 56702 76655
rect 56646 76601 56648 76653
rect 56648 76601 56700 76653
rect 56700 76601 56702 76653
rect 56646 76599 56702 76601
rect 56857 76653 56913 76655
rect 56857 76601 56859 76653
rect 56859 76601 56911 76653
rect 56911 76601 56913 76653
rect 56857 76599 56913 76601
rect 57068 76653 57124 76655
rect 57068 76601 57070 76653
rect 57070 76601 57122 76653
rect 57122 76601 57124 76653
rect 57068 76599 57124 76601
rect 57279 76653 57335 76655
rect 57279 76601 57281 76653
rect 57281 76601 57333 76653
rect 57333 76601 57335 76653
rect 57279 76599 57335 76601
rect 27788 74853 27844 74855
rect 27788 74801 27790 74853
rect 27790 74801 27842 74853
rect 27842 74801 27844 74853
rect 27788 74799 27844 74801
rect 27999 74853 28055 74855
rect 27999 74801 28001 74853
rect 28001 74801 28053 74853
rect 28053 74801 28055 74853
rect 27999 74799 28055 74801
rect 28210 74853 28266 74855
rect 28210 74801 28212 74853
rect 28212 74801 28264 74853
rect 28264 74801 28266 74853
rect 28210 74799 28266 74801
rect 28421 74853 28477 74855
rect 28421 74801 28423 74853
rect 28423 74801 28475 74853
rect 28475 74801 28477 74853
rect 28421 74799 28477 74801
rect 28632 74853 28688 74855
rect 28632 74801 28634 74853
rect 28634 74801 28686 74853
rect 28686 74801 28688 74853
rect 28632 74799 28688 74801
rect 28843 74853 28899 74855
rect 28843 74801 28845 74853
rect 28845 74801 28897 74853
rect 28897 74801 28899 74853
rect 28843 74799 28899 74801
rect 29054 74853 29110 74855
rect 29054 74801 29056 74853
rect 29056 74801 29108 74853
rect 29108 74801 29110 74853
rect 29054 74799 29110 74801
rect 56013 74853 56069 74855
rect 56013 74801 56015 74853
rect 56015 74801 56067 74853
rect 56067 74801 56069 74853
rect 56013 74799 56069 74801
rect 56224 74853 56280 74855
rect 56224 74801 56226 74853
rect 56226 74801 56278 74853
rect 56278 74801 56280 74853
rect 56224 74799 56280 74801
rect 56435 74853 56491 74855
rect 56435 74801 56437 74853
rect 56437 74801 56489 74853
rect 56489 74801 56491 74853
rect 56435 74799 56491 74801
rect 56646 74853 56702 74855
rect 56646 74801 56648 74853
rect 56648 74801 56700 74853
rect 56700 74801 56702 74853
rect 56646 74799 56702 74801
rect 56857 74853 56913 74855
rect 56857 74801 56859 74853
rect 56859 74801 56911 74853
rect 56911 74801 56913 74853
rect 56857 74799 56913 74801
rect 57068 74853 57124 74855
rect 57068 74801 57070 74853
rect 57070 74801 57122 74853
rect 57122 74801 57124 74853
rect 57068 74799 57124 74801
rect 57279 74853 57335 74855
rect 57279 74801 57281 74853
rect 57281 74801 57333 74853
rect 57333 74801 57335 74853
rect 57279 74799 57335 74801
rect 27788 73053 27844 73055
rect 27788 73001 27790 73053
rect 27790 73001 27842 73053
rect 27842 73001 27844 73053
rect 27788 72999 27844 73001
rect 27999 73053 28055 73055
rect 27999 73001 28001 73053
rect 28001 73001 28053 73053
rect 28053 73001 28055 73053
rect 27999 72999 28055 73001
rect 28210 73053 28266 73055
rect 28210 73001 28212 73053
rect 28212 73001 28264 73053
rect 28264 73001 28266 73053
rect 28210 72999 28266 73001
rect 28421 73053 28477 73055
rect 28421 73001 28423 73053
rect 28423 73001 28475 73053
rect 28475 73001 28477 73053
rect 28421 72999 28477 73001
rect 28632 73053 28688 73055
rect 28632 73001 28634 73053
rect 28634 73001 28686 73053
rect 28686 73001 28688 73053
rect 28632 72999 28688 73001
rect 28843 73053 28899 73055
rect 28843 73001 28845 73053
rect 28845 73001 28897 73053
rect 28897 73001 28899 73053
rect 28843 72999 28899 73001
rect 29054 73053 29110 73055
rect 29054 73001 29056 73053
rect 29056 73001 29108 73053
rect 29108 73001 29110 73053
rect 29054 72999 29110 73001
rect 56013 73053 56069 73055
rect 56013 73001 56015 73053
rect 56015 73001 56067 73053
rect 56067 73001 56069 73053
rect 56013 72999 56069 73001
rect 56224 73053 56280 73055
rect 56224 73001 56226 73053
rect 56226 73001 56278 73053
rect 56278 73001 56280 73053
rect 56224 72999 56280 73001
rect 56435 73053 56491 73055
rect 56435 73001 56437 73053
rect 56437 73001 56489 73053
rect 56489 73001 56491 73053
rect 56435 72999 56491 73001
rect 56646 73053 56702 73055
rect 56646 73001 56648 73053
rect 56648 73001 56700 73053
rect 56700 73001 56702 73053
rect 56646 72999 56702 73001
rect 56857 73053 56913 73055
rect 56857 73001 56859 73053
rect 56859 73001 56911 73053
rect 56911 73001 56913 73053
rect 56857 72999 56913 73001
rect 57068 73053 57124 73055
rect 57068 73001 57070 73053
rect 57070 73001 57122 73053
rect 57122 73001 57124 73053
rect 57068 72999 57124 73001
rect 57279 73053 57335 73055
rect 57279 73001 57281 73053
rect 57281 73001 57333 73053
rect 57333 73001 57335 73053
rect 57279 72999 57335 73001
rect 27788 71253 27844 71255
rect 27788 71201 27790 71253
rect 27790 71201 27842 71253
rect 27842 71201 27844 71253
rect 27788 71199 27844 71201
rect 27999 71253 28055 71255
rect 27999 71201 28001 71253
rect 28001 71201 28053 71253
rect 28053 71201 28055 71253
rect 27999 71199 28055 71201
rect 28210 71253 28266 71255
rect 28210 71201 28212 71253
rect 28212 71201 28264 71253
rect 28264 71201 28266 71253
rect 28210 71199 28266 71201
rect 28421 71253 28477 71255
rect 28421 71201 28423 71253
rect 28423 71201 28475 71253
rect 28475 71201 28477 71253
rect 28421 71199 28477 71201
rect 28632 71253 28688 71255
rect 28632 71201 28634 71253
rect 28634 71201 28686 71253
rect 28686 71201 28688 71253
rect 28632 71199 28688 71201
rect 28843 71253 28899 71255
rect 28843 71201 28845 71253
rect 28845 71201 28897 71253
rect 28897 71201 28899 71253
rect 28843 71199 28899 71201
rect 29054 71253 29110 71255
rect 29054 71201 29056 71253
rect 29056 71201 29108 71253
rect 29108 71201 29110 71253
rect 29054 71199 29110 71201
rect 56013 71253 56069 71255
rect 56013 71201 56015 71253
rect 56015 71201 56067 71253
rect 56067 71201 56069 71253
rect 56013 71199 56069 71201
rect 56224 71253 56280 71255
rect 56224 71201 56226 71253
rect 56226 71201 56278 71253
rect 56278 71201 56280 71253
rect 56224 71199 56280 71201
rect 56435 71253 56491 71255
rect 56435 71201 56437 71253
rect 56437 71201 56489 71253
rect 56489 71201 56491 71253
rect 56435 71199 56491 71201
rect 56646 71253 56702 71255
rect 56646 71201 56648 71253
rect 56648 71201 56700 71253
rect 56700 71201 56702 71253
rect 56646 71199 56702 71201
rect 56857 71253 56913 71255
rect 56857 71201 56859 71253
rect 56859 71201 56911 71253
rect 56911 71201 56913 71253
rect 56857 71199 56913 71201
rect 57068 71253 57124 71255
rect 57068 71201 57070 71253
rect 57070 71201 57122 71253
rect 57122 71201 57124 71253
rect 57068 71199 57124 71201
rect 57279 71253 57335 71255
rect 57279 71201 57281 71253
rect 57281 71201 57333 71253
rect 57333 71201 57335 71253
rect 57279 71199 57335 71201
rect 27788 69453 27844 69455
rect 27788 69401 27790 69453
rect 27790 69401 27842 69453
rect 27842 69401 27844 69453
rect 27788 69399 27844 69401
rect 27999 69453 28055 69455
rect 27999 69401 28001 69453
rect 28001 69401 28053 69453
rect 28053 69401 28055 69453
rect 27999 69399 28055 69401
rect 28210 69453 28266 69455
rect 28210 69401 28212 69453
rect 28212 69401 28264 69453
rect 28264 69401 28266 69453
rect 28210 69399 28266 69401
rect 28421 69453 28477 69455
rect 28421 69401 28423 69453
rect 28423 69401 28475 69453
rect 28475 69401 28477 69453
rect 28421 69399 28477 69401
rect 28632 69453 28688 69455
rect 28632 69401 28634 69453
rect 28634 69401 28686 69453
rect 28686 69401 28688 69453
rect 28632 69399 28688 69401
rect 28843 69453 28899 69455
rect 28843 69401 28845 69453
rect 28845 69401 28897 69453
rect 28897 69401 28899 69453
rect 28843 69399 28899 69401
rect 29054 69453 29110 69455
rect 29054 69401 29056 69453
rect 29056 69401 29108 69453
rect 29108 69401 29110 69453
rect 29054 69399 29110 69401
rect 56013 69453 56069 69455
rect 56013 69401 56015 69453
rect 56015 69401 56067 69453
rect 56067 69401 56069 69453
rect 56013 69399 56069 69401
rect 56224 69453 56280 69455
rect 56224 69401 56226 69453
rect 56226 69401 56278 69453
rect 56278 69401 56280 69453
rect 56224 69399 56280 69401
rect 56435 69453 56491 69455
rect 56435 69401 56437 69453
rect 56437 69401 56489 69453
rect 56489 69401 56491 69453
rect 56435 69399 56491 69401
rect 56646 69453 56702 69455
rect 56646 69401 56648 69453
rect 56648 69401 56700 69453
rect 56700 69401 56702 69453
rect 56646 69399 56702 69401
rect 56857 69453 56913 69455
rect 56857 69401 56859 69453
rect 56859 69401 56911 69453
rect 56911 69401 56913 69453
rect 56857 69399 56913 69401
rect 57068 69453 57124 69455
rect 57068 69401 57070 69453
rect 57070 69401 57122 69453
rect 57122 69401 57124 69453
rect 57068 69399 57124 69401
rect 57279 69453 57335 69455
rect 57279 69401 57281 69453
rect 57281 69401 57333 69453
rect 57333 69401 57335 69453
rect 57279 69399 57335 69401
rect 27788 67653 27844 67655
rect 27788 67601 27790 67653
rect 27790 67601 27842 67653
rect 27842 67601 27844 67653
rect 27788 67599 27844 67601
rect 27999 67653 28055 67655
rect 27999 67601 28001 67653
rect 28001 67601 28053 67653
rect 28053 67601 28055 67653
rect 27999 67599 28055 67601
rect 28210 67653 28266 67655
rect 28210 67601 28212 67653
rect 28212 67601 28264 67653
rect 28264 67601 28266 67653
rect 28210 67599 28266 67601
rect 28421 67653 28477 67655
rect 28421 67601 28423 67653
rect 28423 67601 28475 67653
rect 28475 67601 28477 67653
rect 28421 67599 28477 67601
rect 28632 67653 28688 67655
rect 28632 67601 28634 67653
rect 28634 67601 28686 67653
rect 28686 67601 28688 67653
rect 28632 67599 28688 67601
rect 28843 67653 28899 67655
rect 28843 67601 28845 67653
rect 28845 67601 28897 67653
rect 28897 67601 28899 67653
rect 28843 67599 28899 67601
rect 29054 67653 29110 67655
rect 29054 67601 29056 67653
rect 29056 67601 29108 67653
rect 29108 67601 29110 67653
rect 29054 67599 29110 67601
rect 56013 67653 56069 67655
rect 56013 67601 56015 67653
rect 56015 67601 56067 67653
rect 56067 67601 56069 67653
rect 56013 67599 56069 67601
rect 56224 67653 56280 67655
rect 56224 67601 56226 67653
rect 56226 67601 56278 67653
rect 56278 67601 56280 67653
rect 56224 67599 56280 67601
rect 56435 67653 56491 67655
rect 56435 67601 56437 67653
rect 56437 67601 56489 67653
rect 56489 67601 56491 67653
rect 56435 67599 56491 67601
rect 56646 67653 56702 67655
rect 56646 67601 56648 67653
rect 56648 67601 56700 67653
rect 56700 67601 56702 67653
rect 56646 67599 56702 67601
rect 56857 67653 56913 67655
rect 56857 67601 56859 67653
rect 56859 67601 56911 67653
rect 56911 67601 56913 67653
rect 56857 67599 56913 67601
rect 57068 67653 57124 67655
rect 57068 67601 57070 67653
rect 57070 67601 57122 67653
rect 57122 67601 57124 67653
rect 57068 67599 57124 67601
rect 57279 67653 57335 67655
rect 57279 67601 57281 67653
rect 57281 67601 57333 67653
rect 57333 67601 57335 67653
rect 57279 67599 57335 67601
rect 27788 65853 27844 65855
rect 27788 65801 27790 65853
rect 27790 65801 27842 65853
rect 27842 65801 27844 65853
rect 27788 65799 27844 65801
rect 27999 65853 28055 65855
rect 27999 65801 28001 65853
rect 28001 65801 28053 65853
rect 28053 65801 28055 65853
rect 27999 65799 28055 65801
rect 28210 65853 28266 65855
rect 28210 65801 28212 65853
rect 28212 65801 28264 65853
rect 28264 65801 28266 65853
rect 28210 65799 28266 65801
rect 28421 65853 28477 65855
rect 28421 65801 28423 65853
rect 28423 65801 28475 65853
rect 28475 65801 28477 65853
rect 28421 65799 28477 65801
rect 28632 65853 28688 65855
rect 28632 65801 28634 65853
rect 28634 65801 28686 65853
rect 28686 65801 28688 65853
rect 28632 65799 28688 65801
rect 28843 65853 28899 65855
rect 28843 65801 28845 65853
rect 28845 65801 28897 65853
rect 28897 65801 28899 65853
rect 28843 65799 28899 65801
rect 29054 65853 29110 65855
rect 29054 65801 29056 65853
rect 29056 65801 29108 65853
rect 29108 65801 29110 65853
rect 29054 65799 29110 65801
rect 56013 65853 56069 65855
rect 56013 65801 56015 65853
rect 56015 65801 56067 65853
rect 56067 65801 56069 65853
rect 56013 65799 56069 65801
rect 56224 65853 56280 65855
rect 56224 65801 56226 65853
rect 56226 65801 56278 65853
rect 56278 65801 56280 65853
rect 56224 65799 56280 65801
rect 56435 65853 56491 65855
rect 56435 65801 56437 65853
rect 56437 65801 56489 65853
rect 56489 65801 56491 65853
rect 56435 65799 56491 65801
rect 56646 65853 56702 65855
rect 56646 65801 56648 65853
rect 56648 65801 56700 65853
rect 56700 65801 56702 65853
rect 56646 65799 56702 65801
rect 56857 65853 56913 65855
rect 56857 65801 56859 65853
rect 56859 65801 56911 65853
rect 56911 65801 56913 65853
rect 56857 65799 56913 65801
rect 57068 65853 57124 65855
rect 57068 65801 57070 65853
rect 57070 65801 57122 65853
rect 57122 65801 57124 65853
rect 57068 65799 57124 65801
rect 57279 65853 57335 65855
rect 57279 65801 57281 65853
rect 57281 65801 57333 65853
rect 57333 65801 57335 65853
rect 57279 65799 57335 65801
rect 27788 64053 27844 64055
rect 27788 64001 27790 64053
rect 27790 64001 27842 64053
rect 27842 64001 27844 64053
rect 27788 63999 27844 64001
rect 27999 64053 28055 64055
rect 27999 64001 28001 64053
rect 28001 64001 28053 64053
rect 28053 64001 28055 64053
rect 27999 63999 28055 64001
rect 28210 64053 28266 64055
rect 28210 64001 28212 64053
rect 28212 64001 28264 64053
rect 28264 64001 28266 64053
rect 28210 63999 28266 64001
rect 28421 64053 28477 64055
rect 28421 64001 28423 64053
rect 28423 64001 28475 64053
rect 28475 64001 28477 64053
rect 28421 63999 28477 64001
rect 28632 64053 28688 64055
rect 28632 64001 28634 64053
rect 28634 64001 28686 64053
rect 28686 64001 28688 64053
rect 28632 63999 28688 64001
rect 28843 64053 28899 64055
rect 28843 64001 28845 64053
rect 28845 64001 28897 64053
rect 28897 64001 28899 64053
rect 28843 63999 28899 64001
rect 29054 64053 29110 64055
rect 29054 64001 29056 64053
rect 29056 64001 29108 64053
rect 29108 64001 29110 64053
rect 29054 63999 29110 64001
rect 56013 64053 56069 64055
rect 56013 64001 56015 64053
rect 56015 64001 56067 64053
rect 56067 64001 56069 64053
rect 56013 63999 56069 64001
rect 56224 64053 56280 64055
rect 56224 64001 56226 64053
rect 56226 64001 56278 64053
rect 56278 64001 56280 64053
rect 56224 63999 56280 64001
rect 56435 64053 56491 64055
rect 56435 64001 56437 64053
rect 56437 64001 56489 64053
rect 56489 64001 56491 64053
rect 56435 63999 56491 64001
rect 56646 64053 56702 64055
rect 56646 64001 56648 64053
rect 56648 64001 56700 64053
rect 56700 64001 56702 64053
rect 56646 63999 56702 64001
rect 56857 64053 56913 64055
rect 56857 64001 56859 64053
rect 56859 64001 56911 64053
rect 56911 64001 56913 64053
rect 56857 63999 56913 64001
rect 57068 64053 57124 64055
rect 57068 64001 57070 64053
rect 57070 64001 57122 64053
rect 57122 64001 57124 64053
rect 57068 63999 57124 64001
rect 57279 64053 57335 64055
rect 57279 64001 57281 64053
rect 57281 64001 57333 64053
rect 57333 64001 57335 64053
rect 57279 63999 57335 64001
rect 27788 62253 27844 62255
rect 27788 62201 27790 62253
rect 27790 62201 27842 62253
rect 27842 62201 27844 62253
rect 27788 62199 27844 62201
rect 27999 62253 28055 62255
rect 27999 62201 28001 62253
rect 28001 62201 28053 62253
rect 28053 62201 28055 62253
rect 27999 62199 28055 62201
rect 28210 62253 28266 62255
rect 28210 62201 28212 62253
rect 28212 62201 28264 62253
rect 28264 62201 28266 62253
rect 28210 62199 28266 62201
rect 28421 62253 28477 62255
rect 28421 62201 28423 62253
rect 28423 62201 28475 62253
rect 28475 62201 28477 62253
rect 28421 62199 28477 62201
rect 28632 62253 28688 62255
rect 28632 62201 28634 62253
rect 28634 62201 28686 62253
rect 28686 62201 28688 62253
rect 28632 62199 28688 62201
rect 28843 62253 28899 62255
rect 28843 62201 28845 62253
rect 28845 62201 28897 62253
rect 28897 62201 28899 62253
rect 28843 62199 28899 62201
rect 29054 62253 29110 62255
rect 29054 62201 29056 62253
rect 29056 62201 29108 62253
rect 29108 62201 29110 62253
rect 29054 62199 29110 62201
rect 56013 62253 56069 62255
rect 56013 62201 56015 62253
rect 56015 62201 56067 62253
rect 56067 62201 56069 62253
rect 56013 62199 56069 62201
rect 56224 62253 56280 62255
rect 56224 62201 56226 62253
rect 56226 62201 56278 62253
rect 56278 62201 56280 62253
rect 56224 62199 56280 62201
rect 56435 62253 56491 62255
rect 56435 62201 56437 62253
rect 56437 62201 56489 62253
rect 56489 62201 56491 62253
rect 56435 62199 56491 62201
rect 56646 62253 56702 62255
rect 56646 62201 56648 62253
rect 56648 62201 56700 62253
rect 56700 62201 56702 62253
rect 56646 62199 56702 62201
rect 56857 62253 56913 62255
rect 56857 62201 56859 62253
rect 56859 62201 56911 62253
rect 56911 62201 56913 62253
rect 56857 62199 56913 62201
rect 57068 62253 57124 62255
rect 57068 62201 57070 62253
rect 57070 62201 57122 62253
rect 57122 62201 57124 62253
rect 57068 62199 57124 62201
rect 57279 62253 57335 62255
rect 57279 62201 57281 62253
rect 57281 62201 57333 62253
rect 57333 62201 57335 62253
rect 57279 62199 57335 62201
rect 27788 60453 27844 60455
rect 27788 60401 27790 60453
rect 27790 60401 27842 60453
rect 27842 60401 27844 60453
rect 27788 60399 27844 60401
rect 27999 60453 28055 60455
rect 27999 60401 28001 60453
rect 28001 60401 28053 60453
rect 28053 60401 28055 60453
rect 27999 60399 28055 60401
rect 28210 60453 28266 60455
rect 28210 60401 28212 60453
rect 28212 60401 28264 60453
rect 28264 60401 28266 60453
rect 28210 60399 28266 60401
rect 28421 60453 28477 60455
rect 28421 60401 28423 60453
rect 28423 60401 28475 60453
rect 28475 60401 28477 60453
rect 28421 60399 28477 60401
rect 28632 60453 28688 60455
rect 28632 60401 28634 60453
rect 28634 60401 28686 60453
rect 28686 60401 28688 60453
rect 28632 60399 28688 60401
rect 28843 60453 28899 60455
rect 28843 60401 28845 60453
rect 28845 60401 28897 60453
rect 28897 60401 28899 60453
rect 28843 60399 28899 60401
rect 29054 60453 29110 60455
rect 29054 60401 29056 60453
rect 29056 60401 29108 60453
rect 29108 60401 29110 60453
rect 29054 60399 29110 60401
rect 56013 60453 56069 60455
rect 56013 60401 56015 60453
rect 56015 60401 56067 60453
rect 56067 60401 56069 60453
rect 56013 60399 56069 60401
rect 56224 60453 56280 60455
rect 56224 60401 56226 60453
rect 56226 60401 56278 60453
rect 56278 60401 56280 60453
rect 56224 60399 56280 60401
rect 56435 60453 56491 60455
rect 56435 60401 56437 60453
rect 56437 60401 56489 60453
rect 56489 60401 56491 60453
rect 56435 60399 56491 60401
rect 56646 60453 56702 60455
rect 56646 60401 56648 60453
rect 56648 60401 56700 60453
rect 56700 60401 56702 60453
rect 56646 60399 56702 60401
rect 56857 60453 56913 60455
rect 56857 60401 56859 60453
rect 56859 60401 56911 60453
rect 56911 60401 56913 60453
rect 56857 60399 56913 60401
rect 57068 60453 57124 60455
rect 57068 60401 57070 60453
rect 57070 60401 57122 60453
rect 57122 60401 57124 60453
rect 57068 60399 57124 60401
rect 57279 60453 57335 60455
rect 57279 60401 57281 60453
rect 57281 60401 57333 60453
rect 57333 60401 57335 60453
rect 57279 60399 57335 60401
rect 27788 58653 27844 58655
rect 27788 58601 27790 58653
rect 27790 58601 27842 58653
rect 27842 58601 27844 58653
rect 27788 58599 27844 58601
rect 27999 58653 28055 58655
rect 27999 58601 28001 58653
rect 28001 58601 28053 58653
rect 28053 58601 28055 58653
rect 27999 58599 28055 58601
rect 28210 58653 28266 58655
rect 28210 58601 28212 58653
rect 28212 58601 28264 58653
rect 28264 58601 28266 58653
rect 28210 58599 28266 58601
rect 28421 58653 28477 58655
rect 28421 58601 28423 58653
rect 28423 58601 28475 58653
rect 28475 58601 28477 58653
rect 28421 58599 28477 58601
rect 28632 58653 28688 58655
rect 28632 58601 28634 58653
rect 28634 58601 28686 58653
rect 28686 58601 28688 58653
rect 28632 58599 28688 58601
rect 28843 58653 28899 58655
rect 28843 58601 28845 58653
rect 28845 58601 28897 58653
rect 28897 58601 28899 58653
rect 28843 58599 28899 58601
rect 29054 58653 29110 58655
rect 29054 58601 29056 58653
rect 29056 58601 29108 58653
rect 29108 58601 29110 58653
rect 29054 58599 29110 58601
rect 56013 58653 56069 58655
rect 56013 58601 56015 58653
rect 56015 58601 56067 58653
rect 56067 58601 56069 58653
rect 56013 58599 56069 58601
rect 56224 58653 56280 58655
rect 56224 58601 56226 58653
rect 56226 58601 56278 58653
rect 56278 58601 56280 58653
rect 56224 58599 56280 58601
rect 56435 58653 56491 58655
rect 56435 58601 56437 58653
rect 56437 58601 56489 58653
rect 56489 58601 56491 58653
rect 56435 58599 56491 58601
rect 56646 58653 56702 58655
rect 56646 58601 56648 58653
rect 56648 58601 56700 58653
rect 56700 58601 56702 58653
rect 56646 58599 56702 58601
rect 56857 58653 56913 58655
rect 56857 58601 56859 58653
rect 56859 58601 56911 58653
rect 56911 58601 56913 58653
rect 56857 58599 56913 58601
rect 57068 58653 57124 58655
rect 57068 58601 57070 58653
rect 57070 58601 57122 58653
rect 57122 58601 57124 58653
rect 57068 58599 57124 58601
rect 57279 58653 57335 58655
rect 57279 58601 57281 58653
rect 57281 58601 57333 58653
rect 57333 58601 57335 58653
rect 57279 58599 57335 58601
rect 27788 56853 27844 56855
rect 27788 56801 27790 56853
rect 27790 56801 27842 56853
rect 27842 56801 27844 56853
rect 27788 56799 27844 56801
rect 27999 56853 28055 56855
rect 27999 56801 28001 56853
rect 28001 56801 28053 56853
rect 28053 56801 28055 56853
rect 27999 56799 28055 56801
rect 28210 56853 28266 56855
rect 28210 56801 28212 56853
rect 28212 56801 28264 56853
rect 28264 56801 28266 56853
rect 28210 56799 28266 56801
rect 28421 56853 28477 56855
rect 28421 56801 28423 56853
rect 28423 56801 28475 56853
rect 28475 56801 28477 56853
rect 28421 56799 28477 56801
rect 28632 56853 28688 56855
rect 28632 56801 28634 56853
rect 28634 56801 28686 56853
rect 28686 56801 28688 56853
rect 28632 56799 28688 56801
rect 28843 56853 28899 56855
rect 28843 56801 28845 56853
rect 28845 56801 28897 56853
rect 28897 56801 28899 56853
rect 28843 56799 28899 56801
rect 29054 56853 29110 56855
rect 29054 56801 29056 56853
rect 29056 56801 29108 56853
rect 29108 56801 29110 56853
rect 29054 56799 29110 56801
rect 56013 56853 56069 56855
rect 56013 56801 56015 56853
rect 56015 56801 56067 56853
rect 56067 56801 56069 56853
rect 56013 56799 56069 56801
rect 56224 56853 56280 56855
rect 56224 56801 56226 56853
rect 56226 56801 56278 56853
rect 56278 56801 56280 56853
rect 56224 56799 56280 56801
rect 56435 56853 56491 56855
rect 56435 56801 56437 56853
rect 56437 56801 56489 56853
rect 56489 56801 56491 56853
rect 56435 56799 56491 56801
rect 56646 56853 56702 56855
rect 56646 56801 56648 56853
rect 56648 56801 56700 56853
rect 56700 56801 56702 56853
rect 56646 56799 56702 56801
rect 56857 56853 56913 56855
rect 56857 56801 56859 56853
rect 56859 56801 56911 56853
rect 56911 56801 56913 56853
rect 56857 56799 56913 56801
rect 57068 56853 57124 56855
rect 57068 56801 57070 56853
rect 57070 56801 57122 56853
rect 57122 56801 57124 56853
rect 57068 56799 57124 56801
rect 57279 56853 57335 56855
rect 57279 56801 57281 56853
rect 57281 56801 57333 56853
rect 57333 56801 57335 56853
rect 57279 56799 57335 56801
rect 27788 55053 27844 55055
rect 27788 55001 27790 55053
rect 27790 55001 27842 55053
rect 27842 55001 27844 55053
rect 27788 54999 27844 55001
rect 27999 55053 28055 55055
rect 27999 55001 28001 55053
rect 28001 55001 28053 55053
rect 28053 55001 28055 55053
rect 27999 54999 28055 55001
rect 28210 55053 28266 55055
rect 28210 55001 28212 55053
rect 28212 55001 28264 55053
rect 28264 55001 28266 55053
rect 28210 54999 28266 55001
rect 28421 55053 28477 55055
rect 28421 55001 28423 55053
rect 28423 55001 28475 55053
rect 28475 55001 28477 55053
rect 28421 54999 28477 55001
rect 28632 55053 28688 55055
rect 28632 55001 28634 55053
rect 28634 55001 28686 55053
rect 28686 55001 28688 55053
rect 28632 54999 28688 55001
rect 28843 55053 28899 55055
rect 28843 55001 28845 55053
rect 28845 55001 28897 55053
rect 28897 55001 28899 55053
rect 28843 54999 28899 55001
rect 29054 55053 29110 55055
rect 29054 55001 29056 55053
rect 29056 55001 29108 55053
rect 29108 55001 29110 55053
rect 29054 54999 29110 55001
rect 56013 55053 56069 55055
rect 56013 55001 56015 55053
rect 56015 55001 56067 55053
rect 56067 55001 56069 55053
rect 56013 54999 56069 55001
rect 56224 55053 56280 55055
rect 56224 55001 56226 55053
rect 56226 55001 56278 55053
rect 56278 55001 56280 55053
rect 56224 54999 56280 55001
rect 56435 55053 56491 55055
rect 56435 55001 56437 55053
rect 56437 55001 56489 55053
rect 56489 55001 56491 55053
rect 56435 54999 56491 55001
rect 56646 55053 56702 55055
rect 56646 55001 56648 55053
rect 56648 55001 56700 55053
rect 56700 55001 56702 55053
rect 56646 54999 56702 55001
rect 56857 55053 56913 55055
rect 56857 55001 56859 55053
rect 56859 55001 56911 55053
rect 56911 55001 56913 55053
rect 56857 54999 56913 55001
rect 57068 55053 57124 55055
rect 57068 55001 57070 55053
rect 57070 55001 57122 55053
rect 57122 55001 57124 55053
rect 57068 54999 57124 55001
rect 57279 55053 57335 55055
rect 57279 55001 57281 55053
rect 57281 55001 57333 55053
rect 57333 55001 57335 55053
rect 57279 54999 57335 55001
rect 27788 53253 27844 53255
rect 27788 53201 27790 53253
rect 27790 53201 27842 53253
rect 27842 53201 27844 53253
rect 27788 53199 27844 53201
rect 27999 53253 28055 53255
rect 27999 53201 28001 53253
rect 28001 53201 28053 53253
rect 28053 53201 28055 53253
rect 27999 53199 28055 53201
rect 28210 53253 28266 53255
rect 28210 53201 28212 53253
rect 28212 53201 28264 53253
rect 28264 53201 28266 53253
rect 28210 53199 28266 53201
rect 28421 53253 28477 53255
rect 28421 53201 28423 53253
rect 28423 53201 28475 53253
rect 28475 53201 28477 53253
rect 28421 53199 28477 53201
rect 28632 53253 28688 53255
rect 28632 53201 28634 53253
rect 28634 53201 28686 53253
rect 28686 53201 28688 53253
rect 28632 53199 28688 53201
rect 28843 53253 28899 53255
rect 28843 53201 28845 53253
rect 28845 53201 28897 53253
rect 28897 53201 28899 53253
rect 28843 53199 28899 53201
rect 29054 53253 29110 53255
rect 29054 53201 29056 53253
rect 29056 53201 29108 53253
rect 29108 53201 29110 53253
rect 29054 53199 29110 53201
rect 56013 53253 56069 53255
rect 56013 53201 56015 53253
rect 56015 53201 56067 53253
rect 56067 53201 56069 53253
rect 56013 53199 56069 53201
rect 56224 53253 56280 53255
rect 56224 53201 56226 53253
rect 56226 53201 56278 53253
rect 56278 53201 56280 53253
rect 56224 53199 56280 53201
rect 56435 53253 56491 53255
rect 56435 53201 56437 53253
rect 56437 53201 56489 53253
rect 56489 53201 56491 53253
rect 56435 53199 56491 53201
rect 56646 53253 56702 53255
rect 56646 53201 56648 53253
rect 56648 53201 56700 53253
rect 56700 53201 56702 53253
rect 56646 53199 56702 53201
rect 56857 53253 56913 53255
rect 56857 53201 56859 53253
rect 56859 53201 56911 53253
rect 56911 53201 56913 53253
rect 56857 53199 56913 53201
rect 57068 53253 57124 53255
rect 57068 53201 57070 53253
rect 57070 53201 57122 53253
rect 57122 53201 57124 53253
rect 57068 53199 57124 53201
rect 57279 53253 57335 53255
rect 57279 53201 57281 53253
rect 57281 53201 57333 53253
rect 57333 53201 57335 53253
rect 57279 53199 57335 53201
rect 27788 51453 27844 51455
rect 27788 51401 27790 51453
rect 27790 51401 27842 51453
rect 27842 51401 27844 51453
rect 27788 51399 27844 51401
rect 27999 51453 28055 51455
rect 27999 51401 28001 51453
rect 28001 51401 28053 51453
rect 28053 51401 28055 51453
rect 27999 51399 28055 51401
rect 28210 51453 28266 51455
rect 28210 51401 28212 51453
rect 28212 51401 28264 51453
rect 28264 51401 28266 51453
rect 28210 51399 28266 51401
rect 28421 51453 28477 51455
rect 28421 51401 28423 51453
rect 28423 51401 28475 51453
rect 28475 51401 28477 51453
rect 28421 51399 28477 51401
rect 28632 51453 28688 51455
rect 28632 51401 28634 51453
rect 28634 51401 28686 51453
rect 28686 51401 28688 51453
rect 28632 51399 28688 51401
rect 28843 51453 28899 51455
rect 28843 51401 28845 51453
rect 28845 51401 28897 51453
rect 28897 51401 28899 51453
rect 28843 51399 28899 51401
rect 29054 51453 29110 51455
rect 29054 51401 29056 51453
rect 29056 51401 29108 51453
rect 29108 51401 29110 51453
rect 29054 51399 29110 51401
rect 56013 51453 56069 51455
rect 56013 51401 56015 51453
rect 56015 51401 56067 51453
rect 56067 51401 56069 51453
rect 56013 51399 56069 51401
rect 56224 51453 56280 51455
rect 56224 51401 56226 51453
rect 56226 51401 56278 51453
rect 56278 51401 56280 51453
rect 56224 51399 56280 51401
rect 56435 51453 56491 51455
rect 56435 51401 56437 51453
rect 56437 51401 56489 51453
rect 56489 51401 56491 51453
rect 56435 51399 56491 51401
rect 56646 51453 56702 51455
rect 56646 51401 56648 51453
rect 56648 51401 56700 51453
rect 56700 51401 56702 51453
rect 56646 51399 56702 51401
rect 56857 51453 56913 51455
rect 56857 51401 56859 51453
rect 56859 51401 56911 51453
rect 56911 51401 56913 51453
rect 56857 51399 56913 51401
rect 57068 51453 57124 51455
rect 57068 51401 57070 51453
rect 57070 51401 57122 51453
rect 57122 51401 57124 51453
rect 57068 51399 57124 51401
rect 57279 51453 57335 51455
rect 57279 51401 57281 51453
rect 57281 51401 57333 51453
rect 57333 51401 57335 51453
rect 57279 51399 57335 51401
rect 27788 49653 27844 49655
rect 27788 49601 27790 49653
rect 27790 49601 27842 49653
rect 27842 49601 27844 49653
rect 27788 49599 27844 49601
rect 27999 49653 28055 49655
rect 27999 49601 28001 49653
rect 28001 49601 28053 49653
rect 28053 49601 28055 49653
rect 27999 49599 28055 49601
rect 28210 49653 28266 49655
rect 28210 49601 28212 49653
rect 28212 49601 28264 49653
rect 28264 49601 28266 49653
rect 28210 49599 28266 49601
rect 28421 49653 28477 49655
rect 28421 49601 28423 49653
rect 28423 49601 28475 49653
rect 28475 49601 28477 49653
rect 28421 49599 28477 49601
rect 28632 49653 28688 49655
rect 28632 49601 28634 49653
rect 28634 49601 28686 49653
rect 28686 49601 28688 49653
rect 28632 49599 28688 49601
rect 28843 49653 28899 49655
rect 28843 49601 28845 49653
rect 28845 49601 28897 49653
rect 28897 49601 28899 49653
rect 28843 49599 28899 49601
rect 29054 49653 29110 49655
rect 29054 49601 29056 49653
rect 29056 49601 29108 49653
rect 29108 49601 29110 49653
rect 29054 49599 29110 49601
rect 56013 49653 56069 49655
rect 56013 49601 56015 49653
rect 56015 49601 56067 49653
rect 56067 49601 56069 49653
rect 56013 49599 56069 49601
rect 56224 49653 56280 49655
rect 56224 49601 56226 49653
rect 56226 49601 56278 49653
rect 56278 49601 56280 49653
rect 56224 49599 56280 49601
rect 56435 49653 56491 49655
rect 56435 49601 56437 49653
rect 56437 49601 56489 49653
rect 56489 49601 56491 49653
rect 56435 49599 56491 49601
rect 56646 49653 56702 49655
rect 56646 49601 56648 49653
rect 56648 49601 56700 49653
rect 56700 49601 56702 49653
rect 56646 49599 56702 49601
rect 56857 49653 56913 49655
rect 56857 49601 56859 49653
rect 56859 49601 56911 49653
rect 56911 49601 56913 49653
rect 56857 49599 56913 49601
rect 57068 49653 57124 49655
rect 57068 49601 57070 49653
rect 57070 49601 57122 49653
rect 57122 49601 57124 49653
rect 57068 49599 57124 49601
rect 57279 49653 57335 49655
rect 57279 49601 57281 49653
rect 57281 49601 57333 49653
rect 57333 49601 57335 49653
rect 57279 49599 57335 49601
rect 27788 47853 27844 47855
rect 27788 47801 27790 47853
rect 27790 47801 27842 47853
rect 27842 47801 27844 47853
rect 27788 47799 27844 47801
rect 27999 47853 28055 47855
rect 27999 47801 28001 47853
rect 28001 47801 28053 47853
rect 28053 47801 28055 47853
rect 27999 47799 28055 47801
rect 28210 47853 28266 47855
rect 28210 47801 28212 47853
rect 28212 47801 28264 47853
rect 28264 47801 28266 47853
rect 28210 47799 28266 47801
rect 28421 47853 28477 47855
rect 28421 47801 28423 47853
rect 28423 47801 28475 47853
rect 28475 47801 28477 47853
rect 28421 47799 28477 47801
rect 28632 47853 28688 47855
rect 28632 47801 28634 47853
rect 28634 47801 28686 47853
rect 28686 47801 28688 47853
rect 28632 47799 28688 47801
rect 28843 47853 28899 47855
rect 28843 47801 28845 47853
rect 28845 47801 28897 47853
rect 28897 47801 28899 47853
rect 28843 47799 28899 47801
rect 29054 47853 29110 47855
rect 29054 47801 29056 47853
rect 29056 47801 29108 47853
rect 29108 47801 29110 47853
rect 29054 47799 29110 47801
rect 56013 47853 56069 47855
rect 56013 47801 56015 47853
rect 56015 47801 56067 47853
rect 56067 47801 56069 47853
rect 56013 47799 56069 47801
rect 56224 47853 56280 47855
rect 56224 47801 56226 47853
rect 56226 47801 56278 47853
rect 56278 47801 56280 47853
rect 56224 47799 56280 47801
rect 56435 47853 56491 47855
rect 56435 47801 56437 47853
rect 56437 47801 56489 47853
rect 56489 47801 56491 47853
rect 56435 47799 56491 47801
rect 56646 47853 56702 47855
rect 56646 47801 56648 47853
rect 56648 47801 56700 47853
rect 56700 47801 56702 47853
rect 56646 47799 56702 47801
rect 56857 47853 56913 47855
rect 56857 47801 56859 47853
rect 56859 47801 56911 47853
rect 56911 47801 56913 47853
rect 56857 47799 56913 47801
rect 57068 47853 57124 47855
rect 57068 47801 57070 47853
rect 57070 47801 57122 47853
rect 57122 47801 57124 47853
rect 57068 47799 57124 47801
rect 57279 47853 57335 47855
rect 57279 47801 57281 47853
rect 57281 47801 57333 47853
rect 57333 47801 57335 47853
rect 57279 47799 57335 47801
rect 27788 46053 27844 46055
rect 27788 46001 27790 46053
rect 27790 46001 27842 46053
rect 27842 46001 27844 46053
rect 27788 45999 27844 46001
rect 27999 46053 28055 46055
rect 27999 46001 28001 46053
rect 28001 46001 28053 46053
rect 28053 46001 28055 46053
rect 27999 45999 28055 46001
rect 28210 46053 28266 46055
rect 28210 46001 28212 46053
rect 28212 46001 28264 46053
rect 28264 46001 28266 46053
rect 28210 45999 28266 46001
rect 28421 46053 28477 46055
rect 28421 46001 28423 46053
rect 28423 46001 28475 46053
rect 28475 46001 28477 46053
rect 28421 45999 28477 46001
rect 28632 46053 28688 46055
rect 28632 46001 28634 46053
rect 28634 46001 28686 46053
rect 28686 46001 28688 46053
rect 28632 45999 28688 46001
rect 28843 46053 28899 46055
rect 28843 46001 28845 46053
rect 28845 46001 28897 46053
rect 28897 46001 28899 46053
rect 28843 45999 28899 46001
rect 29054 46053 29110 46055
rect 29054 46001 29056 46053
rect 29056 46001 29108 46053
rect 29108 46001 29110 46053
rect 29054 45999 29110 46001
rect 56013 46053 56069 46055
rect 56013 46001 56015 46053
rect 56015 46001 56067 46053
rect 56067 46001 56069 46053
rect 56013 45999 56069 46001
rect 56224 46053 56280 46055
rect 56224 46001 56226 46053
rect 56226 46001 56278 46053
rect 56278 46001 56280 46053
rect 56224 45999 56280 46001
rect 56435 46053 56491 46055
rect 56435 46001 56437 46053
rect 56437 46001 56489 46053
rect 56489 46001 56491 46053
rect 56435 45999 56491 46001
rect 56646 46053 56702 46055
rect 56646 46001 56648 46053
rect 56648 46001 56700 46053
rect 56700 46001 56702 46053
rect 56646 45999 56702 46001
rect 56857 46053 56913 46055
rect 56857 46001 56859 46053
rect 56859 46001 56911 46053
rect 56911 46001 56913 46053
rect 56857 45999 56913 46001
rect 57068 46053 57124 46055
rect 57068 46001 57070 46053
rect 57070 46001 57122 46053
rect 57122 46001 57124 46053
rect 57068 45999 57124 46001
rect 57279 46053 57335 46055
rect 57279 46001 57281 46053
rect 57281 46001 57333 46053
rect 57333 46001 57335 46053
rect 57279 45999 57335 46001
rect 27788 44253 27844 44255
rect 27788 44201 27790 44253
rect 27790 44201 27842 44253
rect 27842 44201 27844 44253
rect 27788 44199 27844 44201
rect 27999 44253 28055 44255
rect 27999 44201 28001 44253
rect 28001 44201 28053 44253
rect 28053 44201 28055 44253
rect 27999 44199 28055 44201
rect 28210 44253 28266 44255
rect 28210 44201 28212 44253
rect 28212 44201 28264 44253
rect 28264 44201 28266 44253
rect 28210 44199 28266 44201
rect 28421 44253 28477 44255
rect 28421 44201 28423 44253
rect 28423 44201 28475 44253
rect 28475 44201 28477 44253
rect 28421 44199 28477 44201
rect 28632 44253 28688 44255
rect 28632 44201 28634 44253
rect 28634 44201 28686 44253
rect 28686 44201 28688 44253
rect 28632 44199 28688 44201
rect 28843 44253 28899 44255
rect 28843 44201 28845 44253
rect 28845 44201 28897 44253
rect 28897 44201 28899 44253
rect 28843 44199 28899 44201
rect 29054 44253 29110 44255
rect 29054 44201 29056 44253
rect 29056 44201 29108 44253
rect 29108 44201 29110 44253
rect 29054 44199 29110 44201
rect 56013 44253 56069 44255
rect 56013 44201 56015 44253
rect 56015 44201 56067 44253
rect 56067 44201 56069 44253
rect 56013 44199 56069 44201
rect 56224 44253 56280 44255
rect 56224 44201 56226 44253
rect 56226 44201 56278 44253
rect 56278 44201 56280 44253
rect 56224 44199 56280 44201
rect 56435 44253 56491 44255
rect 56435 44201 56437 44253
rect 56437 44201 56489 44253
rect 56489 44201 56491 44253
rect 56435 44199 56491 44201
rect 56646 44253 56702 44255
rect 56646 44201 56648 44253
rect 56648 44201 56700 44253
rect 56700 44201 56702 44253
rect 56646 44199 56702 44201
rect 56857 44253 56913 44255
rect 56857 44201 56859 44253
rect 56859 44201 56911 44253
rect 56911 44201 56913 44253
rect 56857 44199 56913 44201
rect 57068 44253 57124 44255
rect 57068 44201 57070 44253
rect 57070 44201 57122 44253
rect 57122 44201 57124 44253
rect 57068 44199 57124 44201
rect 57279 44253 57335 44255
rect 57279 44201 57281 44253
rect 57281 44201 57333 44253
rect 57333 44201 57335 44253
rect 57279 44199 57335 44201
rect 27788 42453 27844 42455
rect 27788 42401 27790 42453
rect 27790 42401 27842 42453
rect 27842 42401 27844 42453
rect 27788 42399 27844 42401
rect 27999 42453 28055 42455
rect 27999 42401 28001 42453
rect 28001 42401 28053 42453
rect 28053 42401 28055 42453
rect 27999 42399 28055 42401
rect 28210 42453 28266 42455
rect 28210 42401 28212 42453
rect 28212 42401 28264 42453
rect 28264 42401 28266 42453
rect 28210 42399 28266 42401
rect 28421 42453 28477 42455
rect 28421 42401 28423 42453
rect 28423 42401 28475 42453
rect 28475 42401 28477 42453
rect 28421 42399 28477 42401
rect 28632 42453 28688 42455
rect 28632 42401 28634 42453
rect 28634 42401 28686 42453
rect 28686 42401 28688 42453
rect 28632 42399 28688 42401
rect 28843 42453 28899 42455
rect 28843 42401 28845 42453
rect 28845 42401 28897 42453
rect 28897 42401 28899 42453
rect 28843 42399 28899 42401
rect 29054 42453 29110 42455
rect 29054 42401 29056 42453
rect 29056 42401 29108 42453
rect 29108 42401 29110 42453
rect 29054 42399 29110 42401
rect 56013 42453 56069 42455
rect 56013 42401 56015 42453
rect 56015 42401 56067 42453
rect 56067 42401 56069 42453
rect 56013 42399 56069 42401
rect 56224 42453 56280 42455
rect 56224 42401 56226 42453
rect 56226 42401 56278 42453
rect 56278 42401 56280 42453
rect 56224 42399 56280 42401
rect 56435 42453 56491 42455
rect 56435 42401 56437 42453
rect 56437 42401 56489 42453
rect 56489 42401 56491 42453
rect 56435 42399 56491 42401
rect 56646 42453 56702 42455
rect 56646 42401 56648 42453
rect 56648 42401 56700 42453
rect 56700 42401 56702 42453
rect 56646 42399 56702 42401
rect 56857 42453 56913 42455
rect 56857 42401 56859 42453
rect 56859 42401 56911 42453
rect 56911 42401 56913 42453
rect 56857 42399 56913 42401
rect 57068 42453 57124 42455
rect 57068 42401 57070 42453
rect 57070 42401 57122 42453
rect 57122 42401 57124 42453
rect 57068 42399 57124 42401
rect 57279 42453 57335 42455
rect 57279 42401 57281 42453
rect 57281 42401 57333 42453
rect 57333 42401 57335 42453
rect 57279 42399 57335 42401
rect 27788 40653 27844 40655
rect 27788 40601 27790 40653
rect 27790 40601 27842 40653
rect 27842 40601 27844 40653
rect 27788 40599 27844 40601
rect 27999 40653 28055 40655
rect 27999 40601 28001 40653
rect 28001 40601 28053 40653
rect 28053 40601 28055 40653
rect 27999 40599 28055 40601
rect 28210 40653 28266 40655
rect 28210 40601 28212 40653
rect 28212 40601 28264 40653
rect 28264 40601 28266 40653
rect 28210 40599 28266 40601
rect 28421 40653 28477 40655
rect 28421 40601 28423 40653
rect 28423 40601 28475 40653
rect 28475 40601 28477 40653
rect 28421 40599 28477 40601
rect 28632 40653 28688 40655
rect 28632 40601 28634 40653
rect 28634 40601 28686 40653
rect 28686 40601 28688 40653
rect 28632 40599 28688 40601
rect 28843 40653 28899 40655
rect 28843 40601 28845 40653
rect 28845 40601 28897 40653
rect 28897 40601 28899 40653
rect 28843 40599 28899 40601
rect 29054 40653 29110 40655
rect 29054 40601 29056 40653
rect 29056 40601 29108 40653
rect 29108 40601 29110 40653
rect 29054 40599 29110 40601
rect 56013 40653 56069 40655
rect 56013 40601 56015 40653
rect 56015 40601 56067 40653
rect 56067 40601 56069 40653
rect 56013 40599 56069 40601
rect 56224 40653 56280 40655
rect 56224 40601 56226 40653
rect 56226 40601 56278 40653
rect 56278 40601 56280 40653
rect 56224 40599 56280 40601
rect 56435 40653 56491 40655
rect 56435 40601 56437 40653
rect 56437 40601 56489 40653
rect 56489 40601 56491 40653
rect 56435 40599 56491 40601
rect 56646 40653 56702 40655
rect 56646 40601 56648 40653
rect 56648 40601 56700 40653
rect 56700 40601 56702 40653
rect 56646 40599 56702 40601
rect 56857 40653 56913 40655
rect 56857 40601 56859 40653
rect 56859 40601 56911 40653
rect 56911 40601 56913 40653
rect 56857 40599 56913 40601
rect 57068 40653 57124 40655
rect 57068 40601 57070 40653
rect 57070 40601 57122 40653
rect 57122 40601 57124 40653
rect 57068 40599 57124 40601
rect 57279 40653 57335 40655
rect 57279 40601 57281 40653
rect 57281 40601 57333 40653
rect 57333 40601 57335 40653
rect 57279 40599 57335 40601
rect 27788 38853 27844 38855
rect 27788 38801 27790 38853
rect 27790 38801 27842 38853
rect 27842 38801 27844 38853
rect 27788 38799 27844 38801
rect 27999 38853 28055 38855
rect 27999 38801 28001 38853
rect 28001 38801 28053 38853
rect 28053 38801 28055 38853
rect 27999 38799 28055 38801
rect 28210 38853 28266 38855
rect 28210 38801 28212 38853
rect 28212 38801 28264 38853
rect 28264 38801 28266 38853
rect 28210 38799 28266 38801
rect 28421 38853 28477 38855
rect 28421 38801 28423 38853
rect 28423 38801 28475 38853
rect 28475 38801 28477 38853
rect 28421 38799 28477 38801
rect 28632 38853 28688 38855
rect 28632 38801 28634 38853
rect 28634 38801 28686 38853
rect 28686 38801 28688 38853
rect 28632 38799 28688 38801
rect 28843 38853 28899 38855
rect 28843 38801 28845 38853
rect 28845 38801 28897 38853
rect 28897 38801 28899 38853
rect 28843 38799 28899 38801
rect 29054 38853 29110 38855
rect 29054 38801 29056 38853
rect 29056 38801 29108 38853
rect 29108 38801 29110 38853
rect 29054 38799 29110 38801
rect 56013 38853 56069 38855
rect 56013 38801 56015 38853
rect 56015 38801 56067 38853
rect 56067 38801 56069 38853
rect 56013 38799 56069 38801
rect 56224 38853 56280 38855
rect 56224 38801 56226 38853
rect 56226 38801 56278 38853
rect 56278 38801 56280 38853
rect 56224 38799 56280 38801
rect 56435 38853 56491 38855
rect 56435 38801 56437 38853
rect 56437 38801 56489 38853
rect 56489 38801 56491 38853
rect 56435 38799 56491 38801
rect 56646 38853 56702 38855
rect 56646 38801 56648 38853
rect 56648 38801 56700 38853
rect 56700 38801 56702 38853
rect 56646 38799 56702 38801
rect 56857 38853 56913 38855
rect 56857 38801 56859 38853
rect 56859 38801 56911 38853
rect 56911 38801 56913 38853
rect 56857 38799 56913 38801
rect 57068 38853 57124 38855
rect 57068 38801 57070 38853
rect 57070 38801 57122 38853
rect 57122 38801 57124 38853
rect 57068 38799 57124 38801
rect 57279 38853 57335 38855
rect 57279 38801 57281 38853
rect 57281 38801 57333 38853
rect 57333 38801 57335 38853
rect 57279 38799 57335 38801
rect 27788 37053 27844 37055
rect 27788 37001 27790 37053
rect 27790 37001 27842 37053
rect 27842 37001 27844 37053
rect 27788 36999 27844 37001
rect 27999 37053 28055 37055
rect 27999 37001 28001 37053
rect 28001 37001 28053 37053
rect 28053 37001 28055 37053
rect 27999 36999 28055 37001
rect 28210 37053 28266 37055
rect 28210 37001 28212 37053
rect 28212 37001 28264 37053
rect 28264 37001 28266 37053
rect 28210 36999 28266 37001
rect 28421 37053 28477 37055
rect 28421 37001 28423 37053
rect 28423 37001 28475 37053
rect 28475 37001 28477 37053
rect 28421 36999 28477 37001
rect 28632 37053 28688 37055
rect 28632 37001 28634 37053
rect 28634 37001 28686 37053
rect 28686 37001 28688 37053
rect 28632 36999 28688 37001
rect 28843 37053 28899 37055
rect 28843 37001 28845 37053
rect 28845 37001 28897 37053
rect 28897 37001 28899 37053
rect 28843 36999 28899 37001
rect 29054 37053 29110 37055
rect 29054 37001 29056 37053
rect 29056 37001 29108 37053
rect 29108 37001 29110 37053
rect 29054 36999 29110 37001
rect 56013 37053 56069 37055
rect 56013 37001 56015 37053
rect 56015 37001 56067 37053
rect 56067 37001 56069 37053
rect 56013 36999 56069 37001
rect 56224 37053 56280 37055
rect 56224 37001 56226 37053
rect 56226 37001 56278 37053
rect 56278 37001 56280 37053
rect 56224 36999 56280 37001
rect 56435 37053 56491 37055
rect 56435 37001 56437 37053
rect 56437 37001 56489 37053
rect 56489 37001 56491 37053
rect 56435 36999 56491 37001
rect 56646 37053 56702 37055
rect 56646 37001 56648 37053
rect 56648 37001 56700 37053
rect 56700 37001 56702 37053
rect 56646 36999 56702 37001
rect 56857 37053 56913 37055
rect 56857 37001 56859 37053
rect 56859 37001 56911 37053
rect 56911 37001 56913 37053
rect 56857 36999 56913 37001
rect 57068 37053 57124 37055
rect 57068 37001 57070 37053
rect 57070 37001 57122 37053
rect 57122 37001 57124 37053
rect 57068 36999 57124 37001
rect 57279 37053 57335 37055
rect 57279 37001 57281 37053
rect 57281 37001 57333 37053
rect 57333 37001 57335 37053
rect 57279 36999 57335 37001
rect 36958 35825 37014 35881
rect 37169 35825 37225 35881
rect 37381 35825 37437 35881
rect 37592 35825 37648 35881
rect 27447 34990 27503 34992
rect 27447 34938 27449 34990
rect 27449 34938 27501 34990
rect 27501 34938 27503 34990
rect 27447 34936 27503 34938
rect 27571 34990 27627 34992
rect 27571 34938 27573 34990
rect 27573 34938 27625 34990
rect 27625 34938 27627 34990
rect 27571 34936 27627 34938
rect 27695 34990 27751 34992
rect 27695 34938 27697 34990
rect 27697 34938 27749 34990
rect 27749 34938 27751 34990
rect 27695 34936 27751 34938
rect 27447 34866 27503 34868
rect 27447 34814 27449 34866
rect 27449 34814 27501 34866
rect 27501 34814 27503 34866
rect 27447 34812 27503 34814
rect 27571 34866 27627 34868
rect 27571 34814 27573 34866
rect 27573 34814 27625 34866
rect 27625 34814 27627 34866
rect 27571 34812 27627 34814
rect 27695 34866 27751 34868
rect 27695 34814 27697 34866
rect 27697 34814 27749 34866
rect 27749 34814 27751 34866
rect 27695 34812 27751 34814
rect 27447 34742 27503 34744
rect 27447 34690 27449 34742
rect 27449 34690 27501 34742
rect 27501 34690 27503 34742
rect 27447 34688 27503 34690
rect 27571 34742 27627 34744
rect 27571 34690 27573 34742
rect 27573 34690 27625 34742
rect 27625 34690 27627 34742
rect 27571 34688 27627 34690
rect 27695 34742 27751 34744
rect 27695 34690 27697 34742
rect 27697 34690 27749 34742
rect 27749 34690 27751 34742
rect 27695 34688 27751 34690
rect 27447 34618 27503 34620
rect 27447 34566 27449 34618
rect 27449 34566 27501 34618
rect 27501 34566 27503 34618
rect 27447 34564 27503 34566
rect 27571 34618 27627 34620
rect 27571 34566 27573 34618
rect 27573 34566 27625 34618
rect 27625 34566 27627 34618
rect 27571 34564 27627 34566
rect 27695 34618 27751 34620
rect 27695 34566 27697 34618
rect 27697 34566 27749 34618
rect 27749 34566 27751 34618
rect 27695 34564 27751 34566
rect 26859 33955 26915 34011
rect 27071 33955 27127 34011
rect 26859 33737 26915 33793
rect 27071 33737 27127 33793
rect 26859 33520 26915 33576
rect 27071 33520 27127 33576
rect 26859 33302 26915 33358
rect 27071 33302 27127 33358
rect 26859 33084 26915 33140
rect 27071 33084 27127 33140
rect 26859 32866 26915 32922
rect 27071 32866 27127 32922
rect 26859 32649 26915 32705
rect 27071 32649 27127 32705
rect 26859 32431 26915 32487
rect 27071 32431 27127 32487
rect 26859 32075 26861 32088
rect 26861 32075 26913 32088
rect 26913 32075 26915 32088
rect 26859 32032 26915 32075
rect 27071 32075 27073 32088
rect 27073 32075 27125 32088
rect 27125 32075 27127 32088
rect 27071 32032 27127 32075
rect 26859 31857 26861 31870
rect 26861 31857 26913 31870
rect 26913 31857 26915 31870
rect 26859 31814 26915 31857
rect 27071 31857 27073 31870
rect 27073 31857 27125 31870
rect 27125 31857 27127 31870
rect 27071 31814 27127 31857
rect 26859 31639 26861 31652
rect 26861 31639 26913 31652
rect 26913 31639 26915 31652
rect 26859 31596 26915 31639
rect 27071 31639 27073 31652
rect 27073 31639 27125 31652
rect 27125 31639 27127 31652
rect 27071 31596 27127 31639
rect 26859 29950 26915 29968
rect 26859 29912 26861 29950
rect 26861 29912 26913 29950
rect 26913 29912 26915 29950
rect 27071 29950 27127 29968
rect 27071 29912 27073 29950
rect 27073 29912 27125 29950
rect 27125 29912 27127 29950
rect 26859 29733 26915 29750
rect 26859 29694 26861 29733
rect 26861 29694 26913 29733
rect 26913 29694 26915 29733
rect 27071 29733 27127 29750
rect 27071 29694 27073 29733
rect 27073 29694 27125 29733
rect 27125 29694 27127 29733
rect 26859 29515 26915 29533
rect 26859 29477 26861 29515
rect 26861 29477 26913 29515
rect 26913 29477 26915 29515
rect 27071 29515 27127 29533
rect 27071 29477 27073 29515
rect 27073 29477 27125 29515
rect 27125 29477 27127 29515
rect 26859 29297 26915 29315
rect 26859 29259 26861 29297
rect 26861 29259 26913 29297
rect 26913 29259 26915 29297
rect 27071 29297 27127 29315
rect 27071 29259 27073 29297
rect 27073 29259 27125 29297
rect 27125 29259 27127 29297
rect 26859 29080 26915 29098
rect 26859 29042 26861 29080
rect 26861 29042 26913 29080
rect 26913 29042 26915 29080
rect 27071 29080 27127 29098
rect 27071 29042 27073 29080
rect 27073 29042 27125 29080
rect 27125 29042 27127 29080
rect 26859 28862 26915 28880
rect 26859 28824 26861 28862
rect 26861 28824 26913 28862
rect 26913 28824 26915 28862
rect 27071 28862 27127 28880
rect 27071 28824 27073 28862
rect 27073 28824 27125 28862
rect 27125 28824 27127 28862
rect 26859 28644 26915 28662
rect 26859 28606 26861 28644
rect 26861 28606 26913 28644
rect 26913 28606 26915 28644
rect 27071 28644 27127 28662
rect 27071 28606 27073 28644
rect 27073 28606 27125 28644
rect 27125 28606 27127 28644
rect 26859 28427 26915 28444
rect 26859 28388 26861 28427
rect 26861 28388 26913 28427
rect 26913 28388 26915 28427
rect 27071 28427 27127 28444
rect 27071 28388 27073 28427
rect 27073 28388 27125 28427
rect 27125 28388 27127 28427
rect 26859 28209 26915 28227
rect 26859 28171 26861 28209
rect 26861 28171 26913 28209
rect 26913 28171 26915 28209
rect 27071 28209 27127 28227
rect 27071 28171 27073 28209
rect 27073 28171 27125 28209
rect 27125 28171 27127 28209
rect 26859 27992 26915 28009
rect 26859 27953 26861 27992
rect 26861 27953 26913 27992
rect 26913 27953 26915 27992
rect 27071 27992 27127 28009
rect 27071 27953 27073 27992
rect 27073 27953 27125 27992
rect 27125 27953 27127 27992
rect 26859 27774 26915 27792
rect 26859 27736 26861 27774
rect 26861 27736 26913 27774
rect 26913 27736 26915 27774
rect 27071 27774 27127 27792
rect 27071 27736 27073 27774
rect 27073 27736 27125 27774
rect 27125 27736 27127 27774
rect 26859 27556 26915 27574
rect 26859 27518 26861 27556
rect 26861 27518 26913 27556
rect 26913 27518 26915 27556
rect 27071 27556 27127 27574
rect 27071 27518 27073 27556
rect 27073 27518 27125 27556
rect 27125 27518 27127 27556
rect 25404 27269 25460 27325
rect 25528 27269 25584 27325
rect 25652 27269 25708 27325
rect 25776 27269 25832 27325
rect 25900 27269 25956 27325
rect 25404 27145 25460 27201
rect 25528 27145 25584 27201
rect 25652 27145 25708 27201
rect 25776 27145 25832 27201
rect 25900 27145 25956 27201
rect 25404 27021 25460 27077
rect 25528 27021 25584 27077
rect 25652 27021 25708 27077
rect 25776 27021 25832 27077
rect 25900 27021 25956 27077
rect 25404 26897 25460 26953
rect 25528 26897 25584 26953
rect 25652 26897 25708 26953
rect 25776 26897 25832 26953
rect 25900 26897 25956 26953
rect 25404 26773 25460 26829
rect 25528 26773 25584 26829
rect 25652 26773 25708 26829
rect 25776 26773 25832 26829
rect 25900 26773 25956 26829
rect 25404 26649 25460 26705
rect 25528 26649 25584 26705
rect 25652 26649 25708 26705
rect 25776 26649 25832 26705
rect 25900 26649 25956 26705
rect 25404 26525 25460 26581
rect 25528 26525 25584 26581
rect 25652 26525 25708 26581
rect 25776 26525 25832 26581
rect 25900 26525 25956 26581
rect 26450 26126 26610 26286
rect 26092 25807 26252 25967
rect 25756 25487 25916 25647
rect 25421 25168 25581 25328
rect 25081 24477 25241 24637
rect 24744 24156 24904 24316
rect 24416 23835 24576 23995
rect 24057 23513 24217 23673
rect 26465 19532 26625 19692
rect 26858 24074 27122 24075
rect 26858 24022 26861 24074
rect 26861 24022 26913 24074
rect 26913 24022 27073 24074
rect 27073 24022 27122 24074
rect 26858 23857 27122 24022
rect 26858 23805 26861 23857
rect 26861 23805 26913 23857
rect 26913 23805 27073 23857
rect 27073 23805 27122 23857
rect 26858 23639 27122 23805
rect 26858 23587 26861 23639
rect 26861 23587 26913 23639
rect 26913 23587 27073 23639
rect 27073 23587 27122 23639
rect 26858 23421 27122 23587
rect 26858 23369 26861 23421
rect 26861 23369 26913 23421
rect 26913 23369 27073 23421
rect 27073 23369 27122 23421
rect 26858 23204 27122 23369
rect 26858 23187 26861 23204
rect 26861 23187 26913 23204
rect 26913 23187 27073 23204
rect 27073 23187 27122 23204
rect 26924 20540 27073 20570
rect 27073 20540 27084 20570
rect 26924 20410 27084 20540
rect 26924 20157 27084 20226
rect 26924 20105 27073 20157
rect 27073 20105 27084 20157
rect 26924 20066 27084 20105
rect 26107 19187 26267 19347
rect 25771 18867 25931 19027
rect 25434 18524 25594 18684
rect 25094 18190 25254 18350
rect 24757 17817 24917 17977
rect 24429 17496 24589 17656
rect 24069 17157 24229 17317
rect 26859 14063 26915 14119
rect 27071 14063 27127 14119
rect 26859 13846 26915 13902
rect 27071 13846 27127 13902
rect 26859 13628 26915 13684
rect 27071 13628 27127 13684
rect 26859 13411 26915 13467
rect 27071 13411 27127 13467
rect 26859 13193 26915 13249
rect 27071 13193 27127 13249
rect 26859 12975 26915 13031
rect 27071 12975 27127 13031
rect 26859 12757 26915 12813
rect 27071 12757 27127 12813
rect 26859 12540 26915 12596
rect 27071 12540 27127 12596
rect 26859 12322 26915 12378
rect 27071 12322 27127 12378
rect 26859 12105 26915 12161
rect 27071 12105 27127 12161
rect 26859 9351 26915 9407
rect 27071 9351 27127 9407
rect 26859 9134 26915 9190
rect 27071 9134 27127 9190
rect 26859 8916 26915 8972
rect 27071 8916 27127 8972
rect 26859 8698 26915 8754
rect 27071 8698 27127 8754
rect 26859 8480 26915 8536
rect 27071 8480 27127 8536
rect 26859 8263 26915 8319
rect 27071 8263 27127 8319
rect 26859 5523 26861 5539
rect 26861 5523 26913 5539
rect 26913 5523 26915 5539
rect 26859 5483 26915 5523
rect 27071 5523 27073 5539
rect 27073 5523 27125 5539
rect 27125 5523 27127 5539
rect 27071 5483 27127 5523
rect 26859 5306 26861 5321
rect 26861 5306 26913 5321
rect 26913 5306 26915 5321
rect 26859 5265 26915 5306
rect 27071 5306 27073 5321
rect 27073 5306 27125 5321
rect 27125 5306 27127 5321
rect 27071 5265 27127 5306
rect 57996 33955 58052 34011
rect 58208 33955 58264 34011
rect 57996 33737 58052 33793
rect 58208 33737 58264 33793
rect 57996 33520 58052 33576
rect 58208 33520 58264 33576
rect 27474 33085 27530 33141
rect 27686 33085 27742 33141
rect 27474 32867 27530 32923
rect 27686 32867 27742 32923
rect 27474 32649 27530 32705
rect 27686 32649 27742 32705
rect 27474 32431 27530 32487
rect 27686 32431 27742 32487
rect 27474 31204 27476 31252
rect 27476 31204 27528 31252
rect 27528 31204 27530 31252
rect 27474 31196 27530 31204
rect 27686 31204 27688 31252
rect 27688 31204 27740 31252
rect 27740 31204 27742 31252
rect 27686 31196 27742 31204
rect 27474 30986 27476 31034
rect 27476 30986 27528 31034
rect 27528 30986 27530 31034
rect 27474 30978 27530 30986
rect 27686 30986 27688 31034
rect 27688 30986 27740 31034
rect 27740 30986 27742 31034
rect 27686 30978 27742 30986
rect 27474 30769 27476 30816
rect 27476 30769 27528 30816
rect 27528 30769 27530 30816
rect 27474 30760 27530 30769
rect 27686 30769 27688 30816
rect 27688 30769 27740 30816
rect 27740 30769 27742 30816
rect 27686 30760 27742 30769
rect 27474 30551 27476 30598
rect 27476 30551 27528 30598
rect 27528 30551 27530 30598
rect 27474 30542 27530 30551
rect 27686 30551 27688 30598
rect 27688 30551 27740 30598
rect 27740 30551 27742 30598
rect 27686 30542 27742 30551
rect 27474 26743 27530 26799
rect 27686 26743 27742 26799
rect 27474 26525 27530 26581
rect 27686 26525 27742 26581
rect 27474 24972 27530 25028
rect 27686 24972 27742 25028
rect 27474 24754 27530 24810
rect 27686 24754 27742 24810
rect 27475 22934 27476 22936
rect 27476 22934 27528 22936
rect 27528 22934 27688 22936
rect 27688 22934 27739 22936
rect 27475 22768 27739 22934
rect 27475 22716 27476 22768
rect 27476 22716 27528 22768
rect 27528 22716 27688 22768
rect 27688 22716 27739 22768
rect 27475 22551 27739 22716
rect 27475 22499 27476 22551
rect 27476 22499 27528 22551
rect 27528 22499 27688 22551
rect 27688 22499 27739 22551
rect 27475 22333 27739 22499
rect 27475 22281 27476 22333
rect 27476 22281 27528 22333
rect 27528 22281 27688 22333
rect 27688 22281 27739 22333
rect 27475 22115 27739 22281
rect 27475 22063 27476 22115
rect 27476 22063 27528 22115
rect 27528 22063 27688 22115
rect 27688 22063 27739 22115
rect 27475 22048 27739 22063
rect 27474 16457 27530 16470
rect 27474 16414 27476 16457
rect 27476 16414 27528 16457
rect 27528 16414 27530 16457
rect 27686 16457 27742 16470
rect 27686 16414 27688 16457
rect 27688 16414 27740 16457
rect 27740 16414 27742 16457
rect 27474 16239 27530 16253
rect 27474 16197 27476 16239
rect 27476 16197 27528 16239
rect 27528 16197 27530 16239
rect 27686 16239 27742 16253
rect 27686 16197 27688 16239
rect 27688 16197 27740 16239
rect 27740 16197 27742 16239
rect 27474 16022 27530 16035
rect 27474 15979 27476 16022
rect 27476 15979 27528 16022
rect 27528 15979 27530 16022
rect 27686 16022 27742 16035
rect 27686 15979 27688 16022
rect 27688 15979 27740 16022
rect 27740 15979 27742 16022
rect 27474 15804 27530 15818
rect 27474 15762 27476 15804
rect 27476 15762 27528 15804
rect 27528 15762 27530 15804
rect 27686 15804 27742 15818
rect 27686 15762 27688 15804
rect 27688 15762 27740 15804
rect 27740 15762 27742 15804
rect 27474 15586 27530 15600
rect 27474 15544 27476 15586
rect 27476 15544 27528 15586
rect 27528 15544 27530 15586
rect 27686 15586 27742 15600
rect 27686 15544 27688 15586
rect 27688 15544 27740 15586
rect 27740 15544 27742 15586
rect 27474 15369 27530 15382
rect 27474 15326 27476 15369
rect 27476 15326 27528 15369
rect 27528 15326 27530 15369
rect 27686 15369 27742 15382
rect 27686 15326 27688 15369
rect 27688 15326 27740 15369
rect 27740 15326 27742 15369
rect 27474 15151 27530 15164
rect 27474 15108 27476 15151
rect 27476 15108 27528 15151
rect 27528 15108 27530 15151
rect 27686 15151 27742 15164
rect 27686 15108 27688 15151
rect 27688 15108 27740 15151
rect 27740 15108 27742 15151
rect 27474 14933 27530 14947
rect 27474 14891 27476 14933
rect 27476 14891 27528 14933
rect 27528 14891 27530 14933
rect 27686 14933 27742 14947
rect 27686 14891 27688 14933
rect 27688 14891 27740 14933
rect 27740 14891 27742 14933
rect 27474 14716 27530 14729
rect 27474 14673 27476 14716
rect 27476 14673 27528 14716
rect 27528 14673 27530 14716
rect 27686 14716 27742 14729
rect 27686 14673 27688 14716
rect 27688 14673 27740 14716
rect 27740 14673 27742 14716
rect 27474 14498 27530 14512
rect 27474 14456 27476 14498
rect 27476 14456 27528 14498
rect 27528 14456 27530 14498
rect 27686 14498 27742 14512
rect 27686 14456 27688 14498
rect 27688 14456 27740 14498
rect 27740 14456 27742 14498
rect 27474 14229 27476 14231
rect 27476 14229 27528 14231
rect 27528 14229 27530 14231
rect 27474 14175 27530 14229
rect 27686 14229 27688 14231
rect 27688 14229 27740 14231
rect 27740 14229 27742 14231
rect 27686 14175 27742 14229
rect 27474 14011 27476 14014
rect 27476 14011 27528 14014
rect 27528 14011 27530 14014
rect 27474 13958 27530 14011
rect 27686 14011 27688 14014
rect 27688 14011 27740 14014
rect 27740 14011 27742 14014
rect 27686 13958 27742 14011
rect 27474 13793 27476 13796
rect 27476 13793 27528 13796
rect 27528 13793 27530 13796
rect 27474 13740 27530 13793
rect 27686 13793 27688 13796
rect 27688 13793 27740 13796
rect 27740 13793 27742 13796
rect 27686 13740 27742 13793
rect 27474 13576 27476 13578
rect 27476 13576 27528 13578
rect 27528 13576 27530 13578
rect 27474 13522 27530 13576
rect 27686 13576 27688 13578
rect 27688 13576 27740 13578
rect 27740 13576 27742 13578
rect 27686 13522 27742 13576
rect 27474 13358 27476 13361
rect 27476 13358 27528 13361
rect 27528 13358 27530 13361
rect 27474 13305 27530 13358
rect 27686 13358 27688 13361
rect 27688 13358 27740 13361
rect 27740 13358 27742 13361
rect 27686 13305 27742 13358
rect 27474 11399 27476 11406
rect 27476 11399 27528 11406
rect 27528 11399 27530 11406
rect 27474 11350 27530 11399
rect 27686 11399 27688 11406
rect 27688 11399 27740 11406
rect 27740 11399 27742 11406
rect 27686 11350 27742 11399
rect 27474 11182 27476 11189
rect 27476 11182 27528 11189
rect 27528 11182 27530 11189
rect 27474 11133 27530 11182
rect 27686 11182 27688 11189
rect 27688 11182 27740 11189
rect 27740 11182 27742 11189
rect 27686 11133 27742 11182
rect 27474 10964 27476 10971
rect 27476 10964 27528 10971
rect 27528 10964 27530 10971
rect 27474 10915 27530 10964
rect 27686 10964 27688 10971
rect 27688 10964 27740 10971
rect 27740 10964 27742 10971
rect 27686 10915 27742 10964
rect 27474 10746 27476 10753
rect 27476 10746 27528 10753
rect 27528 10746 27530 10753
rect 27474 10697 27530 10746
rect 27686 10746 27688 10753
rect 27688 10746 27740 10753
rect 27740 10746 27742 10753
rect 27686 10697 27742 10746
rect 27474 10529 27476 10535
rect 27476 10529 27528 10535
rect 27528 10529 27530 10535
rect 27474 10479 27530 10529
rect 27686 10529 27688 10535
rect 27688 10529 27740 10535
rect 27740 10529 27742 10535
rect 27686 10479 27742 10529
rect 27474 10311 27476 10318
rect 27476 10311 27528 10318
rect 27528 10311 27530 10318
rect 27474 10262 27530 10311
rect 27686 10311 27688 10318
rect 27688 10311 27740 10318
rect 27740 10311 27742 10318
rect 27686 10262 27742 10311
rect 57381 33085 57437 33141
rect 57593 33085 57649 33141
rect 57381 32867 57437 32923
rect 57593 32867 57649 32923
rect 57381 32649 57437 32705
rect 57593 32649 57649 32705
rect 57381 32431 57437 32487
rect 57593 32431 57649 32487
rect 57381 31204 57383 31252
rect 57383 31204 57435 31252
rect 57435 31204 57437 31252
rect 57381 31196 57437 31204
rect 57593 31204 57595 31252
rect 57595 31204 57647 31252
rect 57647 31204 57649 31252
rect 57593 31196 57649 31204
rect 57381 30986 57383 31034
rect 57383 30986 57435 31034
rect 57435 30986 57437 31034
rect 57381 30978 57437 30986
rect 57593 30986 57595 31034
rect 57595 30986 57647 31034
rect 57647 30986 57649 31034
rect 57593 30978 57649 30986
rect 57381 30769 57383 30816
rect 57383 30769 57435 30816
rect 57435 30769 57437 30816
rect 57381 30760 57437 30769
rect 57593 30769 57595 30816
rect 57595 30769 57647 30816
rect 57647 30769 57649 30816
rect 57593 30760 57649 30769
rect 57381 30551 57383 30598
rect 57383 30551 57435 30598
rect 57435 30551 57437 30598
rect 57381 30542 57437 30551
rect 57593 30551 57595 30598
rect 57595 30551 57647 30598
rect 57647 30551 57649 30598
rect 57593 30542 57649 30551
rect 57381 26743 57437 26799
rect 57593 26743 57649 26799
rect 57381 26525 57437 26581
rect 57593 26525 57649 26581
rect 57363 22768 57627 22923
rect 57363 22716 57383 22768
rect 57383 22716 57435 22768
rect 57435 22716 57595 22768
rect 57595 22716 57627 22768
rect 57363 22551 57627 22716
rect 57363 22499 57383 22551
rect 57383 22499 57435 22551
rect 57435 22499 57595 22551
rect 57595 22499 57627 22551
rect 57363 22333 57627 22499
rect 57363 22281 57383 22333
rect 57383 22281 57435 22333
rect 57435 22281 57595 22333
rect 57595 22281 57627 22333
rect 57363 22115 57627 22281
rect 57363 22063 57383 22115
rect 57383 22063 57435 22115
rect 57435 22063 57595 22115
rect 57595 22063 57627 22115
rect 57363 22035 57627 22063
rect 57381 16675 57437 16678
rect 57381 16623 57383 16675
rect 57383 16623 57435 16675
rect 57435 16623 57437 16675
rect 57381 16622 57437 16623
rect 57593 16675 57649 16678
rect 57593 16623 57595 16675
rect 57595 16623 57647 16675
rect 57647 16623 57649 16675
rect 57593 16622 57649 16623
rect 57381 16457 57437 16461
rect 57381 16405 57383 16457
rect 57383 16405 57435 16457
rect 57435 16405 57437 16457
rect 57593 16457 57649 16461
rect 57593 16405 57595 16457
rect 57595 16405 57647 16457
rect 57647 16405 57649 16457
rect 57381 16239 57437 16243
rect 57381 16187 57383 16239
rect 57383 16187 57435 16239
rect 57435 16187 57437 16239
rect 57593 16239 57649 16243
rect 57593 16187 57595 16239
rect 57595 16187 57647 16239
rect 57647 16187 57649 16239
rect 57381 16022 57437 16026
rect 57381 15970 57383 16022
rect 57383 15970 57435 16022
rect 57435 15970 57437 16022
rect 57593 16022 57649 16026
rect 57593 15970 57595 16022
rect 57595 15970 57647 16022
rect 57647 15970 57649 16022
rect 57381 15804 57437 15808
rect 57381 15752 57383 15804
rect 57383 15752 57435 15804
rect 57435 15752 57437 15804
rect 57593 15804 57649 15808
rect 57593 15752 57595 15804
rect 57595 15752 57647 15804
rect 57647 15752 57649 15804
rect 57381 15586 57437 15590
rect 57381 15534 57383 15586
rect 57383 15534 57435 15586
rect 57435 15534 57437 15586
rect 57593 15586 57649 15590
rect 57593 15534 57595 15586
rect 57595 15534 57647 15586
rect 57647 15534 57649 15586
rect 57381 15369 57437 15372
rect 57381 15317 57383 15369
rect 57383 15317 57435 15369
rect 57435 15317 57437 15369
rect 57381 15316 57437 15317
rect 57593 15369 57649 15372
rect 57593 15317 57595 15369
rect 57595 15317 57647 15369
rect 57647 15317 57649 15369
rect 57593 15316 57649 15317
rect 57381 15151 57437 15155
rect 57381 15099 57383 15151
rect 57383 15099 57435 15151
rect 57435 15099 57437 15151
rect 57593 15151 57649 15155
rect 57593 15099 57595 15151
rect 57595 15099 57647 15151
rect 57647 15099 57649 15151
rect 57381 14933 57437 14937
rect 57381 14881 57383 14933
rect 57383 14881 57435 14933
rect 57435 14881 57437 14933
rect 57593 14933 57649 14937
rect 57593 14881 57595 14933
rect 57595 14881 57647 14933
rect 57647 14881 57649 14933
rect 57381 14716 57437 14720
rect 57381 14664 57383 14716
rect 57383 14664 57435 14716
rect 57435 14664 57437 14716
rect 57593 14716 57649 14720
rect 57593 14664 57595 14716
rect 57595 14664 57647 14716
rect 57647 14664 57649 14716
rect 57381 11399 57383 11406
rect 57383 11399 57435 11406
rect 57435 11399 57437 11406
rect 57381 11350 57437 11399
rect 57593 11399 57595 11406
rect 57595 11399 57647 11406
rect 57647 11399 57649 11406
rect 57593 11350 57649 11399
rect 57381 11182 57383 11189
rect 57383 11182 57435 11189
rect 57435 11182 57437 11189
rect 57381 11133 57437 11182
rect 57593 11182 57595 11189
rect 57595 11182 57647 11189
rect 57647 11182 57649 11189
rect 57593 11133 57649 11182
rect 57381 10964 57383 10971
rect 57383 10964 57435 10971
rect 57435 10964 57437 10971
rect 57381 10915 57437 10964
rect 57593 10964 57595 10971
rect 57595 10964 57647 10971
rect 57647 10964 57649 10971
rect 57593 10915 57649 10964
rect 57381 10746 57383 10753
rect 57383 10746 57435 10753
rect 57435 10746 57437 10753
rect 57381 10697 57437 10746
rect 57593 10746 57595 10753
rect 57595 10746 57647 10753
rect 57647 10746 57649 10753
rect 57593 10697 57649 10746
rect 57381 10529 57383 10535
rect 57383 10529 57435 10535
rect 57435 10529 57437 10535
rect 57381 10479 57437 10529
rect 57593 10529 57595 10535
rect 57595 10529 57647 10535
rect 57647 10529 57649 10535
rect 57593 10479 57649 10529
rect 57381 10311 57383 10318
rect 57383 10311 57435 10318
rect 57435 10311 57437 10318
rect 57381 10262 57437 10311
rect 57593 10311 57595 10318
rect 57595 10311 57647 10318
rect 57647 10311 57649 10318
rect 57593 10262 57649 10311
rect 51766 9811 51822 9971
rect 49897 8897 50057 8953
rect 27474 7534 27530 7535
rect 27474 7482 27476 7534
rect 27476 7482 27528 7534
rect 27528 7482 27530 7534
rect 27474 7479 27530 7482
rect 27686 7534 27742 7535
rect 27686 7482 27688 7534
rect 27688 7482 27740 7534
rect 27740 7482 27742 7534
rect 27686 7479 27742 7482
rect 27474 7316 27530 7317
rect 27474 7264 27476 7316
rect 27476 7264 27528 7316
rect 27528 7264 27530 7316
rect 27474 7261 27530 7264
rect 27686 7316 27742 7317
rect 27686 7264 27688 7316
rect 27688 7264 27740 7316
rect 27740 7264 27742 7316
rect 27686 7261 27742 7264
rect 27474 7047 27476 7099
rect 27476 7047 27528 7099
rect 27528 7047 27530 7099
rect 27474 7043 27530 7047
rect 27686 7047 27688 7099
rect 27688 7047 27740 7099
rect 27740 7047 27742 7099
rect 27686 7043 27742 7047
rect 28273 6780 28329 6836
rect 28484 6780 28540 6836
rect 28696 6780 28752 6836
rect 28907 6780 28963 6836
rect 28273 6562 28329 6618
rect 28484 6562 28540 6618
rect 28696 6562 28752 6618
rect 28907 6562 28963 6618
rect 28273 6344 28329 6400
rect 28484 6344 28540 6400
rect 28696 6344 28752 6400
rect 28907 6344 28963 6400
rect 27474 6064 27530 6120
rect 27686 6064 27742 6120
rect 27474 5846 27530 5902
rect 27686 5846 27742 5902
rect 26859 4472 26915 4528
rect 27071 4472 27127 4528
rect 26859 4254 26915 4310
rect 27071 4254 27127 4310
rect 27474 3781 27530 3837
rect 27686 3781 27742 3837
rect 27474 3563 27530 3619
rect 27686 3563 27742 3619
rect 28801 3781 28857 3837
rect 28801 3563 28857 3619
rect 43800 2994 43960 3050
rect 57381 8840 57437 8843
rect 57381 8788 57383 8840
rect 57383 8788 57435 8840
rect 57435 8788 57437 8840
rect 57381 8787 57437 8788
rect 57593 8840 57649 8843
rect 57593 8788 57595 8840
rect 57595 8788 57647 8840
rect 57647 8788 57649 8840
rect 57593 8787 57649 8788
rect 57381 8622 57437 8625
rect 57381 8570 57383 8622
rect 57383 8570 57435 8622
rect 57435 8570 57437 8622
rect 57381 8569 57437 8570
rect 57593 8622 57649 8625
rect 57593 8570 57595 8622
rect 57595 8570 57647 8622
rect 57647 8570 57649 8622
rect 57593 8569 57649 8570
rect 57381 8404 57437 8408
rect 57381 8352 57383 8404
rect 57383 8352 57435 8404
rect 57435 8352 57437 8404
rect 57593 8404 57649 8408
rect 57593 8352 57595 8404
rect 57595 8352 57647 8404
rect 57647 8352 57649 8404
rect 57381 8187 57437 8190
rect 57381 8135 57383 8187
rect 57383 8135 57435 8187
rect 57435 8135 57437 8187
rect 57381 8134 57437 8135
rect 57593 8187 57649 8190
rect 57593 8135 57595 8187
rect 57595 8135 57647 8187
rect 57647 8135 57649 8187
rect 57593 8134 57649 8135
rect 57381 7969 57437 7972
rect 57381 7917 57383 7969
rect 57383 7917 57435 7969
rect 57435 7917 57437 7969
rect 57381 7916 57437 7917
rect 57593 7969 57649 7972
rect 57593 7917 57595 7969
rect 57595 7917 57647 7969
rect 57647 7917 57649 7969
rect 57593 7916 57649 7917
rect 57381 7752 57437 7755
rect 57381 7700 57383 7752
rect 57383 7700 57435 7752
rect 57435 7700 57437 7752
rect 57381 7699 57437 7700
rect 57593 7752 57649 7755
rect 57593 7700 57595 7752
rect 57595 7700 57647 7752
rect 57647 7700 57649 7752
rect 57593 7699 57649 7700
rect 57381 7534 57437 7537
rect 57381 7482 57383 7534
rect 57383 7482 57435 7534
rect 57435 7482 57437 7534
rect 57381 7481 57437 7482
rect 57593 7534 57649 7537
rect 57593 7482 57595 7534
rect 57595 7482 57647 7534
rect 57647 7482 57649 7534
rect 57593 7481 57649 7482
rect 57381 7316 57437 7319
rect 57381 7264 57383 7316
rect 57383 7264 57435 7316
rect 57435 7264 57437 7316
rect 57381 7263 57437 7264
rect 57593 7316 57649 7319
rect 57593 7264 57595 7316
rect 57595 7264 57647 7316
rect 57647 7264 57649 7316
rect 57593 7263 57649 7264
rect 57381 7099 57437 7102
rect 57381 7047 57383 7099
rect 57383 7047 57435 7099
rect 57435 7047 57437 7099
rect 57381 7046 57437 7047
rect 57593 7099 57649 7102
rect 57593 7047 57595 7099
rect 57595 7047 57647 7099
rect 57647 7047 57649 7099
rect 57593 7046 57649 7047
rect 56160 6780 56216 6836
rect 56371 6780 56427 6836
rect 56583 6780 56639 6836
rect 56794 6780 56850 6836
rect 56160 6562 56216 6618
rect 56371 6562 56427 6618
rect 56583 6562 56639 6618
rect 56794 6562 56850 6618
rect 56160 6344 56216 6400
rect 56371 6344 56427 6400
rect 56583 6344 56639 6400
rect 56794 6344 56850 6400
rect 57381 6064 57437 6120
rect 57593 6064 57649 6120
rect 57381 5846 57437 5902
rect 57593 5846 57649 5902
rect 57381 3781 57437 3837
rect 57593 3781 57649 3837
rect 57381 3563 57437 3619
rect 57593 3563 57649 3619
rect 57996 33302 58052 33358
rect 58208 33302 58264 33358
rect 57996 33084 58052 33140
rect 58208 33084 58264 33140
rect 57996 32866 58052 32922
rect 58208 32866 58264 32922
rect 57996 32649 58052 32705
rect 58208 32649 58264 32705
rect 57996 32431 58052 32487
rect 58208 32431 58264 32487
rect 57996 32075 57998 32088
rect 57998 32075 58050 32088
rect 58050 32075 58052 32088
rect 57996 32032 58052 32075
rect 58208 32075 58210 32088
rect 58210 32075 58262 32088
rect 58262 32075 58264 32088
rect 58208 32032 58264 32075
rect 57996 31857 57998 31870
rect 57998 31857 58050 31870
rect 58050 31857 58052 31870
rect 57996 31814 58052 31857
rect 58208 31857 58210 31870
rect 58210 31857 58262 31870
rect 58262 31857 58264 31870
rect 58208 31814 58264 31857
rect 57996 31639 57998 31652
rect 57998 31639 58050 31652
rect 58050 31639 58052 31652
rect 57996 31596 58052 31639
rect 58208 31639 58210 31652
rect 58210 31639 58262 31652
rect 58262 31639 58264 31652
rect 58208 31596 58264 31639
rect 57996 29950 58052 29968
rect 57996 29912 57998 29950
rect 57998 29912 58050 29950
rect 58050 29912 58052 29950
rect 58208 29950 58264 29968
rect 58208 29912 58210 29950
rect 58210 29912 58262 29950
rect 58262 29912 58264 29950
rect 57996 29733 58052 29750
rect 57996 29694 57998 29733
rect 57998 29694 58050 29733
rect 58050 29694 58052 29733
rect 58208 29733 58264 29750
rect 58208 29694 58210 29733
rect 58210 29694 58262 29733
rect 58262 29694 58264 29733
rect 57996 29515 58052 29533
rect 57996 29477 57998 29515
rect 57998 29477 58050 29515
rect 58050 29477 58052 29515
rect 58208 29515 58264 29533
rect 58208 29477 58210 29515
rect 58210 29477 58262 29515
rect 58262 29477 58264 29515
rect 57996 29297 58052 29315
rect 57996 29259 57998 29297
rect 57998 29259 58050 29297
rect 58050 29259 58052 29297
rect 58208 29297 58264 29315
rect 58208 29259 58210 29297
rect 58210 29259 58262 29297
rect 58262 29259 58264 29297
rect 57996 29080 58052 29098
rect 57996 29042 57998 29080
rect 57998 29042 58050 29080
rect 58050 29042 58052 29080
rect 58208 29080 58264 29098
rect 58208 29042 58210 29080
rect 58210 29042 58262 29080
rect 58262 29042 58264 29080
rect 57996 28862 58052 28880
rect 57996 28824 57998 28862
rect 57998 28824 58050 28862
rect 58050 28824 58052 28862
rect 58208 28862 58264 28880
rect 58208 28824 58210 28862
rect 58210 28824 58262 28862
rect 58262 28824 58264 28862
rect 57996 28644 58052 28662
rect 57996 28606 57998 28644
rect 57998 28606 58050 28644
rect 58050 28606 58052 28644
rect 58208 28644 58264 28662
rect 58208 28606 58210 28644
rect 58210 28606 58262 28644
rect 58262 28606 58264 28644
rect 57996 28427 58052 28444
rect 57996 28388 57998 28427
rect 57998 28388 58050 28427
rect 58050 28388 58052 28427
rect 58208 28427 58264 28444
rect 58208 28388 58210 28427
rect 58210 28388 58262 28427
rect 58262 28388 58264 28427
rect 57996 28209 58052 28227
rect 57996 28171 57998 28209
rect 57998 28171 58050 28209
rect 58050 28171 58052 28209
rect 58208 28209 58264 28227
rect 58208 28171 58210 28209
rect 58210 28171 58262 28209
rect 58262 28171 58264 28209
rect 57996 27992 58052 28009
rect 57996 27953 57998 27992
rect 57998 27953 58050 27992
rect 58050 27953 58052 27992
rect 58208 27992 58264 28009
rect 58208 27953 58210 27992
rect 58210 27953 58262 27992
rect 58262 27953 58264 27992
rect 57996 27774 58052 27792
rect 57996 27736 57998 27774
rect 57998 27736 58050 27774
rect 58050 27736 58052 27774
rect 58208 27774 58264 27792
rect 58208 27736 58210 27774
rect 58210 27736 58262 27774
rect 58262 27736 58264 27774
rect 57996 27556 58052 27574
rect 57996 27518 57998 27556
rect 57998 27518 58050 27556
rect 58050 27518 58052 27556
rect 58208 27556 58264 27574
rect 58208 27518 58210 27556
rect 58210 27518 58262 27556
rect 58262 27518 58264 27556
rect 58865 94773 58921 94775
rect 58865 94721 58867 94773
rect 58867 94721 58919 94773
rect 58919 94721 58921 94773
rect 58865 94719 58921 94721
rect 58989 94773 59045 94775
rect 58989 94721 58991 94773
rect 58991 94721 59043 94773
rect 59043 94721 59045 94773
rect 58989 94719 59045 94721
rect 59113 94773 59169 94775
rect 59113 94721 59115 94773
rect 59115 94721 59167 94773
rect 59167 94721 59169 94773
rect 59113 94719 59169 94721
rect 59237 94773 59293 94775
rect 59237 94721 59239 94773
rect 59239 94721 59291 94773
rect 59291 94721 59293 94773
rect 59237 94719 59293 94721
rect 59361 94773 59417 94775
rect 59361 94721 59363 94773
rect 59363 94721 59415 94773
rect 59415 94721 59417 94773
rect 59361 94719 59417 94721
rect 58865 94649 58921 94651
rect 58865 94597 58867 94649
rect 58867 94597 58919 94649
rect 58919 94597 58921 94649
rect 58865 94595 58921 94597
rect 58989 94649 59045 94651
rect 58989 94597 58991 94649
rect 58991 94597 59043 94649
rect 59043 94597 59045 94649
rect 58989 94595 59045 94597
rect 59113 94649 59169 94651
rect 59113 94597 59115 94649
rect 59115 94597 59167 94649
rect 59167 94597 59169 94649
rect 59113 94595 59169 94597
rect 59237 94649 59293 94651
rect 59237 94597 59239 94649
rect 59239 94597 59291 94649
rect 59291 94597 59293 94649
rect 59237 94595 59293 94597
rect 59361 94649 59417 94651
rect 59361 94597 59363 94649
rect 59363 94597 59415 94649
rect 59415 94597 59417 94649
rect 59361 94595 59417 94597
rect 58865 94525 58921 94527
rect 58865 94473 58867 94525
rect 58867 94473 58919 94525
rect 58919 94473 58921 94525
rect 58865 94471 58921 94473
rect 58989 94525 59045 94527
rect 58989 94473 58991 94525
rect 58991 94473 59043 94525
rect 59043 94473 59045 94525
rect 58989 94471 59045 94473
rect 59113 94525 59169 94527
rect 59113 94473 59115 94525
rect 59115 94473 59167 94525
rect 59167 94473 59169 94525
rect 59113 94471 59169 94473
rect 59237 94525 59293 94527
rect 59237 94473 59239 94525
rect 59239 94473 59291 94525
rect 59291 94473 59293 94525
rect 59237 94471 59293 94473
rect 59361 94525 59417 94527
rect 59361 94473 59363 94525
rect 59363 94473 59415 94525
rect 59415 94473 59417 94525
rect 59361 94471 59417 94473
rect 58816 34936 58872 34992
rect 58940 34936 58996 34992
rect 59064 34936 59120 34992
rect 59188 34936 59244 34992
rect 59312 34936 59368 34992
rect 59436 34936 59492 34992
rect 58816 34812 58872 34868
rect 58940 34812 58996 34868
rect 59064 34812 59120 34868
rect 59188 34812 59244 34868
rect 59312 34812 59368 34868
rect 59436 34812 59492 34868
rect 58816 34688 58872 34744
rect 58940 34688 58996 34744
rect 59064 34688 59120 34744
rect 59188 34688 59244 34744
rect 59312 34688 59368 34744
rect 59436 34688 59492 34744
rect 58816 34564 58872 34620
rect 58940 34564 58996 34620
rect 59064 34564 59120 34620
rect 59188 34564 59244 34620
rect 59312 34564 59368 34620
rect 59436 34564 59492 34620
rect 58873 31242 58929 31298
rect 58997 31242 59053 31298
rect 59121 31242 59177 31298
rect 59245 31242 59301 31298
rect 59369 31242 59425 31298
rect 58873 31118 58929 31174
rect 58997 31118 59053 31174
rect 59121 31118 59177 31174
rect 59245 31118 59301 31174
rect 59369 31118 59425 31174
rect 58873 30994 58929 31050
rect 58997 30994 59053 31050
rect 59121 30994 59177 31050
rect 59245 30994 59301 31050
rect 59369 30994 59425 31050
rect 58873 30797 58929 30853
rect 58997 30797 59053 30853
rect 59121 30797 59177 30853
rect 59245 30797 59301 30853
rect 59369 30797 59425 30853
rect 58873 30673 58929 30729
rect 58997 30673 59053 30729
rect 59121 30673 59177 30729
rect 59245 30673 59301 30729
rect 59369 30673 59425 30729
rect 58873 30549 58929 30605
rect 58997 30549 59053 30605
rect 59121 30549 59177 30605
rect 59245 30549 59301 30605
rect 59369 30549 59425 30605
rect 58859 28239 58915 28295
rect 58983 28239 59039 28295
rect 59107 28239 59163 28295
rect 59231 28239 59287 28295
rect 59355 28239 59411 28295
rect 58859 28115 58915 28171
rect 58983 28115 59039 28171
rect 59107 28115 59163 28171
rect 59231 28115 59287 28171
rect 59355 28115 59411 28171
rect 58859 27991 58915 28047
rect 58983 27991 59039 28047
rect 59107 27991 59163 28047
rect 59231 27991 59287 28047
rect 59355 27991 59411 28047
rect 58859 27867 58915 27923
rect 58983 27867 59039 27923
rect 59107 27867 59163 27923
rect 59231 27867 59287 27923
rect 59355 27867 59411 27923
rect 58859 27743 58915 27799
rect 58983 27743 59039 27799
rect 59107 27743 59163 27799
rect 59231 27743 59287 27799
rect 59355 27743 59411 27799
rect 58859 27619 58915 27675
rect 58983 27619 59039 27675
rect 59107 27619 59163 27675
rect 59231 27619 59287 27675
rect 59355 27619 59411 27675
rect 58859 27495 58915 27551
rect 58983 27495 59039 27551
rect 59107 27495 59163 27551
rect 59231 27495 59287 27551
rect 59355 27495 59411 27551
rect 58859 27371 58915 27427
rect 58983 27371 59039 27427
rect 59107 27371 59163 27427
rect 59231 27371 59287 27427
rect 59355 27371 59411 27427
rect 58859 27247 58915 27303
rect 58983 27247 59039 27303
rect 59107 27247 59163 27303
rect 59231 27247 59287 27303
rect 59355 27247 59411 27303
rect 58859 27123 58915 27179
rect 58983 27123 59039 27179
rect 59107 27123 59163 27179
rect 59231 27123 59287 27179
rect 59355 27123 59411 27179
rect 58859 26999 58915 27055
rect 58983 26999 59039 27055
rect 59107 26999 59163 27055
rect 59231 26999 59287 27055
rect 59355 26999 59411 27055
rect 58859 26875 58915 26931
rect 58983 26875 59039 26931
rect 59107 26875 59163 26931
rect 59231 26875 59287 26931
rect 59355 26875 59411 26931
rect 58859 26751 58915 26807
rect 58983 26751 59039 26807
rect 59107 26751 59163 26807
rect 59231 26751 59287 26807
rect 59355 26751 59411 26807
rect 58859 26627 58915 26683
rect 58983 26627 59039 26683
rect 59107 26627 59163 26683
rect 59231 26627 59287 26683
rect 59355 26627 59411 26683
rect 58859 26503 58915 26559
rect 58983 26503 59039 26559
rect 59107 26503 59163 26559
rect 59231 26503 59287 26559
rect 59355 26503 59411 26559
rect 57994 24074 58258 24075
rect 57994 24022 57998 24074
rect 57998 24022 58050 24074
rect 58050 24022 58210 24074
rect 58210 24022 58258 24074
rect 57994 23857 58258 24022
rect 57994 23805 57998 23857
rect 57998 23805 58050 23857
rect 58050 23805 58210 23857
rect 58210 23805 58258 23857
rect 57994 23639 58258 23805
rect 57994 23587 57998 23639
rect 57998 23587 58050 23639
rect 58050 23587 58210 23639
rect 58210 23587 58258 23639
rect 57994 23421 58258 23587
rect 57994 23369 57998 23421
rect 57998 23369 58050 23421
rect 58050 23369 58210 23421
rect 58210 23369 58258 23421
rect 57994 23204 58258 23369
rect 57994 23187 57998 23204
rect 57998 23187 58050 23204
rect 58050 23187 58210 23204
rect 58210 23187 58258 23204
rect 58048 20540 58050 20570
rect 58050 20540 58208 20570
rect 58048 20410 58208 20540
rect 58048 20157 58208 20226
rect 58048 20105 58050 20157
rect 58050 20105 58208 20157
rect 58048 20066 58208 20105
rect 57996 13734 58052 13790
rect 58208 13734 58264 13790
rect 57996 13517 58052 13573
rect 58208 13517 58264 13573
rect 57996 13299 58052 13355
rect 58208 13299 58264 13355
rect 57996 13082 58052 13138
rect 58208 13082 58264 13138
rect 57996 12864 58052 12920
rect 58208 12864 58264 12920
rect 57996 12646 58052 12702
rect 58208 12646 58264 12702
rect 57996 12428 58052 12484
rect 58208 12428 58264 12484
rect 57996 12211 58052 12267
rect 58208 12211 58264 12267
rect 57996 11993 58052 12049
rect 58208 11993 58264 12049
rect 57996 11776 58052 11832
rect 58208 11776 58264 11832
rect 57996 9351 58052 9407
rect 58208 9351 58264 9407
rect 57996 9134 58052 9190
rect 58208 9134 58264 9190
rect 57996 8916 58052 8972
rect 58208 8916 58264 8972
rect 57996 8698 58052 8754
rect 58208 8698 58264 8754
rect 57996 8480 58052 8536
rect 58208 8480 58264 8536
rect 57996 8263 58052 8319
rect 58208 8263 58264 8319
rect 57996 5523 57998 5539
rect 57998 5523 58050 5539
rect 58050 5523 58052 5539
rect 57996 5483 58052 5523
rect 58208 5523 58210 5539
rect 58210 5523 58262 5539
rect 58262 5523 58264 5539
rect 58208 5483 58264 5523
rect 57996 5306 57998 5321
rect 57998 5306 58050 5321
rect 58050 5306 58052 5321
rect 57996 5265 58052 5306
rect 58208 5306 58210 5321
rect 58210 5306 58262 5321
rect 58262 5306 58264 5321
rect 58208 5265 58264 5306
rect 57996 4472 58052 4528
rect 58208 4472 58264 4528
rect 57996 4254 58052 4310
rect 58208 4254 58264 4310
<< metal3 >>
rect 1401 96176 2401 96976
rect 2626 96368 3626 96976
rect 4137 96176 5137 96976
rect 5362 96368 6362 96976
rect 6801 96176 7801 96976
rect 8026 96368 9026 96976
rect 9537 96176 10537 96976
rect 10762 96368 11762 96976
rect 12201 96176 13201 96976
rect 13426 96368 14426 96976
rect 14937 96176 15937 96976
rect 16162 96368 17162 96976
rect 17601 96176 18601 96976
rect 18826 96368 19826 96976
rect 20653 96176 21653 96976
rect 22258 96368 23258 96976
rect 23483 96176 24483 96976
rect 25158 96368 26158 96976
rect 26572 96176 27572 96976
rect 27877 96368 28877 96976
rect 29273 96368 30273 96976
rect 30710 96176 31710 96976
rect 32381 96368 33381 96976
rect 34024 96368 35024 96976
rect 35415 96176 36415 96976
rect 36948 96368 37948 96976
rect 38585 96176 39585 96976
rect 39882 96368 40882 96976
rect 41230 96176 42230 96976
rect 42430 96368 43430 96976
rect 43713 96368 44713 96976
rect 45069 96176 46069 96976
rect 46313 96176 47313 96976
rect 47538 96368 48538 96976
rect 48901 96176 49901 96976
rect 50465 96368 51465 96976
rect 52569 96176 53569 96976
rect 54262 96176 55262 96976
rect 55990 96368 56990 96976
rect 57547 96176 58547 96976
rect 58791 96368 59791 96976
rect 60977 96176 61977 96976
rect 62202 96368 63202 96976
rect 63713 96176 64713 96976
rect 64938 96368 65938 96976
rect 66377 96176 67377 96976
rect 67602 96368 68602 96976
rect 69113 96176 70113 96976
rect 70338 96368 71338 96976
rect 71777 96176 72777 96976
rect 73002 96368 74002 96976
rect 74513 96176 75513 96976
rect 75738 96368 76738 96976
rect 77177 96176 78177 96976
rect 78402 96368 79402 96976
rect 80229 96176 81229 96976
rect 81834 96368 82834 96976
rect 83059 96176 84059 96976
rect 84666 96176 85666 96976
rect 0 95176 86372 96176
rect 0 94776 1014 94976
rect 25376 94776 25948 94785
rect 58855 94776 59427 94785
rect 85358 94776 86372 94976
rect 0 94775 27272 94776
rect 0 94719 25386 94775
rect 25442 94719 25510 94775
rect 25566 94719 25634 94775
rect 25690 94719 25758 94775
rect 25814 94719 25882 94775
rect 25938 94728 27272 94775
rect 58855 94775 86372 94776
rect 58855 94728 58865 94775
rect 25938 94719 58865 94728
rect 58921 94719 58989 94775
rect 59045 94719 59113 94775
rect 59169 94719 59237 94775
rect 59293 94719 59361 94775
rect 59417 94719 86372 94775
rect 0 94655 86372 94719
rect 0 94651 27788 94655
rect 0 94595 25386 94651
rect 25442 94595 25510 94651
rect 25566 94595 25634 94651
rect 25690 94595 25758 94651
rect 25814 94595 25882 94651
rect 25938 94599 27788 94651
rect 27844 94599 27999 94655
rect 28055 94599 28210 94655
rect 28266 94599 28421 94655
rect 28477 94599 28632 94655
rect 28688 94599 28843 94655
rect 28899 94599 29054 94655
rect 29110 94599 56013 94655
rect 56069 94599 56224 94655
rect 56280 94599 56435 94655
rect 56491 94599 56646 94655
rect 56702 94599 56857 94655
rect 56913 94599 57068 94655
rect 57124 94599 57279 94655
rect 57335 94651 86372 94655
rect 57335 94599 58865 94651
rect 25938 94595 58865 94599
rect 58921 94595 58989 94651
rect 59045 94595 59113 94651
rect 59169 94595 59237 94651
rect 59293 94595 59361 94651
rect 59417 94595 86372 94651
rect 0 94527 86372 94595
rect 0 94476 25386 94527
rect 0 94276 1014 94476
rect 25376 94471 25386 94476
rect 25442 94471 25510 94527
rect 25566 94471 25634 94527
rect 25690 94471 25758 94527
rect 25814 94471 25882 94527
rect 25938 94476 27272 94527
rect 30402 94526 54622 94527
rect 25938 94471 25948 94476
rect 25376 94461 25948 94471
rect 58855 94471 58865 94527
rect 58921 94471 58989 94527
rect 59045 94471 59113 94527
rect 59169 94471 59237 94527
rect 59293 94471 59361 94527
rect 59417 94476 86372 94527
rect 59417 94471 59427 94476
rect 58855 94461 59427 94471
rect 85358 94276 86372 94476
rect 0 93376 1706 94076
rect 56271 94066 61644 94268
rect 84666 93376 86372 94076
rect 0 92976 1014 93176
rect 85358 92976 86372 93176
rect 0 92928 27272 92976
rect 59421 92928 86372 92976
rect 0 92855 86372 92928
rect 0 92799 27788 92855
rect 27844 92799 27999 92855
rect 28055 92799 28210 92855
rect 28266 92799 28421 92855
rect 28477 92799 28632 92855
rect 28688 92799 28843 92855
rect 28899 92799 29054 92855
rect 29110 92799 56013 92855
rect 56069 92799 56224 92855
rect 56280 92799 56435 92855
rect 56491 92799 56646 92855
rect 56702 92799 56857 92855
rect 56913 92799 57068 92855
rect 57124 92799 57279 92855
rect 57335 92799 86372 92855
rect 0 92727 86372 92799
rect 0 92676 27272 92727
rect 30403 92726 54622 92727
rect 59421 92676 86372 92727
rect 0 92476 1014 92676
rect 85358 92476 86372 92676
rect 0 91576 1706 92276
rect 84666 91576 86372 92276
rect 0 91176 1014 91376
rect 85358 91176 86372 91376
rect 0 91128 27272 91176
rect 59421 91128 86372 91176
rect 0 91055 86372 91128
rect 0 90999 27788 91055
rect 27844 90999 27999 91055
rect 28055 90999 28210 91055
rect 28266 90999 28421 91055
rect 28477 90999 28632 91055
rect 28688 90999 28843 91055
rect 28899 90999 29054 91055
rect 29110 90999 56013 91055
rect 56069 90999 56224 91055
rect 56280 90999 56435 91055
rect 56491 90999 56646 91055
rect 56702 90999 56857 91055
rect 56913 90999 57068 91055
rect 57124 90999 57279 91055
rect 57335 90999 86372 91055
rect 0 90927 86372 90999
rect 0 90876 27272 90927
rect 30403 90926 54622 90927
rect 59421 90876 86372 90927
rect 0 90676 1014 90876
rect 85358 90676 86372 90876
rect 0 89776 1706 90476
rect 84666 89776 86372 90476
rect 0 89376 1014 89576
rect 85358 89376 86372 89576
rect 0 89328 27272 89376
rect 59421 89328 86372 89376
rect 0 89255 86372 89328
rect 0 89199 27788 89255
rect 27844 89199 27999 89255
rect 28055 89199 28210 89255
rect 28266 89199 28421 89255
rect 28477 89199 28632 89255
rect 28688 89199 28843 89255
rect 28899 89199 29054 89255
rect 29110 89199 56013 89255
rect 56069 89199 56224 89255
rect 56280 89199 56435 89255
rect 56491 89199 56646 89255
rect 56702 89199 56857 89255
rect 56913 89199 57068 89255
rect 57124 89199 57279 89255
rect 57335 89199 86372 89255
rect 0 89127 86372 89199
rect 0 89076 27272 89127
rect 30403 89126 54622 89127
rect 59421 89076 86372 89127
rect 0 88876 1014 89076
rect 85358 88876 86372 89076
rect 0 87976 1706 88676
rect 84666 87976 86372 88676
rect 0 87576 1014 87776
rect 85358 87576 86372 87776
rect 0 87528 27272 87576
rect 59421 87528 86372 87576
rect 0 87455 86372 87528
rect 0 87399 27788 87455
rect 27844 87399 27999 87455
rect 28055 87399 28210 87455
rect 28266 87399 28421 87455
rect 28477 87399 28632 87455
rect 28688 87399 28843 87455
rect 28899 87399 29054 87455
rect 29110 87399 56013 87455
rect 56069 87399 56224 87455
rect 56280 87399 56435 87455
rect 56491 87399 56646 87455
rect 56702 87399 56857 87455
rect 56913 87399 57068 87455
rect 57124 87399 57279 87455
rect 57335 87399 86372 87455
rect 0 87327 86372 87399
rect 0 87276 27272 87327
rect 30403 87326 54622 87327
rect 59421 87276 86372 87327
rect 0 87076 1014 87276
rect 85358 87076 86372 87276
rect 0 86176 1706 86876
rect 84666 86176 86372 86876
rect 0 85776 1014 85976
rect 85358 85776 86372 85976
rect 0 85728 27272 85776
rect 59421 85728 86372 85776
rect 0 85655 86372 85728
rect 0 85599 27788 85655
rect 27844 85599 27999 85655
rect 28055 85599 28210 85655
rect 28266 85599 28421 85655
rect 28477 85599 28632 85655
rect 28688 85599 28843 85655
rect 28899 85599 29054 85655
rect 29110 85599 56013 85655
rect 56069 85599 56224 85655
rect 56280 85599 56435 85655
rect 56491 85599 56646 85655
rect 56702 85599 56857 85655
rect 56913 85599 57068 85655
rect 57124 85599 57279 85655
rect 57335 85599 86372 85655
rect 0 85527 86372 85599
rect 0 85476 27272 85527
rect 30403 85526 54622 85527
rect 59421 85476 86372 85527
rect 0 85276 1014 85476
rect 85358 85276 86372 85476
rect 0 84376 1706 85076
rect 84666 84376 86372 85076
rect 0 83976 1014 84176
rect 85358 83976 86372 84176
rect 0 83928 27272 83976
rect 59421 83928 86372 83976
rect 0 83855 86372 83928
rect 0 83799 27788 83855
rect 27844 83799 27999 83855
rect 28055 83799 28210 83855
rect 28266 83799 28421 83855
rect 28477 83799 28632 83855
rect 28688 83799 28843 83855
rect 28899 83799 29054 83855
rect 29110 83799 56013 83855
rect 56069 83799 56224 83855
rect 56280 83799 56435 83855
rect 56491 83799 56646 83855
rect 56702 83799 56857 83855
rect 56913 83799 57068 83855
rect 57124 83799 57279 83855
rect 57335 83799 86372 83855
rect 0 83727 86372 83799
rect 0 83676 27272 83727
rect 30403 83726 54622 83727
rect 59421 83676 86372 83727
rect 0 83476 1014 83676
rect 85358 83476 86372 83676
rect 0 82576 1706 83276
rect 84666 82576 86372 83276
rect 0 82176 1014 82376
rect 85358 82176 86372 82376
rect 0 82128 27272 82176
rect 59421 82128 86372 82176
rect 0 82055 86372 82128
rect 0 81999 27788 82055
rect 27844 81999 27999 82055
rect 28055 81999 28210 82055
rect 28266 81999 28421 82055
rect 28477 81999 28632 82055
rect 28688 81999 28843 82055
rect 28899 81999 29054 82055
rect 29110 81999 56013 82055
rect 56069 81999 56224 82055
rect 56280 81999 56435 82055
rect 56491 81999 56646 82055
rect 56702 81999 56857 82055
rect 56913 81999 57068 82055
rect 57124 81999 57279 82055
rect 57335 81999 86372 82055
rect 0 81927 86372 81999
rect 0 81876 27272 81927
rect 30403 81926 54622 81927
rect 59421 81876 86372 81927
rect 0 81676 1014 81876
rect 85358 81676 86372 81876
rect 0 80776 1706 81476
rect 84666 80776 86372 81476
rect 0 80376 1014 80576
rect 85358 80376 86372 80576
rect 0 80328 27272 80376
rect 59421 80328 86372 80376
rect 0 80255 86372 80328
rect 0 80199 27788 80255
rect 27844 80199 27999 80255
rect 28055 80199 28210 80255
rect 28266 80199 28421 80255
rect 28477 80199 28632 80255
rect 28688 80199 28843 80255
rect 28899 80199 29054 80255
rect 29110 80199 56013 80255
rect 56069 80199 56224 80255
rect 56280 80199 56435 80255
rect 56491 80199 56646 80255
rect 56702 80199 56857 80255
rect 56913 80199 57068 80255
rect 57124 80199 57279 80255
rect 57335 80199 86372 80255
rect 0 80127 86372 80199
rect 0 80076 27272 80127
rect 30403 80126 54622 80127
rect 59421 80076 86372 80127
rect 0 79876 1014 80076
rect 85358 79876 86372 80076
rect 0 78976 1706 79676
rect 84666 78976 86372 79676
rect 0 78576 1014 78776
rect 85358 78576 86372 78776
rect 0 78528 27272 78576
rect 59421 78528 86372 78576
rect 0 78455 86372 78528
rect 0 78399 27788 78455
rect 27844 78399 27999 78455
rect 28055 78399 28210 78455
rect 28266 78399 28421 78455
rect 28477 78399 28632 78455
rect 28688 78399 28843 78455
rect 28899 78399 29054 78455
rect 29110 78399 56013 78455
rect 56069 78399 56224 78455
rect 56280 78399 56435 78455
rect 56491 78399 56646 78455
rect 56702 78399 56857 78455
rect 56913 78399 57068 78455
rect 57124 78399 57279 78455
rect 57335 78399 86372 78455
rect 0 78327 86372 78399
rect 0 78276 27272 78327
rect 30403 78326 54622 78327
rect 59421 78276 86372 78327
rect 0 78076 1014 78276
rect 85358 78076 86372 78276
rect 0 77176 1706 77876
rect 84666 77176 86372 77876
rect 0 76776 1014 76976
rect 85358 76776 86372 76976
rect 0 76728 27272 76776
rect 59421 76728 86372 76776
rect 0 76655 86372 76728
rect 0 76599 27788 76655
rect 27844 76599 27999 76655
rect 28055 76599 28210 76655
rect 28266 76599 28421 76655
rect 28477 76599 28632 76655
rect 28688 76599 28843 76655
rect 28899 76599 29054 76655
rect 29110 76599 56013 76655
rect 56069 76599 56224 76655
rect 56280 76599 56435 76655
rect 56491 76599 56646 76655
rect 56702 76599 56857 76655
rect 56913 76599 57068 76655
rect 57124 76599 57279 76655
rect 57335 76599 86372 76655
rect 0 76527 86372 76599
rect 0 76476 27272 76527
rect 30403 76526 54622 76527
rect 59421 76476 86372 76527
rect 0 76276 1014 76476
rect 85358 76276 86372 76476
rect 0 75376 1706 76076
rect 84666 75376 86372 76076
rect 0 74976 1014 75176
rect 85358 74976 86372 75176
rect 0 74928 27272 74976
rect 59421 74928 86372 74976
rect 0 74855 86372 74928
rect 0 74799 27788 74855
rect 27844 74799 27999 74855
rect 28055 74799 28210 74855
rect 28266 74799 28421 74855
rect 28477 74799 28632 74855
rect 28688 74799 28843 74855
rect 28899 74799 29054 74855
rect 29110 74799 56013 74855
rect 56069 74799 56224 74855
rect 56280 74799 56435 74855
rect 56491 74799 56646 74855
rect 56702 74799 56857 74855
rect 56913 74799 57068 74855
rect 57124 74799 57279 74855
rect 57335 74799 86372 74855
rect 0 74727 86372 74799
rect 0 74676 27272 74727
rect 30403 74726 54622 74727
rect 59421 74676 86372 74727
rect 0 74476 1014 74676
rect 85358 74476 86372 74676
rect 0 73576 1706 74276
rect 84666 73576 86372 74276
rect 0 73176 1014 73376
rect 85358 73176 86372 73376
rect 0 73128 27272 73176
rect 59421 73128 86372 73176
rect 0 73055 86372 73128
rect 0 72999 27788 73055
rect 27844 72999 27999 73055
rect 28055 72999 28210 73055
rect 28266 72999 28421 73055
rect 28477 72999 28632 73055
rect 28688 72999 28843 73055
rect 28899 72999 29054 73055
rect 29110 72999 56013 73055
rect 56069 72999 56224 73055
rect 56280 72999 56435 73055
rect 56491 72999 56646 73055
rect 56702 72999 56857 73055
rect 56913 72999 57068 73055
rect 57124 72999 57279 73055
rect 57335 72999 86372 73055
rect 0 72927 86372 72999
rect 0 72876 27272 72927
rect 30403 72926 54622 72927
rect 59421 72876 86372 72927
rect 0 72676 1014 72876
rect 85358 72676 86372 72876
rect 0 71776 1706 72476
rect 84666 71776 86372 72476
rect 0 71376 1014 71576
rect 85358 71376 86372 71576
rect 0 71328 27272 71376
rect 59421 71328 86372 71376
rect 0 71255 86372 71328
rect 0 71199 27788 71255
rect 27844 71199 27999 71255
rect 28055 71199 28210 71255
rect 28266 71199 28421 71255
rect 28477 71199 28632 71255
rect 28688 71199 28843 71255
rect 28899 71199 29054 71255
rect 29110 71199 56013 71255
rect 56069 71199 56224 71255
rect 56280 71199 56435 71255
rect 56491 71199 56646 71255
rect 56702 71199 56857 71255
rect 56913 71199 57068 71255
rect 57124 71199 57279 71255
rect 57335 71199 86372 71255
rect 0 71127 86372 71199
rect 0 71076 27272 71127
rect 30403 71126 54622 71127
rect 59421 71076 86372 71127
rect 0 70876 1014 71076
rect 85358 70876 86372 71076
rect 0 69976 1706 70676
rect 84666 69976 86372 70676
rect 0 69576 1014 69776
rect 85358 69576 86372 69776
rect 0 69528 27272 69576
rect 59421 69528 86372 69576
rect 0 69455 86372 69528
rect 0 69399 27788 69455
rect 27844 69399 27999 69455
rect 28055 69399 28210 69455
rect 28266 69399 28421 69455
rect 28477 69399 28632 69455
rect 28688 69399 28843 69455
rect 28899 69399 29054 69455
rect 29110 69399 56013 69455
rect 56069 69399 56224 69455
rect 56280 69399 56435 69455
rect 56491 69399 56646 69455
rect 56702 69399 56857 69455
rect 56913 69399 57068 69455
rect 57124 69399 57279 69455
rect 57335 69399 86372 69455
rect 0 69327 86372 69399
rect 0 69276 27272 69327
rect 30403 69326 54622 69327
rect 59421 69276 86372 69327
rect 0 69076 1014 69276
rect 85358 69076 86372 69276
rect 0 68176 1706 68876
rect 84666 68176 86372 68876
rect 0 67776 1014 67976
rect 85358 67776 86372 67976
rect 0 67728 27272 67776
rect 59421 67728 86372 67776
rect 0 67655 86372 67728
rect 0 67599 27788 67655
rect 27844 67599 27999 67655
rect 28055 67599 28210 67655
rect 28266 67599 28421 67655
rect 28477 67599 28632 67655
rect 28688 67599 28843 67655
rect 28899 67599 29054 67655
rect 29110 67599 56013 67655
rect 56069 67599 56224 67655
rect 56280 67599 56435 67655
rect 56491 67599 56646 67655
rect 56702 67599 56857 67655
rect 56913 67599 57068 67655
rect 57124 67599 57279 67655
rect 57335 67599 86372 67655
rect 0 67527 86372 67599
rect 0 67476 27272 67527
rect 30403 67526 54622 67527
rect 59421 67476 86372 67527
rect 0 67276 1014 67476
rect 85358 67276 86372 67476
rect 0 66376 1706 67076
rect 84666 66376 86372 67076
rect 0 65976 1014 66176
rect 85358 65976 86372 66176
rect 0 65928 27272 65976
rect 59421 65928 86372 65976
rect 0 65855 86372 65928
rect 0 65799 27788 65855
rect 27844 65799 27999 65855
rect 28055 65799 28210 65855
rect 28266 65799 28421 65855
rect 28477 65799 28632 65855
rect 28688 65799 28843 65855
rect 28899 65799 29054 65855
rect 29110 65799 56013 65855
rect 56069 65799 56224 65855
rect 56280 65799 56435 65855
rect 56491 65799 56646 65855
rect 56702 65799 56857 65855
rect 56913 65799 57068 65855
rect 57124 65799 57279 65855
rect 57335 65799 86372 65855
rect 0 65727 86372 65799
rect 0 65676 27272 65727
rect 30403 65726 54622 65727
rect 59421 65676 86372 65727
rect 0 65476 1014 65676
rect 85358 65476 86372 65676
rect 0 64576 1706 65276
rect 84666 64576 86372 65276
rect 0 64176 1014 64376
rect 85358 64176 86372 64376
rect 0 64128 27272 64176
rect 59421 64128 86372 64176
rect 0 64055 86372 64128
rect 0 63999 27788 64055
rect 27844 63999 27999 64055
rect 28055 63999 28210 64055
rect 28266 63999 28421 64055
rect 28477 63999 28632 64055
rect 28688 63999 28843 64055
rect 28899 63999 29054 64055
rect 29110 63999 56013 64055
rect 56069 63999 56224 64055
rect 56280 63999 56435 64055
rect 56491 63999 56646 64055
rect 56702 63999 56857 64055
rect 56913 63999 57068 64055
rect 57124 63999 57279 64055
rect 57335 63999 86372 64055
rect 0 63927 86372 63999
rect 0 63876 27272 63927
rect 30403 63926 54622 63927
rect 59421 63876 86372 63927
rect 0 63676 1014 63876
rect 85358 63676 86372 63876
rect 0 62776 1706 63476
rect 84666 62776 86372 63476
rect 0 62376 1014 62576
rect 85358 62376 86372 62576
rect 0 62328 27272 62376
rect 59421 62328 86372 62376
rect 0 62255 86372 62328
rect 0 62199 27788 62255
rect 27844 62199 27999 62255
rect 28055 62199 28210 62255
rect 28266 62199 28421 62255
rect 28477 62199 28632 62255
rect 28688 62199 28843 62255
rect 28899 62199 29054 62255
rect 29110 62199 56013 62255
rect 56069 62199 56224 62255
rect 56280 62199 56435 62255
rect 56491 62199 56646 62255
rect 56702 62199 56857 62255
rect 56913 62199 57068 62255
rect 57124 62199 57279 62255
rect 57335 62199 86372 62255
rect 0 62127 86372 62199
rect 0 62076 27272 62127
rect 30403 62126 54622 62127
rect 59421 62076 86372 62127
rect 0 61876 1014 62076
rect 85358 61876 86372 62076
rect 0 60976 1706 61676
rect 84666 60976 86372 61676
rect 0 60576 1014 60776
rect 85358 60576 86372 60776
rect 0 60528 27272 60576
rect 59421 60528 86372 60576
rect 0 60455 86372 60528
rect 0 60399 27788 60455
rect 27844 60399 27999 60455
rect 28055 60399 28210 60455
rect 28266 60399 28421 60455
rect 28477 60399 28632 60455
rect 28688 60399 28843 60455
rect 28899 60399 29054 60455
rect 29110 60399 56013 60455
rect 56069 60399 56224 60455
rect 56280 60399 56435 60455
rect 56491 60399 56646 60455
rect 56702 60399 56857 60455
rect 56913 60399 57068 60455
rect 57124 60399 57279 60455
rect 57335 60399 86372 60455
rect 0 60327 86372 60399
rect 0 60276 27272 60327
rect 30403 60326 54622 60327
rect 59421 60276 86372 60327
rect 0 60076 1014 60276
rect 85358 60076 86372 60276
rect 0 59176 1706 59876
rect 84666 59176 86372 59876
rect 0 58776 1014 58976
rect 85358 58776 86372 58976
rect 0 58728 27272 58776
rect 59421 58728 86372 58776
rect 0 58655 86372 58728
rect 0 58599 27788 58655
rect 27844 58599 27999 58655
rect 28055 58599 28210 58655
rect 28266 58599 28421 58655
rect 28477 58599 28632 58655
rect 28688 58599 28843 58655
rect 28899 58599 29054 58655
rect 29110 58599 56013 58655
rect 56069 58599 56224 58655
rect 56280 58599 56435 58655
rect 56491 58599 56646 58655
rect 56702 58599 56857 58655
rect 56913 58599 57068 58655
rect 57124 58599 57279 58655
rect 57335 58599 86372 58655
rect 0 58527 86372 58599
rect 0 58476 27272 58527
rect 30403 58526 54622 58527
rect 59421 58476 86372 58527
rect 0 58276 1014 58476
rect 85358 58276 86372 58476
rect 0 57376 1706 58076
rect 84666 57376 86372 58076
rect 0 56976 1014 57176
rect 85358 56976 86372 57176
rect 0 56928 27272 56976
rect 59421 56928 86372 56976
rect 0 56855 86372 56928
rect 0 56799 27788 56855
rect 27844 56799 27999 56855
rect 28055 56799 28210 56855
rect 28266 56799 28421 56855
rect 28477 56799 28632 56855
rect 28688 56799 28843 56855
rect 28899 56799 29054 56855
rect 29110 56799 56013 56855
rect 56069 56799 56224 56855
rect 56280 56799 56435 56855
rect 56491 56799 56646 56855
rect 56702 56799 56857 56855
rect 56913 56799 57068 56855
rect 57124 56799 57279 56855
rect 57335 56799 86372 56855
rect 0 56727 86372 56799
rect 0 56676 27272 56727
rect 30403 56726 54622 56727
rect 59421 56676 86372 56727
rect 0 56476 1014 56676
rect 85358 56476 86372 56676
rect 0 55576 1706 56276
rect 84666 55576 86372 56276
rect 0 55176 1014 55376
rect 85358 55176 86372 55376
rect 0 55128 27272 55176
rect 59421 55128 86372 55176
rect 0 55055 86372 55128
rect 0 54999 27788 55055
rect 27844 54999 27999 55055
rect 28055 54999 28210 55055
rect 28266 54999 28421 55055
rect 28477 54999 28632 55055
rect 28688 54999 28843 55055
rect 28899 54999 29054 55055
rect 29110 54999 56013 55055
rect 56069 54999 56224 55055
rect 56280 54999 56435 55055
rect 56491 54999 56646 55055
rect 56702 54999 56857 55055
rect 56913 54999 57068 55055
rect 57124 54999 57279 55055
rect 57335 54999 86372 55055
rect 0 54927 86372 54999
rect 0 54876 27272 54927
rect 30403 54926 54622 54927
rect 59421 54876 86372 54927
rect 0 54676 1014 54876
rect 85358 54676 86372 54876
rect 0 53776 1706 54476
rect 84666 53776 86372 54476
rect 0 53376 1014 53576
rect 85358 53376 86372 53576
rect 0 53328 27272 53376
rect 59421 53328 86372 53376
rect 0 53255 86372 53328
rect 0 53199 27788 53255
rect 27844 53199 27999 53255
rect 28055 53199 28210 53255
rect 28266 53199 28421 53255
rect 28477 53199 28632 53255
rect 28688 53199 28843 53255
rect 28899 53199 29054 53255
rect 29110 53199 56013 53255
rect 56069 53199 56224 53255
rect 56280 53199 56435 53255
rect 56491 53199 56646 53255
rect 56702 53199 56857 53255
rect 56913 53199 57068 53255
rect 57124 53199 57279 53255
rect 57335 53199 86372 53255
rect 0 53127 86372 53199
rect 0 53076 27272 53127
rect 30403 53126 54622 53127
rect 59421 53076 86372 53127
rect 0 52876 1014 53076
rect 85358 52876 86372 53076
rect 0 51976 1706 52676
rect 84666 51976 86372 52676
rect 0 51576 1014 51776
rect 85358 51576 86372 51776
rect 0 51528 27272 51576
rect 59421 51528 86372 51576
rect 0 51455 86372 51528
rect 0 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 86372 51455
rect 0 51327 86372 51399
rect 0 51276 27272 51327
rect 30403 51326 54622 51327
rect 59421 51276 86372 51327
rect 0 51076 1014 51276
rect 85358 51076 86372 51276
rect 0 50176 1706 50876
rect 84666 50176 86372 50876
rect 0 49776 1014 49976
rect 85358 49776 86372 49976
rect 0 49728 27272 49776
rect 59421 49728 86372 49776
rect 0 49655 86372 49728
rect 0 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 86372 49655
rect 0 49527 86372 49599
rect 0 49476 27272 49527
rect 30403 49526 54622 49527
rect 59421 49476 86372 49527
rect 0 49276 1014 49476
rect 85358 49276 86372 49476
rect 0 48376 1706 49076
rect 84666 48376 86372 49076
rect 0 47976 1014 48176
rect 85358 47976 86372 48176
rect 0 47928 27272 47976
rect 59421 47928 86372 47976
rect 0 47855 86372 47928
rect 0 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 86372 47855
rect 0 47727 86372 47799
rect 0 47676 27272 47727
rect 30403 47726 54622 47727
rect 59421 47676 86372 47727
rect 0 47476 1014 47676
rect 85358 47476 86372 47676
rect 0 46576 1706 47276
rect 84666 46576 86372 47276
rect 0 46176 1014 46376
rect 85358 46176 86372 46376
rect 0 46128 27272 46176
rect 59421 46128 86372 46176
rect 0 46055 86372 46128
rect 0 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 86372 46055
rect 0 45927 86372 45999
rect 0 45876 27272 45927
rect 30403 45926 54622 45927
rect 59421 45876 86372 45927
rect 0 45676 1014 45876
rect 85358 45676 86372 45876
rect 0 44776 1706 45476
rect 84666 44776 86372 45476
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44328 27272 44376
rect 59421 44328 86372 44376
rect 0 44255 86372 44328
rect 0 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 86372 44255
rect 0 44127 86372 44199
rect 0 44076 27272 44127
rect 30403 44126 54622 44127
rect 59421 44076 86372 44127
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42528 27272 42576
rect 59421 42528 86372 42576
rect 0 42455 86372 42528
rect 0 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 86372 42455
rect 0 42327 86372 42399
rect 0 42276 27272 42327
rect 30403 42326 54622 42327
rect 59421 42276 86372 42327
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40728 27272 40776
rect 59421 40728 86372 40776
rect 0 40655 86372 40728
rect 0 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 86372 40655
rect 0 40527 86372 40599
rect 0 40476 27272 40527
rect 30403 40526 54622 40527
rect 59421 40476 86372 40527
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38928 27272 38976
rect 59421 38928 86372 38976
rect 0 38855 86372 38928
rect 0 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 86372 38855
rect 0 38727 86372 38799
rect 0 38676 27272 38727
rect 30403 38726 54622 38727
rect 59421 38676 86372 38727
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37128 27272 37176
rect 59421 37128 86372 37176
rect 0 37055 86372 37128
rect 0 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 86372 37055
rect 0 36927 86372 36999
rect 0 36876 27272 36927
rect 30403 36926 54622 36927
rect 59421 36876 86372 36927
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 36863 35881 37743 35920
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 0 35126 24917 35326
rect 0 35016 1014 35126
rect 0 34992 27830 35016
rect 0 34936 25386 34992
rect 25442 34936 25510 34992
rect 25566 34936 25634 34992
rect 25690 34936 25758 34992
rect 25814 34936 25882 34992
rect 25938 34936 27447 34992
rect 27503 34936 27571 34992
rect 27627 34936 27695 34992
rect 27751 34936 27830 34992
rect 0 34868 27830 34936
rect 0 34812 25386 34868
rect 25442 34812 25510 34868
rect 25566 34812 25634 34868
rect 25690 34812 25758 34868
rect 25814 34812 25882 34868
rect 25938 34812 27447 34868
rect 27503 34812 27571 34868
rect 27627 34812 27695 34868
rect 27751 34812 27830 34868
rect 0 34744 27830 34812
rect 0 34688 25386 34744
rect 25442 34688 25510 34744
rect 25566 34688 25634 34744
rect 25690 34688 25758 34744
rect 25814 34688 25882 34744
rect 25938 34688 27447 34744
rect 27503 34688 27571 34744
rect 27627 34688 27695 34744
rect 27751 34688 27830 34744
rect 0 34620 27830 34688
rect 0 34564 25386 34620
rect 25442 34564 25510 34620
rect 25566 34564 25634 34620
rect 25690 34564 25758 34620
rect 25814 34564 25882 34620
rect 25938 34564 27447 34620
rect 27503 34564 27571 34620
rect 27627 34564 27695 34620
rect 27751 34564 27830 34620
rect 0 34536 27830 34564
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 34011 27214 34124
rect 0 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27214 34011
rect 0 33793 27214 33955
rect 36863 33927 37743 35825
rect 84666 35776 86372 36476
rect 83360 35298 86372 35326
rect 60460 35158 86372 35298
rect 83360 35126 86372 35158
rect 85358 35016 86372 35126
rect 58791 34992 86372 35016
rect 58791 34936 58816 34992
rect 58872 34936 58940 34992
rect 58996 34936 59064 34992
rect 59120 34936 59188 34992
rect 59244 34936 59312 34992
rect 59368 34936 59436 34992
rect 59492 34936 86372 34992
rect 58791 34868 86372 34936
rect 58791 34812 58816 34868
rect 58872 34812 58940 34868
rect 58996 34812 59064 34868
rect 59120 34812 59188 34868
rect 59244 34812 59312 34868
rect 59368 34812 59436 34868
rect 59492 34812 86372 34868
rect 58791 34744 86372 34812
rect 58791 34688 58816 34744
rect 58872 34688 58940 34744
rect 58996 34688 59064 34744
rect 59120 34688 59188 34744
rect 59244 34688 59312 34744
rect 59368 34688 59436 34744
rect 59492 34688 86372 34744
rect 58791 34620 86372 34688
rect 58791 34564 58816 34620
rect 58872 34564 58940 34620
rect 58996 34564 59064 34620
rect 59120 34564 59188 34620
rect 59244 34564 59312 34620
rect 59368 34564 59436 34620
rect 59492 34564 86372 34620
rect 58791 34536 86372 34564
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 34011 86372 34124
rect 57908 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 86372 34011
rect 0 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27214 33793
rect 0 33576 27214 33737
rect 0 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27214 33576
rect 0 33358 27214 33520
rect 0 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27214 33358
rect 0 33140 27214 33302
rect 57908 33793 86372 33955
rect 57908 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 86372 33793
rect 57908 33576 86372 33737
rect 57908 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 86372 33576
rect 57908 33358 86372 33520
rect 57908 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 86372 33358
rect 0 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27214 33140
rect 0 32922 27214 33084
rect 0 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27214 32922
rect 0 32705 27214 32866
rect 0 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27214 32705
rect 0 32487 27214 32649
rect 0 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27214 32487
rect 0 32318 27214 32431
rect 27387 33141 28929 33263
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 28929 33141
rect 27387 32923 28929 33085
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 28929 32923
rect 27387 32705 28929 32867
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 28929 32705
rect 27387 32487 28929 32649
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 28929 32487
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 27387 32311 28929 32431
rect 56135 33141 57736 33263
rect 56135 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 56135 32923 57736 33085
rect 56135 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 56135 32705 57736 32867
rect 56135 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 56135 32487 57736 32649
rect 56135 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 56135 32311 57736 32431
rect 57908 33140 86372 33302
rect 57908 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 86372 33140
rect 57908 32922 86372 33084
rect 57908 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 86372 32922
rect 57908 32705 86372 32866
rect 57908 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 86372 32705
rect 57908 32487 86372 32649
rect 57908 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 86372 32487
rect 57908 32315 86372 32431
rect 57908 32199 58351 32315
rect 26772 32088 58351 32199
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 26772 31870 58351 32032
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 26772 31652 58351 31814
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 26772 31486 58351 31596
rect 25293 31252 28929 31352
rect 25293 31248 27474 31252
rect 25293 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31196 27474 31248
rect 27530 31196 27686 31252
rect 27742 31196 28929 31252
rect 25950 31192 28929 31196
rect 25293 31124 28929 31192
rect 25293 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 28929 31124
rect 25293 31034 28929 31068
rect 25293 31000 27474 31034
rect 25293 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30978 27474 31000
rect 27530 30978 27686 31034
rect 27742 30978 28929 31034
rect 25950 30944 28929 30978
rect 25293 30816 28929 30944
rect 25293 30793 27474 30816
rect 25293 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30760 27474 30793
rect 27530 30760 27686 30816
rect 27742 30760 28929 30816
rect 25950 30737 28929 30760
rect 25293 30669 28929 30737
rect 25293 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 28929 30669
rect 25293 30598 28929 30613
rect 25293 30545 27474 30598
rect 25293 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30542 27474 30545
rect 27530 30542 27686 30598
rect 27742 30542 28929 30598
rect 25950 30489 28929 30542
rect 25293 30443 28929 30489
rect 56186 31298 59524 31352
rect 56186 31252 58873 31298
rect 56186 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31242 58873 31252
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59524 31298
rect 57649 31196 59524 31242
rect 56186 31174 59524 31196
rect 56186 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59524 31174
rect 56186 31050 59524 31118
rect 56186 31034 58873 31050
rect 56186 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30994 58873 31034
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59524 31050
rect 57649 30978 59524 30994
rect 56186 30853 59524 30978
rect 56186 30816 58873 30853
rect 56186 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30797 58873 30816
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59524 30853
rect 57649 30760 59524 30797
rect 56186 30729 59524 30760
rect 56186 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59524 30729
rect 56186 30605 59524 30673
rect 56186 30598 58873 30605
rect 56186 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30549 58873 30598
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59524 30605
rect 57649 30542 59524 30549
rect 56186 30443 59524 30542
rect 26772 29968 58351 30105
rect 26772 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 26772 29750 58351 29912
rect 26772 29714 26859 29750
rect 0 29694 26859 29714
rect 26915 29694 27071 29750
rect 27127 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29714 58351 29750
rect 84666 29714 86372 32315
rect 58264 29694 86372 29714
rect 0 29533 86372 29694
rect 0 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 86372 29533
rect 0 29430 86372 29477
rect 26772 29315 58351 29430
rect 26772 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 26772 29098 58351 29259
rect 26772 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 26772 28880 58351 29042
rect 26772 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 26772 28662 58351 28824
rect 26772 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 26772 28444 58351 28606
rect 0 28412 3011 28416
rect 0 28317 26070 28412
rect 0 28261 25404 28317
rect 25460 28261 25528 28317
rect 25584 28261 25652 28317
rect 25708 28261 25776 28317
rect 25832 28261 25900 28317
rect 25956 28261 26070 28317
rect 0 28193 26070 28261
rect 0 28137 25404 28193
rect 25460 28137 25528 28193
rect 25584 28137 25652 28193
rect 25708 28137 25776 28193
rect 25832 28137 25900 28193
rect 25956 28137 26070 28193
rect 0 28069 26070 28137
rect 0 28013 25404 28069
rect 25460 28013 25528 28069
rect 25584 28013 25652 28069
rect 25708 28013 25776 28069
rect 25832 28013 25900 28069
rect 25956 28013 26070 28069
rect 0 27945 26070 28013
rect 0 27889 25404 27945
rect 25460 27889 25528 27945
rect 25584 27889 25652 27945
rect 25708 27889 25776 27945
rect 25832 27889 25900 27945
rect 25956 27889 26070 27945
rect 0 27821 26070 27889
rect 0 27765 25404 27821
rect 25460 27765 25528 27821
rect 25584 27765 25652 27821
rect 25708 27765 25776 27821
rect 25832 27765 25900 27821
rect 25956 27765 26070 27821
rect 0 27697 26070 27765
rect 0 27641 25404 27697
rect 25460 27641 25528 27697
rect 25584 27641 25652 27697
rect 25708 27641 25776 27697
rect 25832 27641 25900 27697
rect 25956 27641 26070 27697
rect 0 27573 26070 27641
rect 0 27517 25404 27573
rect 25460 27517 25528 27573
rect 25584 27517 25652 27573
rect 25708 27517 25776 27573
rect 25832 27517 25900 27573
rect 25956 27517 26070 27573
rect 0 27449 26070 27517
rect 0 27393 25404 27449
rect 25460 27393 25528 27449
rect 25584 27393 25652 27449
rect 25708 27393 25776 27449
rect 25832 27393 25900 27449
rect 25956 27393 26070 27449
rect 0 27325 26070 27393
rect 26772 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 83361 28412 86372 28416
rect 26772 28227 58351 28388
rect 26772 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 26772 28009 58351 28171
rect 26772 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 26772 27792 58351 27953
rect 26772 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 26772 27574 58351 27736
rect 26772 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 26772 27382 58351 27518
rect 58785 28295 86372 28412
rect 58785 28239 58859 28295
rect 58915 28239 58983 28295
rect 59039 28239 59107 28295
rect 59163 28239 59231 28295
rect 59287 28239 59355 28295
rect 59411 28239 86372 28295
rect 58785 28171 86372 28239
rect 58785 28115 58859 28171
rect 58915 28115 58983 28171
rect 59039 28115 59107 28171
rect 59163 28115 59231 28171
rect 59287 28115 59355 28171
rect 59411 28115 86372 28171
rect 58785 28047 86372 28115
rect 58785 27991 58859 28047
rect 58915 27991 58983 28047
rect 59039 27991 59107 28047
rect 59163 27991 59231 28047
rect 59287 27991 59355 28047
rect 59411 27991 86372 28047
rect 58785 27923 86372 27991
rect 58785 27867 58859 27923
rect 58915 27867 58983 27923
rect 59039 27867 59107 27923
rect 59163 27867 59231 27923
rect 59287 27867 59355 27923
rect 59411 27867 86372 27923
rect 58785 27799 86372 27867
rect 58785 27743 58859 27799
rect 58915 27743 58983 27799
rect 59039 27743 59107 27799
rect 59163 27743 59231 27799
rect 59287 27743 59355 27799
rect 59411 27743 86372 27799
rect 58785 27675 86372 27743
rect 58785 27619 58859 27675
rect 58915 27619 58983 27675
rect 59039 27619 59107 27675
rect 59163 27619 59231 27675
rect 59287 27619 59355 27675
rect 59411 27619 86372 27675
rect 58785 27551 86372 27619
rect 58785 27495 58859 27551
rect 58915 27495 58983 27551
rect 59039 27495 59107 27551
rect 59163 27495 59231 27551
rect 59287 27495 59355 27551
rect 59411 27495 86372 27551
rect 58785 27427 86372 27495
rect 0 27269 25404 27325
rect 25460 27269 25528 27325
rect 25584 27269 25652 27325
rect 25708 27269 25776 27325
rect 25832 27269 25900 27325
rect 25956 27269 26070 27325
rect 0 27201 26070 27269
rect 0 27145 25404 27201
rect 25460 27145 25528 27201
rect 25584 27145 25652 27201
rect 25708 27145 25776 27201
rect 25832 27145 25900 27201
rect 25956 27145 26070 27201
rect 0 27077 26070 27145
rect 0 27021 25404 27077
rect 25460 27021 25528 27077
rect 25584 27021 25652 27077
rect 25708 27021 25776 27077
rect 25832 27021 25900 27077
rect 25956 27021 26070 27077
rect 0 26953 26070 27021
rect 0 26897 25404 26953
rect 25460 26897 25528 26953
rect 25584 26897 25652 26953
rect 25708 26897 25776 26953
rect 25832 26897 25900 26953
rect 25956 26897 26070 26953
rect 0 26890 26070 26897
rect 58785 27371 58859 27427
rect 58915 27371 58983 27427
rect 59039 27371 59107 27427
rect 59163 27371 59231 27427
rect 59287 27371 59355 27427
rect 59411 27371 86372 27427
rect 58785 27303 86372 27371
rect 58785 27247 58859 27303
rect 58915 27247 58983 27303
rect 59039 27247 59107 27303
rect 59163 27247 59231 27303
rect 59287 27247 59355 27303
rect 59411 27247 86372 27303
rect 58785 27179 86372 27247
rect 58785 27123 58859 27179
rect 58915 27123 58983 27179
rect 59039 27123 59107 27179
rect 59163 27123 59231 27179
rect 59287 27123 59355 27179
rect 59411 27123 86372 27179
rect 58785 27055 86372 27123
rect 58785 26999 58859 27055
rect 58915 26999 58983 27055
rect 59039 26999 59107 27055
rect 59163 26999 59231 27055
rect 59287 26999 59355 27055
rect 59411 26999 86372 27055
rect 58785 26931 86372 26999
rect 58785 26890 58859 26931
rect 0 26829 27828 26890
rect 0 26773 25404 26829
rect 25460 26773 25528 26829
rect 25584 26773 25652 26829
rect 25708 26773 25776 26829
rect 25832 26773 25900 26829
rect 25956 26799 27828 26829
rect 25956 26773 27474 26799
rect 0 26743 27474 26773
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 0 26705 27828 26743
rect 0 26649 25404 26705
rect 25460 26649 25528 26705
rect 25584 26649 25652 26705
rect 25708 26649 25776 26705
rect 25832 26649 25900 26705
rect 25956 26649 27828 26705
rect 0 26581 27828 26649
rect 0 26525 25404 26581
rect 25460 26525 25528 26581
rect 25584 26525 25652 26581
rect 25708 26525 25776 26581
rect 25832 26525 25900 26581
rect 25956 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 0 26435 27828 26525
rect 57295 26875 58859 26890
rect 58915 26875 58983 26931
rect 59039 26875 59107 26931
rect 59163 26875 59231 26931
rect 59287 26875 59355 26931
rect 59411 26875 86372 26931
rect 57295 26807 86372 26875
rect 57295 26799 58859 26807
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26751 58859 26799
rect 58915 26751 58983 26807
rect 59039 26751 59107 26807
rect 59163 26751 59231 26807
rect 59287 26751 59355 26807
rect 59411 26751 86372 26807
rect 57649 26743 86372 26751
rect 57295 26683 86372 26743
rect 57295 26627 58859 26683
rect 58915 26627 58983 26683
rect 59039 26627 59107 26683
rect 59163 26627 59231 26683
rect 59287 26627 59355 26683
rect 59411 26627 86372 26683
rect 57295 26581 86372 26627
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26559 86372 26581
rect 57649 26525 58859 26559
rect 57295 26503 58859 26525
rect 58915 26503 58983 26559
rect 59039 26503 59107 26559
rect 59163 26503 59231 26559
rect 59287 26503 59355 26559
rect 59411 26503 86372 26559
rect 57295 26435 86372 26503
rect 6921 26434 8163 26435
rect 17721 26434 18963 26435
rect 23425 26434 27828 26435
rect 66497 26434 67739 26435
rect 77297 26434 78539 26435
rect 23828 26286 26642 26324
rect 23828 26126 26450 26286
rect 26610 26126 26642 26286
rect 23828 26109 26642 26126
rect 23828 25967 26285 26002
rect 23828 25807 26092 25967
rect 26252 25807 26285 25967
rect 23828 25787 26285 25807
rect 23828 25647 25949 25681
rect 23828 25487 25756 25647
rect 25916 25487 25949 25647
rect 23828 25466 25949 25487
rect 23828 25328 25614 25359
rect 23828 25168 25421 25328
rect 25581 25168 25614 25328
rect 23828 25144 25614 25168
rect 27382 25028 29699 25208
rect 27382 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 29699 25028
rect 27382 24810 29699 24972
rect 27382 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 29699 24810
rect 23828 24637 25274 24667
rect 23828 24477 25081 24637
rect 25241 24477 25274 24637
rect 27382 24526 29699 24754
rect 23828 24452 25274 24477
rect 23828 24316 24935 24345
rect 23828 24156 24744 24316
rect 24904 24156 24935 24316
rect 23828 24130 24935 24156
rect 26770 24075 58348 24278
rect 23828 23995 24607 24024
rect 0 23380 1706 23938
rect 23828 23835 24416 23995
rect 24576 23835 24607 23995
rect 23828 23809 24607 23835
rect 24047 23673 24227 23683
rect 24047 23513 24057 23673
rect 24217 23513 24227 23673
rect 24047 23503 24227 23513
rect 26770 23380 26858 24075
rect 0 23187 26858 23380
rect 27122 23370 57994 24075
rect 27122 23187 27214 23370
rect 0 22938 27214 23187
rect 27387 22936 57681 23199
rect 57908 23187 57994 23370
rect 58258 23380 58348 24075
rect 84666 23380 86372 23938
rect 58258 23187 86372 23380
rect 57908 22938 86372 23187
rect 57908 22937 83763 22938
rect 27387 22282 27475 22936
rect 0 22048 27475 22282
rect 27739 22923 57681 22936
rect 27739 22291 57363 22923
rect 27739 22048 27826 22291
rect 0 21827 27826 22048
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 22035 57363 22291
rect 57627 22282 57681 22923
rect 57627 22035 86372 22282
rect 56078 21827 86372 22035
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 20570 86372 20739
rect 0 20410 26924 20570
rect 27084 20410 58048 20570
rect 58208 20410 86372 20570
rect 0 20226 86372 20410
rect 0 20066 26924 20226
rect 27084 20066 58048 20226
rect 58208 20066 86372 20226
rect 0 19969 86372 20066
rect 0 18016 24250 19969
rect 26435 19692 29403 19731
rect 26435 19532 26465 19692
rect 26625 19532 29403 19692
rect 26435 19502 29403 19532
rect 55720 19502 58817 19731
rect 26077 19347 29403 19391
rect 26077 19187 26107 19347
rect 26267 19187 29403 19347
rect 26077 19162 29403 19187
rect 55720 19162 59177 19391
rect 25742 19027 29403 19051
rect 25742 18867 25771 19027
rect 25931 18867 29403 19027
rect 25742 18822 29403 18867
rect 55720 18822 59515 19051
rect 25406 18684 29403 18711
rect 25406 18524 25434 18684
rect 25594 18524 29403 18684
rect 25406 18482 29403 18524
rect 55720 18482 59846 18711
rect 25066 18350 29403 18371
rect 25066 18190 25094 18350
rect 25254 18190 29403 18350
rect 25066 18142 29403 18190
rect 55720 18142 60184 18371
rect 24730 17977 29403 18031
rect 24730 17817 24757 17977
rect 24917 17817 29403 17977
rect 24730 17802 29403 17817
rect 55720 17802 60525 18031
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 24401 17656 29403 17691
rect 24401 17496 24429 17656
rect 24589 17496 29403 17656
rect 24401 17462 29403 17496
rect 55720 17462 60855 17691
rect 24042 17317 29403 17351
rect 24042 17157 24069 17317
rect 24229 17157 29403 17317
rect 24042 17122 29403 17157
rect 55720 17122 61205 17351
rect 61807 16784 86372 17730
rect 46982 16678 86372 16784
rect 46982 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 86372 16678
rect 24111 16597 27828 16598
rect 0 16470 27828 16597
rect 0 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 0 16253 27828 16414
rect 0 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 0 16035 27828 16197
rect 0 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 0 15818 27828 15979
rect 0 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 0 15600 27828 15762
rect 0 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 0 15382 27828 15544
rect 0 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 0 15164 27828 15326
rect 0 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 0 15015 27828 15108
rect 46982 16461 86372 16622
rect 46982 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 86372 16461
rect 46982 16243 86372 16405
rect 46982 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 86372 16243
rect 46982 16026 86372 16187
rect 46982 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 86372 16026
rect 46982 15808 86372 15970
rect 46982 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 86372 15808
rect 46982 15590 86372 15752
rect 46982 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 86372 15590
rect 46982 15372 86372 15534
rect 46982 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 86372 15372
rect 46982 15155 86372 15316
rect 46982 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 86372 15155
rect 46982 15015 86372 15099
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14947 51760 14966
rect 0 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14936 51760 14947
rect 57295 14937 86372 14968
rect 27742 14891 47683 14936
rect 0 14729 47683 14891
rect 0 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 47683 14729
rect 0 14512 47683 14673
rect 0 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14491 47683 14512
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 86372 14937
rect 57295 14720 86372 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 86372 14720
rect 27742 14456 45977 14491
rect 0 14329 45977 14456
rect 0 14328 24250 14329
rect 27387 14231 45977 14329
rect 57295 14328 86372 14664
rect 57295 14327 83763 14328
rect 24047 14178 27214 14179
rect 0 14119 27214 14178
rect 0 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27214 14119
rect 0 13902 27214 14063
rect 0 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27214 13902
rect 0 13684 27214 13846
rect 0 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27214 13684
rect 0 13467 27214 13628
rect 0 13461 26859 13467
rect 0 12846 1706 13461
rect 24047 13411 26859 13461
rect 26915 13411 27071 13467
rect 27127 13411 27214 13467
rect 24047 13249 27214 13411
rect 24047 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27214 13249
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 45977 14231
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 27387 14014 45977 14175
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 45977 14014
rect 27387 13796 45977 13958
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13760 45977 13796
rect 50228 13790 86372 13866
rect 27742 13740 49775 13760
rect 27387 13578 49775 13740
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 49775 13578
rect 27387 13361 49775 13522
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 49775 13361
rect 27387 13245 49775 13305
rect 29478 13243 49775 13245
rect 24047 13031 27214 13193
rect 41493 13078 49775 13243
rect 50228 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 86372 13790
rect 50228 13573 86372 13734
rect 50228 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 86372 13573
rect 50228 13461 86372 13517
rect 50228 13355 58421 13461
rect 50228 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58421 13355
rect 50228 13138 58421 13299
rect 50228 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58421 13138
rect 24047 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27214 13031
rect 24047 12934 27214 12975
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12813 34761 12846
rect 0 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 34761 12813
rect 0 12596 34761 12757
rect 0 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12570 34761 12596
rect 50228 12920 58421 13082
rect 50228 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58421 12920
rect 50228 12846 58421 12864
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12702 86372 12846
rect 50228 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 86372 12702
rect 50228 12570 86372 12646
rect 27127 12540 86372 12570
rect 0 12484 86372 12540
rect 0 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 86372 12484
rect 0 12378 86372 12428
rect 0 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 86372 12378
rect 0 12267 86372 12322
rect 0 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 86372 12267
rect 0 12161 86372 12211
rect 0 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 86372 12161
rect 0 12049 86372 12105
rect 0 12046 57996 12049
rect 0 12036 24250 12046
rect 26772 11993 57996 12046
rect 58052 11993 58208 12049
rect 58264 12036 86372 12049
rect 58264 12035 84999 12036
rect 58264 11993 58351 12035
rect 26772 11844 58351 11993
rect 29478 11832 58351 11844
rect 29478 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 29478 11697 58351 11776
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 11406 27828 11491
rect 0 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 0 11189 27828 11350
rect 0 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 0 10971 27828 11133
rect 0 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 0 10753 27828 10915
rect 29478 10756 41516 11697
rect 61825 11491 86372 11493
rect 0 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 0 10535 27828 10697
rect 0 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 0 10318 27828 10479
rect 0 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 0 10176 27828 10262
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 23612 9942 29221 10030
rect 34741 9972 41516 10756
rect 42261 11406 86372 11491
rect 42261 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 86372 11406
rect 42261 11189 86372 11350
rect 42261 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 86372 11189
rect 42261 10971 86372 11133
rect 42261 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 86372 10971
rect 42261 10753 86372 10915
rect 42261 10740 57381 10753
rect 57295 10697 57381 10740
rect 57437 10697 57593 10753
rect 57649 10697 86372 10753
rect 57295 10535 86372 10697
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 86372 10535
rect 24047 9515 28729 9516
rect 0 9514 1014 9515
rect 2226 9514 28729 9515
rect 0 9407 28729 9514
rect 0 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 28729 9407
rect 0 9190 28729 9351
rect 29133 9302 29221 9942
rect 41857 9502 51430 10420
rect 57295 10318 86372 10479
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 86372 10318
rect 51750 10097 54952 10185
rect 57295 10176 86372 10262
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 51750 9971 51838 10097
rect 51750 9811 51766 9971
rect 51822 9811 51838 9971
rect 54864 10030 54952 10097
rect 54864 9942 62145 10030
rect 51750 9801 51838 9811
rect 58688 9681 61743 9777
rect 57909 9515 62278 9516
rect 57909 9514 72434 9515
rect 72602 9514 83234 9515
rect 85358 9514 86372 9515
rect 29133 9214 41656 9302
rect 0 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 28729 9190
rect 0 8972 28729 9134
rect 0 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 28729 8972
rect 0 8754 28729 8916
rect 41568 8972 41656 9214
rect 41857 9165 55482 9502
rect 41568 8953 50067 8972
rect 41568 8897 49897 8953
rect 50057 8897 50067 8953
rect 41568 8884 50067 8897
rect 50922 8930 55482 9165
rect 57909 9407 86372 9514
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 86372 9407
rect 57909 9190 86372 9351
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 86372 9190
rect 57909 8972 86372 9134
rect 0 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 28729 8754
rect 0 8536 28729 8698
rect 50922 8843 57736 8930
rect 50922 8787 57381 8843
rect 57437 8787 57593 8843
rect 57649 8787 57736 8843
rect 50922 8625 57736 8787
rect 0 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 28729 8536
rect 0 8319 28729 8480
rect 0 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 28729 8319
rect 0 8154 28729 8263
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 28178 7652 28729 8154
rect 29513 7900 41397 8582
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 7535 27828 7595
rect 0 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 0 7317 27828 7479
rect 0 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 0 7099 27828 7261
rect 0 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 28178 7084 34622 7652
rect 0 6982 27828 7043
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 23625 6836 29058 6875
rect 23625 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 29058 6836
rect 23625 6618 29058 6780
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 8569 57381 8625
rect 57437 8569 57593 8625
rect 57649 8569 57736 8625
rect 50922 8408 57736 8569
rect 50922 8352 57381 8408
rect 57437 8352 57593 8408
rect 57649 8352 57736 8408
rect 50922 8190 57736 8352
rect 50922 8134 57381 8190
rect 57437 8134 57593 8190
rect 57649 8134 57736 8190
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 86372 8972
rect 57909 8754 86372 8916
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 86372 8754
rect 57909 8536 86372 8698
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 86372 8536
rect 57909 8319 86372 8480
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 86372 8319
rect 57909 8154 86372 8263
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7972 57736 8134
rect 50922 7916 57381 7972
rect 57437 7916 57593 7972
rect 57649 7916 57736 7972
rect 50922 7755 57736 7916
rect 50922 7699 57381 7755
rect 57437 7699 57593 7755
rect 57649 7699 57736 7755
rect 50922 7596 57736 7699
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7537 86372 7595
rect 50922 7481 57381 7537
rect 57437 7481 57593 7537
rect 57649 7481 86372 7537
rect 50922 7392 86372 7481
rect 34860 7319 86372 7392
rect 34860 7263 57381 7319
rect 57437 7263 57593 7319
rect 57649 7263 86372 7319
rect 34860 7102 86372 7263
rect 34860 7046 57381 7102
rect 57437 7046 57593 7102
rect 57649 7046 86372 7102
rect 34860 6984 86372 7046
rect 23625 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 29058 6618
rect 34860 6592 55482 6984
rect 61802 6982 86372 6984
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 23625 6400 29058 6562
rect 23625 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 29058 6400
rect 23625 6306 29058 6344
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 50922 6199 55482 6592
rect 56065 6836 62747 6874
rect 56065 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 62747 6836
rect 56065 6618 62747 6780
rect 56065 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 62747 6618
rect 56065 6400 62747 6562
rect 56065 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 62747 6400
rect 56065 6306 62747 6344
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 0 6120 34622 6177
rect 0 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 34622 6120
rect 0 5902 34622 6064
rect 0 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 34622 5902
rect 0 5766 34622 5846
rect 29458 5665 34622 5766
rect 50922 6120 86372 6198
rect 50922 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 86372 6120
rect 50922 5902 86372 6064
rect 50922 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 86372 5902
rect 50922 5766 86372 5846
rect 23687 5629 27214 5630
rect 0 5539 27214 5629
rect 50922 5605 55482 5766
rect 57909 5629 62429 5630
rect 0 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27214 5539
rect 0 5321 27214 5483
rect 0 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27214 5321
rect 0 5175 27214 5265
rect 57909 5539 86372 5629
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 86372 5539
rect 57909 5321 86372 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 86372 5321
rect 57909 5175 86372 5265
rect 0 5174 24250 5175
rect 61802 5174 86372 5175
rect 0 5173 3011 5174
rect 83361 5173 86372 5174
rect 0 4515 1712 5173
rect 57909 4619 62429 4621
rect 23909 4528 62429 4619
rect 23909 4515 26859 4528
rect 0 4472 26859 4515
rect 26915 4472 27071 4528
rect 27127 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4515 62429 4528
rect 84660 4515 86372 5173
rect 58264 4472 86372 4515
rect 0 4310 86372 4472
rect 0 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 86372 4310
rect 0 4166 86372 4254
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3837 61215 3875
rect 23909 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 28801 3837
rect 28857 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 61215 3837
rect 23909 3772 61215 3781
rect 0 3619 86372 3772
rect 0 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 28801 3619
rect 28857 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 86372 3619
rect 0 3524 86372 3563
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 60886 3420 86372 3524
rect 0 2854 1014 3420
rect 24169 3050 62588 3066
rect 24169 2994 43800 3050
rect 43960 2994 62588 3050
rect 24169 2978 62588 2994
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
use 512x8M8W_PWR_512x8m81  512x8M8W_PWR_512x8m81_0
timestamp 1762296095
transform 1 0 0 0 1 0
box 1912 6592 83548 35222
use control_512x8_512x8m81  control_512x8_512x8m81_0
timestamp 1762296095
transform 1 0 27533 0 1 4711
box -3624 -1833 31790 30125
use G_ring_512x8m81  G_ring_512x8m81_0
timestamp 1762296095
transform 1 0 282 0 1 0
box 112 620 85672 96289
use GF018_512x8M8WM1_lef_512x8m81  GF018_512x8M8WM1_lef_512x8m81_0
timestamp 1762296095
transform 1 0 0 0 1 0
box 0 0 86372 96976
use lcol4_512_512x8m81  lcol4_512_512x8m81_0
timestamp 1762296095
transform 1 0 2921 0 1 5019
box -1235 -3394 22810 89707
use M1_PSUB4310591302010_512x8m81  M1_PSUB4310591302010_512x8m81_0
timestamp 1762296095
transform 1 0 53710 0 1 2781
box 0 0 1 1
use M1_PSUB4310591302014_512x8m81  M1_PSUB4310591302014_512x8m81_0
timestamp 1762296095
transform 1 0 34404 0 1 2781
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_0
timestamp 1762296095
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_1
timestamp 1762296095
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_2
timestamp 1762296095
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_3
timestamp 1762296095
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_4
timestamp 1762296095
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_5
timestamp 1762296095
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_6
timestamp 1762296095
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_7
timestamp 1762296095
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_8
timestamp 1762296095
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_9
timestamp 1762296095
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_10
timestamp 1762296095
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_11
timestamp 1762296095
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_12
timestamp 1762296095
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_13
timestamp 1762296095
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_14
timestamp 1762296095
transform 1 0 28449 0 1 92827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_15
timestamp 1762296095
transform 1 0 28449 0 1 91027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_16
timestamp 1762296095
transform 1 0 28449 0 1 89227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_17
timestamp 1762296095
transform 1 0 28449 0 1 87427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_18
timestamp 1762296095
transform 1 0 28449 0 1 85627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_19
timestamp 1762296095
transform 1 0 28449 0 1 83827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_20
timestamp 1762296095
transform 1 0 28449 0 1 82027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_21
timestamp 1762296095
transform 1 0 28449 0 1 80227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_22
timestamp 1762296095
transform 1 0 28449 0 1 78427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_23
timestamp 1762296095
transform 1 0 28449 0 1 76627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_24
timestamp 1762296095
transform 1 0 28449 0 1 74827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_25
timestamp 1762296095
transform 1 0 28449 0 1 73027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_26
timestamp 1762296095
transform 1 0 28449 0 1 71227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_27
timestamp 1762296095
transform 1 0 28449 0 1 69427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_28
timestamp 1762296095
transform 1 0 28449 0 1 67627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_29
timestamp 1762296095
transform 1 0 28449 0 1 65827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_30
timestamp 1762296095
transform 1 0 28449 0 1 64027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_31
timestamp 1762296095
transform 1 0 28449 0 1 62227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_32
timestamp 1762296095
transform 1 0 28449 0 1 60427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_33
timestamp 1762296095
transform 1 0 28449 0 1 58627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_34
timestamp 1762296095
transform 1 0 28449 0 1 56827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_35
timestamp 1762296095
transform 1 0 28449 0 1 55027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_36
timestamp 1762296095
transform 1 0 28449 0 1 53227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_37
timestamp 1762296095
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_38
timestamp 1762296095
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_39
timestamp 1762296095
transform 1 0 28449 0 1 94627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_40
timestamp 1762296095
transform 1 0 56674 0 1 87427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_41
timestamp 1762296095
transform 1 0 56674 0 1 89227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_42
timestamp 1762296095
transform 1 0 56674 0 1 91027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_43
timestamp 1762296095
transform 1 0 56674 0 1 92827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_44
timestamp 1762296095
transform 1 0 56674 0 1 94627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_45
timestamp 1762296095
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_46
timestamp 1762296095
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_47
timestamp 1762296095
transform 1 0 56674 0 1 53227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_48
timestamp 1762296095
transform 1 0 56674 0 1 55027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_49
timestamp 1762296095
transform 1 0 56674 0 1 56827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_50
timestamp 1762296095
transform 1 0 56674 0 1 58627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_51
timestamp 1762296095
transform 1 0 56674 0 1 60427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_52
timestamp 1762296095
transform 1 0 56674 0 1 62227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_53
timestamp 1762296095
transform 1 0 56674 0 1 64027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_54
timestamp 1762296095
transform 1 0 56674 0 1 65827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_55
timestamp 1762296095
transform 1 0 56674 0 1 67627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_56
timestamp 1762296095
transform 1 0 56674 0 1 69427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_57
timestamp 1762296095
transform 1 0 56674 0 1 71227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_58
timestamp 1762296095
transform 1 0 56674 0 1 73027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_59
timestamp 1762296095
transform 1 0 56674 0 1 74827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_60
timestamp 1762296095
transform 1 0 56674 0 1 76627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_61
timestamp 1762296095
transform 1 0 56674 0 1 78427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_62
timestamp 1762296095
transform 1 0 56674 0 1 80227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_63
timestamp 1762296095
transform 1 0 56674 0 1 82027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_64
timestamp 1762296095
transform 1 0 56674 0 1 83827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_65
timestamp 1762296095
transform 1 0 56674 0 1 85627
box 0 0 1 1
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_0
timestamp 1762296095
transform -1 0 57515 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_1
timestamp 1762296095
transform -1 0 58130 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 19369
box 0 0 1 1
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_1
timestamp 1762296095
transform -1 0 57515 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 4126
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1762296095
transform 1 0 62228 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1762296095
transform 1 0 49986 0 1 6323
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1762296095
transform 1 0 82808 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_3
timestamp 1762296095
transform 1 0 51732 0 1 5173
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_4
timestamp 1762296095
transform 1 0 72743 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_5
timestamp 1762296095
transform 1 0 72293 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_6
timestamp 1762296095
transform 1 0 23517 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_7
timestamp 1762296095
transform 1 0 13167 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_8
timestamp 1762296095
transform 1 0 12717 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_9
timestamp 1762296095
transform 1 0 2652 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_10
timestamp 1762296095
transform 1 0 40701 0 1 3256
box 0 0 1 1
use M2_M1431059130203_512x8m81  M2_M1431059130203_512x8m81_0
timestamp 1762296095
transform 1 0 25662 0 1 34778
box 0 0 1 1
use M2_M1431059130204_512x8m81  M2_M1431059130204_512x8m81_0
timestamp 1762296095
transform 1 0 25662 0 1 94623
box 0 0 1 1
use M2_M1431059130204_512x8m81  M2_M1431059130204_512x8m81_1
timestamp 1762296095
transform 1 0 59141 0 1 94623
box 0 0 1 1
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1762296095
transform 1 0 60601 0 1 35416
box 0 0 1 1
use M2_M14310591302012_512x8m81  M2_M14310591302012_512x8m81_0
timestamp 1762296095
transform 1 0 27599 0 1 34778
box 0 0 1 1
use m2m3_512x8m81  m2m3_512x8m81_0
timestamp 1762296095
transform 1 0 58611 0 1 17122
box 0 0 3541 9202
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 12783
box 0 0 1 1
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_1
timestamp 1762296095
transform -1 0 57515 0 1 15671
box 0 0 1 1
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 15463
box 0 0 1 1
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 13112
box 0 0 1 1
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_0
timestamp 1762296095
transform -1 0 57515 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_1
timestamp 1762296095
transform -1 0 58130 0 1 8835
box 0 0 1 1
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 8835
box 0 0 1 1
use M3_M2$$201250860_512x8m81  M3_M2$$201250860_512x8m81_0
timestamp 1762296095
transform -1 0 56505 0 1 6590
box 0 0 1 1
use M3_M2$$201250860_512x8m81  M3_M2$$201250860_512x8m81_1
timestamp 1762296095
transform 1 0 28618 0 1 6590
box 0 0 1 1
use M3_M2$$201251884_512x8m81  M3_M2$$201251884_512x8m81_0
timestamp 1762296095
transform 1 0 37303 0 1 35853
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_0
timestamp 1762296095
transform 1 0 28829 0 1 3700
box 0 0 1 1
use M3_M2$$201253932_512x8m81  M3_M2$$201253932_512x8m81_0
timestamp 1762296095
transform 1 0 57515 0 1 8162
box 0 0 1 1
use M3_M2$$201254956_512x8m81  M3_M2$$201254956_512x8m81_0
timestamp 1762296095
transform 1 0 27608 0 1 13768
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_0
timestamp 1762296095
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_1
timestamp 1762296095
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_2
timestamp 1762296095
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_3
timestamp 1762296095
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_4
timestamp 1762296095
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_5
timestamp 1762296095
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_6
timestamp 1762296095
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_7
timestamp 1762296095
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_8
timestamp 1762296095
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_9
timestamp 1762296095
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_10
timestamp 1762296095
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_11
timestamp 1762296095
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_12
timestamp 1762296095
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_13
timestamp 1762296095
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_14
timestamp 1762296095
transform 1 0 28449 0 1 82027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_15
timestamp 1762296095
transform 1 0 28449 0 1 80227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_16
timestamp 1762296095
transform 1 0 28449 0 1 78427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_17
timestamp 1762296095
transform 1 0 28449 0 1 76627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_18
timestamp 1762296095
transform 1 0 28449 0 1 74827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_19
timestamp 1762296095
transform 1 0 28449 0 1 73027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_20
timestamp 1762296095
transform 1 0 28449 0 1 71227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_21
timestamp 1762296095
transform 1 0 28449 0 1 69427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_22
timestamp 1762296095
transform 1 0 28449 0 1 67627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_23
timestamp 1762296095
transform 1 0 28449 0 1 65827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_24
timestamp 1762296095
transform 1 0 28449 0 1 64027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_25
timestamp 1762296095
transform 1 0 28449 0 1 62227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_26
timestamp 1762296095
transform 1 0 28449 0 1 60427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_27
timestamp 1762296095
transform 1 0 28449 0 1 58627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_28
timestamp 1762296095
transform 1 0 28449 0 1 56827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_29
timestamp 1762296095
transform 1 0 28449 0 1 55027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_30
timestamp 1762296095
transform 1 0 28449 0 1 53227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_31
timestamp 1762296095
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_32
timestamp 1762296095
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_33
timestamp 1762296095
transform 1 0 28449 0 1 94627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_34
timestamp 1762296095
transform 1 0 28449 0 1 92827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_35
timestamp 1762296095
transform 1 0 28449 0 1 91027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_36
timestamp 1762296095
transform 1 0 28449 0 1 89227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_37
timestamp 1762296095
transform 1 0 28449 0 1 87427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_38
timestamp 1762296095
transform 1 0 28449 0 1 85627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_39
timestamp 1762296095
transform 1 0 28449 0 1 83827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_40
timestamp 1762296095
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_41
timestamp 1762296095
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_42
timestamp 1762296095
transform 1 0 56674 0 1 53227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_43
timestamp 1762296095
transform 1 0 56674 0 1 55027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_44
timestamp 1762296095
transform 1 0 56674 0 1 56827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_45
timestamp 1762296095
transform 1 0 56674 0 1 58627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_46
timestamp 1762296095
transform 1 0 56674 0 1 60427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_47
timestamp 1762296095
transform 1 0 56674 0 1 62227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_48
timestamp 1762296095
transform 1 0 56674 0 1 64027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_49
timestamp 1762296095
transform 1 0 56674 0 1 65827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_50
timestamp 1762296095
transform 1 0 56674 0 1 67627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_51
timestamp 1762296095
transform 1 0 56674 0 1 69427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_52
timestamp 1762296095
transform 1 0 56674 0 1 71227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_53
timestamp 1762296095
transform 1 0 56674 0 1 73027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_54
timestamp 1762296095
transform 1 0 56674 0 1 74827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_55
timestamp 1762296095
transform 1 0 56674 0 1 76627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_56
timestamp 1762296095
transform 1 0 56674 0 1 78427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_57
timestamp 1762296095
transform 1 0 56674 0 1 80227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_58
timestamp 1762296095
transform 1 0 56674 0 1 82027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_59
timestamp 1762296095
transform 1 0 56674 0 1 83827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_60
timestamp 1762296095
transform 1 0 56674 0 1 85627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_61
timestamp 1762296095
transform 1 0 56674 0 1 87427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_62
timestamp 1762296095
transform 1 0 56674 0 1 89227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_63
timestamp 1762296095
transform 1 0 56674 0 1 91027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_64
timestamp 1762296095
transform 1 0 56674 0 1 92827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_65
timestamp 1762296095
transform 1 0 56674 0 1 94627
box 0 0 1 1
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_0
timestamp 1762296095
transform -1 0 57515 0 1 30897
box 0 0 1 1
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_1
timestamp 1762296095
transform -1 0 57515 0 1 32786
box 0 0 1 1
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 32786
box 0 0 1 1
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_3
timestamp 1762296095
transform 1 0 27608 0 1 30897
box 0 0 1 1
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_1
timestamp 1762296095
transform 1 0 26993 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 7289
box 0 0 1 1
use M3_M2$$201414700_512x8m81  M3_M2$$201414700_512x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 33221
box 0 0 1 1
use M3_M2$$201414700_512x8m81  M3_M2$$201414700_512x8m81_1
timestamp 1762296095
transform 1 0 26993 0 1 33221
box 0 0 1 1
use M3_M2$$201415724_512x8m81  M3_M2$$201415724_512x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 28743
box 0 0 1 1
use M3_M2$$201415724_512x8m81  M3_M2$$201415724_512x8m81_1
timestamp 1762296095
transform 1 0 26993 0 1 28743
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_0
timestamp 1762296095
transform -1 0 57515 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_1
timestamp 1762296095
transform -1 0 58130 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_2
timestamp 1762296095
transform -1 0 57515 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_3
timestamp 1762296095
transform -1 0 58130 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_4
timestamp 1762296095
transform -1 0 57515 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_5
timestamp 1762296095
transform 1 0 27608 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_6
timestamp 1762296095
transform 1 0 26993 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_7
timestamp 1762296095
transform 1 0 27608 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_8
timestamp 1762296095
transform 1 0 26993 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_9
timestamp 1762296095
transform 1 0 27608 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_10
timestamp 1762296095
transform 1 0 27608 0 1 24891
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_0
timestamp 1762296095
transform 0 -1 49977 1 0 8925
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1762296095
transform 1 0 51794 0 1 9891
box 0 0 1 1
use M3_M2431059130202_512x8m81  M3_M2431059130202_512x8m81_0
timestamp 1762296095
transform 1 0 25662 0 1 34778
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_0
timestamp 1762296095
transform 1 0 58128 0 1 20490
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_1
timestamp 1762296095
transform 1 0 58128 0 1 20146
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_2
timestamp 1762296095
transform 1 0 24149 0 1 17237
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_3
timestamp 1762296095
transform 1 0 24496 0 1 23915
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_4
timestamp 1762296095
transform 1 0 24509 0 1 17576
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_5
timestamp 1762296095
transform 1 0 24824 0 1 24236
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_6
timestamp 1762296095
transform 1 0 24837 0 1 17897
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_7
timestamp 1762296095
transform 1 0 25161 0 1 24557
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_8
timestamp 1762296095
transform 1 0 25174 0 1 18270
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_9
timestamp 1762296095
transform 1 0 25501 0 1 25248
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_10
timestamp 1762296095
transform 1 0 25514 0 1 18604
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_11
timestamp 1762296095
transform 1 0 25836 0 1 25567
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_12
timestamp 1762296095
transform 1 0 25851 0 1 18947
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_13
timestamp 1762296095
transform 1 0 26172 0 1 25887
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_14
timestamp 1762296095
transform 1 0 26187 0 1 19267
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_15
timestamp 1762296095
transform 1 0 26530 0 1 26206
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_16
timestamp 1762296095
transform 1 0 26545 0 1 19612
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_17
timestamp 1762296095
transform 1 0 27004 0 1 20490
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_18
timestamp 1762296095
transform 1 0 27004 0 1 20146
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_19
timestamp 1762296095
transform 1 0 24137 0 1 23593
box 0 0 1 1
use M3_M2431059130206_512x8m81  M3_M2431059130206_512x8m81_0
timestamp 1762296095
transform 1 0 27599 0 1 34778
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1762296095
transform 1 0 43880 0 1 3022
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_0
timestamp 1762296095
transform 1 0 59149 0 1 31146
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_1
timestamp 1762296095
transform 1 0 59149 0 1 30701
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_2
timestamp 1762296095
transform 1 0 25674 0 1 31096
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_3
timestamp 1762296095
transform 1 0 25674 0 1 30641
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_4
timestamp 1762296095
transform 1 0 25662 0 1 94623
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_5
timestamp 1762296095
transform 1 0 59141 0 1 94623
box 0 0 1 1
use M3_M24310591302011_512x8m81  M3_M24310591302011_512x8m81_0
timestamp 1762296095
transform 1 0 59154 0 1 34778
box 0 0 1 1
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_0
timestamp 1762296095
transform 1 0 58126 0 1 23631
box 0 0 1 1
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_1
timestamp 1762296095
transform 1 0 57495 0 1 22479
box 0 0 1 1
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_2
timestamp 1762296095
transform 1 0 26990 0 1 23631
box 0 0 1 1
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_3
timestamp 1762296095
transform 1 0 27607 0 1 22492
box 0 0 1 1
use M3_M24310591302015_512x8m81  M3_M24310591302015_512x8m81_0
timestamp 1762296095
transform 1 0 59135 0 1 27399
box 0 0 1 1
use M3_M24310591302015_512x8m81  M3_M24310591302015_512x8m81_1
timestamp 1762296095
transform 1 0 25680 0 1 27421
box 0 0 1 1
use power_a_512x8m81  power_a_512x8m81_0
timestamp 1762296095
transform -1 0 70018 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_1
timestamp 1762296095
transform -1 0 80818 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_2
timestamp 1762296095
transform 1 0 75018 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_3
timestamp 1762296095
transform 1 0 46033 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_4
timestamp 1762296095
transform 1 0 52478 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_5
timestamp 1762296095
transform 1 0 43633 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_6
timestamp 1762296095
transform 1 0 51233 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_7
timestamp 1762296095
transform 1 0 64218 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_8
timestamp 1762296095
transform -1 0 34022 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_9
timestamp 1762296095
transform -1 0 32324 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_10
timestamp 1762296095
transform -1 0 10442 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_11
timestamp 1762296095
transform -1 0 21242 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_12
timestamp 1762296095
transform 1 0 41233 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_13
timestamp 1762296095
transform 1 0 15442 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_14
timestamp 1762296095
transform 1 0 34831 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_15
timestamp 1762296095
transform 1 0 4642 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_16
timestamp 1762296095
transform 1 0 38028 0 1 282
box 0 -282 1000 1000
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_0
timestamp 1762296095
transform 1 0 15448 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_1
timestamp 1762296095
transform 1 0 10048 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_2
timestamp 1762296095
transform 1 0 4648 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_3
timestamp 1762296095
transform 1 0 75024 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_4
timestamp 1762296095
transform 1 0 69624 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_5
timestamp 1762296095
transform 1 0 64224 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_6
timestamp 1762296095
transform 1 0 46824 0 1 94546
box -511 630 1714 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_0
timestamp 1762296095
transform -1 0 41719 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_1
timestamp 1762296095
transform -1 0 39074 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_2
timestamp 1762296095
transform -1 0 35904 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_3
timestamp 1762296095
transform -1 0 31199 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_4
timestamp 1762296095
transform -1 0 27061 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_5
timestamp 1762296095
transform -1 0 21142 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_6
timestamp 1762296095
transform -1 0 80718 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_7
timestamp 1762296095
transform -1 0 58036 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_8
timestamp 1762296095
transform -1 0 85155 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_9
timestamp 1762296095
transform -1 0 54751 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_10
timestamp 1762296095
transform -1 0 49390 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_11
timestamp 1762296095
transform -1 0 45558 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_12
timestamp 1762296095
transform -1 0 53058 0 1 94546
box -511 630 489 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_0
timestamp 1762296095
transform -1 0 26872 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_1
timestamp 1762296095
transform -1 0 41596 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_2
timestamp 1762296095
transform -1 0 38662 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_3
timestamp 1762296095
transform -1 0 35738 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_4
timestamp 1762296095
transform -1 0 34095 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_5
timestamp 1762296095
transform -1 0 30987 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_6
timestamp 1762296095
transform -1 0 29591 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_7
timestamp 1762296095
transform -1 0 60505 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_8
timestamp 1762296095
transform -1 0 52179 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_9
timestamp 1762296095
transform -1 0 45427 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_10
timestamp 1762296095
transform -1 0 57704 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_11
timestamp 1762296095
transform -1 0 44144 0 1 94546
box 714 1822 1714 2430
use power_route_512x8m81  power_route_512x8m81_0
timestamp 1762296095
transform 1 0 -1921 0 1 -2063
box 1921 2345 88293 99039
use rcol4_512_512x8m81  rcol4_512_512x8m81_0
timestamp 1762296095
transform 1 0 60511 0 1 5019
box -1090 -3394 24835 89717
use xdec64_512x8m81  xdec64_512x8m81_0
timestamp 1762296095
transform 1 0 28677 0 1 36127
box -3364 -228 31133 58748
<< labels >>
flabel metal3 s 0 93376 1706 94076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 91576 1706 92276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 89776 1706 90476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 87976 1706 88676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 86176 1706 86876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 2626 96368 3626 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 4642 0 5642 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 5362 96368 6362 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 8026 96368 9026 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 9442 0 10442 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 10762 96368 11762 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 13426 96368 14426 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 15442 0 16442 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 84376 1706 85076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 82576 1706 83276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 80776 1706 81476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 78976 1706 79676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 77176 1706 77876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 75376 1706 76076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 73576 1706 74276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 71776 1706 72476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 16162 96368 17162 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 18826 96368 19826 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 20242 0 21242 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 22258 96368 23258 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 25158 96368 26158 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 26435 3011 28416 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 6921 26434 8163 28412 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 69976 1706 70676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 68176 1706 68876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 66376 1706 67076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 64576 1706 65276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 62776 1706 63476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 17721 26434 18963 28412 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 60976 1706 61676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 26435 26070 28412 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 59176 1706 59876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 23425 26434 27828 26890 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 10176 3011 11493 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2249 10174 24250 11491 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2229 10175 24250 11491 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 24047 10176 27828 11493 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 34536 1014 35326 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 35126 24917 35326 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 34536 27830 35016 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 27877 96368 28877 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 57376 1706 58076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 55576 1706 56276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 53776 1706 54476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 51976 1706 52676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 50176 1706 50876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 48376 1706 49076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 46576 1706 47276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 44776 1706 45476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 42976 1706 43676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29273 96368 30273 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 31324 0 32324 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 32381 96368 33381 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 33022 0 34022 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 34024 96368 35024 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 34831 0 35831 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 41176 1706 41876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 39376 1706 40076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 37576 1706 38276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 35776 1706 36476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 8152 1014 9515 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 8152 3011 9514 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 36948 96368 37948 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 38028 0 39028 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 39882 96368 40882 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 41233 0 42233 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 42430 96368 43430 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 43633 0 44633 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 43713 96368 44713 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 46033 0 47033 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 47538 96368 48538 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2226 8154 28729 9515 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 8153 24250 9514 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 28178 7084 28729 9516 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 24047 8154 28729 9516 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29537 6744 34622 7652 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 28178 7084 34622 7652 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 1401 95176 2401 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 4137 95176 5137 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 6801 95176 7801 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 9537 95176 10537 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50465 96368 51465 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 51233 0 52233 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 12201 95176 13201 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 52478 0 53478 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 55990 96368 56990 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58791 96368 59791 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 62202 96368 63202 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 14937 95176 15937 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 17601 95176 18601 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 20653 95176 21653 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 23483 95176 24483 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26572 95176 27572 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30710 95176 31710 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 35415 95176 36415 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 38585 95176 39585 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 41230 95176 42230 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 64218 0 65218 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 64938 96368 65938 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 67602 96368 68602 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 69018 0 70018 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 70338 96368 71338 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 73002 96368 74002 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 75018 0 76018 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 75738 96368 76738 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 78402 96368 79402 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 45069 95176 46069 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 46313 95176 47313 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 79818 0 80818 932 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 48901 95176 49901 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 52569 95176 53569 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 81834 96368 82834 96976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 94276 1014 94976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 25376 94461 25948 94785 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 94476 27272 94776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30402 94526 54622 94728 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 94527 86372 94728 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58855 94461 59427 94785 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58855 94476 86372 94776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 94276 86372 94976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 54262 95176 55262 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57547 95176 58547 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 92476 1014 93176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 60977 95176 61977 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 92676 27272 92976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 63713 95176 64713 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 66377 95176 67377 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 69113 95176 70113 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 71777 95176 72777 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 74513 95176 75513 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 77177 95176 78177 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 80229 95176 81229 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 83059 95176 84059 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 92726 54622 92928 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 95176 85666 96976 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 92727 86372 92928 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 95176 86372 96176 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 92676 86372 92976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 93376 86372 94076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 92476 86372 93176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 91576 86372 92276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 90676 1014 91376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 90876 27272 91176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 90926 54622 91128 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 90927 86372 91128 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59421 90876 86372 91176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 90676 86372 91376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 88876 1014 89576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 89776 86372 90476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 87976 86372 88676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 86176 86372 86876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 89076 27272 89376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 89126 54622 89328 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 89127 86372 89328 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59421 89076 86372 89376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 84376 86372 85076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 82576 86372 83276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 80776 86372 81476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 78976 86372 79676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 77176 86372 77876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 75376 86372 76076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 73576 86372 74276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 71776 86372 72476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 69976 86372 70676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 68176 86372 68876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 66376 86372 67076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 64576 86372 65276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 62776 86372 63476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 88876 86372 89576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 60976 86372 61676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 87076 1014 87776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 87276 27272 87576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 59176 86372 59876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 57376 86372 58076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 55576 86372 56276 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 53776 86372 54476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 51976 86372 52676 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 50176 86372 50876 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 48376 86372 49076 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 46576 86372 47276 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 87326 54622 87528 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 44776 86372 45476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 87327 86372 87528 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 42976 86372 43676 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 87276 86372 87576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 41176 86372 41876 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 39376 86372 40076 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 87076 86372 87776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 85276 1014 85976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 37576 86372 38276 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 35776 86372 36476 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 29430 1706 34125 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 85476 27272 85776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 85526 54622 85728 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 85527 86372 85728 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2095 32315 2188 34126 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 32315 3011 34125 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 85476 86372 85776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 85276 86372 85976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 32316 25085 34125 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 32318 27214 34124 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 83476 1014 84176 0 FreeSans 448 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 83676 27272 83976 0 FreeSans 448 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 83726 54622 83928 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 83727 86372 83928 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59421 83676 86372 83976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26772 31486 58351 32199 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26772 27382 58351 30105 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 31486 58351 34124 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61853 32315 72383 34125 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 32315 86372 34124 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 83476 86372 84176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 81676 1014 82376 0 FreeSans 448 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 81876 27272 82176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 81926 54622 82128 0 FreeSans 448 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 29430 86372 29714 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 81927 86372 82128 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 29430 86372 34125 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 72653 32315 86372 34125 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 22938 1706 23938 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 22938 27214 23380 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26770 23370 58348 24278 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 22937 83763 23380 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 22938 86372 23380 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 22938 86372 23938 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 81876 86372 82176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 18016 24250 20739 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 81676 86372 82376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 29513 19969 55645 21625 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 79876 1014 80576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 29521 19969 55645 21707 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 80076 27272 80376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 80126 54622 80328 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 80127 86372 80328 0 FreeSans 448 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 44432 19969 55645 21708 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61825 18015 83763 20739 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61807 18016 86372 20739 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 19969 86372 20739 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 12036 1706 14178 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 23821 12046 34761 12847 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 13461 27214 14178 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 12036 24250 12846 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 24047 12046 27214 14179 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 24047 12046 34761 12934 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 34741 9972 41516 12570 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29478 10756 41516 12570 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29478 11697 58351 12570 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26772 11844 58351 12570 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50228 12035 58421 13866 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59826 12035 60026 14017 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50228 13461 86372 13866 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61807 13461 72429 14178 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61773 13461 86372 14177 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 83169 12035 84221 12847 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 83169 13461 84221 14179 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 80076 86372 80376 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 50228 12036 86372 12846 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 79876 86372 80576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 78076 1014 78776 0 FreeSans 448 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 78276 27272 78576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26772 12035 84999 12570 0 FreeSans 448 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 78326 54622 78528 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 78327 86372 78528 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 12036 86372 14178 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 72607 13461 86372 14178 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 78276 86372 78576 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 61802 8153 86372 9514 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 78076 86372 78776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 57909 8154 62278 9516 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 76276 1014 76976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 57909 8154 72434 9515 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 76476 27272 76776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 72602 8152 83234 9515 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 76526 54622 76728 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 61825 8152 86372 9514 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 76527 86372 76728 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 8152 86372 9515 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 76476 86372 76776 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 76276 86372 76976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 4060 1712 5629 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 74476 1014 75176 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 5173 3011 5629 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 74676 27272 74976 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 5174 24250 5629 0 FreeSans 448 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 74726 54622 74928 0 FreeSans 448 0 0 0 VSS
port 30 nsew ground bidirectional
rlabel metal2 s 27936 0 28160 200 4 CLK
port 11 nsew signal input
rlabel metal2 s 1864 0 2088 200 4 D[0]
port 19 nsew signal input
rlabel metal2 s 29006 0 29230 200 4 A[8]
port 1 nsew signal input
rlabel metal2 s 29705 0 29929 200 4 A[7]
port 2 nsew signal input
rlabel metal2 s 30859 0 31083 200 4 A[2]
port 7 nsew signal input
rlabel metal2 s 32552 0 32776 200 4 A[1]
port 8 nsew signal input
rlabel metal2 s 34243 0 34467 200 4 A[0]
port 9 nsew signal input
rlabel metal2 s 14127 0 14351 200 4 Q[2]
port 26 nsew signal output
rlabel metal2 s 22279 0 22503 200 4 Q[3]
port 25 nsew signal output
rlabel metal2 s 50342 0 50566 200 4 CEN
port 10 nsew signal input
rlabel metal2 s 54417 0 54641 200 4 A[5]
port 4 nsew signal input
rlabel metal2 s 53772 0 53996 200 4 A[6]
port 3 nsew signal input
rlabel metal2 s 55164 0 55388 200 4 A[4]
port 5 nsew signal input
rlabel metal2 s 23404 0 23628 200 4 WEN[3]
port 35 nsew signal input
rlabel metal2 s 83372 0 83596 200 4 D[7]
port 12 nsew signal input
rlabel metal2 s 81855 0 82079 200 4 Q[7]
port 21 nsew signal output
rlabel metal2 s 23795 0 24019 200 4 D[3]
port 16 nsew signal input
rlabel metal2 s 12206 0 12430 200 4 D[1]
port 18 nsew signal input
rlabel metal2 s 13454 0 13678 200 4 D[2]
port 17 nsew signal input
rlabel metal2 s 56265 0 56489 200 4 A[3]
port 6 nsew signal input
rlabel metal2 s 11533 0 11757 200 4 Q[1]
port 27 nsew signal output
rlabel metal2 s 73703 0 73927 200 4 Q[6]
port 22 nsew signal output
rlabel metal2 s 71782 0 72006 200 4 D[5]
port 14 nsew signal input
rlabel metal2 s 62958 0 63182 200 4 Q[4]
port 24 nsew signal output
rlabel metal2 s 72180 0 72404 200 4 WEN[5]
port 33 nsew signal input
rlabel metal2 s 13054 0 13278 200 4 WEN[2]
port 36 nsew signal input
rlabel metal2 s 12604 0 12828 200 4 WEN[1]
port 37 nsew signal input
rlabel metal2 s 62115 0 62339 200 4 WEN[4]
port 34 nsew signal input
rlabel metal2 s 82695 0 82919 200 4 WEN[7]
port 31 nsew signal input
rlabel metal2 s 72630 0 72854 200 4 WEN[6]
port 32 nsew signal input
rlabel metal2 s 61447 0 61671 200 4 D[4]
port 15 nsew signal input
rlabel metal2 s 73030 0 73254 200 4 D[6]
port 13 nsew signal input
rlabel metal2 s 71109 0 71333 200 4 Q[5]
port 23 nsew signal output
rlabel metal2 s 3380 0 3604 200 4 Q[0]
port 28 nsew signal output
rlabel metal2 s 40588 0 40812 200 4 GWEN
port 20 nsew signal input
rlabel metal2 s 2539 0 2763 200 4 WEN[0]
port 38 nsew signal input
rlabel metal3 s 0 4060 24341 4515 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 74727 86372 74928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 74676 86372 74976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 74476 86372 75176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72676 1014 73376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72876 27272 73176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 72926 54622 73128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72927 86372 73128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 72876 86372 73176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 72676 86372 73376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 70876 1014 71576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 71076 27272 71376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 71126 54622 71328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 71127 86372 71328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 71076 86372 71376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 70876 86372 71576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69076 1014 69776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69276 27272 69576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 69326 54622 69528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69327 86372 69528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 69276 86372 69576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 69076 86372 69776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67276 1014 67976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67476 27272 67776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 67526 54622 67728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67527 86372 67728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 67476 86372 67776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 67276 86372 67976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65476 1014 66176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65676 27272 65976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 65726 54622 65928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65727 86372 65928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 65676 86372 65976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 65476 86372 66176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63676 1014 64376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63876 27272 64176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 63926 54622 64128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63927 86372 64128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 63876 86372 64176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 63676 86372 64376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 61876 1014 62576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 62076 27272 62376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 62126 54622 62328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 62127 86372 62328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 62076 86372 62376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 61876 86372 62576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60076 1014 60776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60276 27272 60576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 60326 54622 60528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60327 86372 60528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 60276 86372 60576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 60076 86372 60776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58276 1014 58976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58476 27272 58776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 58526 54622 58728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58527 86372 58728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 58476 86372 58776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 58276 86372 58976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56476 1014 57176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56676 27272 56976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 56726 54622 56928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56727 86372 56928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 56676 86372 56976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 56476 86372 57176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54676 1014 55376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54876 27272 55176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 54926 54622 55128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54927 86372 55128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 54876 86372 55176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 54676 86372 55376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 52876 1014 53576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 53076 27272 53376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 53126 54622 53328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 53127 86372 53328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 53076 86372 53376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 52876 86372 53576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51076 1014 51776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51276 27272 51576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 51326 54622 51528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51327 86372 51528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 51276 86372 51576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 51076 86372 51776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49276 1014 49976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49476 27272 49776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 49526 54622 49728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49527 86372 49728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 49476 86372 49776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 49276 86372 49976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47476 1014 48176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47676 27272 47976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 47726 54622 47928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47727 86372 47928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 47676 86372 47976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 47476 86372 48176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45676 1014 46376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45876 27272 46176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 45926 54622 46128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45927 86372 46128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 45876 86372 46176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 45676 86372 46376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 43876 1014 44576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 44076 27272 44376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 44127 86372 44328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 44076 86372 44376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42327 86372 42528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40527 86372 40728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38727 86372 38928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36927 86372 37128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 60460 35158 86372 35298 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58791 34536 86372 35016 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 34536 86372 35326 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83360 35126 86372 35326 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 66497 26434 67739 28412 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 77297 26434 78539 28412 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28412 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 26435 86372 28416 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21826 57681 23199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 22291 57681 23199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42261 10740 86372 11491 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8930 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 2502 1014 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 1 VSS
port 30 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 96976
string GDS_END 2941248
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2875980
string LEFclass BLOCK
string LEFsymmetry X Y R90
string path 232.665 4.660 232.665 0.000 
<< end >>
