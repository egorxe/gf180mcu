magic
tech gf180mcuD
timestamp 1762296095
<< properties >>
string GDS_END 273530
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 273174
<< end >>
