magic
tech gf180mcuD
timestamp 1759194789
<< properties >>
string GDS_END 7919528
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 7685348
<< end >>
