magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_0
timestamp 1762296095
transform -1 0 85672 0 1 96288
box 0 0 1 1
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_1
timestamp 1762296095
transform -1 0 85672 0 1 620
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_0
timestamp 1762296095
transform 1 0 85474 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_1
timestamp 1762296095
transform 1 0 27139 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_2
timestamp 1762296095
transform 1 0 57047 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_3
timestamp 1762296095
transform 1 0 112 0 1 1140
box 0 0 1 1
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_0
timestamp 1762296095
transform 1 0 56123 0 1 36019
box 0 0 1 1
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_1
timestamp 1762296095
transform 1 0 27563 0 1 36019
box 0 0 1 1
use M1_PSUB4310591302046_512x8m81  M1_PSUB4310591302046_512x8m81_0
timestamp 1762296095
transform 1 0 27563 0 1 34197
box 0 0 1 1
<< properties >>
string GDS_END 2641408
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2640098
string path 4.620 11.160 4.620 0.000 
<< end >>
