magic
tech gf180mcuD
timestamp 1759194789
<< properties >>
string GDS_END 9504374
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 9255474
<< end >>
