magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< psubdiff >>
rect 13097 70975 69968 71000
rect 13097 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69968 70975
rect 13097 70871 69968 70929
rect 13097 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69968 70871
rect 13097 70803 69968 70825
rect 13097 70767 13291 70803
rect 13097 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13291 70767
rect 13097 70663 13291 70721
rect 13097 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13291 70663
rect 13097 70559 13291 70617
rect 13097 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13291 70559
rect 13097 70455 13291 70513
rect 13097 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13291 70455
rect 13097 70351 13291 70409
rect 13097 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13291 70351
rect 13097 70247 13291 70305
rect 13097 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13291 70247
rect 13097 70143 13291 70201
rect 13097 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13291 70143
rect 13097 70039 13291 70097
rect 13097 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13291 70039
rect 13097 69935 13291 69993
rect 13097 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13291 69935
rect 13097 69831 13291 69889
rect 13097 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13291 69831
rect 13097 69727 13291 69785
rect 69774 70720 69968 70803
rect 69774 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69968 70720
rect 69774 70616 69968 70674
rect 69774 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69968 70616
rect 69774 70512 69968 70570
rect 69774 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69968 70512
rect 69774 70408 69968 70466
rect 69774 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69968 70408
rect 69774 70304 69968 70362
rect 69774 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69968 70304
rect 69774 70200 69968 70258
rect 69774 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69968 70200
rect 69774 70096 69968 70154
rect 69774 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69968 70096
rect 69774 69968 69968 70050
rect 69774 69946 71000 69968
rect 69774 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69774 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69774 69842 71000 69862
rect 69774 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69774 69774 70824 69796
rect 13097 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13291 69727
rect 13097 69623 13291 69681
rect 13097 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13291 69623
rect 13097 69519 13291 69577
rect 13097 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13291 69519
rect 13097 69415 13291 69473
rect 13097 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13291 69415
rect 13097 69311 13291 69369
rect 13097 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13291 69311
rect 13097 69207 13291 69265
rect 13097 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13291 69207
rect 13097 69103 13291 69161
rect 13097 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13291 69103
rect 13097 68999 13291 69057
rect 13097 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13291 68999
rect 13097 68895 13291 68953
rect 13097 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13291 68895
rect 13097 68791 13291 68849
rect 13097 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13291 68791
rect 13097 68687 13291 68745
rect 13097 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13291 68687
rect 13097 68583 13291 68641
rect 13097 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13291 68583
rect 13097 68479 13291 68537
rect 13097 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13291 68479
rect 13097 68375 13291 68433
rect 13097 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13291 68375
rect 13097 68271 13291 68329
rect 13097 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13291 68271
rect 13097 68167 13291 68225
rect 13097 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13291 68167
rect 13097 68063 13291 68121
rect 13097 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13291 68063
rect 13097 67959 13291 68017
rect 13097 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13291 67959
rect 13097 67855 13291 67913
rect 13097 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13291 67855
rect 13097 67751 13291 67809
rect 13097 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13291 67751
rect 13097 67647 13291 67705
rect 13097 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13291 67647
rect 13097 67543 13291 67601
rect 13097 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13291 67543
rect 13097 67439 13291 67497
rect 13097 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13291 67439
rect 13097 67335 13291 67393
rect 13097 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13291 67335
rect 13097 67231 13291 67289
rect 13097 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13291 67231
rect 13097 67127 13291 67185
rect 13097 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13291 67127
rect 13097 67023 13291 67081
rect 13097 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13291 67023
rect 13097 66919 13291 66977
rect 13097 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13291 66919
rect 13097 66815 13291 66873
rect 13097 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13291 66815
rect 13097 66711 13291 66769
rect 13097 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13291 66711
rect 13097 66607 13291 66665
rect 13097 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13291 66607
rect 13097 66503 13291 66561
rect 13097 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13291 66503
rect 13097 66399 13291 66457
rect 13097 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13291 66399
rect 13097 66295 13291 66353
rect 13097 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13291 66295
rect 13097 66191 13291 66249
rect 13097 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13291 66191
rect 13097 66087 13291 66145
rect 13097 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13291 66087
rect 13097 65983 13291 66041
rect 13097 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13291 65983
rect 13097 65879 13291 65937
rect 13097 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13291 65879
rect 13097 65775 13291 65833
rect 13097 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13291 65775
rect 13097 65671 13291 65729
rect 13097 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13291 65671
rect 13097 65567 13291 65625
rect 13097 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13291 65567
rect 13097 65463 13291 65521
rect 13097 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13291 65463
rect 13097 65359 13291 65417
rect 13097 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13291 65359
rect 13097 65255 13291 65313
rect 13097 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13291 65255
rect 13097 65151 13291 65209
rect 13097 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13291 65151
rect 13097 65047 13291 65105
rect 13097 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13291 65047
rect 13097 64943 13291 65001
rect 13097 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13291 64943
rect 13097 64839 13291 64897
rect 13097 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13291 64839
rect 13097 64735 13291 64793
rect 13097 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13291 64735
rect 13097 64631 13291 64689
rect 13097 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13291 64631
rect 13097 64527 13291 64585
rect 13097 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13291 64527
rect 13097 64423 13291 64481
rect 13097 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13291 64423
rect 13097 64319 13291 64377
rect 13097 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13291 64319
rect 13097 64215 13291 64273
rect 13097 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13291 64215
rect 13097 64111 13291 64169
rect 13097 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13291 64111
rect 13097 64007 13291 64065
rect 13097 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13291 64007
rect 13097 63903 13291 63961
rect 13097 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13291 63903
rect 13097 63799 13291 63857
rect 13097 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13291 63799
rect 13097 63695 13291 63753
rect 13097 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13291 63695
rect 13097 63591 13291 63649
rect 13097 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13291 63591
rect 13097 63487 13291 63545
rect 13097 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13291 63487
rect 13097 63383 13291 63441
rect 13097 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13291 63383
rect 13097 63279 13291 63337
rect 13097 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13291 63279
rect 13097 63175 13291 63233
rect 13097 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13291 63175
rect 13097 63071 13291 63129
rect 13097 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13291 63071
rect 13097 62967 13291 63025
rect 13097 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13291 62967
rect 13097 62863 13291 62921
rect 13097 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13291 62863
rect 13097 62759 13291 62817
rect 13097 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13291 62759
rect 13097 62655 13291 62713
rect 13097 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13291 62655
rect 13097 62551 13291 62609
rect 13097 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13291 62551
rect 13097 62447 13291 62505
rect 13097 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13291 62447
rect 13097 62343 13291 62401
rect 13097 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13291 62343
rect 13097 62239 13291 62297
rect 13097 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13291 62239
rect 13097 62135 13291 62193
rect 13097 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13291 62135
rect 13097 62031 13291 62089
rect 13097 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13291 62031
rect 13097 61927 13291 61985
rect 13097 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13291 61927
rect 13097 61823 13291 61881
rect 13097 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13291 61823
rect 13097 61719 13291 61777
rect 13097 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13291 61719
rect 13097 61615 13291 61673
rect 13097 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13291 61615
rect 13097 61511 13291 61569
rect 13097 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13291 61511
rect 13097 61407 13291 61465
rect 13097 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13291 61407
rect 13097 61303 13291 61361
rect 13097 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13291 61303
rect 13097 61199 13291 61257
rect 13097 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13291 61199
rect 13097 61095 13291 61153
rect 13097 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13291 61095
rect 13097 60991 13291 61049
rect 13097 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13291 60991
rect 13097 60887 13291 60945
rect 13097 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13291 60887
rect 13097 60783 13291 60841
rect 13097 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13291 60783
rect 13097 60679 13291 60737
rect 13097 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13291 60679
rect 13097 60575 13291 60633
rect 13097 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13291 60575
rect 13097 60471 13291 60529
rect 13097 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13291 60471
rect 13097 60367 13291 60425
rect 13097 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13291 60367
rect 13097 60263 13291 60321
rect 13097 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13291 60263
rect 13097 60159 13291 60217
rect 13097 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13291 60159
rect 13097 60055 13291 60113
rect 13097 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13291 60055
rect 13097 59951 13291 60009
rect 13097 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13291 59951
rect 13097 59847 13291 59905
rect 13097 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13291 59847
rect 13097 59743 13291 59801
rect 13097 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13291 59743
rect 13097 59639 13291 59697
rect 13097 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13291 59639
rect 13097 59535 13291 59593
rect 13097 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13291 59535
rect 13097 59431 13291 59489
rect 13097 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13291 59431
rect 13097 59327 13291 59385
rect 13097 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13291 59327
rect 13097 59223 13291 59281
rect 13097 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13291 59223
rect 13097 59119 13291 59177
rect 13097 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13291 59119
rect 13097 59015 13291 59073
rect 13097 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13291 59015
rect 13097 58911 13291 58969
rect 13097 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13291 58911
rect 13097 58807 13291 58865
rect 13097 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13291 58807
rect 13097 58703 13291 58761
rect 13097 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13291 58703
rect 13097 58599 13291 58657
rect 13097 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13291 58599
rect 13097 58495 13291 58553
rect 13097 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13291 58495
rect 13097 58391 13291 58449
rect 13097 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13291 58391
rect 13097 58287 13291 58345
rect 13097 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13291 58287
rect 13097 58183 13291 58241
rect 13097 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13291 58183
rect 13097 58079 13291 58137
rect 13097 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13291 58079
rect 13097 57975 13291 58033
rect 13097 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13291 57975
rect 13097 57871 13291 57929
rect 13097 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13291 57871
rect 13097 57767 13291 57825
rect 13097 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13291 57767
rect 13097 57663 13291 57721
rect 13097 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13291 57663
rect 13097 57559 13291 57617
rect 13097 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13291 57559
rect 13097 57455 13291 57513
rect 13097 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13291 57455
rect 13097 57351 13291 57409
rect 13097 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13291 57351
rect 13097 57247 13291 57305
rect 13097 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13291 57247
rect 13097 57143 13291 57201
rect 13097 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13291 57143
rect 13097 57039 13291 57097
rect 13097 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13291 57039
rect 13097 56935 13291 56993
rect 13097 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13291 56935
rect 13097 56831 13291 56889
rect 13097 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13291 56831
rect 13097 56727 13291 56785
rect 13097 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13291 56727
rect 13097 56623 13291 56681
rect 13097 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13291 56623
rect 13097 56519 13291 56577
rect 13097 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13291 56519
rect 13097 56415 13291 56473
rect 13097 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13291 56415
rect 13097 56311 13291 56369
rect 13097 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13291 56311
rect 13097 56207 13291 56265
rect 13097 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13291 56207
rect 13097 56103 13291 56161
rect 13097 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13291 56103
rect 13097 55999 13291 56057
rect 13097 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13291 55999
rect 13097 55895 13291 55953
rect 13097 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13291 55895
rect 13097 55791 13291 55849
rect 13097 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13291 55791
rect 13097 55687 13291 55745
rect 13097 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13291 55687
rect 13097 55583 13291 55641
rect 13097 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13291 55583
rect 13097 55479 13291 55537
rect 13097 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13291 55479
rect 13097 55375 13291 55433
rect 13097 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13291 55375
rect 13097 55271 13291 55329
rect 13097 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13291 55271
rect 13097 55167 13291 55225
rect 13097 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13291 55167
rect 13097 55063 13291 55121
rect 13097 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13291 55063
rect 13097 54959 13291 55017
rect 13097 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13291 54959
rect 13097 54855 13291 54913
rect 13097 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13291 54855
rect 13097 54751 13291 54809
rect 13097 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13291 54751
rect 13097 54647 13291 54705
rect 13097 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13291 54647
rect 13097 54543 13291 54601
rect 13097 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13291 54543
rect 13097 54439 13291 54497
rect 13097 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13291 54439
rect 13097 54335 13291 54393
rect 13097 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13291 54335
rect 13097 54231 13291 54289
rect 13097 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13291 54231
rect 13097 54127 13291 54185
rect 13097 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13291 54127
rect 13097 54023 13291 54081
rect 13097 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13291 54023
rect 13097 53919 13291 53977
rect 13097 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13291 53919
rect 13097 53815 13291 53873
rect 13097 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13291 53815
rect 13097 53711 13291 53769
rect 13097 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13291 53711
rect 13097 53607 13291 53665
rect 13097 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13291 53607
rect 13097 53503 13291 53561
rect 13097 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13291 53503
rect 13097 53399 13291 53457
rect 13097 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13291 53399
rect 13097 53295 13291 53353
rect 13097 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13291 53295
rect 13097 53191 13291 53249
rect 13097 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13291 53191
rect 13097 53087 13291 53145
rect 13097 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13291 53087
rect 13097 52983 13291 53041
rect 13097 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13291 52983
rect 13097 52879 13291 52937
rect 13097 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13291 52879
rect 13097 52775 13291 52833
rect 13097 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13291 52775
rect 13097 52671 13291 52729
rect 13097 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13291 52671
rect 13097 52567 13291 52625
rect 13097 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13291 52567
rect 13097 52463 13291 52521
rect 13097 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13291 52463
rect 13097 52359 13291 52417
rect 13097 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13291 52359
rect 13097 52255 13291 52313
rect 13097 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13291 52255
rect 13097 52151 13291 52209
rect 13097 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13291 52151
rect 13097 52047 13291 52105
rect 13097 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13291 52047
rect 13097 51943 13291 52001
rect 13097 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13291 51943
rect 13097 51839 13291 51897
rect 13097 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13291 51839
rect 13097 51735 13291 51793
rect 13097 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13291 51735
rect 13097 51631 13291 51689
rect 13097 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13291 51631
rect 13097 51527 13291 51585
rect 13097 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13291 51527
rect 13097 51423 13291 51481
rect 13097 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13291 51423
rect 13097 51319 13291 51377
rect 13097 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13291 51319
rect 13097 51215 13291 51273
rect 13097 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13291 51215
rect 13097 51111 13291 51169
rect 13097 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13291 51111
rect 13097 51007 13291 51065
rect 13097 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13291 51007
rect 13097 50903 13291 50961
rect 13097 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13291 50903
rect 13097 50799 13291 50857
rect 13097 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13291 50799
rect 13097 50695 13291 50753
rect 13097 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13291 50695
rect 13097 50591 13291 50649
rect 13097 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13291 50591
rect 13097 50487 13291 50545
rect 13097 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13291 50487
rect 13097 50383 13291 50441
rect 13097 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13291 50383
rect 13097 50279 13291 50337
rect 13097 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13291 50279
rect 13097 50175 13291 50233
rect 13097 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13291 50175
rect 13097 50071 13291 50129
rect 13097 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13291 50071
rect 13097 49967 13291 50025
rect 13097 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13291 49967
rect 13097 49863 13291 49921
rect 13097 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13291 49863
rect 13097 49759 13291 49817
rect 13097 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13291 49759
rect 13097 49655 13291 49713
rect 13097 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13291 49655
rect 13097 49551 13291 49609
rect 13097 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13291 49551
rect 13097 49447 13291 49505
rect 13097 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13291 49447
rect 13097 49343 13291 49401
rect 13097 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13291 49343
rect 13097 49239 13291 49297
rect 13097 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13291 49239
rect 13097 49135 13291 49193
rect 13097 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13291 49135
rect 13097 49031 13291 49089
rect 13097 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13291 49031
rect 13097 48927 13291 48985
rect 13097 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13291 48927
rect 13097 48823 13291 48881
rect 13097 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13291 48823
rect 13097 48719 13291 48777
rect 13097 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13291 48719
rect 13097 48615 13291 48673
rect 13097 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13291 48615
rect 13097 48511 13291 48569
rect 13097 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13291 48511
rect 13097 48407 13291 48465
rect 13097 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13291 48407
rect 13097 48303 13291 48361
rect 13097 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13291 48303
rect 13097 48199 13291 48257
rect 13097 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13291 48199
rect 13097 48095 13291 48153
rect 13097 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13291 48095
rect 13097 47991 13291 48049
rect 13097 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13291 47991
rect 13097 47887 13291 47945
rect 13097 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13291 47887
rect 13097 47783 13291 47841
rect 13097 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13291 47783
rect 13097 47679 13291 47737
rect 13097 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13291 47679
rect 13097 47575 13291 47633
rect 13097 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13291 47575
rect 13097 47471 13291 47529
rect 13097 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13291 47471
rect 13097 47367 13291 47425
rect 13097 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13291 47367
rect 13097 47263 13291 47321
rect 13097 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13291 47263
rect 13097 47159 13291 47217
rect 13097 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13291 47159
rect 13097 47055 13291 47113
rect 13097 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13291 47055
rect 13097 46951 13291 47009
rect 13097 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13291 46951
rect 13097 46847 13291 46905
rect 13097 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13291 46847
rect 13097 46743 13291 46801
rect 13097 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13291 46743
rect 13097 46639 13291 46697
rect 13097 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13291 46639
rect 13097 46535 13291 46593
rect 13097 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13291 46535
rect 13097 46431 13291 46489
rect 13097 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13291 46431
rect 13097 46327 13291 46385
rect 13097 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13291 46327
rect 13097 46223 13291 46281
rect 13097 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13291 46223
rect 13097 46119 13291 46177
rect 13097 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13291 46119
rect 13097 46015 13291 46073
rect 13097 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13291 46015
rect 13097 45911 13291 45969
rect 13097 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13291 45911
rect 13097 45807 13291 45865
rect 13097 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13291 45807
rect 13097 45703 13291 45761
rect 13097 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13291 45703
rect 13097 45599 13291 45657
rect 13097 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13291 45599
rect 13097 45495 13291 45553
rect 13097 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13291 45495
rect 13097 45391 13291 45449
rect 13097 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13291 45391
rect 13097 45287 13291 45345
rect 13097 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13291 45287
rect 13097 45183 13291 45241
rect 13097 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13291 45183
rect 13097 45079 13291 45137
rect 13097 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13291 45079
rect 13097 44893 13291 45033
rect 70802 69758 70824 69774
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70802 69700 71000 69758
rect 70802 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70802 69596 71000 69654
rect 70802 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70802 69492 71000 69550
rect 70802 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70802 69388 71000 69446
rect 70802 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70802 69284 71000 69342
rect 70802 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70802 69180 71000 69238
rect 70802 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70802 69076 71000 69134
rect 70802 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70802 68972 71000 69030
rect 70802 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70802 68868 71000 68926
rect 70802 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70802 68764 71000 68822
rect 70802 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70802 68660 71000 68718
rect 70802 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70802 68556 71000 68614
rect 70802 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70802 68452 71000 68510
rect 70802 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70802 68348 71000 68406
rect 70802 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70802 68244 71000 68302
rect 70802 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70802 68140 71000 68198
rect 70802 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70802 68036 71000 68094
rect 70802 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70802 67932 71000 67990
rect 70802 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70802 67828 71000 67886
rect 70802 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70802 67724 71000 67782
rect 70802 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70802 67620 71000 67678
rect 70802 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70802 67516 71000 67574
rect 70802 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70802 67412 71000 67470
rect 70802 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70802 67308 71000 67366
rect 70802 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70802 67204 71000 67262
rect 70802 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70802 67100 71000 67158
rect 70802 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70802 66996 71000 67054
rect 70802 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70802 66892 71000 66950
rect 70802 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70802 66788 71000 66846
rect 70802 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70802 66684 71000 66742
rect 70802 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70802 66580 71000 66638
rect 70802 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70802 66476 71000 66534
rect 70802 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70802 66372 71000 66430
rect 70802 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70802 66268 71000 66326
rect 70802 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70802 66164 71000 66222
rect 70802 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70802 66060 71000 66118
rect 70802 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70802 65956 71000 66014
rect 70802 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70802 65852 71000 65910
rect 70802 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70802 65748 71000 65806
rect 70802 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70802 65644 71000 65702
rect 70802 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70802 65540 71000 65598
rect 70802 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70802 65436 71000 65494
rect 70802 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70802 65332 71000 65390
rect 70802 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70802 65228 71000 65286
rect 70802 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70802 65124 71000 65182
rect 70802 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70802 65020 71000 65078
rect 70802 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70802 64916 71000 64974
rect 70802 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70802 64812 71000 64870
rect 70802 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70802 64708 71000 64766
rect 70802 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70802 64604 71000 64662
rect 70802 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70802 64500 71000 64558
rect 70802 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70802 64396 71000 64454
rect 70802 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70802 64292 71000 64350
rect 70802 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70802 64188 71000 64246
rect 70802 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70802 64084 71000 64142
rect 70802 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70802 63980 71000 64038
rect 70802 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70802 63876 71000 63934
rect 70802 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70802 63772 71000 63830
rect 70802 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70802 63668 71000 63726
rect 70802 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70802 63564 71000 63622
rect 70802 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70802 63460 71000 63518
rect 70802 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70802 63356 71000 63414
rect 70802 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70802 63252 71000 63310
rect 70802 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70802 63148 71000 63206
rect 70802 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70802 63044 71000 63102
rect 70802 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70802 62940 71000 62998
rect 70802 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70802 62836 71000 62894
rect 70802 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70802 62732 71000 62790
rect 70802 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70802 62628 71000 62686
rect 70802 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70802 62524 71000 62582
rect 70802 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70802 62420 71000 62478
rect 70802 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70802 62316 71000 62374
rect 70802 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70802 62212 71000 62270
rect 70802 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70802 62108 71000 62166
rect 70802 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70802 62004 71000 62062
rect 70802 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70802 61900 71000 61958
rect 70802 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70802 61796 71000 61854
rect 70802 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70802 61692 71000 61750
rect 70802 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70802 61588 71000 61646
rect 70802 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70802 61484 71000 61542
rect 70802 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70802 61380 71000 61438
rect 70802 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70802 61276 71000 61334
rect 70802 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70802 61172 71000 61230
rect 70802 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70802 61068 71000 61126
rect 70802 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70802 60964 71000 61022
rect 70802 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70802 60860 71000 60918
rect 70802 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70802 60756 71000 60814
rect 70802 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70802 60652 71000 60710
rect 70802 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70802 60548 71000 60606
rect 70802 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70802 60444 71000 60502
rect 70802 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70802 60340 71000 60398
rect 70802 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70802 60236 71000 60294
rect 70802 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70802 60132 71000 60190
rect 70802 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70802 60028 71000 60086
rect 70802 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70802 59924 71000 59982
rect 70802 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70802 59820 71000 59878
rect 70802 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70802 59716 71000 59774
rect 70802 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70802 59612 71000 59670
rect 70802 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70802 59508 71000 59566
rect 70802 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70802 59404 71000 59462
rect 70802 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70802 59300 71000 59358
rect 70802 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70802 59196 71000 59254
rect 70802 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70802 59092 71000 59150
rect 70802 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70802 58988 71000 59046
rect 70802 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70802 58884 71000 58942
rect 70802 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70802 58780 71000 58838
rect 70802 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70802 58676 71000 58734
rect 70802 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70802 58572 71000 58630
rect 70802 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70802 58468 71000 58526
rect 70802 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70802 58364 71000 58422
rect 70802 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70802 58260 71000 58318
rect 70802 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70802 58156 71000 58214
rect 70802 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70802 58052 71000 58110
rect 70802 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70802 57948 71000 58006
rect 70802 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70802 57844 71000 57902
rect 70802 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70802 57740 71000 57798
rect 70802 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70802 57636 71000 57694
rect 70802 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70802 57532 71000 57590
rect 70802 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70802 57428 71000 57486
rect 70802 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70802 57324 71000 57382
rect 70802 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70802 57220 71000 57278
rect 70802 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70802 57116 71000 57174
rect 70802 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70802 57012 71000 57070
rect 70802 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70802 56908 71000 56966
rect 70802 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70802 56804 71000 56862
rect 70802 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70802 56700 71000 56758
rect 70802 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70802 56596 71000 56654
rect 70802 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70802 56492 71000 56550
rect 70802 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70802 56388 71000 56446
rect 70802 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70802 56284 71000 56342
rect 70802 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70802 56180 71000 56238
rect 70802 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70802 56076 71000 56134
rect 70802 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70802 55972 71000 56030
rect 70802 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70802 55868 71000 55926
rect 70802 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70802 55764 71000 55822
rect 70802 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70802 55660 71000 55718
rect 70802 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70802 55556 71000 55614
rect 70802 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70802 55452 71000 55510
rect 70802 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70802 55348 71000 55406
rect 70802 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70802 55244 71000 55302
rect 70802 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70802 55140 71000 55198
rect 70802 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70802 55036 71000 55094
rect 70802 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70802 54932 71000 54990
rect 70802 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70802 54828 71000 54886
rect 70802 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70802 54724 71000 54782
rect 70802 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70802 54620 71000 54678
rect 70802 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70802 54516 71000 54574
rect 70802 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70802 54412 71000 54470
rect 70802 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70802 54308 71000 54366
rect 70802 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70802 54204 71000 54262
rect 70802 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70802 54100 71000 54158
rect 70802 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70802 53996 71000 54054
rect 70802 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70802 53892 71000 53950
rect 70802 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70802 53788 71000 53846
rect 70802 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70802 53684 71000 53742
rect 70802 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70802 53580 71000 53638
rect 70802 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70802 53476 71000 53534
rect 70802 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70802 53372 71000 53430
rect 70802 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70802 53268 71000 53326
rect 70802 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70802 53164 71000 53222
rect 70802 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70802 53060 71000 53118
rect 70802 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70802 52956 71000 53014
rect 70802 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70802 52852 71000 52910
rect 70802 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70802 52748 71000 52806
rect 70802 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70802 52644 71000 52702
rect 70802 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70802 52540 71000 52598
rect 70802 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70802 52436 71000 52494
rect 70802 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70802 52332 71000 52390
rect 70802 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70802 52228 71000 52286
rect 70802 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70802 52124 71000 52182
rect 70802 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70802 52020 71000 52078
rect 70802 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70802 51916 71000 51974
rect 70802 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70802 51812 71000 51870
rect 70802 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70802 51708 71000 51766
rect 70802 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70802 51604 71000 51662
rect 70802 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70802 51500 71000 51558
rect 70802 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70802 51396 71000 51454
rect 70802 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70802 51292 71000 51350
rect 70802 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70802 51188 71000 51246
rect 70802 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70802 51084 71000 51142
rect 70802 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70802 50980 71000 51038
rect 70802 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70802 50876 71000 50934
rect 70802 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70802 50772 71000 50830
rect 70802 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70802 50668 71000 50726
rect 70802 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70802 50564 71000 50622
rect 70802 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70802 50460 71000 50518
rect 70802 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70802 50356 71000 50414
rect 70802 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70802 50252 71000 50310
rect 70802 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70802 50148 71000 50206
rect 70802 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70802 50044 71000 50102
rect 70802 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70802 49940 71000 49998
rect 70802 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70802 49836 71000 49894
rect 70802 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70802 49732 71000 49790
rect 70802 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70802 49628 71000 49686
rect 70802 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70802 49524 71000 49582
rect 70802 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70802 49420 71000 49478
rect 70802 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70802 49316 71000 49374
rect 70802 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70802 49212 71000 49270
rect 70802 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70802 49108 71000 49166
rect 70802 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70802 49004 71000 49062
rect 70802 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70802 48900 71000 48958
rect 70802 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70802 48796 71000 48854
rect 70802 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70802 48692 71000 48750
rect 70802 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70802 48588 71000 48646
rect 70802 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70802 48484 71000 48542
rect 70802 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70802 48380 71000 48438
rect 70802 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70802 48276 71000 48334
rect 70802 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70802 48172 71000 48230
rect 70802 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70802 48068 71000 48126
rect 70802 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70802 47964 71000 48022
rect 70802 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70802 47860 71000 47918
rect 70802 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70802 47756 71000 47814
rect 70802 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70802 47652 71000 47710
rect 70802 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70802 47548 71000 47606
rect 70802 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70802 47444 71000 47502
rect 70802 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70802 47340 71000 47398
rect 70802 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70802 47236 71000 47294
rect 70802 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70802 47132 71000 47190
rect 70802 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70802 47028 71000 47086
rect 70802 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70802 46924 71000 46982
rect 70802 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70802 46820 71000 46878
rect 70802 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70802 46716 71000 46774
rect 70802 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70802 46612 71000 46670
rect 70802 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70802 46508 71000 46566
rect 70802 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70802 46404 71000 46462
rect 70802 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70802 46300 71000 46358
rect 70802 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70802 46196 71000 46254
rect 70802 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70802 46092 71000 46150
rect 70802 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70802 45988 71000 46046
rect 70802 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70802 45884 71000 45942
rect 70802 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70802 45780 71000 45838
rect 70802 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70802 45676 71000 45734
rect 70802 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70802 45572 71000 45630
rect 70802 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70802 45468 71000 45526
rect 70802 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70802 45364 71000 45422
rect 70802 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70802 45260 71000 45318
rect 70802 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70802 45156 71000 45214
rect 70802 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70802 45052 71000 45110
rect 70802 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70802 44948 71000 45006
tri 13291 44893 13323 44925 sw
rect 70802 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13097 44892 13323 44893
tri 13323 44892 13324 44893 sw
rect 13097 44847 13324 44892
tri 13324 44847 13369 44892 sw
rect 13097 44843 13369 44847
tri 13097 44842 13098 44843 ne
rect 13098 44842 13369 44843
tri 13098 44841 13099 44842 ne
rect 13099 44841 13369 44842
tri 13099 44840 13100 44841 ne
rect 13100 44840 13369 44841
tri 13100 44839 13101 44840 ne
rect 13101 44839 13369 44840
tri 13101 44838 13102 44839 ne
rect 13102 44838 13369 44839
tri 13102 44837 13103 44838 ne
rect 13103 44837 13369 44838
tri 13369 44837 13379 44847 sw
rect 70802 44844 71000 44902
tri 13103 44830 13110 44837 ne
rect 13110 44830 13379 44837
tri 13110 44785 13155 44830 ne
rect 13155 44824 13379 44830
rect 13155 44785 13254 44824
tri 13155 44740 13200 44785 ne
rect 13200 44778 13254 44785
rect 13300 44792 13379 44824
tri 13379 44792 13424 44837 sw
rect 70802 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 13300 44786 13424 44792
tri 13424 44786 13430 44792 sw
rect 13300 44778 13430 44786
rect 13200 44741 13430 44778
tri 13430 44741 13475 44786 sw
rect 13200 44740 13475 44741
tri 13200 44708 13232 44740 ne
rect 13232 44708 13475 44740
tri 13232 44663 13277 44708 ne
rect 13277 44696 13475 44708
tri 13475 44696 13520 44741 sw
rect 70802 44740 71000 44798
rect 13277 44692 13520 44696
rect 13277 44663 13386 44692
tri 13277 44618 13322 44663 ne
rect 13322 44646 13386 44663
rect 13432 44651 13520 44692
tri 13520 44651 13565 44696 sw
rect 70802 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 13432 44646 13565 44651
rect 13322 44618 13565 44646
tri 13565 44618 13598 44651 sw
rect 70802 44636 71000 44694
tri 13322 44573 13367 44618 ne
rect 13367 44573 13598 44618
tri 13598 44573 13643 44618 sw
rect 70802 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13367 44572 13368 44573 ne
rect 13368 44572 13643 44573
tri 13368 44571 13369 44572 ne
rect 13369 44571 13643 44572
tri 13369 44570 13370 44571 ne
rect 13370 44570 13643 44571
tri 13370 44569 13371 44570 ne
rect 13371 44569 13643 44570
tri 13371 44568 13372 44569 ne
rect 13372 44568 13643 44569
tri 13372 44567 13373 44568 ne
rect 13373 44567 13643 44568
tri 13373 44566 13374 44567 ne
rect 13374 44566 13643 44567
tri 13374 44565 13375 44566 ne
rect 13375 44565 13643 44566
tri 13375 44564 13376 44565 ne
rect 13376 44564 13643 44565
tri 13376 44563 13377 44564 ne
rect 13377 44563 13643 44564
tri 13377 44562 13378 44563 ne
rect 13378 44562 13643 44563
tri 13378 44561 13379 44562 ne
rect 13379 44561 13643 44562
tri 13643 44561 13655 44573 sw
tri 13379 44516 13424 44561 ne
rect 13424 44560 13655 44561
rect 13424 44516 13518 44560
tri 13424 44471 13469 44516 ne
rect 13469 44514 13518 44516
rect 13564 44541 13655 44560
tri 13655 44541 13675 44561 sw
rect 13564 44514 13675 44541
rect 13469 44496 13675 44514
tri 13675 44496 13720 44541 sw
rect 70802 44532 71000 44590
rect 13469 44471 13720 44496
tri 13469 44466 13474 44471 ne
rect 13474 44466 13720 44471
tri 13474 44421 13519 44466 ne
rect 13519 44451 13720 44466
tri 13720 44451 13765 44496 sw
rect 70802 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
rect 13519 44428 13765 44451
rect 13519 44421 13650 44428
tri 13519 44376 13564 44421 ne
rect 13564 44382 13650 44421
rect 13696 44406 13765 44428
tri 13765 44406 13810 44451 sw
rect 70802 44428 71000 44486
rect 13696 44382 13810 44406
rect 13564 44376 13810 44382
tri 13564 44331 13609 44376 ne
rect 13609 44375 13810 44376
tri 13810 44375 13841 44406 sw
rect 70802 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
rect 13609 44331 13841 44375
tri 13609 44298 13642 44331 ne
rect 13642 44330 13841 44331
tri 13841 44330 13886 44375 sw
rect 13642 44298 13886 44330
tri 13642 44297 13643 44298 ne
rect 13643 44297 13886 44298
tri 13643 44296 13644 44297 ne
rect 13644 44296 13886 44297
tri 13644 44295 13645 44296 ne
rect 13645 44295 13782 44296
tri 13645 44294 13646 44295 ne
rect 13646 44294 13782 44295
tri 13646 44293 13647 44294 ne
rect 13647 44293 13782 44294
tri 13647 44292 13648 44293 ne
rect 13648 44292 13782 44293
tri 13648 44291 13649 44292 ne
rect 13649 44291 13782 44292
tri 13649 44290 13650 44291 ne
rect 13650 44290 13782 44291
tri 13650 44289 13651 44290 ne
rect 13651 44289 13782 44290
tri 13651 44288 13652 44289 ne
rect 13652 44288 13782 44289
tri 13652 44287 13653 44288 ne
rect 13653 44287 13782 44288
tri 13653 44286 13654 44287 ne
rect 13654 44286 13782 44287
tri 13654 44285 13655 44286 ne
rect 13655 44285 13782 44286
tri 13655 44240 13700 44285 ne
rect 13700 44250 13782 44285
rect 13828 44285 13886 44296
tri 13886 44285 13931 44330 sw
rect 70802 44324 71000 44382
rect 13828 44250 13931 44285
rect 13700 44240 13931 44250
tri 13931 44240 13976 44285 sw
rect 70802 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
tri 13700 44220 13720 44240 ne
rect 13720 44220 13976 44240
tri 13976 44220 13996 44240 sw
rect 70802 44220 71000 44278
tri 13720 44195 13745 44220 ne
rect 13745 44195 13996 44220
tri 13745 44175 13765 44195 ne
rect 13765 44175 13996 44195
tri 13996 44175 14041 44220 sw
tri 13765 44130 13810 44175 ne
rect 13810 44164 14041 44175
rect 13810 44130 13914 44164
tri 13810 44085 13855 44130 ne
rect 13855 44118 13914 44130
rect 13960 44130 14041 44164
tri 14041 44130 14086 44175 sw
rect 70802 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 13960 44118 14086 44130
rect 13855 44085 14086 44118
tri 14086 44085 14131 44130 sw
rect 70802 44116 71000 44174
tri 13855 44069 13871 44085 ne
rect 13871 44069 14131 44085
tri 13871 44024 13916 44069 ne
rect 13916 44054 14131 44069
tri 14131 44054 14162 44085 sw
rect 70802 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 13916 44032 14162 44054
rect 13916 44024 14046 44032
tri 13916 44023 13917 44024 ne
rect 13917 44023 14046 44024
tri 13917 44022 13918 44023 ne
rect 13918 44022 14046 44023
tri 13918 44021 13919 44022 ne
rect 13919 44021 14046 44022
tri 13919 44020 13920 44021 ne
rect 13920 44020 14046 44021
tri 13920 44019 13921 44020 ne
rect 13921 44019 14046 44020
tri 13921 44018 13922 44019 ne
rect 13922 44018 14046 44019
tri 13922 44017 13923 44018 ne
rect 13923 44017 14046 44018
tri 13923 44016 13924 44017 ne
rect 13924 44016 14046 44017
tri 13924 44015 13925 44016 ne
rect 13925 44015 14046 44016
tri 13925 44014 13926 44015 ne
rect 13926 44014 14046 44015
tri 13926 44013 13927 44014 ne
rect 13927 44013 14046 44014
tri 13927 44012 13928 44013 ne
rect 13928 44012 14046 44013
tri 13928 44011 13929 44012 ne
rect 13929 44011 14046 44012
tri 13929 44010 13930 44011 ne
rect 13930 44010 14046 44011
tri 13930 44009 13931 44010 ne
rect 13931 44009 14046 44010
tri 13931 43964 13976 44009 ne
rect 13976 43986 14046 44009
rect 14092 44009 14162 44032
tri 14162 44009 14207 44054 sw
rect 70802 44012 71000 44070
rect 14092 43986 14207 44009
rect 13976 43964 14207 43986
tri 14207 43964 14252 44009 sw
rect 70802 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13976 43919 14021 43964 ne
rect 14021 43919 14252 43964
tri 14252 43919 14297 43964 sw
tri 14021 43874 14066 43919 ne
rect 14066 43900 14297 43919
rect 14066 43874 14178 43900
tri 14066 43854 14086 43874 ne
rect 14086 43854 14178 43874
rect 14224 43899 14297 43900
tri 14297 43899 14317 43919 sw
rect 70802 43908 71000 43966
rect 14224 43854 14317 43899
tri 14317 43854 14362 43899 sw
rect 70802 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
tri 14086 43829 14111 43854 ne
rect 14111 43829 14362 43854
tri 14111 43809 14131 43829 ne
rect 14131 43809 14362 43829
tri 14362 43809 14407 43854 sw
tri 14131 43764 14176 43809 ne
rect 14176 43768 14407 43809
rect 14176 43764 14310 43768
tri 14176 43749 14191 43764 ne
rect 14191 43749 14310 43764
tri 14191 43748 14192 43749 ne
rect 14192 43748 14310 43749
tri 14192 43747 14193 43748 ne
rect 14193 43747 14310 43748
tri 14193 43746 14194 43747 ne
rect 14194 43746 14310 43747
tri 14194 43745 14195 43746 ne
rect 14195 43745 14310 43746
tri 14195 43744 14196 43745 ne
rect 14196 43744 14310 43745
tri 14196 43743 14197 43744 ne
rect 14197 43743 14310 43744
tri 14197 43742 14198 43743 ne
rect 14198 43742 14310 43743
tri 14198 43741 14199 43742 ne
rect 14199 43741 14310 43742
tri 14199 43740 14200 43741 ne
rect 14200 43740 14310 43741
tri 14200 43739 14201 43740 ne
rect 14201 43739 14310 43740
tri 14201 43738 14202 43739 ne
rect 14202 43738 14310 43739
tri 14202 43737 14203 43738 ne
rect 14203 43737 14310 43738
tri 14203 43736 14204 43737 ne
rect 14204 43736 14310 43737
tri 14204 43735 14205 43736 ne
rect 14205 43735 14310 43736
tri 14205 43734 14206 43735 ne
rect 14206 43734 14310 43735
tri 14206 43733 14207 43734 ne
rect 14207 43733 14310 43734
tri 14207 43688 14252 43733 ne
rect 14252 43722 14310 43733
rect 14356 43764 14407 43768
tri 14407 43764 14452 43809 sw
rect 70802 43804 71000 43862
rect 14356 43733 14452 43764
tri 14452 43733 14483 43764 sw
rect 70802 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43722 14483 43733
rect 14252 43688 14483 43722
tri 14483 43688 14528 43733 sw
rect 70802 43700 71000 43758
tri 14252 43646 14294 43688 ne
rect 14294 43646 14528 43688
tri 14294 43601 14339 43646 ne
rect 14339 43643 14528 43646
tri 14528 43643 14573 43688 sw
rect 70802 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14339 43636 14573 43643
rect 14339 43601 14442 43636
tri 14339 43556 14384 43601 ne
rect 14384 43590 14442 43601
rect 14488 43598 14573 43636
tri 14573 43598 14618 43643 sw
rect 14488 43592 14618 43598
tri 14618 43592 14624 43598 sw
rect 70802 43596 71000 43654
rect 14488 43590 14624 43592
rect 14384 43556 14624 43590
tri 14384 43511 14429 43556 ne
rect 14429 43547 14624 43556
tri 14624 43547 14669 43592 sw
rect 70802 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
rect 14429 43511 14669 43547
tri 14429 43488 14452 43511 ne
rect 14452 43504 14669 43511
rect 14452 43488 14574 43504
tri 14452 43475 14465 43488 ne
rect 14465 43475 14574 43488
tri 14465 43474 14466 43475 ne
rect 14466 43474 14574 43475
tri 14466 43473 14467 43474 ne
rect 14467 43473 14574 43474
tri 14467 43472 14468 43473 ne
rect 14468 43472 14574 43473
tri 14468 43471 14469 43472 ne
rect 14469 43471 14574 43472
tri 14469 43470 14470 43471 ne
rect 14470 43470 14574 43471
tri 14470 43469 14471 43470 ne
rect 14471 43469 14574 43470
tri 14471 43468 14472 43469 ne
rect 14472 43468 14574 43469
tri 14472 43467 14473 43468 ne
rect 14473 43467 14574 43468
tri 14473 43466 14474 43467 ne
rect 14474 43466 14574 43467
tri 14474 43465 14475 43466 ne
rect 14475 43465 14574 43466
tri 14475 43464 14476 43465 ne
rect 14476 43464 14574 43465
tri 14476 43463 14477 43464 ne
rect 14477 43463 14574 43464
tri 14477 43462 14478 43463 ne
rect 14478 43462 14574 43463
tri 14478 43461 14479 43462 ne
rect 14479 43461 14574 43462
tri 14479 43460 14480 43461 ne
rect 14480 43460 14574 43461
tri 14480 43459 14481 43460 ne
rect 14481 43459 14574 43460
tri 14481 43458 14482 43459 ne
rect 14482 43458 14574 43459
rect 14620 43502 14669 43504
tri 14669 43502 14714 43547 sw
rect 14620 43458 14714 43502
tri 14482 43457 14483 43458 ne
rect 14483 43457 14714 43458
tri 14714 43457 14759 43502 sw
rect 70802 43492 71000 43550
tri 14483 43443 14497 43457 ne
rect 14497 43443 14759 43457
tri 14759 43443 14773 43457 sw
rect 70802 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14497 43398 14542 43443 ne
rect 14542 43398 14773 43443
tri 14773 43398 14818 43443 sw
tri 14542 43353 14587 43398 ne
rect 14587 43372 14818 43398
rect 14587 43353 14706 43372
tri 14587 43327 14613 43353 ne
rect 14613 43327 14706 43353
tri 14613 43282 14658 43327 ne
rect 14658 43326 14706 43327
rect 14752 43353 14818 43372
tri 14818 43353 14863 43398 sw
rect 70802 43388 71000 43446
rect 14752 43326 14863 43353
rect 14658 43308 14863 43326
tri 14863 43308 14908 43353 sw
rect 70802 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 14658 43282 14908 43308
tri 14658 43237 14703 43282 ne
rect 14703 43271 14908 43282
tri 14908 43271 14945 43308 sw
rect 70802 43284 71000 43342
rect 14703 43240 14945 43271
rect 14703 43237 14838 43240
tri 14703 43201 14739 43237 ne
rect 14739 43201 14838 43237
tri 14739 43200 14740 43201 ne
rect 14740 43200 14838 43201
tri 14740 43199 14741 43200 ne
rect 14741 43199 14838 43200
tri 14741 43198 14742 43199 ne
rect 14742 43198 14838 43199
tri 14742 43197 14743 43198 ne
rect 14743 43197 14838 43198
tri 14743 43196 14744 43197 ne
rect 14744 43196 14838 43197
tri 14744 43195 14745 43196 ne
rect 14745 43195 14838 43196
tri 14745 43194 14746 43195 ne
rect 14746 43194 14838 43195
rect 14884 43226 14945 43240
tri 14945 43226 14990 43271 sw
rect 70802 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43194 14990 43226
tri 14746 43193 14747 43194 ne
rect 14747 43193 14990 43194
tri 14747 43192 14748 43193 ne
rect 14748 43192 14990 43193
tri 14748 43191 14749 43192 ne
rect 14749 43191 14990 43192
tri 14749 43190 14750 43191 ne
rect 14750 43190 14990 43191
tri 14750 43189 14751 43190 ne
rect 14751 43189 14990 43190
tri 14751 43188 14752 43189 ne
rect 14752 43188 14990 43189
tri 14752 43187 14753 43188 ne
rect 14753 43187 14990 43188
tri 14753 43186 14754 43187 ne
rect 14754 43186 14990 43187
tri 14754 43185 14755 43186 ne
rect 14755 43185 14990 43186
tri 14755 43184 14756 43185 ne
rect 14756 43184 14990 43185
tri 14756 43183 14757 43184 ne
rect 14757 43183 14990 43184
tri 14757 43182 14758 43183 ne
rect 14758 43182 14990 43183
tri 14758 43181 14759 43182 ne
rect 14759 43181 14990 43182
tri 14990 43181 15035 43226 sw
tri 14759 43136 14804 43181 ne
rect 14804 43136 15035 43181
tri 15035 43136 15080 43181 sw
rect 70802 43180 71000 43238
tri 14804 43122 14818 43136 ne
rect 14818 43122 15080 43136
tri 15080 43122 15094 43136 sw
rect 70802 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14818 43091 14849 43122 ne
rect 14849 43108 15094 43122
rect 14849 43091 14970 43108
tri 14849 43077 14863 43091 ne
rect 14863 43077 14970 43091
tri 14863 43032 14908 43077 ne
rect 14908 43062 14970 43077
rect 15016 43077 15094 43108
tri 15094 43077 15139 43122 sw
rect 15016 43062 15139 43077
rect 14908 43032 15139 43062
tri 15139 43032 15184 43077 sw
rect 70802 43076 71000 43134
tri 14908 42987 14953 43032 ne
rect 14953 42987 15184 43032
tri 15184 42987 15229 43032 sw
rect 70802 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14953 42971 14969 42987 ne
rect 14969 42976 15229 42987
rect 14969 42971 15102 42976
tri 14969 42926 15014 42971 ne
rect 15014 42930 15102 42971
rect 15148 42950 15229 42976
tri 15229 42950 15266 42987 sw
rect 70802 42972 71000 43030
rect 15148 42930 15266 42950
rect 15014 42926 15266 42930
tri 15014 42925 15015 42926 ne
rect 15015 42925 15266 42926
tri 15015 42924 15016 42925 ne
rect 15016 42924 15266 42925
tri 15016 42923 15017 42924 ne
rect 15017 42923 15266 42924
tri 15017 42922 15018 42923 ne
rect 15018 42922 15266 42923
tri 15018 42921 15019 42922 ne
rect 15019 42921 15266 42922
tri 15019 42920 15020 42921 ne
rect 15020 42920 15266 42921
tri 15020 42919 15021 42920 ne
rect 15021 42919 15266 42920
tri 15021 42918 15022 42919 ne
rect 15022 42918 15266 42919
tri 15022 42917 15023 42918 ne
rect 15023 42917 15266 42918
tri 15023 42916 15024 42917 ne
rect 15024 42916 15266 42917
tri 15024 42915 15025 42916 ne
rect 15025 42915 15266 42916
tri 15025 42914 15026 42915 ne
rect 15026 42914 15266 42915
tri 15026 42913 15027 42914 ne
rect 15027 42913 15266 42914
tri 15027 42912 15028 42913 ne
rect 15028 42912 15266 42913
tri 15028 42911 15029 42912 ne
rect 15029 42911 15266 42912
tri 15029 42910 15030 42911 ne
rect 15030 42910 15266 42911
tri 15030 42909 15031 42910 ne
rect 15031 42909 15266 42910
tri 15031 42908 15032 42909 ne
rect 15032 42908 15266 42909
tri 15032 42907 15033 42908 ne
rect 15033 42907 15266 42908
tri 15033 42906 15034 42907 ne
rect 15034 42906 15266 42907
tri 15034 42905 15035 42906 ne
rect 15035 42905 15266 42906
tri 15266 42905 15311 42950 sw
rect 70802 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15035 42860 15080 42905 ne
rect 15080 42860 15311 42905
tri 15311 42860 15356 42905 sw
rect 70802 42868 71000 42926
tri 15080 42815 15125 42860 ne
rect 15125 42844 15356 42860
rect 15125 42815 15234 42844
tri 15125 42770 15170 42815 ne
rect 15170 42798 15234 42815
rect 15280 42815 15356 42844
tri 15356 42815 15401 42860 sw
rect 70802 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 15280 42801 15401 42815
tri 15401 42801 15415 42815 sw
rect 15280 42798 15415 42801
rect 15170 42770 15415 42798
tri 15170 42756 15184 42770 ne
rect 15184 42756 15415 42770
tri 15415 42756 15460 42801 sw
rect 70802 42764 71000 42822
tri 15184 42725 15215 42756 ne
rect 15215 42725 15460 42756
tri 15215 42711 15229 42725 ne
rect 15229 42712 15460 42725
rect 15229 42711 15366 42712
tri 15229 42666 15274 42711 ne
rect 15274 42666 15366 42711
rect 15412 42711 15460 42712
tri 15460 42711 15505 42756 sw
rect 70802 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 15412 42666 15505 42711
tri 15505 42666 15550 42711 sw
tri 15274 42652 15288 42666 ne
rect 15288 42652 15550 42666
tri 15288 42651 15289 42652 ne
rect 15289 42651 15550 42652
tri 15289 42650 15290 42651 ne
rect 15290 42650 15550 42651
tri 15290 42649 15291 42650 ne
rect 15291 42649 15550 42650
tri 15291 42648 15292 42649 ne
rect 15292 42648 15550 42649
tri 15292 42647 15293 42648 ne
rect 15293 42647 15550 42648
tri 15293 42646 15294 42647 ne
rect 15294 42646 15550 42647
tri 15294 42645 15295 42646 ne
rect 15295 42645 15550 42646
tri 15295 42644 15296 42645 ne
rect 15296 42644 15550 42645
tri 15296 42643 15297 42644 ne
rect 15297 42643 15550 42644
tri 15297 42642 15298 42643 ne
rect 15298 42642 15550 42643
tri 15298 42641 15299 42642 ne
rect 15299 42641 15550 42642
tri 15299 42640 15300 42641 ne
rect 15300 42640 15550 42641
tri 15300 42639 15301 42640 ne
rect 15301 42639 15550 42640
tri 15301 42638 15302 42639 ne
rect 15302 42638 15550 42639
tri 15302 42637 15303 42638 ne
rect 15303 42637 15550 42638
tri 15303 42636 15304 42637 ne
rect 15304 42636 15550 42637
tri 15304 42635 15305 42636 ne
rect 15305 42635 15550 42636
tri 15305 42634 15306 42635 ne
rect 15306 42634 15550 42635
tri 15306 42633 15307 42634 ne
rect 15307 42633 15550 42634
tri 15307 42632 15308 42633 ne
rect 15308 42632 15550 42633
tri 15308 42631 15309 42632 ne
rect 15309 42631 15550 42632
tri 15309 42630 15310 42631 ne
rect 15310 42630 15550 42631
tri 15310 42629 15311 42630 ne
rect 15311 42629 15550 42630
tri 15550 42629 15587 42666 sw
rect 70802 42660 71000 42718
tri 15311 42584 15356 42629 ne
rect 15356 42584 15587 42629
tri 15587 42584 15632 42629 sw
rect 70802 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15356 42552 15388 42584 ne
rect 15388 42580 15632 42584
rect 15388 42552 15498 42580
tri 15388 42507 15433 42552 ne
rect 15433 42534 15498 42552
rect 15544 42539 15632 42580
tri 15632 42539 15677 42584 sw
rect 70802 42556 71000 42614
rect 15544 42534 15677 42539
rect 15433 42507 15677 42534
tri 15433 42462 15478 42507 ne
rect 15478 42494 15677 42507
tri 15677 42494 15722 42539 sw
rect 70802 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 15478 42488 15722 42494
tri 15722 42488 15728 42494 sw
rect 15478 42462 15728 42488
tri 15478 42417 15523 42462 ne
rect 15523 42448 15728 42462
rect 15523 42417 15630 42448
tri 15523 42390 15550 42417 ne
rect 15550 42402 15630 42417
rect 15676 42443 15728 42448
tri 15728 42443 15773 42488 sw
rect 70802 42452 71000 42510
rect 15676 42402 15773 42443
rect 15550 42398 15773 42402
tri 15773 42398 15818 42443 sw
rect 70802 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 15550 42390 15818 42398
tri 15550 42377 15563 42390 ne
rect 15563 42377 15818 42390
tri 15563 42376 15564 42377 ne
rect 15564 42376 15818 42377
tri 15564 42375 15565 42376 ne
rect 15565 42375 15818 42376
tri 15565 42374 15566 42375 ne
rect 15566 42374 15818 42375
tri 15566 42373 15567 42374 ne
rect 15567 42373 15818 42374
tri 15567 42372 15568 42373 ne
rect 15568 42372 15818 42373
tri 15568 42371 15569 42372 ne
rect 15569 42371 15818 42372
tri 15569 42370 15570 42371 ne
rect 15570 42370 15818 42371
tri 15570 42369 15571 42370 ne
rect 15571 42369 15818 42370
tri 15571 42368 15572 42369 ne
rect 15572 42368 15818 42369
tri 15572 42367 15573 42368 ne
rect 15573 42367 15818 42368
tri 15573 42366 15574 42367 ne
rect 15574 42366 15818 42367
tri 15574 42365 15575 42366 ne
rect 15575 42365 15818 42366
tri 15575 42364 15576 42365 ne
rect 15576 42364 15818 42365
tri 15576 42363 15577 42364 ne
rect 15577 42363 15818 42364
tri 15577 42362 15578 42363 ne
rect 15578 42362 15818 42363
tri 15578 42361 15579 42362 ne
rect 15579 42361 15818 42362
tri 15579 42360 15580 42361 ne
rect 15580 42360 15818 42361
tri 15580 42359 15581 42360 ne
rect 15581 42359 15818 42360
tri 15581 42358 15582 42359 ne
rect 15582 42358 15818 42359
tri 15582 42357 15583 42358 ne
rect 15583 42357 15818 42358
tri 15583 42356 15584 42357 ne
rect 15584 42356 15818 42357
tri 15584 42355 15585 42356 ne
rect 15585 42355 15818 42356
tri 15585 42354 15586 42355 ne
rect 15586 42354 15818 42355
tri 15586 42353 15587 42354 ne
rect 15587 42353 15818 42354
tri 15818 42353 15863 42398 sw
tri 15587 42345 15595 42353 ne
rect 15595 42345 15863 42353
tri 15863 42345 15871 42353 sw
rect 70802 42348 71000 42406
tri 15595 42300 15640 42345 ne
rect 15640 42316 15871 42345
rect 15640 42300 15762 42316
tri 15640 42255 15685 42300 ne
rect 15685 42270 15762 42300
rect 15808 42300 15871 42316
tri 15871 42300 15916 42345 sw
rect 70802 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42270 15916 42300
rect 15685 42255 15916 42270
tri 15916 42255 15961 42300 sw
tri 15685 42232 15708 42255 ne
rect 15708 42232 15961 42255
tri 15708 42187 15753 42232 ne
rect 15753 42210 15961 42232
tri 15961 42210 16006 42255 sw
rect 70802 42244 71000 42302
rect 15753 42187 16006 42210
tri 15753 42142 15798 42187 ne
rect 15798 42184 16006 42187
rect 15798 42142 15894 42184
tri 15798 42103 15837 42142 ne
rect 15837 42138 15894 42142
rect 15940 42167 16006 42184
tri 16006 42167 16049 42210 sw
rect 70802 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
rect 15940 42138 16049 42167
rect 15837 42122 16049 42138
tri 16049 42122 16094 42167 sw
rect 70802 42140 71000 42198
rect 15837 42103 16094 42122
tri 15837 42102 15838 42103 ne
rect 15838 42102 16094 42103
tri 15838 42101 15839 42102 ne
rect 15839 42101 16094 42102
tri 15839 42100 15840 42101 ne
rect 15840 42100 16094 42101
tri 15840 42099 15841 42100 ne
rect 15841 42099 16094 42100
tri 15841 42098 15842 42099 ne
rect 15842 42098 16094 42099
tri 15842 42097 15843 42098 ne
rect 15843 42097 16094 42098
tri 15843 42096 15844 42097 ne
rect 15844 42096 16094 42097
tri 15844 42095 15845 42096 ne
rect 15845 42095 16094 42096
tri 15845 42094 15846 42095 ne
rect 15846 42094 16094 42095
tri 15846 42093 15847 42094 ne
rect 15847 42093 16094 42094
tri 15847 42092 15848 42093 ne
rect 15848 42092 16094 42093
tri 15848 42091 15849 42092 ne
rect 15849 42091 16094 42092
tri 15849 42090 15850 42091 ne
rect 15850 42090 16094 42091
tri 15850 42089 15851 42090 ne
rect 15851 42089 16094 42090
tri 15851 42088 15852 42089 ne
rect 15852 42088 16094 42089
tri 15852 42087 15853 42088 ne
rect 15853 42087 16094 42088
tri 15853 42086 15854 42087 ne
rect 15854 42086 16094 42087
tri 15854 42085 15855 42086 ne
rect 15855 42085 16094 42086
tri 15855 42084 15856 42085 ne
rect 15856 42084 16094 42085
tri 15856 42083 15857 42084 ne
rect 15857 42083 16094 42084
tri 15857 42082 15858 42083 ne
rect 15858 42082 16094 42083
tri 15858 42081 15859 42082 ne
rect 15859 42081 16094 42082
tri 15859 42080 15860 42081 ne
rect 15860 42080 16094 42081
tri 15860 42079 15861 42080 ne
rect 15861 42079 16094 42080
tri 15861 42078 15862 42079 ne
rect 15862 42078 16094 42079
tri 15862 42077 15863 42078 ne
rect 15863 42077 16094 42078
tri 16094 42077 16139 42122 sw
rect 70802 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15863 42032 15908 42077 ne
rect 15908 42052 16139 42077
rect 15908 42032 16026 42052
tri 15908 42024 15916 42032 ne
rect 15916 42024 16026 42032
tri 15916 41987 15953 42024 ne
rect 15953 42006 16026 42024
rect 16072 42032 16139 42052
tri 16139 42032 16184 42077 sw
rect 70802 42036 71000 42094
rect 16072 42024 16184 42032
tri 16184 42024 16192 42032 sw
rect 16072 42006 16192 42024
rect 15953 41987 16192 42006
tri 15953 41979 15961 41987 ne
rect 15961 41979 16192 41987
tri 16192 41979 16237 42024 sw
rect 70802 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15961 41934 16006 41979 ne
rect 16006 41934 16237 41979
tri 16237 41934 16282 41979 sw
tri 16006 41889 16051 41934 ne
rect 16051 41920 16282 41934
rect 16051 41889 16158 41920
tri 16051 41874 16066 41889 ne
rect 16066 41874 16158 41889
rect 16204 41889 16282 41920
tri 16282 41889 16327 41934 sw
rect 70802 41932 71000 41990
rect 16204 41874 16327 41889
tri 16066 41829 16111 41874 ne
rect 16111 41846 16327 41874
tri 16327 41846 16370 41889 sw
rect 70802 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 16111 41829 16370 41846
tri 16111 41828 16112 41829 ne
rect 16112 41828 16370 41829
tri 16112 41827 16113 41828 ne
rect 16113 41827 16370 41828
tri 16113 41826 16114 41827 ne
rect 16114 41826 16370 41827
tri 16114 41825 16115 41826 ne
rect 16115 41825 16370 41826
tri 16115 41824 16116 41825 ne
rect 16116 41824 16370 41825
tri 16116 41823 16117 41824 ne
rect 16117 41823 16370 41824
tri 16117 41822 16118 41823 ne
rect 16118 41822 16370 41823
tri 16118 41821 16119 41822 ne
rect 16119 41821 16370 41822
tri 16119 41820 16120 41821 ne
rect 16120 41820 16370 41821
tri 16120 41819 16121 41820 ne
rect 16121 41819 16370 41820
tri 16121 41818 16122 41819 ne
rect 16122 41818 16370 41819
tri 16122 41817 16123 41818 ne
rect 16123 41817 16370 41818
tri 16123 41816 16124 41817 ne
rect 16124 41816 16370 41817
tri 16124 41815 16125 41816 ne
rect 16125 41815 16370 41816
tri 16125 41814 16126 41815 ne
rect 16126 41814 16370 41815
tri 16126 41813 16127 41814 ne
rect 16127 41813 16370 41814
tri 16127 41812 16128 41813 ne
rect 16128 41812 16370 41813
tri 16128 41811 16129 41812 ne
rect 16129 41811 16370 41812
tri 16129 41810 16130 41811 ne
rect 16130 41810 16370 41811
tri 16130 41809 16131 41810 ne
rect 16131 41809 16370 41810
tri 16131 41808 16132 41809 ne
rect 16132 41808 16370 41809
tri 16132 41807 16133 41808 ne
rect 16133 41807 16370 41808
tri 16133 41806 16134 41807 ne
rect 16134 41806 16370 41807
tri 16134 41805 16135 41806 ne
rect 16135 41805 16370 41806
tri 16135 41804 16136 41805 ne
rect 16136 41804 16370 41805
tri 16136 41803 16137 41804 ne
rect 16137 41803 16370 41804
tri 16137 41802 16138 41803 ne
rect 16138 41802 16370 41803
tri 16138 41801 16139 41802 ne
rect 16139 41801 16370 41802
tri 16370 41801 16415 41846 sw
rect 70802 41828 71000 41886
tri 16139 41756 16184 41801 ne
rect 16184 41788 16415 41801
rect 16184 41756 16290 41788
tri 16184 41711 16229 41756 ne
rect 16229 41742 16290 41756
rect 16336 41756 16415 41788
tri 16415 41756 16460 41801 sw
rect 70802 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41742 16460 41756
rect 16229 41711 16460 41742
tri 16460 41711 16505 41756 sw
rect 70802 41724 71000 41782
tri 16229 41666 16274 41711 ne
rect 16274 41703 16505 41711
tri 16505 41703 16513 41711 sw
rect 16274 41666 16513 41703
tri 16274 41658 16282 41666 ne
rect 16282 41658 16513 41666
tri 16513 41658 16558 41703 sw
rect 70802 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
tri 16282 41621 16319 41658 ne
rect 16319 41656 16558 41658
rect 16319 41621 16422 41656
tri 16319 41613 16327 41621 ne
rect 16327 41613 16422 41621
tri 16327 41568 16372 41613 ne
rect 16372 41610 16422 41613
rect 16468 41613 16558 41656
tri 16558 41613 16603 41658 sw
rect 70802 41620 71000 41678
rect 16468 41610 16603 41613
rect 16372 41568 16603 41610
tri 16603 41568 16648 41613 sw
rect 70802 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16372 41554 16386 41568 ne
rect 16386 41554 16648 41568
tri 16386 41553 16387 41554 ne
rect 16387 41553 16648 41554
tri 16387 41552 16388 41553 ne
rect 16388 41552 16648 41553
tri 16388 41551 16389 41552 ne
rect 16389 41551 16648 41552
tri 16389 41550 16390 41551 ne
rect 16390 41550 16648 41551
tri 16390 41549 16391 41550 ne
rect 16391 41549 16648 41550
tri 16391 41548 16392 41549 ne
rect 16392 41548 16648 41549
tri 16392 41547 16393 41548 ne
rect 16393 41547 16648 41548
tri 16393 41546 16394 41547 ne
rect 16394 41546 16648 41547
tri 16394 41545 16395 41546 ne
rect 16395 41545 16648 41546
tri 16395 41544 16396 41545 ne
rect 16396 41544 16648 41545
tri 16396 41543 16397 41544 ne
rect 16397 41543 16648 41544
tri 16397 41542 16398 41543 ne
rect 16398 41542 16648 41543
tri 16398 41541 16399 41542 ne
rect 16399 41541 16648 41542
tri 16399 41540 16400 41541 ne
rect 16400 41540 16648 41541
tri 16400 41539 16401 41540 ne
rect 16401 41539 16648 41540
tri 16401 41538 16402 41539 ne
rect 16402 41538 16648 41539
tri 16402 41537 16403 41538 ne
rect 16403 41537 16648 41538
tri 16403 41536 16404 41537 ne
rect 16404 41536 16648 41537
tri 16404 41535 16405 41536 ne
rect 16405 41535 16648 41536
tri 16405 41534 16406 41535 ne
rect 16406 41534 16648 41535
tri 16406 41533 16407 41534 ne
rect 16407 41533 16648 41534
tri 16407 41532 16408 41533 ne
rect 16408 41532 16648 41533
tri 16408 41531 16409 41532 ne
rect 16409 41531 16648 41532
tri 16409 41530 16410 41531 ne
rect 16410 41530 16648 41531
tri 16410 41529 16411 41530 ne
rect 16411 41529 16648 41530
tri 16411 41528 16412 41529 ne
rect 16412 41528 16648 41529
tri 16412 41527 16413 41528 ne
rect 16413 41527 16648 41528
tri 16413 41526 16414 41527 ne
rect 16414 41526 16648 41527
tri 16414 41525 16415 41526 ne
rect 16415 41525 16648 41526
tri 16648 41525 16691 41568 sw
tri 16415 41480 16460 41525 ne
rect 16460 41524 16691 41525
rect 16460 41480 16554 41524
tri 16460 41458 16482 41480 ne
rect 16482 41478 16554 41480
rect 16600 41480 16691 41524
tri 16691 41480 16736 41525 sw
rect 70802 41516 71000 41574
rect 16600 41478 16736 41480
rect 16482 41458 16736 41478
tri 16482 41413 16527 41458 ne
rect 16527 41435 16736 41458
tri 16736 41435 16781 41480 sw
rect 70802 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 16527 41413 16781 41435
tri 16527 41368 16572 41413 ne
rect 16572 41392 16781 41413
rect 16572 41368 16686 41392
tri 16572 41323 16617 41368 ne
rect 16617 41346 16686 41368
rect 16732 41390 16781 41392
tri 16781 41390 16826 41435 sw
rect 70802 41412 71000 41470
rect 16732 41384 16826 41390
tri 16826 41384 16832 41390 sw
rect 16732 41346 16832 41384
rect 16617 41339 16832 41346
tri 16832 41339 16877 41384 sw
rect 70802 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 16617 41323 16877 41339
tri 16617 41292 16648 41323 ne
rect 16648 41294 16877 41323
tri 16877 41294 16922 41339 sw
rect 70802 41308 71000 41366
rect 16648 41292 16922 41294
tri 16648 41280 16660 41292 ne
rect 16660 41280 16922 41292
tri 16660 41279 16661 41280 ne
rect 16661 41279 16922 41280
tri 16661 41278 16662 41279 ne
rect 16662 41278 16922 41279
tri 16662 41277 16663 41278 ne
rect 16663 41277 16922 41278
tri 16663 41276 16664 41277 ne
rect 16664 41276 16922 41277
tri 16664 41275 16665 41276 ne
rect 16665 41275 16922 41276
tri 16665 41274 16666 41275 ne
rect 16666 41274 16922 41275
tri 16666 41273 16667 41274 ne
rect 16667 41273 16922 41274
tri 16667 41272 16668 41273 ne
rect 16668 41272 16922 41273
tri 16668 41271 16669 41272 ne
rect 16669 41271 16922 41272
tri 16669 41270 16670 41271 ne
rect 16670 41270 16922 41271
tri 16670 41269 16671 41270 ne
rect 16671 41269 16922 41270
tri 16671 41268 16672 41269 ne
rect 16672 41268 16922 41269
tri 16672 41267 16673 41268 ne
rect 16673 41267 16922 41268
tri 16673 41266 16674 41267 ne
rect 16674 41266 16922 41267
tri 16674 41265 16675 41266 ne
rect 16675 41265 16922 41266
tri 16675 41264 16676 41265 ne
rect 16676 41264 16922 41265
tri 16676 41263 16677 41264 ne
rect 16677 41263 16922 41264
tri 16677 41262 16678 41263 ne
rect 16678 41262 16922 41263
tri 16678 41261 16679 41262 ne
rect 16679 41261 16922 41262
tri 16679 41260 16680 41261 ne
rect 16680 41260 16922 41261
tri 16680 41259 16681 41260 ne
rect 16681 41259 16818 41260
tri 16681 41258 16682 41259 ne
rect 16682 41258 16818 41259
tri 16682 41257 16683 41258 ne
rect 16683 41257 16818 41258
tri 16683 41256 16684 41257 ne
rect 16684 41256 16818 41257
tri 16684 41255 16685 41256 ne
rect 16685 41255 16818 41256
tri 16685 41254 16686 41255 ne
rect 16686 41254 16818 41255
tri 16686 41253 16687 41254 ne
rect 16687 41253 16818 41254
tri 16687 41252 16688 41253 ne
rect 16688 41252 16818 41253
tri 16688 41251 16689 41252 ne
rect 16689 41251 16818 41252
tri 16689 41250 16690 41251 ne
rect 16690 41250 16818 41251
tri 16690 41249 16691 41250 ne
rect 16691 41249 16818 41250
tri 16691 41247 16693 41249 ne
rect 16693 41247 16818 41249
tri 16693 41202 16738 41247 ne
rect 16738 41214 16818 41247
rect 16864 41249 16922 41260
tri 16922 41249 16967 41294 sw
rect 70802 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 16864 41247 16967 41249
tri 16967 41247 16969 41249 sw
rect 16864 41214 16969 41247
rect 16738 41202 16969 41214
tri 16969 41202 17014 41247 sw
rect 70802 41204 71000 41262
tri 16738 41157 16783 41202 ne
rect 16783 41157 17014 41202
tri 17014 41157 17059 41202 sw
rect 70802 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
tri 16783 41138 16802 41157 ne
rect 16802 41138 17059 41157
tri 16802 41093 16847 41138 ne
rect 16847 41128 17059 41138
rect 16847 41093 16950 41128
tri 16847 41048 16892 41093 ne
rect 16892 41082 16950 41093
rect 16996 41112 17059 41128
tri 17059 41112 17104 41157 sw
rect 16996 41108 17104 41112
tri 17104 41108 17108 41112 sw
rect 16996 41082 17108 41108
rect 16892 41063 17108 41082
tri 17108 41063 17153 41108 sw
rect 70802 41100 71000 41158
rect 16892 41048 17153 41063
tri 16892 41005 16935 41048 ne
rect 16935 41018 17153 41048
tri 17153 41018 17198 41063 sw
rect 70802 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 16935 41005 17198 41018
tri 16935 41004 16936 41005 ne
rect 16936 41004 17198 41005
tri 16936 41003 16937 41004 ne
rect 16937 41003 17198 41004
tri 16937 41002 16938 41003 ne
rect 16938 41002 17198 41003
tri 16938 41001 16939 41002 ne
rect 16939 41001 17198 41002
tri 16939 41000 16940 41001 ne
rect 16940 41000 17198 41001
tri 16940 40999 16941 41000 ne
rect 16941 40999 17198 41000
tri 16941 40998 16942 40999 ne
rect 16942 40998 17198 40999
tri 16942 40997 16943 40998 ne
rect 16943 40997 17198 40998
tri 16943 40996 16944 40997 ne
rect 16944 40996 17198 40997
tri 16944 40995 16945 40996 ne
rect 16945 40995 17082 40996
tri 16945 40994 16946 40995 ne
rect 16946 40994 17082 40995
tri 16946 40993 16947 40994 ne
rect 16947 40993 17082 40994
tri 16947 40992 16948 40993 ne
rect 16948 40992 17082 40993
tri 16948 40991 16949 40992 ne
rect 16949 40991 17082 40992
tri 16949 40990 16950 40991 ne
rect 16950 40990 17082 40991
tri 16950 40989 16951 40990 ne
rect 16951 40989 17082 40990
tri 16951 40988 16952 40989 ne
rect 16952 40988 17082 40989
tri 16952 40987 16953 40988 ne
rect 16953 40987 17082 40988
tri 16953 40986 16954 40987 ne
rect 16954 40986 17082 40987
tri 16954 40985 16955 40986 ne
rect 16955 40985 17082 40986
tri 16955 40984 16956 40985 ne
rect 16956 40984 17082 40985
tri 16956 40983 16957 40984 ne
rect 16957 40983 17082 40984
tri 16957 40982 16958 40983 ne
rect 16958 40982 17082 40983
tri 16958 40981 16959 40982 ne
rect 16959 40981 17082 40982
tri 16959 40980 16960 40981 ne
rect 16960 40980 17082 40981
tri 16960 40979 16961 40980 ne
rect 16961 40979 17082 40980
tri 16961 40978 16962 40979 ne
rect 16962 40978 17082 40979
tri 16962 40977 16963 40978 ne
rect 16963 40977 17082 40978
tri 16963 40976 16964 40977 ne
rect 16964 40976 17082 40977
tri 16964 40975 16965 40976 ne
rect 16965 40975 17082 40976
tri 16965 40974 16966 40975 ne
rect 16966 40974 17082 40975
tri 16966 40973 16967 40974 ne
rect 16967 40973 17082 40974
tri 16967 40928 17012 40973 ne
rect 17012 40950 17082 40973
rect 17128 40973 17198 40996
tri 17198 40973 17243 41018 sw
rect 70802 40996 71000 41054
rect 17128 40950 17243 40973
rect 17012 40928 17243 40950
tri 17243 40928 17288 40973 sw
rect 70802 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
tri 17012 40926 17014 40928 ne
rect 17014 40926 17288 40928
tri 17288 40926 17290 40928 sw
tri 17014 40883 17057 40926 ne
rect 17057 40883 17290 40926
tri 17057 40881 17059 40883 ne
rect 17059 40881 17290 40883
tri 17290 40881 17335 40926 sw
rect 70802 40892 71000 40950
tri 17059 40836 17104 40881 ne
rect 17104 40864 17335 40881
rect 17104 40836 17214 40864
tri 17104 40791 17149 40836 ne
rect 17149 40818 17214 40836
rect 17260 40836 17335 40864
tri 17335 40836 17380 40881 sw
rect 70802 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40818 17380 40836
rect 17149 40791 17380 40818
tri 17380 40791 17425 40836 sw
tri 17149 40776 17164 40791 ne
rect 17164 40787 17425 40791
tri 17425 40787 17429 40791 sw
rect 70802 40788 71000 40846
rect 17164 40776 17429 40787
tri 17164 40731 17209 40776 ne
rect 17209 40742 17429 40776
tri 17429 40742 17474 40787 sw
rect 70802 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17209 40732 17474 40742
rect 17209 40731 17346 40732
tri 17209 40730 17210 40731 ne
rect 17210 40730 17346 40731
tri 17210 40729 17211 40730 ne
rect 17211 40729 17346 40730
tri 17211 40728 17212 40729 ne
rect 17212 40728 17346 40729
tri 17212 40727 17213 40728 ne
rect 17213 40727 17346 40728
tri 17213 40726 17214 40727 ne
rect 17214 40726 17346 40727
tri 17214 40725 17215 40726 ne
rect 17215 40725 17346 40726
tri 17215 40724 17216 40725 ne
rect 17216 40724 17346 40725
tri 17216 40723 17217 40724 ne
rect 17217 40723 17346 40724
tri 17217 40722 17218 40723 ne
rect 17218 40722 17346 40723
tri 17218 40721 17219 40722 ne
rect 17219 40721 17346 40722
tri 17219 40720 17220 40721 ne
rect 17220 40720 17346 40721
tri 17220 40719 17221 40720 ne
rect 17221 40719 17346 40720
tri 17221 40718 17222 40719 ne
rect 17222 40718 17346 40719
tri 17222 40717 17223 40718 ne
rect 17223 40717 17346 40718
tri 17223 40716 17224 40717 ne
rect 17224 40716 17346 40717
tri 17224 40715 17225 40716 ne
rect 17225 40715 17346 40716
tri 17225 40714 17226 40715 ne
rect 17226 40714 17346 40715
tri 17226 40713 17227 40714 ne
rect 17227 40713 17346 40714
tri 17227 40712 17228 40713 ne
rect 17228 40712 17346 40713
tri 17228 40711 17229 40712 ne
rect 17229 40711 17346 40712
tri 17229 40710 17230 40711 ne
rect 17230 40710 17346 40711
tri 17230 40709 17231 40710 ne
rect 17231 40709 17346 40710
tri 17231 40708 17232 40709 ne
rect 17232 40708 17346 40709
tri 17232 40707 17233 40708 ne
rect 17233 40707 17346 40708
tri 17233 40706 17234 40707 ne
rect 17234 40706 17346 40707
tri 17234 40705 17235 40706 ne
rect 17235 40705 17346 40706
tri 17235 40704 17236 40705 ne
rect 17236 40704 17346 40705
tri 17236 40703 17237 40704 ne
rect 17237 40703 17346 40704
tri 17237 40702 17238 40703 ne
rect 17238 40702 17346 40703
tri 17238 40701 17239 40702 ne
rect 17239 40701 17346 40702
tri 17239 40700 17240 40701 ne
rect 17240 40700 17346 40701
tri 17240 40699 17241 40700 ne
rect 17241 40699 17346 40700
tri 17241 40698 17242 40699 ne
rect 17242 40698 17346 40699
tri 17242 40697 17243 40698 ne
rect 17243 40697 17346 40698
tri 17243 40652 17288 40697 ne
rect 17288 40686 17346 40697
rect 17392 40697 17474 40732
tri 17474 40697 17519 40742 sw
rect 17392 40686 17519 40697
rect 17288 40652 17519 40686
tri 17519 40652 17564 40697 sw
rect 70802 40684 71000 40742
tri 17288 40607 17333 40652 ne
rect 17333 40607 17564 40652
tri 17564 40607 17609 40652 sw
rect 70802 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17333 40562 17378 40607 ne
rect 17378 40605 17609 40607
tri 17609 40605 17611 40607 sw
rect 17378 40600 17611 40605
rect 17378 40562 17478 40600
tri 17378 40560 17380 40562 ne
rect 17380 40560 17478 40562
tri 17380 40517 17423 40560 ne
rect 17423 40554 17478 40560
rect 17524 40560 17611 40600
tri 17611 40560 17656 40605 sw
rect 70802 40580 71000 40638
rect 17524 40554 17656 40560
rect 17423 40517 17656 40554
tri 17423 40515 17425 40517 ne
rect 17425 40515 17656 40517
tri 17656 40515 17701 40560 sw
rect 70802 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17425 40470 17470 40515 ne
rect 17470 40470 17701 40515
tri 17701 40470 17746 40515 sw
rect 70802 40476 71000 40534
tri 17470 40457 17483 40470 ne
rect 17483 40468 17746 40470
rect 17483 40457 17610 40468
tri 17483 40456 17484 40457 ne
rect 17484 40456 17610 40457
tri 17484 40455 17485 40456 ne
rect 17485 40455 17610 40456
tri 17485 40454 17486 40455 ne
rect 17486 40454 17610 40455
tri 17486 40453 17487 40454 ne
rect 17487 40453 17610 40454
tri 17487 40452 17488 40453 ne
rect 17488 40452 17610 40453
tri 17488 40451 17489 40452 ne
rect 17489 40451 17610 40452
tri 17489 40450 17490 40451 ne
rect 17490 40450 17610 40451
tri 17490 40449 17491 40450 ne
rect 17491 40449 17610 40450
tri 17491 40448 17492 40449 ne
rect 17492 40448 17610 40449
tri 17492 40447 17493 40448 ne
rect 17493 40447 17610 40448
tri 17493 40446 17494 40447 ne
rect 17494 40446 17610 40447
tri 17494 40445 17495 40446 ne
rect 17495 40445 17610 40446
tri 17495 40444 17496 40445 ne
rect 17496 40444 17610 40445
tri 17496 40443 17497 40444 ne
rect 17497 40443 17610 40444
tri 17497 40442 17498 40443 ne
rect 17498 40442 17610 40443
tri 17498 40441 17499 40442 ne
rect 17499 40441 17610 40442
tri 17499 40440 17500 40441 ne
rect 17500 40440 17610 40441
tri 17500 40439 17501 40440 ne
rect 17501 40439 17610 40440
tri 17501 40438 17502 40439 ne
rect 17502 40438 17610 40439
tri 17502 40437 17503 40438 ne
rect 17503 40437 17610 40438
tri 17503 40436 17504 40437 ne
rect 17504 40436 17610 40437
tri 17504 40435 17505 40436 ne
rect 17505 40435 17610 40436
tri 17505 40434 17506 40435 ne
rect 17506 40434 17610 40435
tri 17506 40433 17507 40434 ne
rect 17507 40433 17610 40434
tri 17507 40432 17508 40433 ne
rect 17508 40432 17610 40433
tri 17508 40431 17509 40432 ne
rect 17509 40431 17610 40432
tri 17509 40430 17510 40431 ne
rect 17510 40430 17610 40431
tri 17510 40429 17511 40430 ne
rect 17511 40429 17610 40430
tri 17511 40428 17512 40429 ne
rect 17512 40428 17610 40429
tri 17512 40427 17513 40428 ne
rect 17513 40427 17610 40428
tri 17513 40426 17514 40427 ne
rect 17514 40426 17610 40427
tri 17514 40425 17515 40426 ne
rect 17515 40425 17610 40426
tri 17515 40424 17516 40425 ne
rect 17516 40424 17610 40425
tri 17516 40423 17517 40424 ne
rect 17517 40423 17610 40424
tri 17517 40422 17518 40423 ne
rect 17518 40422 17610 40423
rect 17656 40466 17746 40468
tri 17746 40466 17750 40470 sw
rect 17656 40422 17750 40466
tri 17518 40421 17519 40422 ne
rect 17519 40421 17750 40422
tri 17750 40421 17795 40466 sw
rect 70802 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
tri 17519 40376 17564 40421 ne
rect 17564 40376 17795 40421
tri 17795 40376 17840 40421 sw
tri 17564 40363 17577 40376 ne
rect 17577 40363 17840 40376
tri 17577 40318 17622 40363 ne
rect 17622 40336 17840 40363
rect 17622 40318 17742 40336
tri 17622 40273 17667 40318 ne
rect 17667 40290 17742 40318
rect 17788 40331 17840 40336
tri 17840 40331 17885 40376 sw
rect 70802 40372 71000 40430
rect 17788 40290 17885 40331
rect 17667 40286 17885 40290
tri 17885 40286 17930 40331 sw
rect 70802 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17667 40284 17930 40286
tri 17930 40284 17932 40286 sw
rect 17667 40273 17932 40284
tri 17667 40228 17712 40273 ne
rect 17712 40239 17932 40273
tri 17932 40239 17977 40284 sw
rect 70802 40268 71000 40326
rect 17712 40228 17977 40239
tri 17712 40194 17746 40228 ne
rect 17746 40204 17977 40228
rect 17746 40194 17874 40204
tri 17746 40183 17757 40194 ne
rect 17757 40183 17874 40194
tri 17757 40182 17758 40183 ne
rect 17758 40182 17874 40183
tri 17758 40181 17759 40182 ne
rect 17759 40181 17874 40182
tri 17759 40180 17760 40181 ne
rect 17760 40180 17874 40181
tri 17760 40179 17761 40180 ne
rect 17761 40179 17874 40180
tri 17761 40178 17762 40179 ne
rect 17762 40178 17874 40179
tri 17762 40177 17763 40178 ne
rect 17763 40177 17874 40178
tri 17763 40176 17764 40177 ne
rect 17764 40176 17874 40177
tri 17764 40175 17765 40176 ne
rect 17765 40175 17874 40176
tri 17765 40174 17766 40175 ne
rect 17766 40174 17874 40175
tri 17766 40173 17767 40174 ne
rect 17767 40173 17874 40174
tri 17767 40172 17768 40173 ne
rect 17768 40172 17874 40173
tri 17768 40171 17769 40172 ne
rect 17769 40171 17874 40172
tri 17769 40170 17770 40171 ne
rect 17770 40170 17874 40171
tri 17770 40169 17771 40170 ne
rect 17771 40169 17874 40170
tri 17771 40168 17772 40169 ne
rect 17772 40168 17874 40169
tri 17772 40167 17773 40168 ne
rect 17773 40167 17874 40168
tri 17773 40166 17774 40167 ne
rect 17774 40166 17874 40167
tri 17774 40165 17775 40166 ne
rect 17775 40165 17874 40166
tri 17775 40164 17776 40165 ne
rect 17776 40164 17874 40165
tri 17776 40163 17777 40164 ne
rect 17777 40163 17874 40164
tri 17777 40162 17778 40163 ne
rect 17778 40162 17874 40163
tri 17778 40161 17779 40162 ne
rect 17779 40161 17874 40162
tri 17779 40160 17780 40161 ne
rect 17780 40160 17874 40161
tri 17780 40159 17781 40160 ne
rect 17781 40159 17874 40160
tri 17781 40158 17782 40159 ne
rect 17782 40158 17874 40159
rect 17920 40194 17977 40204
tri 17977 40194 18022 40239 sw
rect 70802 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17920 40158 18022 40194
tri 17782 40157 17783 40158 ne
rect 17783 40157 18022 40158
tri 17783 40156 17784 40157 ne
rect 17784 40156 18022 40157
tri 17784 40155 17785 40156 ne
rect 17785 40155 18022 40156
tri 17785 40154 17786 40155 ne
rect 17786 40154 18022 40155
tri 17786 40153 17787 40154 ne
rect 17787 40153 18022 40154
tri 17787 40152 17788 40153 ne
rect 17788 40152 18022 40153
tri 17788 40151 17789 40152 ne
rect 17789 40151 18022 40152
tri 17789 40150 17790 40151 ne
rect 17790 40150 18022 40151
tri 17790 40149 17791 40150 ne
rect 17791 40149 18022 40150
tri 18022 40149 18067 40194 sw
rect 70802 40164 71000 40222
tri 17791 40148 17792 40149 ne
rect 17792 40148 18067 40149
tri 17792 40147 17793 40148 ne
rect 17793 40147 18067 40148
tri 17793 40146 17794 40147 ne
rect 17794 40146 18067 40147
tri 17794 40145 17795 40146 ne
rect 17795 40145 18067 40146
tri 18067 40145 18071 40149 sw
tri 17795 40100 17840 40145 ne
rect 17840 40104 18071 40145
tri 18071 40104 18112 40145 sw
rect 70802 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
rect 17840 40100 18112 40104
tri 17840 40055 17885 40100 ne
rect 17885 40072 18112 40100
rect 17885 40055 18006 40072
tri 17885 40043 17897 40055 ne
rect 17897 40043 18006 40055
tri 17897 39998 17942 40043 ne
rect 17942 40026 18006 40043
rect 18052 40059 18112 40072
tri 18112 40059 18157 40104 sw
rect 70802 40060 71000 40118
rect 18052 40026 18157 40059
rect 17942 40014 18157 40026
tri 18157 40014 18202 40059 sw
rect 70802 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 17942 40004 18202 40014
tri 18202 40004 18212 40014 sw
rect 17942 39998 18212 40004
tri 17942 39953 17987 39998 ne
rect 17987 39959 18212 39998
tri 18212 39959 18257 40004 sw
rect 17987 39953 18257 39959
tri 17987 39908 18032 39953 ne
rect 18032 39940 18257 39953
rect 18032 39908 18138 39940
tri 18032 39907 18033 39908 ne
rect 18033 39907 18138 39908
tri 18033 39906 18034 39907 ne
rect 18034 39906 18138 39907
tri 18034 39905 18035 39906 ne
rect 18035 39905 18138 39906
tri 18035 39904 18036 39905 ne
rect 18036 39904 18138 39905
tri 18036 39903 18037 39904 ne
rect 18037 39903 18138 39904
tri 18037 39902 18038 39903 ne
rect 18038 39902 18138 39903
tri 18038 39901 18039 39902 ne
rect 18039 39901 18138 39902
tri 18039 39900 18040 39901 ne
rect 18040 39900 18138 39901
tri 18040 39899 18041 39900 ne
rect 18041 39899 18138 39900
tri 18041 39898 18042 39899 ne
rect 18042 39898 18138 39899
tri 18042 39897 18043 39898 ne
rect 18043 39897 18138 39898
tri 18043 39896 18044 39897 ne
rect 18044 39896 18138 39897
tri 18044 39895 18045 39896 ne
rect 18045 39895 18138 39896
tri 18045 39894 18046 39895 ne
rect 18046 39894 18138 39895
rect 18184 39914 18257 39940
tri 18257 39914 18302 39959 sw
rect 70802 39956 71000 40014
rect 18184 39894 18302 39914
tri 18046 39893 18047 39894 ne
rect 18047 39893 18302 39894
tri 18047 39892 18048 39893 ne
rect 18048 39892 18302 39893
tri 18048 39891 18049 39892 ne
rect 18049 39891 18302 39892
tri 18049 39890 18050 39891 ne
rect 18050 39890 18302 39891
tri 18050 39889 18051 39890 ne
rect 18051 39889 18302 39890
tri 18051 39888 18052 39889 ne
rect 18052 39888 18302 39889
tri 18052 39887 18053 39888 ne
rect 18053 39887 18302 39888
tri 18053 39886 18054 39887 ne
rect 18054 39886 18302 39887
tri 18054 39885 18055 39886 ne
rect 18055 39885 18302 39886
tri 18055 39884 18056 39885 ne
rect 18056 39884 18302 39885
tri 18056 39883 18057 39884 ne
rect 18057 39883 18302 39884
tri 18057 39882 18058 39883 ne
rect 18058 39882 18302 39883
tri 18058 39881 18059 39882 ne
rect 18059 39881 18302 39882
tri 18059 39880 18060 39881 ne
rect 18060 39880 18302 39881
tri 18060 39879 18061 39880 ne
rect 18061 39879 18302 39880
tri 18061 39878 18062 39879 ne
rect 18062 39878 18302 39879
tri 18062 39877 18063 39878 ne
rect 18063 39877 18302 39878
tri 18063 39876 18064 39877 ne
rect 18064 39876 18302 39877
tri 18064 39875 18065 39876 ne
rect 18065 39875 18302 39876
tri 18065 39874 18066 39875 ne
rect 18066 39874 18302 39875
tri 18066 39873 18067 39874 ne
rect 18067 39873 18302 39874
tri 18067 39872 18068 39873 ne
rect 18068 39872 18302 39873
tri 18068 39871 18069 39872 ne
rect 18069 39871 18302 39872
tri 18069 39870 18070 39871 ne
rect 18070 39870 18302 39871
tri 18070 39869 18071 39870 ne
rect 18071 39869 18302 39870
tri 18302 39869 18347 39914 sw
rect 70802 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
tri 18071 39828 18112 39869 ne
rect 18112 39828 18347 39869
tri 18347 39828 18388 39869 sw
rect 70802 39852 71000 39910
tri 18112 39824 18116 39828 ne
rect 18116 39824 18388 39828
tri 18116 39783 18157 39824 ne
rect 18157 39808 18388 39824
rect 18157 39783 18270 39808
tri 18157 39738 18202 39783 ne
rect 18202 39762 18270 39783
rect 18316 39783 18388 39808
tri 18388 39783 18433 39828 sw
rect 70802 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39762 18433 39783
rect 18202 39738 18433 39762
tri 18433 39738 18478 39783 sw
rect 70802 39748 71000 39806
tri 18202 39693 18247 39738 ne
rect 18247 39693 18478 39738
tri 18478 39693 18523 39738 sw
rect 70802 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
tri 18247 39679 18261 39693 ne
rect 18261 39683 18523 39693
tri 18523 39683 18533 39693 sw
rect 18261 39679 18533 39683
tri 18261 39634 18306 39679 ne
rect 18306 39676 18533 39679
rect 18306 39634 18402 39676
tri 18306 39633 18307 39634 ne
rect 18307 39633 18402 39634
tri 18307 39632 18308 39633 ne
rect 18308 39632 18402 39633
tri 18308 39631 18309 39632 ne
rect 18309 39631 18402 39632
tri 18309 39630 18310 39631 ne
rect 18310 39630 18402 39631
rect 18448 39638 18533 39676
tri 18533 39638 18578 39683 sw
rect 70802 39644 71000 39702
rect 18448 39630 18578 39638
tri 18310 39629 18311 39630 ne
rect 18311 39629 18578 39630
tri 18311 39628 18312 39629 ne
rect 18312 39628 18578 39629
tri 18312 39627 18313 39628 ne
rect 18313 39627 18578 39628
tri 18313 39626 18314 39627 ne
rect 18314 39626 18578 39627
tri 18314 39625 18315 39626 ne
rect 18315 39625 18578 39626
tri 18315 39624 18316 39625 ne
rect 18316 39624 18578 39625
tri 18316 39623 18317 39624 ne
rect 18317 39623 18578 39624
tri 18317 39622 18318 39623 ne
rect 18318 39622 18578 39623
tri 18318 39621 18319 39622 ne
rect 18319 39621 18578 39622
tri 18319 39620 18320 39621 ne
rect 18320 39620 18578 39621
tri 18320 39619 18321 39620 ne
rect 18321 39619 18578 39620
tri 18321 39618 18322 39619 ne
rect 18322 39618 18578 39619
tri 18322 39617 18323 39618 ne
rect 18323 39617 18578 39618
tri 18323 39616 18324 39617 ne
rect 18324 39616 18578 39617
tri 18324 39615 18325 39616 ne
rect 18325 39615 18578 39616
tri 18325 39614 18326 39615 ne
rect 18326 39614 18578 39615
tri 18326 39613 18327 39614 ne
rect 18327 39613 18578 39614
tri 18327 39612 18328 39613 ne
rect 18328 39612 18578 39613
tri 18328 39611 18329 39612 ne
rect 18329 39611 18578 39612
tri 18329 39610 18330 39611 ne
rect 18330 39610 18578 39611
tri 18330 39609 18331 39610 ne
rect 18331 39609 18578 39610
tri 18331 39608 18332 39609 ne
rect 18332 39608 18578 39609
tri 18332 39607 18333 39608 ne
rect 18333 39607 18578 39608
tri 18333 39606 18334 39607 ne
rect 18334 39606 18578 39607
tri 18334 39605 18335 39606 ne
rect 18335 39605 18578 39606
tri 18335 39604 18336 39605 ne
rect 18336 39604 18578 39605
tri 18336 39603 18337 39604 ne
rect 18337 39603 18578 39604
tri 18337 39602 18338 39603 ne
rect 18338 39602 18578 39603
tri 18338 39601 18339 39602 ne
rect 18339 39601 18578 39602
tri 18339 39600 18340 39601 ne
rect 18340 39600 18578 39601
tri 18340 39599 18341 39600 ne
rect 18341 39599 18578 39600
tri 18341 39598 18342 39599 ne
rect 18342 39598 18578 39599
tri 18342 39597 18343 39598 ne
rect 18343 39597 18578 39598
tri 18343 39596 18344 39597 ne
rect 18344 39596 18578 39597
tri 18344 39595 18345 39596 ne
rect 18345 39595 18578 39596
tri 18345 39594 18346 39595 ne
rect 18346 39594 18578 39595
tri 18346 39593 18347 39594 ne
rect 18347 39593 18578 39594
tri 18578 39593 18623 39638 sw
rect 70802 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18347 39548 18392 39593 ne
rect 18392 39548 18623 39593
tri 18623 39548 18668 39593 sw
tri 18392 39503 18437 39548 ne
rect 18437 39544 18668 39548
rect 18437 39503 18534 39544
tri 18437 39462 18478 39503 ne
rect 18478 39498 18534 39503
rect 18580 39507 18668 39544
tri 18668 39507 18709 39548 sw
rect 70802 39540 71000 39598
rect 18580 39498 18709 39507
rect 18478 39462 18709 39498
tri 18709 39462 18754 39507 sw
rect 70802 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18478 39458 18482 39462 ne
rect 18482 39458 18754 39462
tri 18482 39417 18523 39458 ne
rect 18523 39417 18754 39458
tri 18754 39417 18799 39462 sw
rect 70802 39436 71000 39494
tri 18523 39372 18568 39417 ne
rect 18568 39412 18799 39417
rect 18568 39372 18666 39412
tri 18568 39359 18581 39372 ne
rect 18581 39366 18666 39372
rect 18712 39372 18799 39412
tri 18799 39372 18844 39417 sw
rect 70802 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 18712 39366 18844 39372
rect 18581 39362 18844 39366
tri 18844 39362 18854 39372 sw
rect 18581 39359 18854 39362
tri 18581 39358 18582 39359 ne
rect 18582 39358 18854 39359
tri 18582 39357 18583 39358 ne
rect 18583 39357 18854 39358
tri 18583 39356 18584 39357 ne
rect 18584 39356 18854 39357
tri 18584 39355 18585 39356 ne
rect 18585 39355 18854 39356
tri 18585 39354 18586 39355 ne
rect 18586 39354 18854 39355
tri 18586 39353 18587 39354 ne
rect 18587 39353 18854 39354
tri 18587 39352 18588 39353 ne
rect 18588 39352 18854 39353
tri 18588 39351 18589 39352 ne
rect 18589 39351 18854 39352
tri 18589 39350 18590 39351 ne
rect 18590 39350 18854 39351
tri 18590 39349 18591 39350 ne
rect 18591 39349 18854 39350
tri 18591 39348 18592 39349 ne
rect 18592 39348 18854 39349
tri 18592 39347 18593 39348 ne
rect 18593 39347 18854 39348
tri 18593 39346 18594 39347 ne
rect 18594 39346 18854 39347
tri 18594 39345 18595 39346 ne
rect 18595 39345 18854 39346
tri 18595 39344 18596 39345 ne
rect 18596 39344 18854 39345
tri 18596 39343 18597 39344 ne
rect 18597 39343 18854 39344
tri 18597 39342 18598 39343 ne
rect 18598 39342 18854 39343
tri 18598 39341 18599 39342 ne
rect 18599 39341 18854 39342
tri 18599 39340 18600 39341 ne
rect 18600 39340 18854 39341
tri 18600 39339 18601 39340 ne
rect 18601 39339 18854 39340
tri 18601 39338 18602 39339 ne
rect 18602 39338 18854 39339
tri 18602 39337 18603 39338 ne
rect 18603 39337 18854 39338
tri 18603 39336 18604 39337 ne
rect 18604 39336 18854 39337
tri 18604 39335 18605 39336 ne
rect 18605 39335 18854 39336
tri 18605 39334 18606 39335 ne
rect 18606 39334 18854 39335
tri 18606 39333 18607 39334 ne
rect 18607 39333 18854 39334
tri 18607 39332 18608 39333 ne
rect 18608 39332 18854 39333
tri 18608 39331 18609 39332 ne
rect 18609 39331 18854 39332
tri 18609 39330 18610 39331 ne
rect 18610 39330 18854 39331
tri 18610 39329 18611 39330 ne
rect 18611 39329 18854 39330
tri 18611 39328 18612 39329 ne
rect 18612 39328 18854 39329
tri 18612 39327 18613 39328 ne
rect 18613 39327 18854 39328
tri 18613 39326 18614 39327 ne
rect 18614 39326 18854 39327
tri 18614 39325 18615 39326 ne
rect 18615 39325 18854 39326
tri 18615 39324 18616 39325 ne
rect 18616 39324 18854 39325
tri 18616 39323 18617 39324 ne
rect 18617 39323 18854 39324
tri 18617 39322 18618 39323 ne
rect 18618 39322 18854 39323
tri 18618 39321 18619 39322 ne
rect 18619 39321 18854 39322
tri 18619 39320 18620 39321 ne
rect 18620 39320 18854 39321
tri 18620 39319 18621 39320 ne
rect 18621 39319 18854 39320
tri 18621 39318 18622 39319 ne
rect 18622 39318 18854 39319
tri 18622 39317 18623 39318 ne
rect 18623 39317 18854 39318
tri 18854 39317 18899 39362 sw
rect 70802 39332 71000 39390
tri 18623 39272 18668 39317 ne
rect 18668 39280 18899 39317
rect 18668 39272 18798 39280
tri 18668 39269 18671 39272 ne
rect 18671 39269 18798 39272
tri 18671 39224 18716 39269 ne
rect 18716 39234 18798 39269
rect 18844 39272 18899 39280
tri 18899 39272 18944 39317 sw
rect 70802 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 18844 39234 18944 39272
rect 18716 39227 18944 39234
tri 18944 39227 18989 39272 sw
rect 70802 39228 71000 39286
rect 18716 39224 18989 39227
tri 18716 39179 18761 39224 ne
rect 18761 39186 18989 39224
tri 18989 39186 19030 39227 sw
rect 18761 39179 19030 39186
tri 18761 39134 18806 39179 ne
rect 18806 39148 19030 39179
rect 18806 39134 18930 39148
tri 18806 39096 18844 39134 ne
rect 18844 39102 18930 39134
rect 18976 39141 19030 39148
tri 19030 39141 19075 39186 sw
rect 70802 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 18976 39102 19075 39141
rect 18844 39096 19075 39102
tri 19075 39096 19120 39141 sw
rect 70802 39124 71000 39182
tri 18844 39089 18851 39096 ne
rect 18851 39089 19120 39096
tri 18851 39085 18855 39089 ne
rect 18855 39085 19120 39089
tri 18855 39084 18856 39085 ne
rect 18856 39084 19120 39085
tri 18856 39083 18857 39084 ne
rect 18857 39083 19120 39084
tri 18857 39082 18858 39083 ne
rect 18858 39082 19120 39083
tri 18858 39081 18859 39082 ne
rect 18859 39081 19120 39082
tri 18859 39080 18860 39081 ne
rect 18860 39080 19120 39081
tri 18860 39079 18861 39080 ne
rect 18861 39079 19120 39080
tri 18861 39078 18862 39079 ne
rect 18862 39078 19120 39079
tri 18862 39077 18863 39078 ne
rect 18863 39077 19120 39078
tri 18863 39076 18864 39077 ne
rect 18864 39076 19120 39077
tri 18864 39075 18865 39076 ne
rect 18865 39075 19120 39076
tri 18865 39074 18866 39075 ne
rect 18866 39074 19120 39075
tri 18866 39073 18867 39074 ne
rect 18867 39073 19120 39074
tri 18867 39072 18868 39073 ne
rect 18868 39072 19120 39073
tri 18868 39071 18869 39072 ne
rect 18869 39071 19120 39072
tri 18869 39070 18870 39071 ne
rect 18870 39070 19120 39071
tri 18870 39069 18871 39070 ne
rect 18871 39069 19120 39070
tri 18871 39068 18872 39069 ne
rect 18872 39068 19120 39069
tri 18872 39067 18873 39068 ne
rect 18873 39067 19120 39068
tri 18873 39066 18874 39067 ne
rect 18874 39066 19120 39067
tri 18874 39065 18875 39066 ne
rect 18875 39065 19120 39066
tri 18875 39064 18876 39065 ne
rect 18876 39064 19120 39065
tri 18876 39063 18877 39064 ne
rect 18877 39063 19120 39064
tri 18877 39062 18878 39063 ne
rect 18878 39062 19120 39063
tri 18878 39061 18879 39062 ne
rect 18879 39061 19120 39062
tri 18879 39060 18880 39061 ne
rect 18880 39060 19120 39061
tri 18880 39059 18881 39060 ne
rect 18881 39059 19120 39060
tri 18881 39058 18882 39059 ne
rect 18882 39058 19120 39059
tri 18882 39057 18883 39058 ne
rect 18883 39057 19120 39058
tri 18883 39056 18884 39057 ne
rect 18884 39056 19120 39057
tri 18884 39055 18885 39056 ne
rect 18885 39055 19120 39056
tri 18885 39054 18886 39055 ne
rect 18886 39054 19120 39055
tri 18886 39053 18887 39054 ne
rect 18887 39053 19120 39054
tri 18887 39052 18888 39053 ne
rect 18888 39052 19120 39053
tri 18888 39051 18889 39052 ne
rect 18889 39051 19120 39052
tri 19120 39051 19165 39096 sw
rect 70802 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18889 39050 18890 39051 ne
rect 18890 39050 19165 39051
tri 18890 39049 18891 39050 ne
rect 18891 39049 19165 39050
tri 18891 39048 18892 39049 ne
rect 18892 39048 19165 39049
tri 18892 39047 18893 39048 ne
rect 18893 39047 19165 39048
tri 18893 39046 18894 39047 ne
rect 18894 39046 19165 39047
tri 18894 39045 18895 39046 ne
rect 18895 39045 19165 39046
tri 18895 39044 18896 39045 ne
rect 18896 39044 19165 39045
tri 18896 39043 18897 39044 ne
rect 18897 39043 19165 39044
tri 18897 39042 18898 39043 ne
rect 18898 39042 19165 39043
tri 18898 39041 18899 39042 ne
rect 18899 39041 19165 39042
tri 19165 39041 19175 39051 sw
tri 18899 38996 18944 39041 ne
rect 18944 39016 19175 39041
rect 18944 38996 19062 39016
tri 18944 38951 18989 38996 ne
rect 18989 38970 19062 38996
rect 19108 39006 19175 39016
tri 19175 39006 19210 39041 sw
rect 70802 39020 71000 39078
rect 19108 38970 19210 39006
rect 18989 38961 19210 38970
tri 19210 38961 19255 39006 sw
rect 70802 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 18989 38951 19255 38961
tri 18989 38949 18991 38951 ne
rect 18991 38949 19255 38951
tri 18991 38904 19036 38949 ne
rect 19036 38916 19255 38949
tri 19255 38916 19300 38961 sw
rect 70802 38916 71000 38974
rect 19036 38904 19300 38916
tri 19036 38859 19081 38904 ne
rect 19081 38900 19300 38904
tri 19300 38900 19316 38916 sw
rect 19081 38884 19316 38900
rect 19081 38859 19194 38884
tri 19081 38814 19126 38859 ne
rect 19126 38838 19194 38859
rect 19240 38855 19316 38884
tri 19316 38855 19361 38900 sw
rect 70802 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38838 19361 38855
rect 19126 38814 19361 38838
tri 19126 38810 19130 38814 ne
rect 19130 38810 19361 38814
tri 19361 38810 19406 38855 sw
rect 70802 38812 71000 38870
tri 19130 38809 19131 38810 ne
rect 19131 38809 19406 38810
tri 19131 38808 19132 38809 ne
rect 19132 38808 19406 38809
tri 19132 38807 19133 38808 ne
rect 19133 38807 19406 38808
tri 19133 38806 19134 38807 ne
rect 19134 38806 19406 38807
tri 19134 38805 19135 38806 ne
rect 19135 38805 19406 38806
tri 19135 38804 19136 38805 ne
rect 19136 38804 19406 38805
tri 19136 38803 19137 38804 ne
rect 19137 38803 19406 38804
tri 19137 38802 19138 38803 ne
rect 19138 38802 19406 38803
tri 19138 38801 19139 38802 ne
rect 19139 38801 19406 38802
tri 19139 38800 19140 38801 ne
rect 19140 38800 19406 38801
tri 19140 38799 19141 38800 ne
rect 19141 38799 19406 38800
tri 19141 38798 19142 38799 ne
rect 19142 38798 19406 38799
tri 19142 38797 19143 38798 ne
rect 19143 38797 19406 38798
tri 19143 38796 19144 38797 ne
rect 19144 38796 19406 38797
tri 19144 38795 19145 38796 ne
rect 19145 38795 19406 38796
tri 19145 38794 19146 38795 ne
rect 19146 38794 19406 38795
tri 19146 38793 19147 38794 ne
rect 19147 38793 19406 38794
tri 19147 38792 19148 38793 ne
rect 19148 38792 19406 38793
tri 19148 38791 19149 38792 ne
rect 19149 38791 19406 38792
tri 19149 38790 19150 38791 ne
rect 19150 38790 19406 38791
tri 19150 38789 19151 38790 ne
rect 19151 38789 19406 38790
tri 19151 38788 19152 38789 ne
rect 19152 38788 19406 38789
tri 19152 38787 19153 38788 ne
rect 19153 38787 19406 38788
tri 19153 38786 19154 38787 ne
rect 19154 38786 19406 38787
tri 19154 38785 19155 38786 ne
rect 19155 38785 19406 38786
tri 19155 38784 19156 38785 ne
rect 19156 38784 19406 38785
tri 19156 38783 19157 38784 ne
rect 19157 38783 19406 38784
tri 19157 38782 19158 38783 ne
rect 19158 38782 19406 38783
tri 19158 38781 19159 38782 ne
rect 19159 38781 19406 38782
tri 19159 38780 19160 38781 ne
rect 19160 38780 19406 38781
tri 19160 38779 19161 38780 ne
rect 19161 38779 19406 38780
tri 19161 38778 19162 38779 ne
rect 19162 38778 19406 38779
tri 19162 38777 19163 38778 ne
rect 19163 38777 19406 38778
tri 19163 38776 19164 38777 ne
rect 19164 38776 19406 38777
tri 19164 38775 19165 38776 ne
rect 19165 38775 19406 38776
tri 19165 38774 19166 38775 ne
rect 19166 38774 19406 38775
tri 19166 38773 19167 38774 ne
rect 19167 38773 19406 38774
tri 19167 38772 19168 38773 ne
rect 19168 38772 19406 38773
tri 19168 38771 19169 38772 ne
rect 19169 38771 19406 38772
tri 19169 38770 19170 38771 ne
rect 19170 38770 19406 38771
tri 19170 38769 19171 38770 ne
rect 19171 38769 19406 38770
tri 19171 38768 19172 38769 ne
rect 19172 38768 19406 38769
tri 19172 38767 19173 38768 ne
rect 19173 38767 19406 38768
tri 19173 38766 19174 38767 ne
rect 19174 38766 19406 38767
tri 19174 38765 19175 38766 ne
rect 19175 38765 19406 38766
tri 19406 38765 19451 38810 sw
rect 70802 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19175 38730 19210 38765 ne
rect 19210 38752 19451 38765
rect 19210 38730 19326 38752
tri 19210 38720 19220 38730 ne
rect 19220 38720 19326 38730
tri 19220 38685 19255 38720 ne
rect 19255 38706 19326 38720
rect 19372 38730 19451 38752
tri 19451 38730 19486 38765 sw
rect 19372 38706 19486 38730
rect 19255 38685 19486 38706
tri 19486 38685 19531 38730 sw
rect 70802 38708 71000 38766
tri 19255 38640 19300 38685 ne
rect 19300 38640 19531 38685
tri 19531 38640 19576 38685 sw
rect 70802 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19300 38595 19345 38640 ne
rect 19345 38620 19576 38640
rect 19345 38595 19458 38620
tri 19345 38584 19356 38595 ne
rect 19356 38584 19458 38595
tri 19356 38539 19401 38584 ne
rect 19401 38574 19458 38584
rect 19504 38595 19576 38620
tri 19576 38595 19621 38640 sw
rect 70802 38604 71000 38662
rect 19504 38579 19621 38595
tri 19621 38579 19637 38595 sw
rect 19504 38574 19637 38579
rect 19401 38539 19637 38574
tri 19401 38536 19404 38539 ne
rect 19404 38536 19637 38539
tri 19404 38535 19405 38536 ne
rect 19405 38535 19637 38536
tri 19405 38534 19406 38535 ne
rect 19406 38534 19637 38535
tri 19637 38534 19682 38579 sw
rect 70802 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
tri 19406 38533 19407 38534 ne
rect 19407 38533 19682 38534
tri 19407 38532 19408 38533 ne
rect 19408 38532 19682 38533
tri 19408 38531 19409 38532 ne
rect 19409 38531 19682 38532
tri 19409 38530 19410 38531 ne
rect 19410 38530 19682 38531
tri 19410 38529 19411 38530 ne
rect 19411 38529 19682 38530
tri 19411 38528 19412 38529 ne
rect 19412 38528 19682 38529
tri 19412 38527 19413 38528 ne
rect 19413 38527 19682 38528
tri 19413 38526 19414 38527 ne
rect 19414 38526 19682 38527
tri 19414 38525 19415 38526 ne
rect 19415 38525 19682 38526
tri 19415 38524 19416 38525 ne
rect 19416 38524 19682 38525
tri 19416 38523 19417 38524 ne
rect 19417 38523 19682 38524
tri 19417 38522 19418 38523 ne
rect 19418 38522 19682 38523
tri 19418 38521 19419 38522 ne
rect 19419 38521 19682 38522
tri 19419 38520 19420 38521 ne
rect 19420 38520 19682 38521
tri 19420 38519 19421 38520 ne
rect 19421 38519 19682 38520
tri 19421 38518 19422 38519 ne
rect 19422 38518 19682 38519
tri 19422 38517 19423 38518 ne
rect 19423 38517 19682 38518
tri 19423 38516 19424 38517 ne
rect 19424 38516 19682 38517
tri 19424 38515 19425 38516 ne
rect 19425 38515 19682 38516
tri 19425 38514 19426 38515 ne
rect 19426 38514 19682 38515
tri 19426 38513 19427 38514 ne
rect 19427 38513 19682 38514
tri 19427 38512 19428 38513 ne
rect 19428 38512 19682 38513
tri 19428 38511 19429 38512 ne
rect 19429 38511 19682 38512
tri 19429 38510 19430 38511 ne
rect 19430 38510 19682 38511
tri 19430 38509 19431 38510 ne
rect 19431 38509 19682 38510
tri 19431 38508 19432 38509 ne
rect 19432 38508 19682 38509
tri 19432 38507 19433 38508 ne
rect 19433 38507 19682 38508
tri 19433 38506 19434 38507 ne
rect 19434 38506 19682 38507
tri 19434 38505 19435 38506 ne
rect 19435 38505 19682 38506
tri 19435 38504 19436 38505 ne
rect 19436 38504 19682 38505
tri 19436 38503 19437 38504 ne
rect 19437 38503 19682 38504
tri 19437 38502 19438 38503 ne
rect 19438 38502 19682 38503
tri 19438 38501 19439 38502 ne
rect 19439 38501 19682 38502
tri 19439 38500 19440 38501 ne
rect 19440 38500 19682 38501
tri 19440 38499 19441 38500 ne
rect 19441 38499 19682 38500
tri 19441 38498 19442 38499 ne
rect 19442 38498 19682 38499
tri 19442 38497 19443 38498 ne
rect 19443 38497 19682 38498
tri 19443 38496 19444 38497 ne
rect 19444 38496 19682 38497
tri 19444 38495 19445 38496 ne
rect 19445 38495 19682 38496
tri 19445 38494 19446 38495 ne
rect 19446 38494 19682 38495
tri 19446 38493 19447 38494 ne
rect 19447 38493 19682 38494
tri 19447 38492 19448 38493 ne
rect 19448 38492 19682 38493
tri 19448 38491 19449 38492 ne
rect 19449 38491 19682 38492
tri 19449 38490 19450 38491 ne
rect 19450 38490 19682 38491
tri 19450 38489 19451 38490 ne
rect 19451 38489 19682 38490
tri 19682 38489 19727 38534 sw
rect 70802 38500 71000 38558
tri 19451 38444 19496 38489 ne
rect 19496 38488 19727 38489
rect 19496 38444 19590 38488
tri 19496 38399 19541 38444 ne
rect 19541 38442 19590 38444
rect 19636 38444 19727 38488
tri 19727 38444 19772 38489 sw
rect 70802 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19772 38444
rect 19541 38409 19772 38442
tri 19772 38409 19807 38444 sw
rect 19541 38399 19807 38409
tri 19541 38364 19576 38399 ne
rect 19576 38364 19807 38399
tri 19807 38364 19852 38409 sw
rect 70802 38396 71000 38454
tri 19576 38354 19586 38364 ne
rect 19586 38356 19852 38364
rect 19586 38354 19722 38356
tri 19586 38319 19621 38354 ne
rect 19621 38319 19722 38354
tri 19621 38274 19666 38319 ne
rect 19666 38310 19722 38319
rect 19768 38319 19852 38356
tri 19852 38319 19897 38364 sw
rect 70802 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 19768 38310 19897 38319
rect 19666 38274 19897 38310
tri 19897 38274 19942 38319 sw
rect 70802 38292 71000 38350
tri 19666 38261 19679 38274 ne
rect 19679 38261 19942 38274
tri 19679 38260 19680 38261 ne
rect 19680 38260 19942 38261
tri 19680 38259 19681 38260 ne
rect 19681 38259 19942 38260
tri 19681 38258 19682 38259 ne
rect 19682 38258 19942 38259
tri 19942 38258 19958 38274 sw
tri 19682 38257 19683 38258 ne
rect 19683 38257 19958 38258
tri 19683 38256 19684 38257 ne
rect 19684 38256 19958 38257
tri 19684 38255 19685 38256 ne
rect 19685 38255 19958 38256
tri 19685 38254 19686 38255 ne
rect 19686 38254 19958 38255
tri 19686 38253 19687 38254 ne
rect 19687 38253 19958 38254
tri 19687 38252 19688 38253 ne
rect 19688 38252 19958 38253
tri 19688 38251 19689 38252 ne
rect 19689 38251 19958 38252
tri 19689 38250 19690 38251 ne
rect 19690 38250 19958 38251
tri 19690 38249 19691 38250 ne
rect 19691 38249 19958 38250
tri 19691 38248 19692 38249 ne
rect 19692 38248 19958 38249
tri 19692 38247 19693 38248 ne
rect 19693 38247 19958 38248
tri 19693 38246 19694 38247 ne
rect 19694 38246 19958 38247
tri 19694 38245 19695 38246 ne
rect 19695 38245 19958 38246
tri 19695 38244 19696 38245 ne
rect 19696 38244 19958 38245
tri 19696 38243 19697 38244 ne
rect 19697 38243 19958 38244
tri 19697 38242 19698 38243 ne
rect 19698 38242 19958 38243
tri 19698 38241 19699 38242 ne
rect 19699 38241 19958 38242
tri 19699 38240 19700 38241 ne
rect 19700 38240 19958 38241
tri 19700 38239 19701 38240 ne
rect 19701 38239 19958 38240
tri 19701 38238 19702 38239 ne
rect 19702 38238 19958 38239
tri 19702 38237 19703 38238 ne
rect 19703 38237 19958 38238
tri 19703 38236 19704 38237 ne
rect 19704 38236 19958 38237
tri 19704 38235 19705 38236 ne
rect 19705 38235 19958 38236
tri 19705 38234 19706 38235 ne
rect 19706 38234 19958 38235
tri 19706 38233 19707 38234 ne
rect 19707 38233 19958 38234
tri 19707 38232 19708 38233 ne
rect 19708 38232 19958 38233
tri 19708 38231 19709 38232 ne
rect 19709 38231 19958 38232
tri 19709 38230 19710 38231 ne
rect 19710 38230 19958 38231
tri 19710 38229 19711 38230 ne
rect 19711 38229 19958 38230
tri 19711 38228 19712 38229 ne
rect 19712 38228 19958 38229
tri 19712 38227 19713 38228 ne
rect 19713 38227 19958 38228
tri 19713 38226 19714 38227 ne
rect 19714 38226 19958 38227
tri 19714 38225 19715 38226 ne
rect 19715 38225 19958 38226
tri 19715 38224 19716 38225 ne
rect 19716 38224 19958 38225
tri 19716 38223 19717 38224 ne
rect 19717 38223 19854 38224
tri 19717 38222 19718 38223 ne
rect 19718 38222 19854 38223
tri 19718 38221 19719 38222 ne
rect 19719 38221 19854 38222
tri 19719 38220 19720 38221 ne
rect 19720 38220 19854 38221
tri 19720 38219 19721 38220 ne
rect 19721 38219 19854 38220
tri 19721 38218 19722 38219 ne
rect 19722 38218 19854 38219
tri 19722 38217 19723 38218 ne
rect 19723 38217 19854 38218
tri 19723 38216 19724 38217 ne
rect 19724 38216 19854 38217
tri 19724 38215 19725 38216 ne
rect 19725 38215 19854 38216
tri 19725 38214 19726 38215 ne
rect 19726 38214 19854 38215
tri 19726 38213 19727 38214 ne
rect 19727 38213 19854 38214
tri 19727 38174 19766 38213 ne
rect 19766 38178 19854 38213
rect 19900 38213 19958 38224
tri 19958 38213 20003 38258 sw
rect 70802 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 19900 38178 20003 38213
rect 19766 38174 20003 38178
tri 19766 38129 19811 38174 ne
rect 19811 38168 20003 38174
tri 20003 38168 20048 38213 sw
rect 70802 38188 71000 38246
rect 19811 38129 20048 38168
tri 19811 38084 19856 38129 ne
rect 19856 38123 20048 38129
tri 20048 38123 20093 38168 sw
rect 70802 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
rect 19856 38092 20093 38123
rect 19856 38084 19986 38092
tri 19856 38039 19901 38084 ne
rect 19901 38046 19986 38084
rect 20032 38088 20093 38092
tri 20093 38088 20128 38123 sw
rect 20032 38046 20128 38088
rect 19901 38043 20128 38046
tri 20128 38043 20173 38088 sw
rect 70802 38084 71000 38142
rect 19901 38039 20173 38043
tri 19901 37998 19942 38039 ne
rect 19942 37998 20173 38039
tri 20173 37998 20218 38043 sw
rect 70802 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
tri 19942 37994 19946 37998 ne
rect 19946 37994 20218 37998
tri 19946 37987 19953 37994 ne
rect 19953 37987 20218 37994
tri 19953 37986 19954 37987 ne
rect 19954 37986 20218 37987
tri 19954 37985 19955 37986 ne
rect 19955 37985 20218 37986
tri 19955 37984 19956 37985 ne
rect 19956 37984 20218 37985
tri 19956 37983 19957 37984 ne
rect 19957 37983 20218 37984
tri 19957 37982 19958 37983 ne
rect 19958 37982 20218 37983
tri 19958 37981 19959 37982 ne
rect 19959 37981 20218 37982
tri 19959 37980 19960 37981 ne
rect 19960 37980 20218 37981
tri 19960 37979 19961 37980 ne
rect 19961 37979 20218 37980
tri 19961 37978 19962 37979 ne
rect 19962 37978 20218 37979
tri 19962 37977 19963 37978 ne
rect 19963 37977 20218 37978
tri 19963 37976 19964 37977 ne
rect 19964 37976 20218 37977
tri 19964 37975 19965 37976 ne
rect 19965 37975 20218 37976
tri 19965 37974 19966 37975 ne
rect 19966 37974 20218 37975
tri 19966 37973 19967 37974 ne
rect 19967 37973 20218 37974
tri 19967 37972 19968 37973 ne
rect 19968 37972 20218 37973
tri 19968 37971 19969 37972 ne
rect 19969 37971 20218 37972
tri 19969 37970 19970 37971 ne
rect 19970 37970 20218 37971
tri 19970 37969 19971 37970 ne
rect 19971 37969 20218 37970
tri 19971 37968 19972 37969 ne
rect 19972 37968 20218 37969
tri 19972 37967 19973 37968 ne
rect 19973 37967 20218 37968
tri 19973 37966 19974 37967 ne
rect 19974 37966 20218 37967
tri 19974 37965 19975 37966 ne
rect 19975 37965 20218 37966
tri 19975 37964 19976 37965 ne
rect 19976 37964 20218 37965
tri 19976 37963 19977 37964 ne
rect 19977 37963 20218 37964
tri 19977 37962 19978 37963 ne
rect 19978 37962 20218 37963
tri 19978 37961 19979 37962 ne
rect 19979 37961 20218 37962
tri 19979 37960 19980 37961 ne
rect 19980 37960 20218 37961
tri 19980 37959 19981 37960 ne
rect 19981 37959 20118 37960
tri 19981 37958 19982 37959 ne
rect 19982 37958 20118 37959
tri 19982 37957 19983 37958 ne
rect 19983 37957 20118 37958
tri 19983 37956 19984 37957 ne
rect 19984 37956 20118 37957
tri 19984 37955 19985 37956 ne
rect 19985 37955 20118 37956
tri 19985 37954 19986 37955 ne
rect 19986 37954 20118 37955
tri 19986 37953 19987 37954 ne
rect 19987 37953 20118 37954
tri 19987 37952 19988 37953 ne
rect 19988 37952 20118 37953
tri 19988 37951 19989 37952 ne
rect 19989 37951 20118 37952
tri 19989 37950 19990 37951 ne
rect 19990 37950 20118 37951
tri 19990 37949 19991 37950 ne
rect 19991 37949 20118 37950
tri 19991 37948 19992 37949 ne
rect 19992 37948 20118 37949
tri 19992 37947 19993 37948 ne
rect 19993 37947 20118 37948
tri 19993 37946 19994 37947 ne
rect 19994 37946 20118 37947
tri 19994 37945 19995 37946 ne
rect 19995 37945 20118 37946
tri 19995 37944 19996 37945 ne
rect 19996 37944 20118 37945
tri 19996 37943 19997 37944 ne
rect 19997 37943 20118 37944
tri 19997 37942 19998 37943 ne
rect 19998 37942 20118 37943
tri 19998 37941 19999 37942 ne
rect 19999 37941 20118 37942
tri 19999 37940 20000 37941 ne
rect 20000 37940 20118 37941
tri 20000 37939 20001 37940 ne
rect 20001 37939 20118 37940
tri 20001 37938 20002 37939 ne
rect 20002 37938 20118 37939
tri 20002 37937 20003 37938 ne
rect 20003 37937 20118 37938
tri 20003 37892 20048 37937 ne
rect 20048 37914 20118 37937
rect 20164 37953 20218 37960
tri 20218 37953 20263 37998 sw
rect 70802 37980 71000 38038
rect 20164 37937 20263 37953
tri 20263 37937 20279 37953 sw
rect 20164 37914 20279 37937
rect 20048 37908 20279 37914
tri 20279 37908 20308 37937 sw
rect 70802 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 20048 37892 20308 37908
tri 20048 37855 20085 37892 ne
rect 20085 37863 20308 37892
tri 20308 37863 20353 37908 sw
rect 70802 37876 71000 37934
rect 20085 37855 20353 37863
tri 20085 37810 20130 37855 ne
rect 20130 37828 20353 37855
rect 20130 37810 20250 37828
tri 20130 37765 20175 37810 ne
rect 20175 37782 20250 37810
rect 20296 37818 20353 37828
tri 20353 37818 20398 37863 sw
rect 70802 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 20296 37796 20398 37818
tri 20398 37796 20420 37818 sw
rect 20296 37782 20420 37796
rect 20175 37765 20420 37782
tri 20175 37720 20220 37765 ne
rect 20220 37751 20420 37765
tri 20420 37751 20465 37796 sw
rect 70802 37772 71000 37830
rect 20220 37720 20465 37751
tri 20220 37713 20227 37720 ne
rect 20227 37713 20465 37720
tri 20227 37712 20228 37713 ne
rect 20228 37712 20465 37713
tri 20228 37711 20229 37712 ne
rect 20229 37711 20465 37712
tri 20229 37710 20230 37711 ne
rect 20230 37710 20465 37711
tri 20230 37709 20231 37710 ne
rect 20231 37709 20465 37710
tri 20231 37708 20232 37709 ne
rect 20232 37708 20465 37709
tri 20232 37707 20233 37708 ne
rect 20233 37707 20465 37708
tri 20233 37706 20234 37707 ne
rect 20234 37706 20465 37707
tri 20465 37706 20510 37751 sw
rect 70802 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
tri 20234 37705 20235 37706 ne
rect 20235 37705 20510 37706
tri 20235 37704 20236 37705 ne
rect 20236 37704 20510 37705
tri 20236 37703 20237 37704 ne
rect 20237 37703 20510 37704
tri 20237 37702 20238 37703 ne
rect 20238 37702 20510 37703
tri 20238 37701 20239 37702 ne
rect 20239 37701 20510 37702
tri 20239 37700 20240 37701 ne
rect 20240 37700 20510 37701
tri 20240 37699 20241 37700 ne
rect 20241 37699 20510 37700
tri 20241 37698 20242 37699 ne
rect 20242 37698 20510 37699
tri 20242 37697 20243 37698 ne
rect 20243 37697 20510 37698
tri 20243 37696 20244 37697 ne
rect 20244 37696 20510 37697
tri 20244 37695 20245 37696 ne
rect 20245 37695 20382 37696
tri 20245 37694 20246 37695 ne
rect 20246 37694 20382 37695
tri 20246 37693 20247 37694 ne
rect 20247 37693 20382 37694
tri 20247 37692 20248 37693 ne
rect 20248 37692 20382 37693
tri 20248 37691 20249 37692 ne
rect 20249 37691 20382 37692
tri 20249 37690 20250 37691 ne
rect 20250 37690 20382 37691
tri 20250 37689 20251 37690 ne
rect 20251 37689 20382 37690
tri 20251 37688 20252 37689 ne
rect 20252 37688 20382 37689
tri 20252 37687 20253 37688 ne
rect 20253 37687 20382 37688
tri 20253 37686 20254 37687 ne
rect 20254 37686 20382 37687
tri 20254 37685 20255 37686 ne
rect 20255 37685 20382 37686
tri 20255 37684 20256 37685 ne
rect 20256 37684 20382 37685
tri 20256 37683 20257 37684 ne
rect 20257 37683 20382 37684
tri 20257 37682 20258 37683 ne
rect 20258 37682 20382 37683
tri 20258 37681 20259 37682 ne
rect 20259 37681 20382 37682
tri 20259 37680 20260 37681 ne
rect 20260 37680 20382 37681
tri 20260 37679 20261 37680 ne
rect 20261 37679 20382 37680
tri 20261 37678 20262 37679 ne
rect 20262 37678 20382 37679
tri 20262 37677 20263 37678 ne
rect 20263 37677 20382 37678
tri 20263 37676 20264 37677 ne
rect 20264 37676 20382 37677
tri 20264 37675 20265 37676 ne
rect 20265 37675 20382 37676
tri 20265 37674 20266 37675 ne
rect 20266 37674 20382 37675
tri 20266 37673 20267 37674 ne
rect 20267 37673 20382 37674
tri 20267 37672 20268 37673 ne
rect 20268 37672 20382 37673
tri 20268 37671 20269 37672 ne
rect 20269 37671 20382 37672
tri 20269 37670 20270 37671 ne
rect 20270 37670 20382 37671
tri 20270 37669 20271 37670 ne
rect 20271 37669 20382 37670
tri 20271 37668 20272 37669 ne
rect 20272 37668 20382 37669
tri 20272 37667 20273 37668 ne
rect 20273 37667 20382 37668
tri 20273 37666 20274 37667 ne
rect 20274 37666 20382 37667
tri 20274 37665 20275 37666 ne
rect 20275 37665 20382 37666
tri 20275 37664 20276 37665 ne
rect 20276 37664 20382 37665
tri 20276 37663 20277 37664 ne
rect 20277 37663 20382 37664
tri 20277 37662 20278 37663 ne
rect 20278 37662 20382 37663
tri 20278 37661 20279 37662 ne
rect 20279 37661 20382 37662
tri 20279 37632 20308 37661 ne
rect 20308 37650 20382 37661
rect 20428 37661 20510 37696
tri 20510 37661 20555 37706 sw
rect 70802 37668 71000 37726
rect 20428 37650 20555 37661
rect 20308 37632 20555 37650
tri 20555 37632 20584 37661 sw
tri 20308 37616 20324 37632 ne
rect 20324 37616 20584 37632
tri 20324 37587 20353 37616 ne
rect 20353 37587 20584 37616
tri 20584 37587 20629 37632 sw
rect 70802 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20353 37542 20398 37587 ne
rect 20398 37564 20629 37587
rect 20398 37542 20514 37564
tri 20398 37497 20443 37542 ne
rect 20443 37518 20514 37542
rect 20560 37542 20629 37564
tri 20629 37542 20674 37587 sw
rect 70802 37564 71000 37622
rect 20560 37518 20674 37542
rect 20443 37497 20674 37518
tri 20674 37497 20719 37542 sw
rect 70802 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
tri 20443 37490 20450 37497 ne
rect 20450 37490 20719 37497
tri 20450 37445 20495 37490 ne
rect 20495 37475 20719 37490
tri 20719 37475 20741 37497 sw
rect 20495 37445 20741 37475
tri 20495 37438 20502 37445 ne
rect 20502 37438 20741 37445
tri 20502 37437 20503 37438 ne
rect 20503 37437 20741 37438
tri 20503 37436 20504 37437 ne
rect 20504 37436 20741 37437
tri 20504 37435 20505 37436 ne
rect 20505 37435 20741 37436
tri 20505 37434 20506 37435 ne
rect 20506 37434 20741 37435
tri 20506 37433 20507 37434 ne
rect 20507 37433 20741 37434
tri 20507 37432 20508 37433 ne
rect 20508 37432 20741 37433
tri 20508 37431 20509 37432 ne
rect 20509 37431 20646 37432
tri 20509 37430 20510 37431 ne
rect 20510 37430 20646 37431
tri 20510 37429 20511 37430 ne
rect 20511 37429 20646 37430
tri 20511 37428 20512 37429 ne
rect 20512 37428 20646 37429
tri 20512 37427 20513 37428 ne
rect 20513 37427 20646 37428
tri 20513 37426 20514 37427 ne
rect 20514 37426 20646 37427
tri 20514 37425 20515 37426 ne
rect 20515 37425 20646 37426
tri 20515 37424 20516 37425 ne
rect 20516 37424 20646 37425
tri 20516 37423 20517 37424 ne
rect 20517 37423 20646 37424
tri 20517 37422 20518 37423 ne
rect 20518 37422 20646 37423
tri 20518 37421 20519 37422 ne
rect 20519 37421 20646 37422
tri 20519 37420 20520 37421 ne
rect 20520 37420 20646 37421
tri 20520 37419 20521 37420 ne
rect 20521 37419 20646 37420
tri 20521 37418 20522 37419 ne
rect 20522 37418 20646 37419
tri 20522 37417 20523 37418 ne
rect 20523 37417 20646 37418
tri 20523 37416 20524 37417 ne
rect 20524 37416 20646 37417
tri 20524 37415 20525 37416 ne
rect 20525 37415 20646 37416
tri 20525 37414 20526 37415 ne
rect 20526 37414 20646 37415
tri 20526 37413 20527 37414 ne
rect 20527 37413 20646 37414
tri 20527 37412 20528 37413 ne
rect 20528 37412 20646 37413
tri 20528 37411 20529 37412 ne
rect 20529 37411 20646 37412
tri 20529 37410 20530 37411 ne
rect 20530 37410 20646 37411
tri 20530 37409 20531 37410 ne
rect 20531 37409 20646 37410
tri 20531 37408 20532 37409 ne
rect 20532 37408 20646 37409
tri 20532 37407 20533 37408 ne
rect 20533 37407 20646 37408
tri 20533 37406 20534 37407 ne
rect 20534 37406 20646 37407
tri 20534 37405 20535 37406 ne
rect 20535 37405 20646 37406
tri 20535 37404 20536 37405 ne
rect 20536 37404 20646 37405
tri 20536 37403 20537 37404 ne
rect 20537 37403 20646 37404
tri 20537 37402 20538 37403 ne
rect 20538 37402 20646 37403
tri 20538 37401 20539 37402 ne
rect 20539 37401 20646 37402
tri 20539 37400 20540 37401 ne
rect 20540 37400 20646 37401
tri 20540 37399 20541 37400 ne
rect 20541 37399 20646 37400
tri 20541 37398 20542 37399 ne
rect 20542 37398 20646 37399
tri 20542 37397 20543 37398 ne
rect 20543 37397 20646 37398
tri 20543 37396 20544 37397 ne
rect 20544 37396 20646 37397
tri 20544 37395 20545 37396 ne
rect 20545 37395 20646 37396
tri 20545 37394 20546 37395 ne
rect 20546 37394 20646 37395
tri 20546 37393 20547 37394 ne
rect 20547 37393 20646 37394
tri 20547 37392 20548 37393 ne
rect 20548 37392 20646 37393
tri 20548 37391 20549 37392 ne
rect 20549 37391 20646 37392
tri 20549 37390 20550 37391 ne
rect 20550 37390 20646 37391
tri 20550 37389 20551 37390 ne
rect 20551 37389 20646 37390
tri 20551 37388 20552 37389 ne
rect 20552 37388 20646 37389
tri 20552 37387 20553 37388 ne
rect 20553 37387 20646 37388
tri 20553 37386 20554 37387 ne
rect 20554 37386 20646 37387
rect 20692 37430 20741 37432
tri 20741 37430 20786 37475 sw
rect 70802 37460 71000 37518
rect 20692 37386 20786 37430
tri 20554 37385 20555 37386 ne
rect 20555 37385 20786 37386
tri 20786 37385 20831 37430 sw
rect 70802 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
tri 20555 37340 20600 37385 ne
rect 20600 37340 20831 37385
tri 20831 37340 20876 37385 sw
rect 70802 37356 71000 37414
tri 20600 37295 20645 37340 ne
rect 20645 37311 20876 37340
tri 20876 37311 20905 37340 sw
rect 20645 37300 20905 37311
rect 20645 37295 20778 37300
tri 20645 37266 20674 37295 ne
rect 20674 37266 20778 37295
tri 20674 37250 20690 37266 ne
rect 20690 37254 20778 37266
rect 20824 37266 20905 37300
tri 20905 37266 20950 37311 sw
rect 70802 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 20824 37254 20950 37266
rect 20690 37250 20950 37254
tri 20690 37221 20719 37250 ne
rect 20719 37221 20950 37250
tri 20950 37221 20995 37266 sw
rect 70802 37252 71000 37310
tri 20719 37176 20764 37221 ne
rect 20764 37176 20995 37221
tri 20995 37176 21040 37221 sw
rect 70802 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
tri 20764 37164 20776 37176 ne
rect 20776 37168 21040 37176
rect 20776 37164 20910 37168
tri 20776 37163 20777 37164 ne
rect 20777 37163 20910 37164
tri 20777 37162 20778 37163 ne
rect 20778 37162 20910 37163
tri 20778 37161 20779 37162 ne
rect 20779 37161 20910 37162
tri 20779 37160 20780 37161 ne
rect 20780 37160 20910 37161
tri 20780 37159 20781 37160 ne
rect 20781 37159 20910 37160
tri 20781 37158 20782 37159 ne
rect 20782 37158 20910 37159
tri 20782 37157 20783 37158 ne
rect 20783 37157 20910 37158
tri 20783 37156 20784 37157 ne
rect 20784 37156 20910 37157
tri 20784 37155 20785 37156 ne
rect 20785 37155 20910 37156
tri 20785 37154 20786 37155 ne
rect 20786 37154 20910 37155
tri 20786 37153 20787 37154 ne
rect 20787 37153 20910 37154
tri 20787 37152 20788 37153 ne
rect 20788 37152 20910 37153
tri 20788 37151 20789 37152 ne
rect 20789 37151 20910 37152
tri 20789 37150 20790 37151 ne
rect 20790 37150 20910 37151
tri 20790 37149 20791 37150 ne
rect 20791 37149 20910 37150
tri 20791 37148 20792 37149 ne
rect 20792 37148 20910 37149
tri 20792 37147 20793 37148 ne
rect 20793 37147 20910 37148
tri 20793 37146 20794 37147 ne
rect 20794 37146 20910 37147
tri 20794 37145 20795 37146 ne
rect 20795 37145 20910 37146
tri 20795 37144 20796 37145 ne
rect 20796 37144 20910 37145
tri 20796 37143 20797 37144 ne
rect 20797 37143 20910 37144
tri 20797 37142 20798 37143 ne
rect 20798 37142 20910 37143
tri 20798 37141 20799 37142 ne
rect 20799 37141 20910 37142
tri 20799 37140 20800 37141 ne
rect 20800 37140 20910 37141
tri 20800 37139 20801 37140 ne
rect 20801 37139 20910 37140
tri 20801 37138 20802 37139 ne
rect 20802 37138 20910 37139
tri 20802 37137 20803 37138 ne
rect 20803 37137 20910 37138
tri 20803 37136 20804 37137 ne
rect 20804 37136 20910 37137
tri 20804 37135 20805 37136 ne
rect 20805 37135 20910 37136
tri 20805 37134 20806 37135 ne
rect 20806 37134 20910 37135
tri 20806 37133 20807 37134 ne
rect 20807 37133 20910 37134
tri 20807 37132 20808 37133 ne
rect 20808 37132 20910 37133
tri 20808 37131 20809 37132 ne
rect 20809 37131 20910 37132
tri 20809 37130 20810 37131 ne
rect 20810 37130 20910 37131
tri 20810 37129 20811 37130 ne
rect 20811 37129 20910 37130
tri 20811 37128 20812 37129 ne
rect 20812 37128 20910 37129
tri 20812 37127 20813 37128 ne
rect 20813 37127 20910 37128
tri 20813 37126 20814 37127 ne
rect 20814 37126 20910 37127
tri 20814 37125 20815 37126 ne
rect 20815 37125 20910 37126
tri 20815 37124 20816 37125 ne
rect 20816 37124 20910 37125
tri 20816 37123 20817 37124 ne
rect 20817 37123 20910 37124
tri 20817 37122 20818 37123 ne
rect 20818 37122 20910 37123
rect 20956 37154 21040 37168
tri 21040 37154 21062 37176 sw
rect 20956 37122 21062 37154
tri 20818 37121 20819 37122 ne
rect 20819 37121 21062 37122
tri 20819 37120 20820 37121 ne
rect 20820 37120 21062 37121
tri 20820 37119 20821 37120 ne
rect 20821 37119 21062 37120
tri 20821 37118 20822 37119 ne
rect 20822 37118 21062 37119
tri 20822 37117 20823 37118 ne
rect 20823 37117 21062 37118
tri 20823 37116 20824 37117 ne
rect 20824 37116 21062 37117
tri 20824 37115 20825 37116 ne
rect 20825 37115 21062 37116
tri 20825 37114 20826 37115 ne
rect 20826 37114 21062 37115
tri 20826 37113 20827 37114 ne
rect 20827 37113 21062 37114
tri 20827 37112 20828 37113 ne
rect 20828 37112 21062 37113
tri 20828 37111 20829 37112 ne
rect 20829 37111 21062 37112
tri 20829 37110 20830 37111 ne
rect 20830 37110 21062 37111
tri 20830 37109 20831 37110 ne
rect 20831 37109 21062 37110
tri 21062 37109 21107 37154 sw
rect 70802 37148 71000 37206
tri 20831 37080 20860 37109 ne
rect 20860 37080 21107 37109
tri 20860 37035 20905 37080 ne
rect 20905 37064 21107 37080
tri 21107 37064 21152 37109 sw
rect 70802 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
rect 20905 37036 21152 37064
rect 20905 37035 21042 37036
tri 20905 36990 20950 37035 ne
rect 20950 36990 21042 37035
rect 21088 37019 21152 37036
tri 21152 37019 21197 37064 sw
rect 70802 37044 71000 37102
rect 21088 36990 21197 37019
tri 21197 36990 21226 37019 sw
rect 70802 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
tri 20950 36945 20995 36990 ne
rect 20995 36945 21226 36990
tri 21226 36945 21271 36990 sw
tri 20995 36900 21040 36945 ne
rect 21040 36904 21271 36945
rect 21040 36900 21174 36904
tri 21040 36889 21051 36900 ne
rect 21051 36889 21174 36900
tri 21051 36888 21052 36889 ne
rect 21052 36888 21174 36889
tri 21052 36887 21053 36888 ne
rect 21053 36887 21174 36888
tri 21053 36886 21054 36887 ne
rect 21054 36886 21174 36887
tri 21054 36885 21055 36886 ne
rect 21055 36885 21174 36886
tri 21055 36884 21056 36885 ne
rect 21056 36884 21174 36885
tri 21056 36883 21057 36884 ne
rect 21057 36883 21174 36884
tri 21057 36882 21058 36883 ne
rect 21058 36882 21174 36883
tri 21058 36881 21059 36882 ne
rect 21059 36881 21174 36882
tri 21059 36880 21060 36881 ne
rect 21060 36880 21174 36881
tri 21060 36879 21061 36880 ne
rect 21061 36879 21174 36880
tri 21061 36878 21062 36879 ne
rect 21062 36878 21174 36879
tri 21062 36877 21063 36878 ne
rect 21063 36877 21174 36878
tri 21063 36876 21064 36877 ne
rect 21064 36876 21174 36877
tri 21064 36875 21065 36876 ne
rect 21065 36875 21174 36876
tri 21065 36874 21066 36875 ne
rect 21066 36874 21174 36875
tri 21066 36873 21067 36874 ne
rect 21067 36873 21174 36874
tri 21067 36872 21068 36873 ne
rect 21068 36872 21174 36873
tri 21068 36871 21069 36872 ne
rect 21069 36871 21174 36872
tri 21069 36870 21070 36871 ne
rect 21070 36870 21174 36871
tri 21070 36869 21071 36870 ne
rect 21071 36869 21174 36870
tri 21071 36868 21072 36869 ne
rect 21072 36868 21174 36869
tri 21072 36867 21073 36868 ne
rect 21073 36867 21174 36868
tri 21073 36866 21074 36867 ne
rect 21074 36866 21174 36867
tri 21074 36865 21075 36866 ne
rect 21075 36865 21174 36866
tri 21075 36864 21076 36865 ne
rect 21076 36864 21174 36865
tri 21076 36863 21077 36864 ne
rect 21077 36863 21174 36864
tri 21077 36862 21078 36863 ne
rect 21078 36862 21174 36863
tri 21078 36861 21079 36862 ne
rect 21079 36861 21174 36862
tri 21079 36860 21080 36861 ne
rect 21080 36860 21174 36861
tri 21080 36859 21081 36860 ne
rect 21081 36859 21174 36860
tri 21081 36858 21082 36859 ne
rect 21082 36858 21174 36859
rect 21220 36900 21271 36904
tri 21271 36900 21316 36945 sw
rect 70802 36940 71000 36998
rect 21220 36858 21316 36900
tri 21082 36857 21083 36858 ne
rect 21083 36857 21316 36858
tri 21083 36856 21084 36857 ne
rect 21084 36856 21316 36857
tri 21084 36855 21085 36856 ne
rect 21085 36855 21316 36856
tri 21316 36855 21361 36900 sw
rect 70802 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
tri 21085 36854 21086 36855 ne
rect 21086 36854 21361 36855
tri 21086 36853 21087 36854 ne
rect 21087 36853 21361 36854
tri 21087 36852 21088 36853 ne
rect 21088 36852 21361 36853
tri 21088 36851 21089 36852 ne
rect 21089 36851 21361 36852
tri 21089 36850 21090 36851 ne
rect 21090 36850 21361 36851
tri 21090 36849 21091 36850 ne
rect 21091 36849 21361 36850
tri 21091 36848 21092 36849 ne
rect 21092 36848 21361 36849
tri 21092 36847 21093 36848 ne
rect 21093 36847 21361 36848
tri 21093 36846 21094 36847 ne
rect 21094 36846 21361 36847
tri 21094 36845 21095 36846 ne
rect 21095 36845 21361 36846
tri 21095 36844 21096 36845 ne
rect 21096 36844 21361 36845
tri 21096 36843 21097 36844 ne
rect 21097 36843 21361 36844
tri 21097 36842 21098 36843 ne
rect 21098 36842 21361 36843
tri 21098 36841 21099 36842 ne
rect 21099 36841 21361 36842
tri 21099 36840 21100 36841 ne
rect 21100 36840 21361 36841
tri 21100 36839 21101 36840 ne
rect 21101 36839 21361 36840
tri 21101 36838 21102 36839 ne
rect 21102 36838 21361 36839
tri 21102 36837 21103 36838 ne
rect 21103 36837 21361 36838
tri 21103 36836 21104 36837 ne
rect 21104 36836 21361 36837
tri 21104 36835 21105 36836 ne
rect 21105 36835 21361 36836
tri 21105 36834 21106 36835 ne
rect 21106 36834 21361 36835
tri 21106 36833 21107 36834 ne
rect 21107 36833 21361 36834
tri 21361 36833 21383 36855 sw
rect 70802 36836 71000 36894
tri 21107 36788 21152 36833 ne
rect 21152 36810 21383 36833
tri 21383 36810 21406 36833 sw
rect 21152 36788 21406 36810
tri 21152 36760 21180 36788 ne
rect 21180 36772 21406 36788
rect 21180 36760 21306 36772
tri 21180 36715 21225 36760 ne
rect 21225 36726 21306 36760
rect 21352 36765 21406 36772
tri 21406 36765 21451 36810 sw
rect 70802 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21352 36726 21451 36765
rect 21225 36720 21451 36726
tri 21451 36720 21496 36765 sw
rect 70802 36732 71000 36790
rect 21225 36715 21496 36720
tri 21225 36670 21270 36715 ne
rect 21270 36692 21496 36715
tri 21496 36692 21524 36720 sw
rect 21270 36670 21524 36692
tri 21270 36625 21315 36670 ne
rect 21315 36647 21524 36670
tri 21524 36647 21569 36692 sw
rect 70802 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21315 36640 21569 36647
rect 21315 36625 21438 36640
tri 21315 36615 21325 36625 ne
rect 21325 36615 21438 36625
tri 21325 36614 21326 36615 ne
rect 21326 36614 21438 36615
tri 21326 36613 21327 36614 ne
rect 21327 36613 21438 36614
tri 21327 36612 21328 36613 ne
rect 21328 36612 21438 36613
tri 21328 36611 21329 36612 ne
rect 21329 36611 21438 36612
tri 21329 36610 21330 36611 ne
rect 21330 36610 21438 36611
tri 21330 36609 21331 36610 ne
rect 21331 36609 21438 36610
tri 21331 36608 21332 36609 ne
rect 21332 36608 21438 36609
tri 21332 36607 21333 36608 ne
rect 21333 36607 21438 36608
tri 21333 36606 21334 36607 ne
rect 21334 36606 21438 36607
tri 21334 36605 21335 36606 ne
rect 21335 36605 21438 36606
tri 21335 36604 21336 36605 ne
rect 21336 36604 21438 36605
tri 21336 36603 21337 36604 ne
rect 21337 36603 21438 36604
tri 21337 36602 21338 36603 ne
rect 21338 36602 21438 36603
tri 21338 36601 21339 36602 ne
rect 21339 36601 21438 36602
tri 21339 36600 21340 36601 ne
rect 21340 36600 21438 36601
tri 21340 36599 21341 36600 ne
rect 21341 36599 21438 36600
tri 21341 36598 21342 36599 ne
rect 21342 36598 21438 36599
tri 21342 36597 21343 36598 ne
rect 21343 36597 21438 36598
tri 21343 36596 21344 36597 ne
rect 21344 36596 21438 36597
tri 21344 36595 21345 36596 ne
rect 21345 36595 21438 36596
tri 21345 36594 21346 36595 ne
rect 21346 36594 21438 36595
rect 21484 36602 21569 36640
tri 21569 36602 21614 36647 sw
rect 70802 36628 71000 36686
rect 21484 36594 21614 36602
tri 21346 36593 21347 36594 ne
rect 21347 36593 21614 36594
tri 21347 36592 21348 36593 ne
rect 21348 36592 21614 36593
tri 21348 36591 21349 36592 ne
rect 21349 36591 21614 36592
tri 21349 36590 21350 36591 ne
rect 21350 36590 21614 36591
tri 21350 36589 21351 36590 ne
rect 21351 36589 21614 36590
tri 21351 36588 21352 36589 ne
rect 21352 36588 21614 36589
tri 21352 36587 21353 36588 ne
rect 21353 36587 21614 36588
tri 21353 36586 21354 36587 ne
rect 21354 36586 21614 36587
tri 21354 36585 21355 36586 ne
rect 21355 36585 21614 36586
tri 21355 36584 21356 36585 ne
rect 21356 36584 21614 36585
tri 21356 36583 21357 36584 ne
rect 21357 36583 21614 36584
tri 21357 36582 21358 36583 ne
rect 21358 36582 21614 36583
tri 21358 36581 21359 36582 ne
rect 21359 36581 21614 36582
tri 21359 36580 21360 36581 ne
rect 21360 36580 21614 36581
tri 21360 36579 21361 36580 ne
rect 21361 36579 21614 36580
tri 21361 36578 21362 36579 ne
rect 21362 36578 21614 36579
tri 21362 36577 21363 36578 ne
rect 21363 36577 21614 36578
tri 21363 36576 21364 36577 ne
rect 21364 36576 21614 36577
tri 21364 36575 21365 36576 ne
rect 21365 36575 21614 36576
tri 21365 36574 21366 36575 ne
rect 21366 36574 21614 36575
tri 21366 36573 21367 36574 ne
rect 21367 36573 21614 36574
tri 21367 36572 21368 36573 ne
rect 21368 36572 21614 36573
tri 21368 36571 21369 36572 ne
rect 21369 36571 21614 36572
tri 21369 36570 21370 36571 ne
rect 21370 36570 21614 36571
tri 21370 36569 21371 36570 ne
rect 21371 36569 21614 36570
tri 21371 36568 21372 36569 ne
rect 21372 36568 21614 36569
tri 21372 36567 21373 36568 ne
rect 21373 36567 21614 36568
tri 21373 36566 21374 36567 ne
rect 21374 36566 21614 36567
tri 21374 36565 21375 36566 ne
rect 21375 36565 21614 36566
tri 21375 36564 21376 36565 ne
rect 21376 36564 21614 36565
tri 21376 36563 21377 36564 ne
rect 21377 36563 21614 36564
tri 21377 36562 21378 36563 ne
rect 21378 36562 21614 36563
tri 21378 36561 21379 36562 ne
rect 21379 36561 21614 36562
tri 21379 36560 21380 36561 ne
rect 21380 36560 21614 36561
tri 21380 36559 21381 36560 ne
rect 21381 36559 21614 36560
tri 21381 36558 21382 36559 ne
rect 21382 36558 21614 36559
tri 21382 36557 21383 36558 ne
rect 21383 36557 21614 36558
tri 21614 36557 21659 36602 sw
rect 70802 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21383 36534 21406 36557 ne
rect 21406 36534 21659 36557
tri 21659 36534 21682 36557 sw
tri 21406 36512 21428 36534 ne
rect 21428 36512 21682 36534
tri 21428 36489 21451 36512 ne
rect 21451 36508 21682 36512
rect 21451 36489 21570 36508
tri 21451 36444 21496 36489 ne
rect 21496 36462 21570 36489
rect 21616 36489 21682 36508
tri 21682 36489 21727 36534 sw
rect 70802 36524 71000 36582
rect 21616 36462 21727 36489
rect 21496 36444 21727 36462
tri 21727 36444 21772 36489 sw
rect 70802 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
tri 21496 36399 21541 36444 ne
rect 21541 36399 21772 36444
tri 21772 36399 21817 36444 sw
rect 70802 36420 71000 36478
tri 21541 36395 21545 36399 ne
rect 21545 36395 21817 36399
tri 21545 36350 21590 36395 ne
rect 21590 36376 21817 36395
rect 21590 36350 21702 36376
tri 21590 36341 21599 36350 ne
rect 21599 36341 21702 36350
tri 21599 36340 21600 36341 ne
rect 21600 36340 21702 36341
tri 21600 36339 21601 36340 ne
rect 21601 36339 21702 36340
tri 21601 36338 21602 36339 ne
rect 21602 36338 21702 36339
tri 21602 36337 21603 36338 ne
rect 21603 36337 21702 36338
tri 21603 36336 21604 36337 ne
rect 21604 36336 21702 36337
tri 21604 36335 21605 36336 ne
rect 21605 36335 21702 36336
tri 21605 36334 21606 36335 ne
rect 21606 36334 21702 36335
tri 21606 36333 21607 36334 ne
rect 21607 36333 21702 36334
tri 21607 36332 21608 36333 ne
rect 21608 36332 21702 36333
tri 21608 36331 21609 36332 ne
rect 21609 36331 21702 36332
tri 21609 36330 21610 36331 ne
rect 21610 36330 21702 36331
rect 21748 36371 21817 36376
tri 21817 36371 21845 36399 sw
rect 70802 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36330 21845 36371
tri 21610 36329 21611 36330 ne
rect 21611 36329 21845 36330
tri 21611 36328 21612 36329 ne
rect 21612 36328 21845 36329
tri 21612 36327 21613 36328 ne
rect 21613 36327 21845 36328
tri 21613 36326 21614 36327 ne
rect 21614 36326 21845 36327
tri 21845 36326 21890 36371 sw
tri 21614 36325 21615 36326 ne
rect 21615 36325 21890 36326
tri 21615 36324 21616 36325 ne
rect 21616 36324 21890 36325
tri 21616 36323 21617 36324 ne
rect 21617 36323 21890 36324
tri 21617 36322 21618 36323 ne
rect 21618 36322 21890 36323
tri 21618 36321 21619 36322 ne
rect 21619 36321 21890 36322
tri 21619 36320 21620 36321 ne
rect 21620 36320 21890 36321
tri 21620 36319 21621 36320 ne
rect 21621 36319 21890 36320
tri 21621 36318 21622 36319 ne
rect 21622 36318 21890 36319
tri 21622 36317 21623 36318 ne
rect 21623 36317 21890 36318
tri 21623 36316 21624 36317 ne
rect 21624 36316 21890 36317
tri 21624 36315 21625 36316 ne
rect 21625 36315 21890 36316
tri 21625 36314 21626 36315 ne
rect 21626 36314 21890 36315
tri 21626 36313 21627 36314 ne
rect 21627 36313 21890 36314
tri 21627 36312 21628 36313 ne
rect 21628 36312 21890 36313
tri 21628 36311 21629 36312 ne
rect 21629 36311 21890 36312
tri 21629 36310 21630 36311 ne
rect 21630 36310 21890 36311
tri 21630 36309 21631 36310 ne
rect 21631 36309 21890 36310
tri 21631 36308 21632 36309 ne
rect 21632 36308 21890 36309
tri 21632 36307 21633 36308 ne
rect 21633 36307 21890 36308
tri 21633 36306 21634 36307 ne
rect 21634 36306 21890 36307
tri 21634 36305 21635 36306 ne
rect 21635 36305 21890 36306
tri 21635 36304 21636 36305 ne
rect 21636 36304 21890 36305
tri 21636 36303 21637 36304 ne
rect 21637 36303 21890 36304
tri 21637 36302 21638 36303 ne
rect 21638 36302 21890 36303
tri 21638 36301 21639 36302 ne
rect 21639 36301 21890 36302
tri 21639 36300 21640 36301 ne
rect 21640 36300 21890 36301
tri 21640 36299 21641 36300 ne
rect 21641 36299 21890 36300
tri 21641 36298 21642 36299 ne
rect 21642 36298 21890 36299
tri 21642 36297 21643 36298 ne
rect 21643 36297 21890 36298
tri 21643 36296 21644 36297 ne
rect 21644 36296 21890 36297
tri 21644 36295 21645 36296 ne
rect 21645 36295 21890 36296
tri 21645 36294 21646 36295 ne
rect 21646 36294 21890 36295
tri 21646 36293 21647 36294 ne
rect 21647 36293 21890 36294
tri 21647 36292 21648 36293 ne
rect 21648 36292 21890 36293
tri 21648 36291 21649 36292 ne
rect 21649 36291 21890 36292
tri 21649 36290 21650 36291 ne
rect 21650 36290 21890 36291
tri 21650 36289 21651 36290 ne
rect 21651 36289 21890 36290
tri 21651 36288 21652 36289 ne
rect 21652 36288 21890 36289
tri 21652 36287 21653 36288 ne
rect 21653 36287 21890 36288
tri 21653 36286 21654 36287 ne
rect 21654 36286 21890 36287
tri 21654 36285 21655 36286 ne
rect 21655 36285 21890 36286
tri 21655 36284 21656 36285 ne
rect 21656 36284 21890 36285
tri 21656 36283 21657 36284 ne
rect 21657 36283 21890 36284
tri 21657 36282 21658 36283 ne
rect 21658 36282 21890 36283
tri 21658 36281 21659 36282 ne
rect 21659 36281 21890 36282
tri 21890 36281 21935 36326 sw
rect 70802 36316 71000 36374
tri 21659 36236 21704 36281 ne
rect 21704 36244 21935 36281
rect 21704 36236 21834 36244
tri 21704 36191 21749 36236 ne
rect 21749 36198 21834 36236
rect 21880 36236 21935 36244
tri 21935 36236 21980 36281 sw
rect 70802 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
rect 21880 36213 21980 36236
tri 21980 36213 22003 36236 sw
rect 21880 36198 22003 36213
rect 21749 36191 22003 36198
tri 21749 36168 21772 36191 ne
rect 21772 36168 22003 36191
tri 22003 36168 22048 36213 sw
rect 70802 36212 71000 36270
tri 21772 36146 21794 36168 ne
rect 21794 36146 22048 36168
tri 21794 36123 21817 36146 ne
rect 21817 36123 22048 36146
tri 22048 36123 22093 36168 sw
rect 70802 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21817 36078 21862 36123 ne
rect 21862 36112 22093 36123
rect 21862 36078 21966 36112
tri 21862 36066 21874 36078 ne
rect 21874 36066 21966 36078
rect 22012 36078 22093 36112
tri 22093 36078 22138 36123 sw
rect 70802 36108 71000 36166
rect 22012 36066 22138 36078
tri 21874 36065 21875 36066 ne
rect 21875 36065 22138 36066
tri 21875 36064 21876 36065 ne
rect 21876 36064 22138 36065
tri 21876 36063 21877 36064 ne
rect 21877 36063 22138 36064
tri 21877 36062 21878 36063 ne
rect 21878 36062 22138 36063
tri 21878 36061 21879 36062 ne
rect 21879 36061 22138 36062
tri 21879 36060 21880 36061 ne
rect 21880 36060 22138 36061
tri 21880 36059 21881 36060 ne
rect 21881 36059 22138 36060
tri 21881 36058 21882 36059 ne
rect 21882 36058 22138 36059
tri 21882 36057 21883 36058 ne
rect 21883 36057 22138 36058
tri 21883 36056 21884 36057 ne
rect 21884 36056 22138 36057
tri 21884 36055 21885 36056 ne
rect 21885 36055 22138 36056
tri 21885 36054 21886 36055 ne
rect 21886 36054 22138 36055
tri 21886 36053 21887 36054 ne
rect 21887 36053 22138 36054
tri 21887 36052 21888 36053 ne
rect 21888 36052 22138 36053
tri 21888 36051 21889 36052 ne
rect 21889 36051 22138 36052
tri 21889 36050 21890 36051 ne
rect 21890 36050 22138 36051
tri 22138 36050 22166 36078 sw
rect 70802 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
tri 21890 36049 21891 36050 ne
rect 21891 36049 22166 36050
tri 21891 36048 21892 36049 ne
rect 21892 36048 22166 36049
tri 21892 36047 21893 36048 ne
rect 21893 36047 22166 36048
tri 21893 36046 21894 36047 ne
rect 21894 36046 22166 36047
tri 21894 36045 21895 36046 ne
rect 21895 36045 22166 36046
tri 21895 36044 21896 36045 ne
rect 21896 36044 22166 36045
tri 21896 36043 21897 36044 ne
rect 21897 36043 22166 36044
tri 21897 36042 21898 36043 ne
rect 21898 36042 22166 36043
tri 21898 36041 21899 36042 ne
rect 21899 36041 22166 36042
tri 21899 36040 21900 36041 ne
rect 21900 36040 22166 36041
tri 21900 36039 21901 36040 ne
rect 21901 36039 22166 36040
tri 21901 36038 21902 36039 ne
rect 21902 36038 22166 36039
tri 21902 36037 21903 36038 ne
rect 21903 36037 22166 36038
tri 21903 36036 21904 36037 ne
rect 21904 36036 22166 36037
tri 21904 36035 21905 36036 ne
rect 21905 36035 22166 36036
tri 21905 36034 21906 36035 ne
rect 21906 36034 22166 36035
tri 21906 36033 21907 36034 ne
rect 21907 36033 22166 36034
tri 21907 36032 21908 36033 ne
rect 21908 36032 22166 36033
tri 21908 36031 21909 36032 ne
rect 21909 36031 22166 36032
tri 21909 36030 21910 36031 ne
rect 21910 36030 22166 36031
tri 21910 36029 21911 36030 ne
rect 21911 36029 22166 36030
tri 21911 36028 21912 36029 ne
rect 21912 36028 22166 36029
tri 21912 36027 21913 36028 ne
rect 21913 36027 22166 36028
tri 21913 36026 21914 36027 ne
rect 21914 36026 22166 36027
tri 21914 36025 21915 36026 ne
rect 21915 36025 22166 36026
tri 21915 36024 21916 36025 ne
rect 21916 36024 22166 36025
tri 21916 36023 21917 36024 ne
rect 21917 36023 22166 36024
tri 21917 36022 21918 36023 ne
rect 21918 36022 22166 36023
tri 21918 36021 21919 36022 ne
rect 21919 36021 22166 36022
tri 21919 36020 21920 36021 ne
rect 21920 36020 22166 36021
tri 21920 36019 21921 36020 ne
rect 21921 36019 22166 36020
tri 21921 36018 21922 36019 ne
rect 21922 36018 22166 36019
tri 21922 36017 21923 36018 ne
rect 21923 36017 22166 36018
tri 21923 36016 21924 36017 ne
rect 21924 36016 22166 36017
tri 21924 36015 21925 36016 ne
rect 21925 36015 22166 36016
tri 21925 36014 21926 36015 ne
rect 21926 36014 22166 36015
tri 21926 36013 21927 36014 ne
rect 21927 36013 22166 36014
tri 21927 36012 21928 36013 ne
rect 21928 36012 22166 36013
tri 21928 36011 21929 36012 ne
rect 21929 36011 22166 36012
tri 21929 36010 21930 36011 ne
rect 21930 36010 22166 36011
tri 21930 36009 21931 36010 ne
rect 21931 36009 22166 36010
tri 21931 36008 21932 36009 ne
rect 21932 36008 22166 36009
tri 21932 36007 21933 36008 ne
rect 21933 36007 22166 36008
tri 21933 36006 21934 36007 ne
rect 21934 36006 22166 36007
tri 21934 36005 21935 36006 ne
rect 21935 36005 22166 36006
tri 22166 36005 22211 36050 sw
tri 21935 35986 21954 36005 ne
rect 21954 35986 22211 36005
tri 21954 35941 21999 35986 ne
rect 21999 35980 22211 35986
rect 21999 35941 22098 35980
tri 21999 35896 22044 35941 ne
rect 22044 35934 22098 35941
rect 22144 35960 22211 35980
tri 22211 35960 22256 36005 sw
rect 70802 36004 71000 36062
rect 22144 35934 22256 35960
rect 22044 35915 22256 35934
tri 22256 35915 22301 35960 sw
rect 70802 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22044 35896 22301 35915
tri 22044 35851 22089 35896 ne
rect 22089 35892 22301 35896
tri 22301 35892 22324 35915 sw
rect 70802 35900 71000 35958
rect 22089 35851 22324 35892
tri 22089 35806 22134 35851 ne
rect 22134 35848 22324 35851
rect 22134 35806 22230 35848
tri 22134 35802 22138 35806 ne
rect 22138 35802 22230 35806
rect 22276 35847 22324 35848
tri 22324 35847 22369 35892 sw
rect 70802 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 22276 35802 22369 35847
tri 22369 35802 22414 35847 sw
tri 22138 35792 22148 35802 ne
rect 22148 35792 22414 35802
tri 22148 35791 22149 35792 ne
rect 22149 35791 22414 35792
tri 22149 35790 22150 35791 ne
rect 22150 35790 22414 35791
tri 22150 35789 22151 35790 ne
rect 22151 35789 22414 35790
tri 22151 35788 22152 35789 ne
rect 22152 35788 22414 35789
tri 22152 35787 22153 35788 ne
rect 22153 35787 22414 35788
tri 22153 35786 22154 35787 ne
rect 22154 35786 22414 35787
tri 22154 35785 22155 35786 ne
rect 22155 35785 22414 35786
tri 22155 35784 22156 35785 ne
rect 22156 35784 22414 35785
tri 22156 35783 22157 35784 ne
rect 22157 35783 22414 35784
tri 22157 35782 22158 35783 ne
rect 22158 35782 22414 35783
tri 22158 35781 22159 35782 ne
rect 22159 35781 22414 35782
tri 22159 35780 22160 35781 ne
rect 22160 35780 22414 35781
tri 22160 35779 22161 35780 ne
rect 22161 35779 22414 35780
tri 22161 35778 22162 35779 ne
rect 22162 35778 22414 35779
tri 22162 35777 22163 35778 ne
rect 22163 35777 22414 35778
tri 22163 35776 22164 35777 ne
rect 22164 35776 22414 35777
tri 22164 35775 22165 35776 ne
rect 22165 35775 22414 35776
tri 22165 35774 22166 35775 ne
rect 22166 35774 22414 35775
tri 22166 35773 22167 35774 ne
rect 22167 35773 22414 35774
tri 22167 35772 22168 35773 ne
rect 22168 35772 22414 35773
tri 22168 35771 22169 35772 ne
rect 22169 35771 22414 35772
tri 22169 35770 22170 35771 ne
rect 22170 35770 22414 35771
tri 22170 35769 22171 35770 ne
rect 22171 35769 22414 35770
tri 22171 35768 22172 35769 ne
rect 22172 35768 22414 35769
tri 22172 35767 22173 35768 ne
rect 22173 35767 22414 35768
tri 22173 35766 22174 35767 ne
rect 22174 35766 22414 35767
tri 22174 35765 22175 35766 ne
rect 22175 35765 22414 35766
tri 22175 35764 22176 35765 ne
rect 22176 35764 22414 35765
tri 22176 35763 22177 35764 ne
rect 22177 35763 22414 35764
tri 22177 35762 22178 35763 ne
rect 22178 35762 22414 35763
tri 22178 35761 22179 35762 ne
rect 22179 35761 22414 35762
tri 22179 35760 22180 35761 ne
rect 22180 35760 22414 35761
tri 22180 35759 22181 35760 ne
rect 22181 35759 22414 35760
tri 22181 35758 22182 35759 ne
rect 22182 35758 22414 35759
tri 22182 35757 22183 35758 ne
rect 22183 35757 22414 35758
tri 22414 35757 22459 35802 sw
rect 70802 35796 71000 35854
tri 22183 35756 22184 35757 ne
rect 22184 35756 22459 35757
tri 22184 35755 22185 35756 ne
rect 22185 35755 22459 35756
tri 22185 35754 22186 35755 ne
rect 22186 35754 22459 35755
tri 22186 35753 22187 35754 ne
rect 22187 35753 22459 35754
tri 22187 35752 22188 35753 ne
rect 22188 35752 22459 35753
tri 22188 35751 22189 35752 ne
rect 22189 35751 22459 35752
tri 22189 35750 22190 35751 ne
rect 22190 35750 22459 35751
tri 22190 35749 22191 35750 ne
rect 22191 35749 22459 35750
tri 22191 35748 22192 35749 ne
rect 22192 35748 22459 35749
tri 22192 35747 22193 35748 ne
rect 22193 35747 22459 35748
tri 22193 35746 22194 35747 ne
rect 22194 35746 22459 35747
tri 22194 35745 22195 35746 ne
rect 22195 35745 22459 35746
tri 22195 35744 22196 35745 ne
rect 22196 35744 22459 35745
tri 22196 35743 22197 35744 ne
rect 22197 35743 22459 35744
tri 22197 35742 22198 35743 ne
rect 22198 35742 22459 35743
tri 22198 35741 22199 35742 ne
rect 22199 35741 22459 35742
tri 22199 35740 22200 35741 ne
rect 22200 35740 22459 35741
tri 22200 35739 22201 35740 ne
rect 22201 35739 22459 35740
tri 22201 35738 22202 35739 ne
rect 22202 35738 22459 35739
tri 22202 35737 22203 35738 ne
rect 22203 35737 22459 35738
tri 22203 35736 22204 35737 ne
rect 22204 35736 22459 35737
tri 22204 35735 22205 35736 ne
rect 22205 35735 22459 35736
tri 22205 35734 22206 35735 ne
rect 22206 35734 22459 35735
tri 22206 35733 22207 35734 ne
rect 22207 35733 22459 35734
tri 22207 35732 22208 35733 ne
rect 22208 35732 22459 35733
tri 22208 35731 22209 35732 ne
rect 22209 35731 22459 35732
tri 22209 35730 22210 35731 ne
rect 22210 35730 22459 35731
tri 22210 35729 22211 35730 ne
rect 22211 35729 22459 35730
tri 22459 35729 22487 35757 sw
rect 70802 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22211 35684 22256 35729 ne
rect 22256 35716 22487 35729
rect 22256 35684 22362 35716
tri 22256 35666 22274 35684 ne
rect 22274 35670 22362 35684
rect 22408 35712 22487 35716
tri 22487 35712 22504 35729 sw
rect 22408 35670 22504 35712
rect 22274 35667 22504 35670
tri 22504 35667 22549 35712 sw
rect 70802 35692 71000 35750
rect 22274 35666 22549 35667
tri 22274 35621 22319 35666 ne
rect 22319 35622 22549 35666
tri 22549 35622 22594 35667 sw
rect 70802 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 22319 35621 22594 35622
tri 22319 35576 22364 35621 ne
rect 22364 35588 22594 35621
tri 22594 35588 22628 35622 sw
rect 70802 35588 71000 35646
rect 22364 35584 22628 35588
rect 22364 35576 22494 35584
tri 22364 35531 22409 35576 ne
rect 22409 35538 22494 35576
rect 22540 35543 22628 35584
tri 22628 35543 22673 35588 sw
rect 22540 35538 22673 35543
rect 22409 35531 22673 35538
tri 22409 35517 22423 35531 ne
rect 22423 35517 22673 35531
tri 22423 35516 22424 35517 ne
rect 22424 35516 22673 35517
tri 22424 35515 22425 35516 ne
rect 22425 35515 22673 35516
tri 22425 35514 22426 35515 ne
rect 22426 35514 22673 35515
tri 22426 35513 22427 35514 ne
rect 22427 35513 22673 35514
tri 22427 35512 22428 35513 ne
rect 22428 35512 22673 35513
tri 22428 35511 22429 35512 ne
rect 22429 35511 22673 35512
tri 22429 35510 22430 35511 ne
rect 22430 35510 22673 35511
tri 22430 35509 22431 35510 ne
rect 22431 35509 22673 35510
tri 22431 35508 22432 35509 ne
rect 22432 35508 22673 35509
tri 22432 35507 22433 35508 ne
rect 22433 35507 22673 35508
tri 22433 35506 22434 35507 ne
rect 22434 35506 22673 35507
tri 22434 35505 22435 35506 ne
rect 22435 35505 22673 35506
tri 22435 35504 22436 35505 ne
rect 22436 35504 22673 35505
tri 22436 35503 22437 35504 ne
rect 22437 35503 22673 35504
tri 22437 35502 22438 35503 ne
rect 22438 35502 22673 35503
tri 22438 35501 22439 35502 ne
rect 22439 35501 22673 35502
tri 22439 35500 22440 35501 ne
rect 22440 35500 22673 35501
tri 22440 35499 22441 35500 ne
rect 22441 35499 22673 35500
tri 22441 35498 22442 35499 ne
rect 22442 35498 22673 35499
tri 22673 35498 22718 35543 sw
rect 70802 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
tri 22442 35497 22443 35498 ne
rect 22443 35497 22718 35498
tri 22443 35496 22444 35497 ne
rect 22444 35496 22718 35497
tri 22444 35495 22445 35496 ne
rect 22445 35495 22718 35496
tri 22445 35494 22446 35495 ne
rect 22446 35494 22718 35495
tri 22446 35493 22447 35494 ne
rect 22447 35493 22718 35494
tri 22447 35492 22448 35493 ne
rect 22448 35492 22718 35493
tri 22448 35491 22449 35492 ne
rect 22449 35491 22718 35492
tri 22449 35490 22450 35491 ne
rect 22450 35490 22718 35491
tri 22450 35489 22451 35490 ne
rect 22451 35489 22718 35490
tri 22451 35488 22452 35489 ne
rect 22452 35488 22718 35489
tri 22452 35487 22453 35488 ne
rect 22453 35487 22718 35488
tri 22453 35486 22454 35487 ne
rect 22454 35486 22718 35487
tri 22454 35485 22455 35486 ne
rect 22455 35485 22718 35486
tri 22455 35484 22456 35485 ne
rect 22456 35484 22718 35485
tri 22456 35483 22457 35484 ne
rect 22457 35483 22718 35484
tri 22457 35482 22458 35483 ne
rect 22458 35482 22718 35483
tri 22458 35481 22459 35482 ne
rect 22459 35481 22718 35482
tri 22459 35480 22460 35481 ne
rect 22460 35480 22718 35481
tri 22460 35479 22461 35480 ne
rect 22461 35479 22718 35480
tri 22461 35478 22462 35479 ne
rect 22462 35478 22718 35479
tri 22462 35477 22463 35478 ne
rect 22463 35477 22718 35478
tri 22463 35476 22464 35477 ne
rect 22464 35476 22718 35477
tri 22464 35475 22465 35476 ne
rect 22465 35475 22718 35476
tri 22465 35474 22466 35475 ne
rect 22466 35474 22718 35475
tri 22466 35473 22467 35474 ne
rect 22467 35473 22718 35474
tri 22467 35472 22468 35473 ne
rect 22468 35472 22718 35473
tri 22468 35471 22469 35472 ne
rect 22469 35471 22718 35472
tri 22469 35470 22470 35471 ne
rect 22470 35470 22718 35471
tri 22470 35469 22471 35470 ne
rect 22471 35469 22718 35470
tri 22471 35468 22472 35469 ne
rect 22472 35468 22718 35469
tri 22472 35467 22473 35468 ne
rect 22473 35467 22718 35468
tri 22473 35466 22474 35467 ne
rect 22474 35466 22718 35467
tri 22474 35465 22475 35466 ne
rect 22475 35465 22718 35466
tri 22475 35464 22476 35465 ne
rect 22476 35464 22718 35465
tri 22476 35463 22477 35464 ne
rect 22477 35463 22718 35464
tri 22477 35462 22478 35463 ne
rect 22478 35462 22718 35463
tri 22478 35461 22479 35462 ne
rect 22479 35461 22718 35462
tri 22479 35460 22480 35461 ne
rect 22480 35460 22718 35461
tri 22480 35459 22481 35460 ne
rect 22481 35459 22718 35460
tri 22481 35458 22482 35459 ne
rect 22482 35458 22718 35459
tri 22482 35457 22483 35458 ne
rect 22483 35457 22718 35458
tri 22483 35456 22484 35457 ne
rect 22484 35456 22718 35457
tri 22484 35455 22485 35456 ne
rect 22485 35455 22718 35456
tri 22485 35454 22486 35455 ne
rect 22486 35454 22718 35455
tri 22486 35453 22487 35454 ne
rect 22487 35453 22718 35454
tri 22718 35453 22763 35498 sw
rect 70802 35484 71000 35542
tri 22487 35436 22504 35453 ne
rect 22504 35452 22763 35453
rect 22504 35436 22626 35452
tri 22504 35408 22532 35436 ne
rect 22532 35408 22626 35436
tri 22532 35391 22549 35408 ne
rect 22549 35406 22626 35408
rect 22672 35436 22763 35452
tri 22763 35436 22780 35453 sw
rect 70802 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35406 22780 35436
rect 22549 35391 22780 35406
tri 22780 35391 22825 35436 sw
tri 22549 35346 22594 35391 ne
rect 22594 35346 22825 35391
tri 22825 35346 22870 35391 sw
rect 70802 35380 71000 35438
tri 22594 35301 22639 35346 ne
rect 22639 35320 22870 35346
rect 22639 35301 22758 35320
tri 22639 35256 22684 35301 ne
rect 22684 35274 22758 35301
rect 22804 35301 22870 35320
tri 22870 35301 22915 35346 sw
rect 70802 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22804 35274 22915 35301
rect 22684 35267 22915 35274
tri 22915 35267 22949 35301 sw
rect 70802 35276 71000 35334
rect 22684 35256 22949 35267
tri 22684 35243 22697 35256 ne
rect 22697 35243 22949 35256
tri 22697 35242 22698 35243 ne
rect 22698 35242 22949 35243
tri 22698 35241 22699 35242 ne
rect 22699 35241 22949 35242
tri 22699 35240 22700 35241 ne
rect 22700 35240 22949 35241
tri 22700 35239 22701 35240 ne
rect 22701 35239 22949 35240
tri 22701 35238 22702 35239 ne
rect 22702 35238 22949 35239
tri 22702 35237 22703 35238 ne
rect 22703 35237 22949 35238
tri 22703 35236 22704 35237 ne
rect 22704 35236 22949 35237
tri 22704 35235 22705 35236 ne
rect 22705 35235 22949 35236
tri 22705 35234 22706 35235 ne
rect 22706 35234 22949 35235
tri 22706 35233 22707 35234 ne
rect 22707 35233 22949 35234
tri 22707 35232 22708 35233 ne
rect 22708 35232 22949 35233
tri 22708 35231 22709 35232 ne
rect 22709 35231 22949 35232
tri 22709 35230 22710 35231 ne
rect 22710 35230 22949 35231
tri 22710 35229 22711 35230 ne
rect 22711 35229 22949 35230
tri 22711 35228 22712 35229 ne
rect 22712 35228 22949 35229
tri 22712 35227 22713 35228 ne
rect 22713 35227 22949 35228
tri 22713 35226 22714 35227 ne
rect 22714 35226 22949 35227
tri 22714 35225 22715 35226 ne
rect 22715 35225 22949 35226
tri 22715 35224 22716 35225 ne
rect 22716 35224 22949 35225
tri 22716 35223 22717 35224 ne
rect 22717 35223 22949 35224
tri 22717 35222 22718 35223 ne
rect 22718 35222 22949 35223
tri 22949 35222 22994 35267 sw
rect 70802 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22718 35221 22719 35222 ne
rect 22719 35221 22994 35222
tri 22719 35220 22720 35221 ne
rect 22720 35220 22994 35221
tri 22720 35219 22721 35220 ne
rect 22721 35219 22994 35220
tri 22721 35218 22722 35219 ne
rect 22722 35218 22994 35219
tri 22722 35217 22723 35218 ne
rect 22723 35217 22994 35218
tri 22723 35216 22724 35217 ne
rect 22724 35216 22994 35217
tri 22724 35215 22725 35216 ne
rect 22725 35215 22994 35216
tri 22725 35214 22726 35215 ne
rect 22726 35214 22994 35215
tri 22726 35213 22727 35214 ne
rect 22727 35213 22994 35214
tri 22727 35212 22728 35213 ne
rect 22728 35212 22994 35213
tri 22728 35211 22729 35212 ne
rect 22729 35211 22994 35212
tri 22729 35210 22730 35211 ne
rect 22730 35210 22994 35211
tri 22730 35209 22731 35210 ne
rect 22731 35209 22994 35210
tri 22731 35208 22732 35209 ne
rect 22732 35208 22994 35209
tri 22732 35207 22733 35208 ne
rect 22733 35207 22994 35208
tri 22733 35206 22734 35207 ne
rect 22734 35206 22994 35207
tri 22734 35205 22735 35206 ne
rect 22735 35205 22994 35206
tri 22735 35204 22736 35205 ne
rect 22736 35204 22994 35205
tri 22736 35203 22737 35204 ne
rect 22737 35203 22994 35204
tri 22737 35202 22738 35203 ne
rect 22738 35202 22994 35203
tri 22738 35201 22739 35202 ne
rect 22739 35201 22994 35202
tri 22739 35200 22740 35201 ne
rect 22740 35200 22994 35201
tri 22740 35199 22741 35200 ne
rect 22741 35199 22994 35200
tri 22741 35198 22742 35199 ne
rect 22742 35198 22994 35199
tri 22742 35197 22743 35198 ne
rect 22743 35197 22994 35198
tri 22743 35196 22744 35197 ne
rect 22744 35196 22994 35197
tri 22744 35195 22745 35196 ne
rect 22745 35195 22994 35196
tri 22745 35194 22746 35195 ne
rect 22746 35194 22994 35195
tri 22746 35193 22747 35194 ne
rect 22747 35193 22994 35194
tri 22747 35192 22748 35193 ne
rect 22748 35192 22994 35193
tri 22748 35191 22749 35192 ne
rect 22749 35191 22994 35192
tri 22749 35190 22750 35191 ne
rect 22750 35190 22994 35191
tri 22750 35189 22751 35190 ne
rect 22751 35189 22994 35190
tri 22751 35188 22752 35189 ne
rect 22752 35188 22994 35189
tri 22752 35187 22753 35188 ne
rect 22753 35187 22890 35188
tri 22753 35186 22754 35187 ne
rect 22754 35186 22890 35187
tri 22754 35185 22755 35186 ne
rect 22755 35185 22890 35186
tri 22755 35184 22756 35185 ne
rect 22756 35184 22890 35185
tri 22756 35183 22757 35184 ne
rect 22757 35183 22890 35184
tri 22757 35182 22758 35183 ne
rect 22758 35182 22890 35183
tri 22758 35181 22759 35182 ne
rect 22759 35181 22890 35182
tri 22759 35180 22760 35181 ne
rect 22760 35180 22890 35181
tri 22760 35179 22761 35180 ne
rect 22761 35179 22890 35180
tri 22761 35178 22762 35179 ne
rect 22762 35178 22890 35179
tri 22762 35177 22763 35178 ne
rect 22763 35177 22890 35178
tri 22763 35132 22808 35177 ne
rect 22808 35142 22890 35177
rect 22936 35177 22994 35188
tri 22994 35177 23039 35222 sw
rect 22936 35142 23039 35177
rect 22808 35132 23039 35142
tri 23039 35132 23084 35177 sw
rect 70802 35172 71000 35230
tri 22808 35087 22853 35132 ne
rect 22853 35115 23084 35132
tri 23084 35115 23101 35132 sw
rect 70802 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
rect 22853 35087 23101 35115
tri 22853 35070 22870 35087 ne
rect 22870 35070 23101 35087
tri 23101 35070 23146 35115 sw
tri 22870 35042 22898 35070 ne
rect 22898 35056 23146 35070
rect 22898 35042 23022 35056
tri 22898 35025 22915 35042 ne
rect 22915 35025 23022 35042
tri 22915 34980 22960 35025 ne
rect 22960 35010 23022 35025
rect 23068 35025 23146 35056
tri 23146 35025 23191 35070 sw
rect 70802 35068 71000 35126
rect 23068 35010 23191 35025
rect 22960 34980 23191 35010
tri 23191 34980 23236 35025 sw
rect 70802 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
tri 22960 34969 22971 34980 ne
rect 22971 34969 23236 34980
tri 22971 34968 22972 34969 ne
rect 22972 34968 23236 34969
tri 22972 34967 22973 34968 ne
rect 22973 34967 23236 34968
tri 22973 34966 22974 34967 ne
rect 22974 34966 23236 34967
tri 22974 34965 22975 34966 ne
rect 22975 34965 23236 34966
tri 22975 34964 22976 34965 ne
rect 22976 34964 23236 34965
tri 22976 34963 22977 34964 ne
rect 22977 34963 23236 34964
tri 22977 34962 22978 34963 ne
rect 22978 34962 23236 34963
tri 22978 34961 22979 34962 ne
rect 22979 34961 23236 34962
tri 22979 34960 22980 34961 ne
rect 22980 34960 23236 34961
tri 22980 34959 22981 34960 ne
rect 22981 34959 23236 34960
tri 22981 34958 22982 34959 ne
rect 22982 34958 23236 34959
tri 22982 34957 22983 34958 ne
rect 22983 34957 23236 34958
tri 22983 34956 22984 34957 ne
rect 22984 34956 23236 34957
tri 22984 34955 22985 34956 ne
rect 22985 34955 23236 34956
tri 22985 34954 22986 34955 ne
rect 22986 34954 23236 34955
tri 22986 34953 22987 34954 ne
rect 22987 34953 23236 34954
tri 22987 34952 22988 34953 ne
rect 22988 34952 23236 34953
tri 22988 34951 22989 34952 ne
rect 22989 34951 23236 34952
tri 22989 34950 22990 34951 ne
rect 22990 34950 23236 34951
tri 22990 34949 22991 34950 ne
rect 22991 34949 23236 34950
tri 22991 34948 22992 34949 ne
rect 22992 34948 23236 34949
tri 22992 34947 22993 34948 ne
rect 22993 34947 23236 34948
tri 22993 34946 22994 34947 ne
rect 22994 34946 23236 34947
tri 23236 34946 23270 34980 sw
rect 70802 34964 71000 35022
tri 22994 34945 22995 34946 ne
rect 22995 34945 23270 34946
tri 22995 34944 22996 34945 ne
rect 22996 34944 23270 34945
tri 22996 34943 22997 34944 ne
rect 22997 34943 23270 34944
tri 22997 34942 22998 34943 ne
rect 22998 34942 23270 34943
tri 22998 34941 22999 34942 ne
rect 22999 34941 23270 34942
tri 22999 34940 23000 34941 ne
rect 23000 34940 23270 34941
tri 23000 34939 23001 34940 ne
rect 23001 34939 23270 34940
tri 23001 34938 23002 34939 ne
rect 23002 34938 23270 34939
tri 23002 34937 23003 34938 ne
rect 23003 34937 23270 34938
tri 23003 34936 23004 34937 ne
rect 23004 34936 23270 34937
tri 23004 34935 23005 34936 ne
rect 23005 34935 23270 34936
tri 23005 34934 23006 34935 ne
rect 23006 34934 23270 34935
tri 23006 34933 23007 34934 ne
rect 23007 34933 23270 34934
tri 23007 34932 23008 34933 ne
rect 23008 34932 23270 34933
tri 23008 34931 23009 34932 ne
rect 23009 34931 23270 34932
tri 23009 34930 23010 34931 ne
rect 23010 34930 23270 34931
tri 23010 34929 23011 34930 ne
rect 23011 34929 23270 34930
tri 23011 34928 23012 34929 ne
rect 23012 34928 23270 34929
tri 23012 34927 23013 34928 ne
rect 23013 34927 23270 34928
tri 23013 34926 23014 34927 ne
rect 23014 34926 23270 34927
tri 23014 34925 23015 34926 ne
rect 23015 34925 23270 34926
tri 23015 34924 23016 34925 ne
rect 23016 34924 23270 34925
tri 23016 34923 23017 34924 ne
rect 23017 34923 23154 34924
tri 23017 34922 23018 34923 ne
rect 23018 34922 23154 34923
tri 23018 34921 23019 34922 ne
rect 23019 34921 23154 34922
tri 23019 34920 23020 34921 ne
rect 23020 34920 23154 34921
tri 23020 34919 23021 34920 ne
rect 23021 34919 23154 34920
tri 23021 34918 23022 34919 ne
rect 23022 34918 23154 34919
tri 23022 34917 23023 34918 ne
rect 23023 34917 23154 34918
tri 23023 34916 23024 34917 ne
rect 23024 34916 23154 34917
tri 23024 34915 23025 34916 ne
rect 23025 34915 23154 34916
tri 23025 34914 23026 34915 ne
rect 23026 34914 23154 34915
tri 23026 34913 23027 34914 ne
rect 23027 34913 23154 34914
tri 23027 34912 23028 34913 ne
rect 23028 34912 23154 34913
tri 23028 34911 23029 34912 ne
rect 23029 34911 23154 34912
tri 23029 34910 23030 34911 ne
rect 23030 34910 23154 34911
tri 23030 34909 23031 34910 ne
rect 23031 34909 23154 34910
tri 23031 34908 23032 34909 ne
rect 23032 34908 23154 34909
tri 23032 34907 23033 34908 ne
rect 23033 34907 23154 34908
tri 23033 34906 23034 34907 ne
rect 23034 34906 23154 34907
tri 23034 34905 23035 34906 ne
rect 23035 34905 23154 34906
tri 23035 34904 23036 34905 ne
rect 23036 34904 23154 34905
tri 23036 34903 23037 34904 ne
rect 23037 34903 23154 34904
tri 23037 34902 23038 34903 ne
rect 23038 34902 23154 34903
tri 23038 34901 23039 34902 ne
rect 23039 34901 23154 34902
tri 23039 34891 23049 34901 ne
rect 23049 34891 23154 34901
tri 23049 34846 23094 34891 ne
rect 23094 34878 23154 34891
rect 23200 34901 23270 34924
tri 23270 34901 23315 34946 sw
rect 70802 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34878 23315 34901
rect 23094 34856 23315 34878
tri 23315 34856 23360 34901 sw
rect 70802 34860 71000 34918
rect 23094 34846 23360 34856
tri 23094 34801 23139 34846 ne
rect 23139 34811 23360 34846
tri 23360 34811 23405 34856 sw
rect 70802 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23139 34801 23405 34811
tri 23139 34756 23184 34801 ne
rect 23184 34794 23405 34801
tri 23405 34794 23422 34811 sw
rect 23184 34792 23422 34794
rect 23184 34756 23286 34792
tri 23184 34711 23229 34756 ne
rect 23229 34746 23286 34756
rect 23332 34749 23422 34792
tri 23422 34749 23467 34794 sw
rect 70802 34756 71000 34814
rect 23332 34746 23467 34749
rect 23229 34711 23467 34746
tri 23229 34704 23236 34711 ne
rect 23236 34704 23467 34711
tri 23467 34704 23512 34749 sw
rect 70802 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23236 34694 23246 34704 ne
rect 23246 34694 23512 34704
tri 23246 34693 23247 34694 ne
rect 23247 34693 23512 34694
tri 23247 34692 23248 34693 ne
rect 23248 34692 23512 34693
tri 23248 34691 23249 34692 ne
rect 23249 34691 23512 34692
tri 23249 34690 23250 34691 ne
rect 23250 34690 23512 34691
tri 23250 34689 23251 34690 ne
rect 23251 34689 23512 34690
tri 23251 34688 23252 34689 ne
rect 23252 34688 23512 34689
tri 23252 34687 23253 34688 ne
rect 23253 34687 23512 34688
tri 23253 34686 23254 34687 ne
rect 23254 34686 23512 34687
tri 23254 34685 23255 34686 ne
rect 23255 34685 23512 34686
tri 23255 34684 23256 34685 ne
rect 23256 34684 23512 34685
tri 23256 34683 23257 34684 ne
rect 23257 34683 23512 34684
tri 23257 34682 23258 34683 ne
rect 23258 34682 23512 34683
tri 23258 34681 23259 34682 ne
rect 23259 34681 23512 34682
tri 23259 34680 23260 34681 ne
rect 23260 34680 23512 34681
tri 23260 34679 23261 34680 ne
rect 23261 34679 23512 34680
tri 23261 34678 23262 34679 ne
rect 23262 34678 23512 34679
tri 23262 34677 23263 34678 ne
rect 23263 34677 23512 34678
tri 23263 34676 23264 34677 ne
rect 23264 34676 23512 34677
tri 23264 34675 23265 34676 ne
rect 23265 34675 23512 34676
tri 23265 34674 23266 34675 ne
rect 23266 34674 23512 34675
tri 23266 34673 23267 34674 ne
rect 23267 34673 23512 34674
tri 23267 34672 23268 34673 ne
rect 23268 34672 23512 34673
tri 23268 34671 23269 34672 ne
rect 23269 34671 23512 34672
tri 23269 34670 23270 34671 ne
rect 23270 34670 23512 34671
tri 23270 34669 23271 34670 ne
rect 23271 34669 23512 34670
tri 23271 34668 23272 34669 ne
rect 23272 34668 23512 34669
tri 23272 34667 23273 34668 ne
rect 23273 34667 23512 34668
tri 23273 34666 23274 34667 ne
rect 23274 34666 23512 34667
tri 23274 34665 23275 34666 ne
rect 23275 34665 23512 34666
tri 23275 34664 23276 34665 ne
rect 23276 34664 23512 34665
tri 23276 34663 23277 34664 ne
rect 23277 34663 23512 34664
tri 23277 34662 23278 34663 ne
rect 23278 34662 23512 34663
tri 23278 34661 23279 34662 ne
rect 23279 34661 23512 34662
tri 23279 34660 23280 34661 ne
rect 23280 34660 23512 34661
tri 23280 34659 23281 34660 ne
rect 23281 34659 23418 34660
tri 23281 34658 23282 34659 ne
rect 23282 34658 23418 34659
tri 23282 34657 23283 34658 ne
rect 23283 34657 23418 34658
tri 23283 34656 23284 34657 ne
rect 23284 34656 23418 34657
tri 23284 34655 23285 34656 ne
rect 23285 34655 23418 34656
tri 23285 34654 23286 34655 ne
rect 23286 34654 23418 34655
tri 23286 34653 23287 34654 ne
rect 23287 34653 23418 34654
tri 23287 34652 23288 34653 ne
rect 23288 34652 23418 34653
tri 23288 34651 23289 34652 ne
rect 23289 34651 23418 34652
tri 23289 34650 23290 34651 ne
rect 23290 34650 23418 34651
tri 23290 34649 23291 34650 ne
rect 23291 34649 23418 34650
tri 23291 34648 23292 34649 ne
rect 23292 34648 23418 34649
tri 23292 34647 23293 34648 ne
rect 23293 34647 23418 34648
tri 23293 34646 23294 34647 ne
rect 23294 34646 23418 34647
tri 23294 34645 23295 34646 ne
rect 23295 34645 23418 34646
tri 23295 34644 23296 34645 ne
rect 23296 34644 23418 34645
tri 23296 34643 23297 34644 ne
rect 23297 34643 23418 34644
tri 23297 34642 23298 34643 ne
rect 23298 34642 23418 34643
tri 23298 34641 23299 34642 ne
rect 23299 34641 23418 34642
tri 23299 34640 23300 34641 ne
rect 23300 34640 23418 34641
tri 23300 34639 23301 34640 ne
rect 23301 34639 23418 34640
tri 23301 34638 23302 34639 ne
rect 23302 34638 23418 34639
tri 23302 34637 23303 34638 ne
rect 23303 34637 23418 34638
tri 23303 34636 23304 34637 ne
rect 23304 34636 23418 34637
tri 23304 34635 23305 34636 ne
rect 23305 34635 23418 34636
tri 23305 34634 23306 34635 ne
rect 23306 34634 23418 34635
tri 23306 34633 23307 34634 ne
rect 23307 34633 23418 34634
tri 23307 34632 23308 34633 ne
rect 23308 34632 23418 34633
tri 23308 34631 23309 34632 ne
rect 23309 34631 23418 34632
tri 23309 34630 23310 34631 ne
rect 23310 34630 23418 34631
tri 23310 34629 23311 34630 ne
rect 23311 34629 23418 34630
tri 23311 34628 23312 34629 ne
rect 23312 34628 23418 34629
tri 23312 34627 23313 34628 ne
rect 23313 34627 23418 34628
tri 23313 34626 23314 34627 ne
rect 23314 34626 23418 34627
tri 23314 34625 23315 34626 ne
rect 23315 34625 23418 34626
tri 23315 34580 23360 34625 ne
rect 23360 34614 23418 34625
rect 23464 34659 23512 34660
tri 23512 34659 23557 34704 sw
rect 23464 34625 23557 34659
tri 23557 34625 23591 34659 sw
rect 70802 34652 71000 34710
rect 23464 34614 23591 34625
tri 23591 34614 23602 34625 sw
rect 23360 34580 23602 34614
tri 23360 34571 23369 34580 ne
rect 23369 34571 23602 34580
tri 23369 34526 23414 34571 ne
rect 23414 34569 23602 34571
tri 23602 34569 23647 34614 sw
rect 70802 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 23414 34528 23647 34569
rect 23414 34526 23550 34528
tri 23414 34481 23459 34526 ne
rect 23459 34482 23550 34526
rect 23596 34524 23647 34528
tri 23647 34524 23692 34569 sw
rect 70802 34548 71000 34606
rect 23596 34484 23692 34524
tri 23692 34484 23732 34524 sw
rect 70802 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 23596 34482 23732 34484
rect 23459 34481 23732 34482
tri 23459 34436 23504 34481 ne
rect 23504 34439 23732 34481
tri 23732 34439 23777 34484 sw
rect 70802 34444 71000 34502
rect 23504 34436 23777 34439
tri 23504 34420 23520 34436 ne
rect 23520 34420 23777 34436
tri 23520 34419 23521 34420 ne
rect 23521 34419 23777 34420
tri 23521 34418 23522 34419 ne
rect 23522 34418 23777 34419
tri 23522 34417 23523 34418 ne
rect 23523 34417 23777 34418
tri 23523 34416 23524 34417 ne
rect 23524 34416 23777 34417
tri 23524 34415 23525 34416 ne
rect 23525 34415 23777 34416
tri 23525 34414 23526 34415 ne
rect 23526 34414 23777 34415
tri 23526 34413 23527 34414 ne
rect 23527 34413 23777 34414
tri 23527 34412 23528 34413 ne
rect 23528 34412 23777 34413
tri 23528 34411 23529 34412 ne
rect 23529 34411 23777 34412
tri 23529 34410 23530 34411 ne
rect 23530 34410 23777 34411
tri 23530 34409 23531 34410 ne
rect 23531 34409 23777 34410
tri 23531 34408 23532 34409 ne
rect 23532 34408 23777 34409
tri 23532 34407 23533 34408 ne
rect 23533 34407 23777 34408
tri 23533 34406 23534 34407 ne
rect 23534 34406 23777 34407
tri 23534 34405 23535 34406 ne
rect 23535 34405 23777 34406
tri 23535 34404 23536 34405 ne
rect 23536 34404 23777 34405
tri 23536 34403 23537 34404 ne
rect 23537 34403 23777 34404
tri 23537 34402 23538 34403 ne
rect 23538 34402 23777 34403
tri 23538 34401 23539 34402 ne
rect 23539 34401 23777 34402
tri 23539 34400 23540 34401 ne
rect 23540 34400 23777 34401
tri 23540 34399 23541 34400 ne
rect 23541 34399 23777 34400
tri 23541 34398 23542 34399 ne
rect 23542 34398 23777 34399
tri 23542 34397 23543 34398 ne
rect 23543 34397 23777 34398
tri 23543 34396 23544 34397 ne
rect 23544 34396 23777 34397
tri 23544 34395 23545 34396 ne
rect 23545 34395 23682 34396
tri 23545 34394 23546 34395 ne
rect 23546 34394 23682 34395
tri 23546 34393 23547 34394 ne
rect 23547 34393 23682 34394
tri 23547 34392 23548 34393 ne
rect 23548 34392 23682 34393
tri 23548 34391 23549 34392 ne
rect 23549 34391 23682 34392
tri 23549 34390 23550 34391 ne
rect 23550 34390 23682 34391
tri 23550 34389 23551 34390 ne
rect 23551 34389 23682 34390
tri 23551 34388 23552 34389 ne
rect 23552 34388 23682 34389
tri 23552 34387 23553 34388 ne
rect 23553 34387 23682 34388
tri 23553 34386 23554 34387 ne
rect 23554 34386 23682 34387
tri 23554 34385 23555 34386 ne
rect 23555 34385 23682 34386
tri 23555 34384 23556 34385 ne
rect 23556 34384 23682 34385
tri 23556 34383 23557 34384 ne
rect 23557 34383 23682 34384
tri 23557 34382 23558 34383 ne
rect 23558 34382 23682 34383
tri 23558 34381 23559 34382 ne
rect 23559 34381 23682 34382
tri 23559 34380 23560 34381 ne
rect 23560 34380 23682 34381
tri 23560 34379 23561 34380 ne
rect 23561 34379 23682 34380
tri 23561 34378 23562 34379 ne
rect 23562 34378 23682 34379
tri 23562 34377 23563 34378 ne
rect 23563 34377 23682 34378
tri 23563 34376 23564 34377 ne
rect 23564 34376 23682 34377
tri 23564 34375 23565 34376 ne
rect 23565 34375 23682 34376
tri 23565 34374 23566 34375 ne
rect 23566 34374 23682 34375
tri 23566 34373 23567 34374 ne
rect 23567 34373 23682 34374
tri 23567 34372 23568 34373 ne
rect 23568 34372 23682 34373
tri 23568 34371 23569 34372 ne
rect 23569 34371 23682 34372
tri 23569 34370 23570 34371 ne
rect 23570 34370 23682 34371
tri 23570 34369 23571 34370 ne
rect 23571 34369 23682 34370
tri 23571 34368 23572 34369 ne
rect 23572 34368 23682 34369
tri 23572 34367 23573 34368 ne
rect 23573 34367 23682 34368
tri 23573 34366 23574 34367 ne
rect 23574 34366 23682 34367
tri 23574 34365 23575 34366 ne
rect 23575 34365 23682 34366
tri 23575 34364 23576 34365 ne
rect 23576 34364 23682 34365
tri 23576 34363 23577 34364 ne
rect 23577 34363 23682 34364
tri 23577 34362 23578 34363 ne
rect 23578 34362 23682 34363
tri 23578 34361 23579 34362 ne
rect 23579 34361 23682 34362
tri 23579 34360 23580 34361 ne
rect 23580 34360 23682 34361
tri 23580 34359 23581 34360 ne
rect 23581 34359 23682 34360
tri 23581 34358 23582 34359 ne
rect 23582 34358 23682 34359
tri 23582 34357 23583 34358 ne
rect 23583 34357 23682 34358
tri 23583 34356 23584 34357 ne
rect 23584 34356 23682 34357
tri 23584 34355 23585 34356 ne
rect 23585 34355 23682 34356
tri 23585 34354 23586 34355 ne
rect 23586 34354 23682 34355
tri 23586 34353 23587 34354 ne
rect 23587 34353 23682 34354
tri 23587 34352 23588 34353 ne
rect 23588 34352 23682 34353
tri 23588 34351 23589 34352 ne
rect 23589 34351 23682 34352
tri 23589 34350 23590 34351 ne
rect 23590 34350 23682 34351
rect 23728 34394 23777 34396
tri 23777 34394 23822 34439 sw
rect 70802 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 23728 34350 23822 34394
tri 23590 34349 23591 34350 ne
rect 23591 34349 23822 34350
tri 23822 34349 23867 34394 sw
tri 23591 34338 23602 34349 ne
rect 23602 34338 23867 34349
tri 23867 34338 23878 34349 sw
rect 70802 34340 71000 34398
tri 23602 34304 23636 34338 ne
rect 23636 34304 23878 34338
tri 23636 34293 23647 34304 ne
rect 23647 34293 23878 34304
tri 23878 34293 23923 34338 sw
rect 70802 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23647 34248 23692 34293 ne
rect 23692 34264 23923 34293
rect 23692 34248 23814 34264
tri 23692 34207 23733 34248 ne
rect 23733 34218 23814 34248
rect 23860 34248 23923 34264
tri 23923 34248 23968 34293 sw
rect 23860 34218 23968 34248
rect 23733 34207 23968 34218
tri 23733 34162 23778 34207 ne
rect 23778 34203 23968 34207
tri 23968 34203 24013 34248 sw
rect 70802 34236 71000 34294
rect 23778 34163 24013 34203
tri 24013 34163 24053 34203 sw
rect 70802 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 23778 34162 24053 34163
tri 23778 34145 23795 34162 ne
rect 23795 34145 24053 34162
tri 23795 34144 23796 34145 ne
rect 23796 34144 24053 34145
tri 23796 34143 23797 34144 ne
rect 23797 34143 24053 34144
tri 23797 34142 23798 34143 ne
rect 23798 34142 24053 34143
tri 23798 34141 23799 34142 ne
rect 23799 34141 24053 34142
tri 23799 34140 23800 34141 ne
rect 23800 34140 24053 34141
tri 23800 34139 23801 34140 ne
rect 23801 34139 24053 34140
tri 23801 34138 23802 34139 ne
rect 23802 34138 24053 34139
tri 23802 34137 23803 34138 ne
rect 23803 34137 24053 34138
tri 23803 34136 23804 34137 ne
rect 23804 34136 24053 34137
tri 23804 34135 23805 34136 ne
rect 23805 34135 24053 34136
tri 23805 34134 23806 34135 ne
rect 23806 34134 24053 34135
tri 23806 34133 23807 34134 ne
rect 23807 34133 24053 34134
tri 23807 34132 23808 34133 ne
rect 23808 34132 24053 34133
tri 23808 34131 23809 34132 ne
rect 23809 34131 23946 34132
tri 23809 34130 23810 34131 ne
rect 23810 34130 23946 34131
tri 23810 34129 23811 34130 ne
rect 23811 34129 23946 34130
tri 23811 34128 23812 34129 ne
rect 23812 34128 23946 34129
tri 23812 34127 23813 34128 ne
rect 23813 34127 23946 34128
tri 23813 34126 23814 34127 ne
rect 23814 34126 23946 34127
tri 23814 34125 23815 34126 ne
rect 23815 34125 23946 34126
tri 23815 34124 23816 34125 ne
rect 23816 34124 23946 34125
tri 23816 34123 23817 34124 ne
rect 23817 34123 23946 34124
tri 23817 34122 23818 34123 ne
rect 23818 34122 23946 34123
tri 23818 34121 23819 34122 ne
rect 23819 34121 23946 34122
tri 23819 34120 23820 34121 ne
rect 23820 34120 23946 34121
tri 23820 34119 23821 34120 ne
rect 23821 34119 23946 34120
tri 23821 34118 23822 34119 ne
rect 23822 34118 23946 34119
tri 23822 34117 23823 34118 ne
rect 23823 34117 23946 34118
tri 23823 34116 23824 34117 ne
rect 23824 34116 23946 34117
tri 23824 34115 23825 34116 ne
rect 23825 34115 23946 34116
tri 23825 34114 23826 34115 ne
rect 23826 34114 23946 34115
tri 23826 34113 23827 34114 ne
rect 23827 34113 23946 34114
tri 23827 34112 23828 34113 ne
rect 23828 34112 23946 34113
tri 23828 34111 23829 34112 ne
rect 23829 34111 23946 34112
tri 23829 34110 23830 34111 ne
rect 23830 34110 23946 34111
tri 23830 34109 23831 34110 ne
rect 23831 34109 23946 34110
tri 23831 34108 23832 34109 ne
rect 23832 34108 23946 34109
tri 23832 34107 23833 34108 ne
rect 23833 34107 23946 34108
tri 23833 34106 23834 34107 ne
rect 23834 34106 23946 34107
tri 23834 34105 23835 34106 ne
rect 23835 34105 23946 34106
tri 23835 34104 23836 34105 ne
rect 23836 34104 23946 34105
tri 23836 34103 23837 34104 ne
rect 23837 34103 23946 34104
tri 23837 34102 23838 34103 ne
rect 23838 34102 23946 34103
tri 23838 34101 23839 34102 ne
rect 23839 34101 23946 34102
tri 23839 34100 23840 34101 ne
rect 23840 34100 23946 34101
tri 23840 34099 23841 34100 ne
rect 23841 34099 23946 34100
tri 23841 34098 23842 34099 ne
rect 23842 34098 23946 34099
tri 23842 34097 23843 34098 ne
rect 23843 34097 23946 34098
tri 23843 34096 23844 34097 ne
rect 23844 34096 23946 34097
tri 23844 34095 23845 34096 ne
rect 23845 34095 23946 34096
tri 23845 34094 23846 34095 ne
rect 23846 34094 23946 34095
tri 23846 34093 23847 34094 ne
rect 23847 34093 23946 34094
tri 23847 34092 23848 34093 ne
rect 23848 34092 23946 34093
tri 23848 34091 23849 34092 ne
rect 23849 34091 23946 34092
tri 23849 34090 23850 34091 ne
rect 23850 34090 23946 34091
tri 23850 34089 23851 34090 ne
rect 23851 34089 23946 34090
tri 23851 34088 23852 34089 ne
rect 23852 34088 23946 34089
tri 23852 34087 23853 34088 ne
rect 23853 34087 23946 34088
tri 23853 34086 23854 34087 ne
rect 23854 34086 23946 34087
rect 23992 34118 24053 34132
tri 24053 34118 24098 34163 sw
rect 70802 34132 71000 34190
rect 23992 34086 24098 34118
tri 23854 34085 23855 34086 ne
rect 23855 34085 24098 34086
tri 23855 34084 23856 34085 ne
rect 23856 34084 24098 34085
tri 23856 34083 23857 34084 ne
rect 23857 34083 24098 34084
tri 23857 34082 23858 34083 ne
rect 23858 34082 24098 34083
tri 23858 34081 23859 34082 ne
rect 23859 34081 24098 34082
tri 23859 34080 23860 34081 ne
rect 23860 34080 24098 34081
tri 23860 34079 23861 34080 ne
rect 23861 34079 24098 34080
tri 23861 34078 23862 34079 ne
rect 23862 34078 24098 34079
tri 23862 34077 23863 34078 ne
rect 23863 34077 24098 34078
tri 23863 34076 23864 34077 ne
rect 23864 34076 24098 34077
tri 23864 34075 23865 34076 ne
rect 23865 34075 24098 34076
tri 23865 34074 23866 34075 ne
rect 23866 34074 24098 34075
tri 23866 34073 23867 34074 ne
rect 23867 34073 24098 34074
tri 24098 34073 24143 34118 sw
rect 70802 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
tri 23867 34028 23912 34073 ne
rect 23912 34028 24143 34073
tri 24143 34028 24188 34073 sw
rect 70802 34028 71000 34086
tri 23912 33983 23957 34028 ne
rect 23957 34017 24188 34028
tri 24188 34017 24199 34028 sw
rect 23957 34000 24199 34017
rect 23957 33983 24078 34000
tri 23957 33972 23968 33983 ne
rect 23968 33972 24078 33983
tri 23968 33938 24002 33972 ne
rect 24002 33954 24078 33972
rect 24124 33972 24199 34000
tri 24199 33972 24244 34017 sw
rect 70802 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33954 24244 33972
rect 24002 33938 24244 33954
tri 24002 33927 24013 33938 ne
rect 24013 33927 24244 33938
tri 24244 33927 24289 33972 sw
tri 24013 33882 24058 33927 ne
rect 24058 33882 24289 33927
tri 24289 33882 24334 33927 sw
rect 70802 33924 71000 33982
tri 24058 33871 24069 33882 ne
rect 24069 33871 24334 33882
tri 24069 33870 24070 33871 ne
rect 24070 33870 24334 33871
tri 24070 33869 24071 33870 ne
rect 24071 33869 24334 33870
tri 24071 33868 24072 33869 ne
rect 24072 33868 24334 33869
tri 24072 33867 24073 33868 ne
rect 24073 33867 24210 33868
tri 24073 33866 24074 33867 ne
rect 24074 33866 24210 33867
tri 24074 33865 24075 33866 ne
rect 24075 33865 24210 33866
tri 24075 33864 24076 33865 ne
rect 24076 33864 24210 33865
tri 24076 33863 24077 33864 ne
rect 24077 33863 24210 33864
tri 24077 33862 24078 33863 ne
rect 24078 33862 24210 33863
tri 24078 33861 24079 33862 ne
rect 24079 33861 24210 33862
tri 24079 33860 24080 33861 ne
rect 24080 33860 24210 33861
tri 24080 33859 24081 33860 ne
rect 24081 33859 24210 33860
tri 24081 33858 24082 33859 ne
rect 24082 33858 24210 33859
tri 24082 33857 24083 33858 ne
rect 24083 33857 24210 33858
tri 24083 33856 24084 33857 ne
rect 24084 33856 24210 33857
tri 24084 33855 24085 33856 ne
rect 24085 33855 24210 33856
tri 24085 33854 24086 33855 ne
rect 24086 33854 24210 33855
tri 24086 33853 24087 33854 ne
rect 24087 33853 24210 33854
tri 24087 33852 24088 33853 ne
rect 24088 33852 24210 33853
tri 24088 33851 24089 33852 ne
rect 24089 33851 24210 33852
tri 24089 33850 24090 33851 ne
rect 24090 33850 24210 33851
tri 24090 33849 24091 33850 ne
rect 24091 33849 24210 33850
tri 24091 33848 24092 33849 ne
rect 24092 33848 24210 33849
tri 24092 33847 24093 33848 ne
rect 24093 33847 24210 33848
tri 24093 33846 24094 33847 ne
rect 24094 33846 24210 33847
tri 24094 33845 24095 33846 ne
rect 24095 33845 24210 33846
tri 24095 33844 24096 33845 ne
rect 24096 33844 24210 33845
tri 24096 33843 24097 33844 ne
rect 24097 33843 24210 33844
tri 24097 33842 24098 33843 ne
rect 24098 33842 24210 33843
tri 24098 33841 24099 33842 ne
rect 24099 33841 24210 33842
tri 24099 33840 24100 33841 ne
rect 24100 33840 24210 33841
tri 24100 33839 24101 33840 ne
rect 24101 33839 24210 33840
tri 24101 33838 24102 33839 ne
rect 24102 33838 24210 33839
tri 24102 33837 24103 33838 ne
rect 24103 33837 24210 33838
tri 24103 33836 24104 33837 ne
rect 24104 33836 24210 33837
tri 24104 33835 24105 33836 ne
rect 24105 33835 24210 33836
tri 24105 33834 24106 33835 ne
rect 24106 33834 24210 33835
tri 24106 33833 24107 33834 ne
rect 24107 33833 24210 33834
tri 24107 33832 24108 33833 ne
rect 24108 33832 24210 33833
tri 24108 33831 24109 33832 ne
rect 24109 33831 24210 33832
tri 24109 33830 24110 33831 ne
rect 24110 33830 24210 33831
tri 24110 33829 24111 33830 ne
rect 24111 33829 24210 33830
tri 24111 33828 24112 33829 ne
rect 24112 33828 24210 33829
tri 24112 33827 24113 33828 ne
rect 24113 33827 24210 33828
tri 24113 33826 24114 33827 ne
rect 24114 33826 24210 33827
tri 24114 33825 24115 33826 ne
rect 24115 33825 24210 33826
tri 24115 33824 24116 33825 ne
rect 24116 33824 24210 33825
tri 24116 33823 24117 33824 ne
rect 24117 33823 24210 33824
tri 24117 33822 24118 33823 ne
rect 24118 33822 24210 33823
rect 24256 33842 24334 33868
tri 24334 33842 24374 33882 sw
rect 70802 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 24256 33822 24374 33842
tri 24118 33821 24119 33822 ne
rect 24119 33821 24374 33822
tri 24119 33820 24120 33821 ne
rect 24120 33820 24374 33821
tri 24120 33819 24121 33820 ne
rect 24121 33819 24374 33820
tri 24121 33818 24122 33819 ne
rect 24122 33818 24374 33819
tri 24122 33817 24123 33818 ne
rect 24123 33817 24374 33818
tri 24123 33816 24124 33817 ne
rect 24124 33816 24374 33817
tri 24124 33815 24125 33816 ne
rect 24125 33815 24374 33816
tri 24125 33814 24126 33815 ne
rect 24126 33814 24374 33815
tri 24126 33813 24127 33814 ne
rect 24127 33813 24374 33814
tri 24127 33812 24128 33813 ne
rect 24128 33812 24374 33813
tri 24128 33811 24129 33812 ne
rect 24129 33811 24374 33812
tri 24129 33810 24130 33811 ne
rect 24130 33810 24374 33811
tri 24130 33809 24131 33810 ne
rect 24131 33809 24374 33810
tri 24131 33808 24132 33809 ne
rect 24132 33808 24374 33809
tri 24132 33807 24133 33808 ne
rect 24133 33807 24374 33808
tri 24133 33806 24134 33807 ne
rect 24134 33806 24374 33807
tri 24134 33805 24135 33806 ne
rect 24135 33805 24374 33806
tri 24135 33804 24136 33805 ne
rect 24136 33804 24374 33805
tri 24136 33803 24137 33804 ne
rect 24137 33803 24374 33804
tri 24137 33802 24138 33803 ne
rect 24138 33802 24374 33803
tri 24138 33801 24139 33802 ne
rect 24139 33801 24374 33802
tri 24139 33800 24140 33801 ne
rect 24140 33800 24374 33801
tri 24140 33799 24141 33800 ne
rect 24141 33799 24374 33800
tri 24141 33798 24142 33799 ne
rect 24142 33798 24374 33799
tri 24142 33797 24143 33798 ne
rect 24143 33797 24374 33798
tri 24374 33797 24419 33842 sw
rect 70802 33820 71000 33878
tri 24143 33752 24188 33797 ne
rect 24188 33752 24419 33797
tri 24419 33752 24464 33797 sw
rect 70802 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24188 33707 24233 33752 ne
rect 24233 33736 24464 33752
rect 24233 33707 24342 33736
tri 24233 33662 24278 33707 ne
rect 24278 33690 24342 33707
rect 24388 33707 24464 33736
tri 24464 33707 24509 33752 sw
rect 70802 33716 71000 33774
rect 24388 33696 24509 33707
tri 24509 33696 24520 33707 sw
rect 24388 33690 24520 33696
rect 24278 33662 24520 33690
tri 24278 33617 24323 33662 ne
rect 24323 33651 24520 33662
tri 24520 33651 24565 33696 sw
rect 70802 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
rect 24323 33617 24565 33651
tri 24323 33606 24334 33617 ne
rect 24334 33606 24565 33617
tri 24565 33606 24610 33651 sw
rect 70802 33612 71000 33670
tri 24334 33597 24343 33606 ne
rect 24343 33604 24610 33606
rect 24343 33597 24474 33604
tri 24343 33596 24344 33597 ne
rect 24344 33596 24474 33597
tri 24344 33595 24345 33596 ne
rect 24345 33595 24474 33596
tri 24345 33594 24346 33595 ne
rect 24346 33594 24474 33595
tri 24346 33593 24347 33594 ne
rect 24347 33593 24474 33594
tri 24347 33592 24348 33593 ne
rect 24348 33592 24474 33593
tri 24348 33591 24349 33592 ne
rect 24349 33591 24474 33592
tri 24349 33590 24350 33591 ne
rect 24350 33590 24474 33591
tri 24350 33589 24351 33590 ne
rect 24351 33589 24474 33590
tri 24351 33588 24352 33589 ne
rect 24352 33588 24474 33589
tri 24352 33587 24353 33588 ne
rect 24353 33587 24474 33588
tri 24353 33586 24354 33587 ne
rect 24354 33586 24474 33587
tri 24354 33585 24355 33586 ne
rect 24355 33585 24474 33586
tri 24355 33584 24356 33585 ne
rect 24356 33584 24474 33585
tri 24356 33583 24357 33584 ne
rect 24357 33583 24474 33584
tri 24357 33582 24358 33583 ne
rect 24358 33582 24474 33583
tri 24358 33581 24359 33582 ne
rect 24359 33581 24474 33582
tri 24359 33580 24360 33581 ne
rect 24360 33580 24474 33581
tri 24360 33579 24361 33580 ne
rect 24361 33579 24474 33580
tri 24361 33578 24362 33579 ne
rect 24362 33578 24474 33579
tri 24362 33577 24363 33578 ne
rect 24363 33577 24474 33578
tri 24363 33576 24364 33577 ne
rect 24364 33576 24474 33577
tri 24364 33575 24365 33576 ne
rect 24365 33575 24474 33576
tri 24365 33574 24366 33575 ne
rect 24366 33574 24474 33575
tri 24366 33573 24367 33574 ne
rect 24367 33573 24474 33574
tri 24367 33572 24368 33573 ne
rect 24368 33572 24474 33573
tri 24368 33571 24369 33572 ne
rect 24369 33571 24474 33572
tri 24369 33570 24370 33571 ne
rect 24370 33570 24474 33571
tri 24370 33569 24371 33570 ne
rect 24371 33569 24474 33570
tri 24371 33568 24372 33569 ne
rect 24372 33568 24474 33569
tri 24372 33567 24373 33568 ne
rect 24373 33567 24474 33568
tri 24373 33566 24374 33567 ne
rect 24374 33566 24474 33567
tri 24374 33565 24375 33566 ne
rect 24375 33565 24474 33566
tri 24375 33564 24376 33565 ne
rect 24376 33564 24474 33565
tri 24376 33563 24377 33564 ne
rect 24377 33563 24474 33564
tri 24377 33562 24378 33563 ne
rect 24378 33562 24474 33563
tri 24378 33561 24379 33562 ne
rect 24379 33561 24474 33562
tri 24379 33560 24380 33561 ne
rect 24380 33560 24474 33561
tri 24380 33559 24381 33560 ne
rect 24381 33559 24474 33560
tri 24381 33558 24382 33559 ne
rect 24382 33558 24474 33559
rect 24520 33561 24610 33604
tri 24610 33561 24655 33606 sw
rect 70802 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 24520 33558 24655 33561
tri 24382 33557 24383 33558 ne
rect 24383 33557 24655 33558
tri 24383 33556 24384 33557 ne
rect 24384 33556 24655 33557
tri 24384 33555 24385 33556 ne
rect 24385 33555 24655 33556
tri 24385 33554 24386 33555 ne
rect 24386 33554 24655 33555
tri 24386 33553 24387 33554 ne
rect 24387 33553 24655 33554
tri 24387 33552 24388 33553 ne
rect 24388 33552 24655 33553
tri 24388 33551 24389 33552 ne
rect 24389 33551 24655 33552
tri 24389 33550 24390 33551 ne
rect 24390 33550 24655 33551
tri 24390 33549 24391 33550 ne
rect 24391 33549 24655 33550
tri 24391 33548 24392 33549 ne
rect 24392 33548 24655 33549
tri 24392 33547 24393 33548 ne
rect 24393 33547 24655 33548
tri 24393 33546 24394 33547 ne
rect 24394 33546 24655 33547
tri 24394 33545 24395 33546 ne
rect 24395 33545 24655 33546
tri 24395 33544 24396 33545 ne
rect 24396 33544 24655 33545
tri 24396 33543 24397 33544 ne
rect 24397 33543 24655 33544
tri 24397 33542 24398 33543 ne
rect 24398 33542 24655 33543
tri 24398 33541 24399 33542 ne
rect 24399 33541 24655 33542
tri 24399 33540 24400 33541 ne
rect 24400 33540 24655 33541
tri 24400 33539 24401 33540 ne
rect 24401 33539 24655 33540
tri 24401 33538 24402 33539 ne
rect 24402 33538 24655 33539
tri 24402 33537 24403 33538 ne
rect 24403 33537 24655 33538
tri 24403 33536 24404 33537 ne
rect 24404 33536 24655 33537
tri 24404 33535 24405 33536 ne
rect 24405 33535 24655 33536
tri 24405 33534 24406 33535 ne
rect 24406 33534 24655 33535
tri 24406 33533 24407 33534 ne
rect 24407 33533 24655 33534
tri 24407 33532 24408 33533 ne
rect 24408 33532 24655 33533
tri 24408 33531 24409 33532 ne
rect 24409 33531 24655 33532
tri 24409 33530 24410 33531 ne
rect 24410 33530 24655 33531
tri 24410 33529 24411 33530 ne
rect 24411 33529 24655 33530
tri 24411 33528 24412 33529 ne
rect 24412 33528 24655 33529
tri 24412 33527 24413 33528 ne
rect 24413 33527 24655 33528
tri 24413 33526 24414 33527 ne
rect 24414 33526 24655 33527
tri 24414 33525 24415 33526 ne
rect 24415 33525 24655 33526
tri 24415 33524 24416 33525 ne
rect 24416 33524 24655 33525
tri 24416 33523 24417 33524 ne
rect 24417 33523 24655 33524
tri 24417 33522 24418 33523 ne
rect 24418 33522 24655 33523
tri 24418 33521 24419 33522 ne
rect 24419 33521 24655 33522
tri 24655 33521 24695 33561 sw
tri 24419 33476 24464 33521 ne
rect 24464 33516 24695 33521
tri 24695 33516 24700 33521 sw
rect 24464 33476 24700 33516
tri 24464 33432 24508 33476 ne
rect 24508 33472 24700 33476
rect 24508 33432 24606 33472
tri 24508 33387 24553 33432 ne
rect 24553 33426 24606 33432
rect 24652 33471 24700 33472
tri 24700 33471 24745 33516 sw
rect 70802 33508 71000 33566
rect 24652 33426 24745 33471
tri 24745 33426 24790 33471 sw
rect 70802 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24553 33387 24790 33426
tri 24553 33342 24598 33387 ne
rect 24598 33381 24790 33387
tri 24790 33381 24835 33426 sw
rect 70802 33404 71000 33462
rect 24598 33380 24835 33381
tri 24835 33380 24836 33381 sw
rect 24598 33342 24836 33380
tri 24598 33322 24618 33342 ne
rect 24618 33340 24836 33342
rect 24618 33322 24738 33340
tri 24618 33321 24619 33322 ne
rect 24619 33321 24738 33322
tri 24619 33320 24620 33321 ne
rect 24620 33320 24738 33321
tri 24620 33319 24621 33320 ne
rect 24621 33319 24738 33320
tri 24621 33318 24622 33319 ne
rect 24622 33318 24738 33319
tri 24622 33317 24623 33318 ne
rect 24623 33317 24738 33318
tri 24623 33316 24624 33317 ne
rect 24624 33316 24738 33317
tri 24624 33315 24625 33316 ne
rect 24625 33315 24738 33316
tri 24625 33314 24626 33315 ne
rect 24626 33314 24738 33315
tri 24626 33313 24627 33314 ne
rect 24627 33313 24738 33314
tri 24627 33312 24628 33313 ne
rect 24628 33312 24738 33313
tri 24628 33311 24629 33312 ne
rect 24629 33311 24738 33312
tri 24629 33310 24630 33311 ne
rect 24630 33310 24738 33311
tri 24630 33309 24631 33310 ne
rect 24631 33309 24738 33310
tri 24631 33308 24632 33309 ne
rect 24632 33308 24738 33309
tri 24632 33307 24633 33308 ne
rect 24633 33307 24738 33308
tri 24633 33306 24634 33307 ne
rect 24634 33306 24738 33307
tri 24634 33305 24635 33306 ne
rect 24635 33305 24738 33306
tri 24635 33304 24636 33305 ne
rect 24636 33304 24738 33305
tri 24636 33303 24637 33304 ne
rect 24637 33303 24738 33304
tri 24637 33302 24638 33303 ne
rect 24638 33302 24738 33303
tri 24638 33301 24639 33302 ne
rect 24639 33301 24738 33302
tri 24639 33300 24640 33301 ne
rect 24640 33300 24738 33301
tri 24640 33299 24641 33300 ne
rect 24641 33299 24738 33300
tri 24641 33298 24642 33299 ne
rect 24642 33298 24738 33299
tri 24642 33297 24643 33298 ne
rect 24643 33297 24738 33298
tri 24643 33296 24644 33297 ne
rect 24644 33296 24738 33297
tri 24644 33295 24645 33296 ne
rect 24645 33295 24738 33296
tri 24645 33294 24646 33295 ne
rect 24646 33294 24738 33295
rect 24784 33335 24836 33340
tri 24836 33335 24881 33380 sw
rect 70802 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 24784 33294 24881 33335
tri 24646 33293 24647 33294 ne
rect 24647 33293 24881 33294
tri 24647 33292 24648 33293 ne
rect 24648 33292 24881 33293
tri 24648 33291 24649 33292 ne
rect 24649 33291 24881 33292
tri 24649 33290 24650 33291 ne
rect 24650 33290 24881 33291
tri 24881 33290 24926 33335 sw
rect 70802 33300 71000 33358
tri 24650 33289 24651 33290 ne
rect 24651 33289 24926 33290
tri 24651 33288 24652 33289 ne
rect 24652 33288 24926 33289
tri 24652 33287 24653 33288 ne
rect 24653 33287 24926 33288
tri 24653 33286 24654 33287 ne
rect 24654 33286 24926 33287
tri 24654 33285 24655 33286 ne
rect 24655 33285 24926 33286
tri 24655 33284 24656 33285 ne
rect 24656 33284 24926 33285
tri 24656 33283 24657 33284 ne
rect 24657 33283 24926 33284
tri 24657 33282 24658 33283 ne
rect 24658 33282 24926 33283
tri 24658 33281 24659 33282 ne
rect 24659 33281 24926 33282
tri 24659 33280 24660 33281 ne
rect 24660 33280 24926 33281
tri 24660 33279 24661 33280 ne
rect 24661 33279 24926 33280
tri 24661 33278 24662 33279 ne
rect 24662 33278 24926 33279
tri 24662 33277 24663 33278 ne
rect 24663 33277 24926 33278
tri 24663 33276 24664 33277 ne
rect 24664 33276 24926 33277
tri 24664 33275 24665 33276 ne
rect 24665 33275 24926 33276
tri 24665 33274 24666 33275 ne
rect 24666 33274 24926 33275
tri 24666 33273 24667 33274 ne
rect 24667 33273 24926 33274
tri 24667 33272 24668 33273 ne
rect 24668 33272 24926 33273
tri 24668 33271 24669 33272 ne
rect 24669 33271 24926 33272
tri 24669 33270 24670 33271 ne
rect 24670 33270 24926 33271
tri 24670 33269 24671 33270 ne
rect 24671 33269 24926 33270
tri 24671 33268 24672 33269 ne
rect 24672 33268 24926 33269
tri 24672 33267 24673 33268 ne
rect 24673 33267 24926 33268
tri 24673 33266 24674 33267 ne
rect 24674 33266 24926 33267
tri 24674 33265 24675 33266 ne
rect 24675 33265 24926 33266
tri 24675 33264 24676 33265 ne
rect 24676 33264 24926 33265
tri 24676 33263 24677 33264 ne
rect 24677 33263 24926 33264
tri 24677 33262 24678 33263 ne
rect 24678 33262 24926 33263
tri 24678 33261 24679 33262 ne
rect 24679 33261 24926 33262
tri 24679 33260 24680 33261 ne
rect 24680 33260 24926 33261
tri 24680 33259 24681 33260 ne
rect 24681 33259 24926 33260
tri 24681 33258 24682 33259 ne
rect 24682 33258 24926 33259
tri 24682 33257 24683 33258 ne
rect 24683 33257 24926 33258
tri 24683 33256 24684 33257 ne
rect 24684 33256 24926 33257
tri 24684 33255 24685 33256 ne
rect 24685 33255 24926 33256
tri 24685 33254 24686 33255 ne
rect 24686 33254 24926 33255
tri 24686 33253 24687 33254 ne
rect 24687 33253 24926 33254
tri 24687 33252 24688 33253 ne
rect 24688 33252 24926 33253
tri 24688 33251 24689 33252 ne
rect 24689 33251 24926 33252
tri 24689 33250 24690 33251 ne
rect 24690 33250 24926 33251
tri 24690 33249 24691 33250 ne
rect 24691 33249 24926 33250
tri 24691 33248 24692 33249 ne
rect 24692 33248 24926 33249
tri 24692 33247 24693 33248 ne
rect 24693 33247 24926 33248
tri 24693 33246 24694 33247 ne
rect 24694 33246 24926 33247
tri 24694 33245 24695 33246 ne
rect 24695 33245 24926 33246
tri 24926 33245 24971 33290 sw
rect 70802 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24695 33240 24700 33245 ne
rect 24700 33240 24971 33245
tri 24971 33240 24976 33245 sw
tri 24700 33200 24740 33240 ne
rect 24740 33208 24976 33240
rect 24740 33200 24870 33208
tri 24740 33195 24745 33200 ne
rect 24745 33195 24870 33200
tri 24745 33150 24790 33195 ne
rect 24790 33162 24870 33195
rect 24916 33195 24976 33208
tri 24976 33195 25021 33240 sw
rect 70802 33196 71000 33254
rect 24916 33162 25021 33195
rect 24790 33150 25021 33162
tri 25021 33150 25066 33195 sw
rect 70802 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
tri 24790 33112 24828 33150 ne
rect 24828 33112 25066 33150
tri 24828 33067 24873 33112 ne
rect 24873 33105 25066 33112
tri 25066 33105 25111 33150 sw
rect 24873 33076 25111 33105
rect 24873 33067 25002 33076
tri 24873 33048 24892 33067 ne
rect 24892 33048 25002 33067
tri 24892 33047 24893 33048 ne
rect 24893 33047 25002 33048
tri 24893 33046 24894 33047 ne
rect 24894 33046 25002 33047
tri 24894 33045 24895 33046 ne
rect 24895 33045 25002 33046
tri 24895 33044 24896 33045 ne
rect 24896 33044 25002 33045
tri 24896 33043 24897 33044 ne
rect 24897 33043 25002 33044
tri 24897 33042 24898 33043 ne
rect 24898 33042 25002 33043
tri 24898 33041 24899 33042 ne
rect 24899 33041 25002 33042
tri 24899 33040 24900 33041 ne
rect 24900 33040 25002 33041
tri 24900 33039 24901 33040 ne
rect 24901 33039 25002 33040
tri 24901 33038 24902 33039 ne
rect 24902 33038 25002 33039
tri 24902 33037 24903 33038 ne
rect 24903 33037 25002 33038
tri 24903 33036 24904 33037 ne
rect 24904 33036 25002 33037
tri 24904 33035 24905 33036 ne
rect 24905 33035 25002 33036
tri 24905 33034 24906 33035 ne
rect 24906 33034 25002 33035
tri 24906 33033 24907 33034 ne
rect 24907 33033 25002 33034
tri 24907 33032 24908 33033 ne
rect 24908 33032 25002 33033
tri 24908 33031 24909 33032 ne
rect 24909 33031 25002 33032
tri 24909 33030 24910 33031 ne
rect 24910 33030 25002 33031
rect 25048 33060 25111 33076
tri 25111 33060 25156 33105 sw
rect 70802 33092 71000 33150
rect 25048 33059 25156 33060
tri 25156 33059 25157 33060 sw
rect 25048 33030 25157 33059
tri 24910 33029 24911 33030 ne
rect 24911 33029 25157 33030
tri 24911 33028 24912 33029 ne
rect 24912 33028 25157 33029
tri 24912 33027 24913 33028 ne
rect 24913 33027 25157 33028
tri 24913 33026 24914 33027 ne
rect 24914 33026 25157 33027
tri 24914 33025 24915 33026 ne
rect 24915 33025 25157 33026
tri 24915 33024 24916 33025 ne
rect 24916 33024 25157 33025
tri 24916 33023 24917 33024 ne
rect 24917 33023 25157 33024
tri 24917 33022 24918 33023 ne
rect 24918 33022 25157 33023
tri 24918 33021 24919 33022 ne
rect 24919 33021 25157 33022
tri 24919 33020 24920 33021 ne
rect 24920 33020 25157 33021
tri 24920 33019 24921 33020 ne
rect 24921 33019 25157 33020
tri 24921 33018 24922 33019 ne
rect 24922 33018 25157 33019
tri 24922 33017 24923 33018 ne
rect 24923 33017 25157 33018
tri 24923 33016 24924 33017 ne
rect 24924 33016 25157 33017
tri 24924 33015 24925 33016 ne
rect 24925 33015 25157 33016
tri 24925 33014 24926 33015 ne
rect 24926 33014 25157 33015
tri 25157 33014 25202 33059 sw
rect 70802 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
tri 24926 33013 24927 33014 ne
rect 24927 33013 25202 33014
tri 24927 33012 24928 33013 ne
rect 24928 33012 25202 33013
tri 24928 33011 24929 33012 ne
rect 24929 33011 25202 33012
tri 24929 33010 24930 33011 ne
rect 24930 33010 25202 33011
tri 24930 33009 24931 33010 ne
rect 24931 33009 25202 33010
tri 24931 33008 24932 33009 ne
rect 24932 33008 25202 33009
tri 24932 33007 24933 33008 ne
rect 24933 33007 25202 33008
tri 24933 33006 24934 33007 ne
rect 24934 33006 25202 33007
tri 24934 33005 24935 33006 ne
rect 24935 33005 25202 33006
tri 24935 33004 24936 33005 ne
rect 24936 33004 25202 33005
tri 24936 33003 24937 33004 ne
rect 24937 33003 25202 33004
tri 24937 33002 24938 33003 ne
rect 24938 33002 25202 33003
tri 24938 33001 24939 33002 ne
rect 24939 33001 25202 33002
tri 24939 33000 24940 33001 ne
rect 24940 33000 25202 33001
tri 24940 32999 24941 33000 ne
rect 24941 32999 25202 33000
tri 24941 32998 24942 32999 ne
rect 24942 32998 25202 32999
tri 24942 32997 24943 32998 ne
rect 24943 32997 25202 32998
tri 24943 32996 24944 32997 ne
rect 24944 32996 25202 32997
tri 24944 32995 24945 32996 ne
rect 24945 32995 25202 32996
tri 24945 32994 24946 32995 ne
rect 24946 32994 25202 32995
tri 24946 32993 24947 32994 ne
rect 24947 32993 25202 32994
tri 24947 32992 24948 32993 ne
rect 24948 32992 25202 32993
tri 24948 32991 24949 32992 ne
rect 24949 32991 25202 32992
tri 24949 32990 24950 32991 ne
rect 24950 32990 25202 32991
tri 24950 32989 24951 32990 ne
rect 24951 32989 25202 32990
tri 24951 32988 24952 32989 ne
rect 24952 32988 25202 32989
tri 24952 32987 24953 32988 ne
rect 24953 32987 25202 32988
tri 24953 32986 24954 32987 ne
rect 24954 32986 25202 32987
tri 24954 32985 24955 32986 ne
rect 24955 32985 25202 32986
tri 24955 32984 24956 32985 ne
rect 24956 32984 25202 32985
tri 24956 32983 24957 32984 ne
rect 24957 32983 25202 32984
tri 24957 32982 24958 32983 ne
rect 24958 32982 25202 32983
tri 24958 32981 24959 32982 ne
rect 24959 32981 25202 32982
tri 24959 32980 24960 32981 ne
rect 24960 32980 25202 32981
tri 24960 32979 24961 32980 ne
rect 24961 32979 25202 32980
tri 24961 32978 24962 32979 ne
rect 24962 32978 25202 32979
tri 24962 32977 24963 32978 ne
rect 24963 32977 25202 32978
tri 24963 32976 24964 32977 ne
rect 24964 32976 25202 32977
tri 24964 32975 24965 32976 ne
rect 24965 32975 25202 32976
tri 24965 32974 24966 32975 ne
rect 24966 32974 25202 32975
tri 24966 32973 24967 32974 ne
rect 24967 32973 25202 32974
tri 24967 32972 24968 32973 ne
rect 24968 32972 25202 32973
tri 24968 32971 24969 32972 ne
rect 24969 32971 25202 32972
tri 24969 32970 24970 32971 ne
rect 24970 32970 25202 32971
tri 24970 32969 24971 32970 ne
rect 24971 32969 25202 32970
tri 25202 32969 25247 33014 sw
rect 70802 32988 71000 33046
tri 24971 32924 25016 32969 ne
rect 25016 32944 25247 32969
rect 25016 32924 25134 32944
tri 25016 32879 25061 32924 ne
rect 25061 32898 25134 32924
rect 25180 32924 25247 32944
tri 25247 32924 25292 32969 sw
rect 70802 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32919 25292 32924
tri 25292 32919 25297 32924 sw
rect 25180 32898 25297 32919
rect 25061 32879 25297 32898
tri 25061 32874 25066 32879 ne
rect 25066 32874 25297 32879
tri 25297 32874 25342 32919 sw
rect 70802 32884 71000 32942
tri 25066 32834 25106 32874 ne
rect 25106 32834 25342 32874
tri 25106 32829 25111 32834 ne
rect 25111 32829 25342 32834
tri 25342 32829 25387 32874 sw
rect 70802 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
tri 25111 32784 25156 32829 ne
rect 25156 32812 25387 32829
rect 25156 32784 25266 32812
tri 25156 32773 25167 32784 ne
rect 25167 32773 25266 32784
tri 25167 32772 25168 32773 ne
rect 25168 32772 25266 32773
tri 25168 32771 25169 32772 ne
rect 25169 32771 25266 32772
tri 25169 32770 25170 32771 ne
rect 25170 32770 25266 32771
tri 25170 32769 25171 32770 ne
rect 25171 32769 25266 32770
tri 25171 32768 25172 32769 ne
rect 25172 32768 25266 32769
tri 25172 32767 25173 32768 ne
rect 25173 32767 25266 32768
tri 25173 32766 25174 32767 ne
rect 25174 32766 25266 32767
rect 25312 32784 25387 32812
tri 25387 32784 25432 32829 sw
rect 25312 32766 25432 32784
tri 25174 32765 25175 32766 ne
rect 25175 32765 25432 32766
tri 25175 32764 25176 32765 ne
rect 25176 32764 25432 32765
tri 25176 32763 25177 32764 ne
rect 25177 32763 25432 32764
tri 25177 32762 25178 32763 ne
rect 25178 32762 25432 32763
tri 25178 32761 25179 32762 ne
rect 25179 32761 25432 32762
tri 25179 32760 25180 32761 ne
rect 25180 32760 25432 32761
tri 25180 32759 25181 32760 ne
rect 25181 32759 25432 32760
tri 25181 32758 25182 32759 ne
rect 25182 32758 25432 32759
tri 25182 32757 25183 32758 ne
rect 25183 32757 25432 32758
tri 25183 32756 25184 32757 ne
rect 25184 32756 25432 32757
tri 25184 32755 25185 32756 ne
rect 25185 32755 25432 32756
tri 25185 32754 25186 32755 ne
rect 25186 32754 25432 32755
tri 25186 32753 25187 32754 ne
rect 25187 32753 25432 32754
tri 25187 32752 25188 32753 ne
rect 25188 32752 25432 32753
tri 25188 32751 25189 32752 ne
rect 25189 32751 25432 32752
tri 25189 32750 25190 32751 ne
rect 25190 32750 25432 32751
tri 25190 32749 25191 32750 ne
rect 25191 32749 25432 32750
tri 25191 32748 25192 32749 ne
rect 25192 32748 25432 32749
tri 25192 32747 25193 32748 ne
rect 25193 32747 25432 32748
tri 25193 32746 25194 32747 ne
rect 25194 32746 25432 32747
tri 25194 32745 25195 32746 ne
rect 25195 32745 25432 32746
tri 25195 32744 25196 32745 ne
rect 25196 32744 25432 32745
tri 25196 32743 25197 32744 ne
rect 25197 32743 25432 32744
tri 25197 32742 25198 32743 ne
rect 25198 32742 25432 32743
tri 25198 32741 25199 32742 ne
rect 25199 32741 25432 32742
tri 25199 32740 25200 32741 ne
rect 25200 32740 25432 32741
tri 25200 32739 25201 32740 ne
rect 25201 32739 25432 32740
tri 25432 32739 25477 32784 sw
rect 70802 32780 71000 32838
tri 25201 32738 25202 32739 ne
rect 25202 32738 25477 32739
tri 25477 32738 25478 32739 sw
tri 25202 32737 25203 32738 ne
rect 25203 32737 25478 32738
tri 25203 32736 25204 32737 ne
rect 25204 32736 25478 32737
tri 25204 32735 25205 32736 ne
rect 25205 32735 25478 32736
tri 25205 32734 25206 32735 ne
rect 25206 32734 25478 32735
tri 25206 32733 25207 32734 ne
rect 25207 32733 25478 32734
tri 25207 32732 25208 32733 ne
rect 25208 32732 25478 32733
tri 25208 32731 25209 32732 ne
rect 25209 32731 25478 32732
tri 25209 32730 25210 32731 ne
rect 25210 32730 25478 32731
tri 25210 32729 25211 32730 ne
rect 25211 32729 25478 32730
tri 25211 32728 25212 32729 ne
rect 25212 32728 25478 32729
tri 25212 32727 25213 32728 ne
rect 25213 32727 25478 32728
tri 25213 32726 25214 32727 ne
rect 25214 32726 25478 32727
tri 25214 32725 25215 32726 ne
rect 25215 32725 25478 32726
tri 25215 32724 25216 32725 ne
rect 25216 32724 25478 32725
tri 25216 32723 25217 32724 ne
rect 25217 32723 25478 32724
tri 25217 32722 25218 32723 ne
rect 25218 32722 25478 32723
tri 25218 32721 25219 32722 ne
rect 25219 32721 25478 32722
tri 25219 32720 25220 32721 ne
rect 25220 32720 25478 32721
tri 25220 32719 25221 32720 ne
rect 25221 32719 25478 32720
tri 25221 32718 25222 32719 ne
rect 25222 32718 25478 32719
tri 25222 32717 25223 32718 ne
rect 25223 32717 25478 32718
tri 25223 32716 25224 32717 ne
rect 25224 32716 25478 32717
tri 25224 32715 25225 32716 ne
rect 25225 32715 25478 32716
tri 25225 32714 25226 32715 ne
rect 25226 32714 25478 32715
tri 25226 32713 25227 32714 ne
rect 25227 32713 25478 32714
tri 25227 32712 25228 32713 ne
rect 25228 32712 25478 32713
tri 25228 32711 25229 32712 ne
rect 25229 32711 25478 32712
tri 25229 32710 25230 32711 ne
rect 25230 32710 25478 32711
tri 25230 32709 25231 32710 ne
rect 25231 32709 25478 32710
tri 25231 32708 25232 32709 ne
rect 25232 32708 25478 32709
tri 25232 32707 25233 32708 ne
rect 25233 32707 25478 32708
tri 25233 32706 25234 32707 ne
rect 25234 32706 25478 32707
tri 25234 32705 25235 32706 ne
rect 25235 32705 25478 32706
tri 25235 32704 25236 32705 ne
rect 25236 32704 25478 32705
tri 25236 32703 25237 32704 ne
rect 25237 32703 25478 32704
tri 25237 32702 25238 32703 ne
rect 25238 32702 25478 32703
tri 25238 32701 25239 32702 ne
rect 25239 32701 25478 32702
tri 25239 32700 25240 32701 ne
rect 25240 32700 25478 32701
tri 25240 32699 25241 32700 ne
rect 25241 32699 25478 32700
tri 25241 32698 25242 32699 ne
rect 25242 32698 25478 32699
tri 25242 32697 25243 32698 ne
rect 25243 32697 25478 32698
tri 25243 32696 25244 32697 ne
rect 25244 32696 25478 32697
tri 25244 32695 25245 32696 ne
rect 25245 32695 25478 32696
tri 25245 32694 25246 32695 ne
rect 25246 32694 25478 32695
tri 25246 32693 25247 32694 ne
rect 25247 32693 25478 32694
tri 25478 32693 25523 32738 sw
rect 70802 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25247 32648 25292 32693 ne
rect 25292 32680 25523 32693
rect 25292 32648 25398 32680
tri 25292 32603 25337 32648 ne
rect 25337 32634 25398 32648
rect 25444 32648 25523 32680
tri 25523 32648 25568 32693 sw
rect 70802 32676 71000 32734
rect 25444 32634 25568 32648
rect 25337 32603 25568 32634
tri 25568 32603 25613 32648 sw
rect 70802 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25337 32558 25382 32603 ne
rect 25382 32598 25613 32603
tri 25613 32598 25618 32603 sw
rect 25382 32558 25618 32598
tri 25382 32513 25427 32558 ne
rect 25427 32553 25618 32558
tri 25618 32553 25663 32598 sw
rect 70802 32572 71000 32630
rect 25427 32548 25663 32553
rect 25427 32513 25530 32548
tri 25427 32508 25432 32513 ne
rect 25432 32508 25530 32513
tri 25432 32499 25441 32508 ne
rect 25441 32502 25530 32508
rect 25576 32508 25663 32548
tri 25663 32508 25708 32553 sw
rect 70802 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 25576 32502 25708 32508
rect 25441 32499 25708 32502
tri 25441 32498 25442 32499 ne
rect 25442 32498 25708 32499
tri 25442 32497 25443 32498 ne
rect 25443 32497 25708 32498
tri 25443 32496 25444 32497 ne
rect 25444 32496 25708 32497
tri 25444 32495 25445 32496 ne
rect 25445 32495 25708 32496
tri 25445 32494 25446 32495 ne
rect 25446 32494 25708 32495
tri 25446 32493 25447 32494 ne
rect 25447 32493 25708 32494
tri 25447 32492 25448 32493 ne
rect 25448 32492 25708 32493
tri 25448 32491 25449 32492 ne
rect 25449 32491 25708 32492
tri 25449 32490 25450 32491 ne
rect 25450 32490 25708 32491
tri 25450 32489 25451 32490 ne
rect 25451 32489 25708 32490
tri 25451 32488 25452 32489 ne
rect 25452 32488 25708 32489
tri 25452 32487 25453 32488 ne
rect 25453 32487 25708 32488
tri 25453 32486 25454 32487 ne
rect 25454 32486 25708 32487
tri 25454 32485 25455 32486 ne
rect 25455 32485 25708 32486
tri 25455 32484 25456 32485 ne
rect 25456 32484 25708 32485
tri 25456 32483 25457 32484 ne
rect 25457 32483 25708 32484
tri 25457 32482 25458 32483 ne
rect 25458 32482 25708 32483
tri 25458 32481 25459 32482 ne
rect 25459 32481 25708 32482
tri 25459 32480 25460 32481 ne
rect 25460 32480 25708 32481
tri 25460 32479 25461 32480 ne
rect 25461 32479 25708 32480
tri 25461 32478 25462 32479 ne
rect 25462 32478 25708 32479
tri 25462 32477 25463 32478 ne
rect 25463 32477 25708 32478
tri 25463 32476 25464 32477 ne
rect 25464 32476 25708 32477
tri 25464 32475 25465 32476 ne
rect 25465 32475 25708 32476
tri 25465 32474 25466 32475 ne
rect 25466 32474 25708 32475
tri 25466 32473 25467 32474 ne
rect 25467 32473 25708 32474
tri 25467 32472 25468 32473 ne
rect 25468 32472 25708 32473
tri 25468 32471 25469 32472 ne
rect 25469 32471 25708 32472
tri 25469 32470 25470 32471 ne
rect 25470 32470 25708 32471
tri 25470 32469 25471 32470 ne
rect 25471 32469 25708 32470
tri 25471 32468 25472 32469 ne
rect 25472 32468 25708 32469
tri 25472 32467 25473 32468 ne
rect 25473 32467 25708 32468
tri 25473 32466 25474 32467 ne
rect 25474 32466 25708 32467
tri 25474 32465 25475 32466 ne
rect 25475 32465 25708 32466
tri 25475 32464 25476 32465 ne
rect 25476 32464 25708 32465
tri 25476 32463 25477 32464 ne
rect 25477 32463 25708 32464
tri 25708 32463 25753 32508 sw
rect 70802 32468 71000 32526
tri 25477 32462 25478 32463 ne
rect 25478 32462 25753 32463
tri 25478 32461 25479 32462 ne
rect 25479 32461 25753 32462
tri 25479 32460 25480 32461 ne
rect 25480 32460 25753 32461
tri 25480 32459 25481 32460 ne
rect 25481 32459 25753 32460
tri 25481 32458 25482 32459 ne
rect 25482 32458 25753 32459
tri 25482 32457 25483 32458 ne
rect 25483 32457 25753 32458
tri 25483 32456 25484 32457 ne
rect 25484 32456 25753 32457
tri 25484 32455 25485 32456 ne
rect 25485 32455 25753 32456
tri 25485 32454 25486 32455 ne
rect 25486 32454 25753 32455
tri 25486 32453 25487 32454 ne
rect 25487 32453 25753 32454
tri 25487 32452 25488 32453 ne
rect 25488 32452 25753 32453
tri 25488 32451 25489 32452 ne
rect 25489 32451 25753 32452
tri 25489 32450 25490 32451 ne
rect 25490 32450 25753 32451
tri 25490 32449 25491 32450 ne
rect 25491 32449 25753 32450
tri 25491 32448 25492 32449 ne
rect 25492 32448 25753 32449
tri 25492 32447 25493 32448 ne
rect 25493 32447 25753 32448
tri 25493 32446 25494 32447 ne
rect 25494 32446 25753 32447
tri 25494 32445 25495 32446 ne
rect 25495 32445 25753 32446
tri 25495 32444 25496 32445 ne
rect 25496 32444 25753 32445
tri 25496 32443 25497 32444 ne
rect 25497 32443 25753 32444
tri 25497 32442 25498 32443 ne
rect 25498 32442 25753 32443
tri 25498 32441 25499 32442 ne
rect 25499 32441 25753 32442
tri 25499 32440 25500 32441 ne
rect 25500 32440 25753 32441
tri 25500 32439 25501 32440 ne
rect 25501 32439 25753 32440
tri 25501 32438 25502 32439 ne
rect 25502 32438 25753 32439
tri 25502 32437 25503 32438 ne
rect 25503 32437 25753 32438
tri 25503 32436 25504 32437 ne
rect 25504 32436 25753 32437
tri 25504 32435 25505 32436 ne
rect 25505 32435 25753 32436
tri 25505 32434 25506 32435 ne
rect 25506 32434 25753 32435
tri 25506 32433 25507 32434 ne
rect 25507 32433 25753 32434
tri 25507 32432 25508 32433 ne
rect 25508 32432 25753 32433
tri 25508 32431 25509 32432 ne
rect 25509 32431 25753 32432
tri 25509 32430 25510 32431 ne
rect 25510 32430 25753 32431
tri 25510 32429 25511 32430 ne
rect 25511 32429 25753 32430
tri 25511 32428 25512 32429 ne
rect 25512 32428 25753 32429
tri 25512 32427 25513 32428 ne
rect 25513 32427 25753 32428
tri 25513 32426 25514 32427 ne
rect 25514 32426 25753 32427
tri 25514 32425 25515 32426 ne
rect 25515 32425 25753 32426
tri 25515 32424 25516 32425 ne
rect 25516 32424 25753 32425
tri 25516 32423 25517 32424 ne
rect 25517 32423 25753 32424
tri 25517 32422 25518 32423 ne
rect 25518 32422 25753 32423
tri 25518 32421 25519 32422 ne
rect 25519 32421 25753 32422
tri 25519 32420 25520 32421 ne
rect 25520 32420 25753 32421
tri 25520 32419 25521 32420 ne
rect 25521 32419 25753 32420
tri 25521 32418 25522 32419 ne
rect 25522 32418 25753 32419
tri 25753 32418 25798 32463 sw
rect 70802 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
tri 25522 32417 25523 32418 ne
rect 25523 32417 25798 32418
tri 25798 32417 25799 32418 sw
tri 25523 32372 25568 32417 ne
rect 25568 32416 25799 32417
rect 25568 32372 25662 32416
tri 25568 32338 25602 32372 ne
rect 25602 32370 25662 32372
rect 25708 32372 25799 32416
tri 25799 32372 25844 32417 sw
rect 25708 32370 25844 32372
rect 25602 32338 25844 32370
tri 25602 32293 25647 32338 ne
rect 25647 32327 25844 32338
tri 25844 32327 25889 32372 sw
rect 70802 32364 71000 32422
rect 25647 32293 25889 32327
tri 25647 32248 25692 32293 ne
rect 25692 32284 25889 32293
rect 25692 32248 25794 32284
tri 25692 32225 25715 32248 ne
rect 25715 32238 25794 32248
rect 25840 32282 25889 32284
tri 25889 32282 25934 32327 sw
rect 70802 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
rect 25840 32276 25934 32282
tri 25934 32276 25940 32282 sw
rect 25840 32238 25940 32276
rect 25715 32231 25940 32238
tri 25940 32231 25985 32276 sw
rect 70802 32260 71000 32318
rect 25715 32225 25985 32231
tri 25715 32224 25716 32225 ne
rect 25716 32224 25985 32225
tri 25716 32223 25717 32224 ne
rect 25717 32223 25985 32224
tri 25717 32222 25718 32223 ne
rect 25718 32222 25985 32223
tri 25718 32221 25719 32222 ne
rect 25719 32221 25985 32222
tri 25719 32220 25720 32221 ne
rect 25720 32220 25985 32221
tri 25720 32219 25721 32220 ne
rect 25721 32219 25985 32220
tri 25721 32218 25722 32219 ne
rect 25722 32218 25985 32219
tri 25722 32217 25723 32218 ne
rect 25723 32217 25985 32218
tri 25723 32216 25724 32217 ne
rect 25724 32216 25985 32217
tri 25724 32215 25725 32216 ne
rect 25725 32215 25985 32216
tri 25725 32214 25726 32215 ne
rect 25726 32214 25985 32215
tri 25726 32213 25727 32214 ne
rect 25727 32213 25985 32214
tri 25727 32212 25728 32213 ne
rect 25728 32212 25985 32213
tri 25728 32211 25729 32212 ne
rect 25729 32211 25985 32212
tri 25729 32210 25730 32211 ne
rect 25730 32210 25985 32211
tri 25730 32209 25731 32210 ne
rect 25731 32209 25985 32210
tri 25731 32208 25732 32209 ne
rect 25732 32208 25985 32209
tri 25732 32207 25733 32208 ne
rect 25733 32207 25985 32208
tri 25733 32206 25734 32207 ne
rect 25734 32206 25985 32207
tri 25734 32205 25735 32206 ne
rect 25735 32205 25985 32206
tri 25735 32204 25736 32205 ne
rect 25736 32204 25985 32205
tri 25736 32203 25737 32204 ne
rect 25737 32203 25985 32204
tri 25737 32202 25738 32203 ne
rect 25738 32202 25985 32203
tri 25738 32201 25739 32202 ne
rect 25739 32201 25985 32202
tri 25739 32200 25740 32201 ne
rect 25740 32200 25985 32201
tri 25740 32199 25741 32200 ne
rect 25741 32199 25985 32200
tri 25741 32198 25742 32199 ne
rect 25742 32198 25985 32199
tri 25742 32197 25743 32198 ne
rect 25743 32197 25985 32198
tri 25743 32196 25744 32197 ne
rect 25744 32196 25985 32197
tri 25744 32195 25745 32196 ne
rect 25745 32195 25985 32196
tri 25745 32194 25746 32195 ne
rect 25746 32194 25985 32195
tri 25746 32193 25747 32194 ne
rect 25747 32193 25985 32194
tri 25747 32192 25748 32193 ne
rect 25748 32192 25985 32193
tri 25748 32191 25749 32192 ne
rect 25749 32191 25985 32192
tri 25749 32190 25750 32191 ne
rect 25750 32190 25985 32191
tri 25750 32189 25751 32190 ne
rect 25751 32189 25985 32190
tri 25751 32188 25752 32189 ne
rect 25752 32188 25985 32189
tri 25752 32187 25753 32188 ne
rect 25753 32187 25985 32188
tri 25753 32186 25754 32187 ne
rect 25754 32186 25985 32187
tri 25985 32186 26030 32231 sw
rect 70802 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25754 32185 25755 32186 ne
rect 25755 32185 26030 32186
tri 25755 32184 25756 32185 ne
rect 25756 32184 26030 32185
tri 25756 32183 25757 32184 ne
rect 25757 32183 26030 32184
tri 25757 32182 25758 32183 ne
rect 25758 32182 26030 32183
tri 25758 32181 25759 32182 ne
rect 25759 32181 26030 32182
tri 25759 32180 25760 32181 ne
rect 25760 32180 26030 32181
tri 25760 32179 25761 32180 ne
rect 25761 32179 26030 32180
tri 25761 32178 25762 32179 ne
rect 25762 32178 26030 32179
tri 25762 32177 25763 32178 ne
rect 25763 32177 26030 32178
tri 25763 32176 25764 32177 ne
rect 25764 32176 26030 32177
tri 25764 32175 25765 32176 ne
rect 25765 32175 26030 32176
tri 25765 32174 25766 32175 ne
rect 25766 32174 26030 32175
tri 25766 32173 25767 32174 ne
rect 25767 32173 26030 32174
tri 25767 32172 25768 32173 ne
rect 25768 32172 26030 32173
tri 25768 32171 25769 32172 ne
rect 25769 32171 26030 32172
tri 25769 32170 25770 32171 ne
rect 25770 32170 26030 32171
tri 25770 32169 25771 32170 ne
rect 25771 32169 26030 32170
tri 25771 32168 25772 32169 ne
rect 25772 32168 26030 32169
tri 25772 32167 25773 32168 ne
rect 25773 32167 26030 32168
tri 25773 32166 25774 32167 ne
rect 25774 32166 26030 32167
tri 25774 32165 25775 32166 ne
rect 25775 32165 26030 32166
tri 25775 32164 25776 32165 ne
rect 25776 32164 26030 32165
tri 25776 32163 25777 32164 ne
rect 25777 32163 26030 32164
tri 25777 32162 25778 32163 ne
rect 25778 32162 26030 32163
tri 25778 32161 25779 32162 ne
rect 25779 32161 26030 32162
tri 25779 32160 25780 32161 ne
rect 25780 32160 26030 32161
tri 25780 32159 25781 32160 ne
rect 25781 32159 26030 32160
tri 25781 32158 25782 32159 ne
rect 25782 32158 26030 32159
tri 25782 32157 25783 32158 ne
rect 25783 32157 26030 32158
tri 25783 32156 25784 32157 ne
rect 25784 32156 26030 32157
tri 25784 32155 25785 32156 ne
rect 25785 32155 26030 32156
tri 25785 32154 25786 32155 ne
rect 25786 32154 26030 32155
tri 25786 32153 25787 32154 ne
rect 25787 32153 26030 32154
tri 25787 32152 25788 32153 ne
rect 25788 32152 26030 32153
tri 25788 32151 25789 32152 ne
rect 25789 32151 25926 32152
tri 25789 32150 25790 32151 ne
rect 25790 32150 25926 32151
tri 25790 32149 25791 32150 ne
rect 25791 32149 25926 32150
tri 25791 32148 25792 32149 ne
rect 25792 32148 25926 32149
tri 25792 32147 25793 32148 ne
rect 25793 32147 25926 32148
tri 25793 32146 25794 32147 ne
rect 25794 32146 25926 32147
tri 25794 32145 25795 32146 ne
rect 25795 32145 25926 32146
tri 25795 32144 25796 32145 ne
rect 25796 32144 25926 32145
tri 25796 32143 25797 32144 ne
rect 25797 32143 25926 32144
tri 25797 32142 25798 32143 ne
rect 25798 32142 25926 32143
tri 25798 32141 25799 32142 ne
rect 25799 32141 25926 32142
tri 25799 32097 25843 32141 ne
rect 25843 32106 25926 32141
rect 25972 32141 26030 32152
tri 26030 32141 26075 32186 sw
rect 70802 32156 71000 32214
rect 25972 32106 26075 32141
rect 25843 32097 26075 32106
tri 26075 32097 26119 32141 sw
rect 70802 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
tri 25843 32052 25888 32097 ne
rect 25888 32052 26119 32097
tri 26119 32052 26164 32097 sw
rect 70802 32052 71000 32110
tri 25888 32018 25922 32052 ne
rect 25922 32020 26164 32052
rect 25922 32018 26058 32020
tri 25922 31973 25967 32018 ne
rect 25967 31974 26058 32018
rect 26104 32007 26164 32020
tri 26164 32007 26209 32052 sw
rect 26104 31974 26209 32007
rect 25967 31973 26209 31974
tri 25967 31950 25990 31973 ne
rect 25990 31962 26209 31973
tri 26209 31962 26254 32007 sw
rect 70802 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 25990 31955 26254 31962
tri 26254 31955 26261 31962 sw
rect 25990 31950 26261 31955
tri 25990 31949 25991 31950 ne
rect 25991 31949 26261 31950
tri 25991 31948 25992 31949 ne
rect 25992 31948 26261 31949
tri 25992 31947 25993 31948 ne
rect 25993 31947 26261 31948
tri 25993 31946 25994 31947 ne
rect 25994 31946 26261 31947
tri 25994 31945 25995 31946 ne
rect 25995 31945 26261 31946
tri 25995 31944 25996 31945 ne
rect 25996 31944 26261 31945
tri 25996 31943 25997 31944 ne
rect 25997 31943 26261 31944
tri 25997 31942 25998 31943 ne
rect 25998 31942 26261 31943
tri 25998 31941 25999 31942 ne
rect 25999 31941 26261 31942
tri 25999 31940 26000 31941 ne
rect 26000 31940 26261 31941
tri 26000 31939 26001 31940 ne
rect 26001 31939 26261 31940
tri 26001 31938 26002 31939 ne
rect 26002 31938 26261 31939
tri 26002 31937 26003 31938 ne
rect 26003 31937 26261 31938
tri 26003 31936 26004 31937 ne
rect 26004 31936 26261 31937
tri 26004 31935 26005 31936 ne
rect 26005 31935 26261 31936
tri 26005 31934 26006 31935 ne
rect 26006 31934 26261 31935
tri 26006 31933 26007 31934 ne
rect 26007 31933 26261 31934
tri 26007 31932 26008 31933 ne
rect 26008 31932 26261 31933
tri 26008 31931 26009 31932 ne
rect 26009 31931 26261 31932
tri 26009 31930 26010 31931 ne
rect 26010 31930 26261 31931
tri 26010 31929 26011 31930 ne
rect 26011 31929 26261 31930
tri 26011 31928 26012 31929 ne
rect 26012 31928 26261 31929
tri 26012 31927 26013 31928 ne
rect 26013 31927 26261 31928
tri 26013 31926 26014 31927 ne
rect 26014 31926 26261 31927
tri 26014 31925 26015 31926 ne
rect 26015 31925 26261 31926
tri 26015 31924 26016 31925 ne
rect 26016 31924 26261 31925
tri 26016 31923 26017 31924 ne
rect 26017 31923 26261 31924
tri 26017 31922 26018 31923 ne
rect 26018 31922 26261 31923
tri 26018 31921 26019 31922 ne
rect 26019 31921 26261 31922
tri 26019 31920 26020 31921 ne
rect 26020 31920 26261 31921
tri 26020 31919 26021 31920 ne
rect 26021 31919 26261 31920
tri 26021 31918 26022 31919 ne
rect 26022 31918 26261 31919
tri 26022 31917 26023 31918 ne
rect 26023 31917 26261 31918
tri 26023 31916 26024 31917 ne
rect 26024 31916 26261 31917
tri 26024 31915 26025 31916 ne
rect 26025 31915 26261 31916
tri 26025 31914 26026 31915 ne
rect 26026 31914 26261 31915
tri 26026 31913 26027 31914 ne
rect 26027 31913 26261 31914
tri 26027 31912 26028 31913 ne
rect 26028 31912 26261 31913
tri 26028 31911 26029 31912 ne
rect 26029 31911 26261 31912
tri 26029 31910 26030 31911 ne
rect 26030 31910 26261 31911
tri 26261 31910 26306 31955 sw
rect 70802 31948 71000 32006
tri 26030 31909 26031 31910 ne
rect 26031 31909 26306 31910
tri 26031 31908 26032 31909 ne
rect 26032 31908 26306 31909
tri 26032 31907 26033 31908 ne
rect 26033 31907 26306 31908
tri 26033 31906 26034 31907 ne
rect 26034 31906 26306 31907
tri 26034 31905 26035 31906 ne
rect 26035 31905 26306 31906
tri 26035 31904 26036 31905 ne
rect 26036 31904 26306 31905
tri 26036 31903 26037 31904 ne
rect 26037 31903 26306 31904
tri 26037 31902 26038 31903 ne
rect 26038 31902 26306 31903
tri 26038 31901 26039 31902 ne
rect 26039 31901 26306 31902
tri 26039 31900 26040 31901 ne
rect 26040 31900 26306 31901
tri 26040 31899 26041 31900 ne
rect 26041 31899 26306 31900
tri 26041 31898 26042 31899 ne
rect 26042 31898 26306 31899
tri 26042 31897 26043 31898 ne
rect 26043 31897 26306 31898
tri 26043 31896 26044 31897 ne
rect 26044 31896 26306 31897
tri 26044 31895 26045 31896 ne
rect 26045 31895 26306 31896
tri 26045 31894 26046 31895 ne
rect 26046 31894 26306 31895
tri 26046 31893 26047 31894 ne
rect 26047 31893 26306 31894
tri 26047 31892 26048 31893 ne
rect 26048 31892 26306 31893
tri 26048 31891 26049 31892 ne
rect 26049 31891 26306 31892
tri 26049 31890 26050 31891 ne
rect 26050 31890 26306 31891
tri 26050 31889 26051 31890 ne
rect 26051 31889 26306 31890
tri 26051 31888 26052 31889 ne
rect 26052 31888 26306 31889
tri 26052 31887 26053 31888 ne
rect 26053 31887 26190 31888
tri 26053 31886 26054 31887 ne
rect 26054 31886 26190 31887
tri 26054 31885 26055 31886 ne
rect 26055 31885 26190 31886
tri 26055 31884 26056 31885 ne
rect 26056 31884 26190 31885
tri 26056 31883 26057 31884 ne
rect 26057 31883 26190 31884
tri 26057 31882 26058 31883 ne
rect 26058 31882 26190 31883
tri 26058 31881 26059 31882 ne
rect 26059 31881 26190 31882
tri 26059 31880 26060 31881 ne
rect 26060 31880 26190 31881
tri 26060 31879 26061 31880 ne
rect 26061 31879 26190 31880
tri 26061 31878 26062 31879 ne
rect 26062 31878 26190 31879
tri 26062 31877 26063 31878 ne
rect 26063 31877 26190 31878
tri 26063 31876 26064 31877 ne
rect 26064 31876 26190 31877
tri 26064 31875 26065 31876 ne
rect 26065 31875 26190 31876
tri 26065 31874 26066 31875 ne
rect 26066 31874 26190 31875
tri 26066 31873 26067 31874 ne
rect 26067 31873 26190 31874
tri 26067 31872 26068 31873 ne
rect 26068 31872 26190 31873
tri 26068 31871 26069 31872 ne
rect 26069 31871 26190 31872
tri 26069 31870 26070 31871 ne
rect 26070 31870 26190 31871
tri 26070 31869 26071 31870 ne
rect 26071 31869 26190 31870
tri 26071 31868 26072 31869 ne
rect 26072 31868 26190 31869
tri 26072 31867 26073 31868 ne
rect 26073 31867 26190 31868
tri 26073 31866 26074 31867 ne
rect 26074 31866 26190 31867
tri 26074 31865 26075 31866 ne
rect 26075 31865 26190 31866
tri 26075 31820 26120 31865 ne
rect 26120 31842 26190 31865
rect 26236 31865 26306 31888
tri 26306 31865 26351 31910 sw
rect 70802 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26236 31842 26351 31865
rect 26120 31820 26351 31842
tri 26351 31820 26396 31865 sw
rect 70802 31844 71000 31902
tri 26120 31776 26164 31820 ne
rect 26164 31776 26396 31820
tri 26396 31776 26440 31820 sw
rect 70802 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
tri 26164 31775 26165 31776 ne
rect 26165 31775 26440 31776
tri 26165 31731 26209 31775 ne
rect 26209 31756 26440 31775
rect 26209 31731 26322 31756
tri 26209 31686 26254 31731 ne
rect 26254 31710 26322 31731
rect 26368 31731 26440 31756
tri 26440 31731 26485 31776 sw
rect 70802 31740 71000 31798
rect 26368 31710 26485 31731
rect 26254 31686 26485 31710
tri 26485 31686 26530 31731 sw
rect 70802 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
tri 26254 31676 26264 31686 ne
rect 26264 31676 26530 31686
tri 26264 31675 26265 31676 ne
rect 26265 31675 26530 31676
tri 26265 31674 26266 31675 ne
rect 26266 31674 26530 31675
tri 26266 31673 26267 31674 ne
rect 26267 31673 26530 31674
tri 26267 31672 26268 31673 ne
rect 26268 31672 26530 31673
tri 26268 31671 26269 31672 ne
rect 26269 31671 26530 31672
tri 26269 31670 26270 31671 ne
rect 26270 31670 26530 31671
tri 26270 31669 26271 31670 ne
rect 26271 31669 26530 31670
tri 26271 31668 26272 31669 ne
rect 26272 31668 26530 31669
tri 26272 31667 26273 31668 ne
rect 26273 31667 26530 31668
tri 26273 31666 26274 31667 ne
rect 26274 31666 26530 31667
tri 26274 31665 26275 31666 ne
rect 26275 31665 26530 31666
tri 26275 31664 26276 31665 ne
rect 26276 31664 26530 31665
tri 26276 31663 26277 31664 ne
rect 26277 31663 26530 31664
tri 26277 31662 26278 31663 ne
rect 26278 31662 26530 31663
tri 26278 31661 26279 31662 ne
rect 26279 31661 26530 31662
tri 26279 31660 26280 31661 ne
rect 26280 31660 26530 31661
tri 26280 31659 26281 31660 ne
rect 26281 31659 26530 31660
tri 26281 31658 26282 31659 ne
rect 26282 31658 26530 31659
tri 26282 31657 26283 31658 ne
rect 26283 31657 26530 31658
tri 26283 31656 26284 31657 ne
rect 26284 31656 26530 31657
tri 26284 31655 26285 31656 ne
rect 26285 31655 26530 31656
tri 26285 31654 26286 31655 ne
rect 26286 31654 26530 31655
tri 26286 31653 26287 31654 ne
rect 26287 31653 26530 31654
tri 26287 31652 26288 31653 ne
rect 26288 31652 26530 31653
tri 26288 31651 26289 31652 ne
rect 26289 31651 26530 31652
tri 26289 31650 26290 31651 ne
rect 26290 31650 26530 31651
tri 26290 31649 26291 31650 ne
rect 26291 31649 26530 31650
tri 26291 31648 26292 31649 ne
rect 26292 31648 26530 31649
tri 26292 31647 26293 31648 ne
rect 26293 31647 26530 31648
tri 26293 31646 26294 31647 ne
rect 26294 31646 26530 31647
tri 26294 31645 26295 31646 ne
rect 26295 31645 26530 31646
tri 26295 31644 26296 31645 ne
rect 26296 31644 26530 31645
tri 26296 31643 26297 31644 ne
rect 26297 31643 26530 31644
tri 26297 31642 26298 31643 ne
rect 26298 31642 26530 31643
tri 26298 31641 26299 31642 ne
rect 26299 31641 26530 31642
tri 26530 31641 26575 31686 sw
tri 26299 31640 26300 31641 ne
rect 26300 31640 26575 31641
tri 26300 31639 26301 31640 ne
rect 26301 31639 26575 31640
tri 26301 31638 26302 31639 ne
rect 26302 31638 26575 31639
tri 26302 31637 26303 31638 ne
rect 26303 31637 26575 31638
tri 26303 31636 26304 31637 ne
rect 26304 31636 26575 31637
tri 26304 31635 26305 31636 ne
rect 26305 31635 26575 31636
tri 26305 31634 26306 31635 ne
rect 26306 31634 26575 31635
tri 26575 31634 26582 31641 sw
rect 70802 31636 71000 31694
tri 26306 31633 26307 31634 ne
rect 26307 31633 26582 31634
tri 26307 31632 26308 31633 ne
rect 26308 31632 26582 31633
tri 26308 31631 26309 31632 ne
rect 26309 31631 26582 31632
tri 26309 31630 26310 31631 ne
rect 26310 31630 26582 31631
tri 26310 31629 26311 31630 ne
rect 26311 31629 26582 31630
tri 26311 31628 26312 31629 ne
rect 26312 31628 26582 31629
tri 26312 31627 26313 31628 ne
rect 26313 31627 26582 31628
tri 26313 31626 26314 31627 ne
rect 26314 31626 26582 31627
tri 26314 31625 26315 31626 ne
rect 26315 31625 26582 31626
tri 26315 31624 26316 31625 ne
rect 26316 31624 26582 31625
tri 26316 31623 26317 31624 ne
rect 26317 31623 26454 31624
tri 26317 31622 26318 31623 ne
rect 26318 31622 26454 31623
tri 26318 31621 26319 31622 ne
rect 26319 31621 26454 31622
tri 26319 31620 26320 31621 ne
rect 26320 31620 26454 31621
tri 26320 31619 26321 31620 ne
rect 26321 31619 26454 31620
tri 26321 31618 26322 31619 ne
rect 26322 31618 26454 31619
tri 26322 31617 26323 31618 ne
rect 26323 31617 26454 31618
tri 26323 31616 26324 31617 ne
rect 26324 31616 26454 31617
tri 26324 31615 26325 31616 ne
rect 26325 31615 26454 31616
tri 26325 31614 26326 31615 ne
rect 26326 31614 26454 31615
tri 26326 31613 26327 31614 ne
rect 26327 31613 26454 31614
tri 26327 31612 26328 31613 ne
rect 26328 31612 26454 31613
tri 26328 31611 26329 31612 ne
rect 26329 31611 26454 31612
tri 26329 31610 26330 31611 ne
rect 26330 31610 26454 31611
tri 26330 31609 26331 31610 ne
rect 26331 31609 26454 31610
tri 26331 31608 26332 31609 ne
rect 26332 31608 26454 31609
tri 26332 31607 26333 31608 ne
rect 26333 31607 26454 31608
tri 26333 31606 26334 31607 ne
rect 26334 31606 26454 31607
tri 26334 31605 26335 31606 ne
rect 26335 31605 26454 31606
tri 26335 31604 26336 31605 ne
rect 26336 31604 26454 31605
tri 26336 31603 26337 31604 ne
rect 26337 31603 26454 31604
tri 26337 31602 26338 31603 ne
rect 26338 31602 26454 31603
tri 26338 31601 26339 31602 ne
rect 26339 31601 26454 31602
tri 26339 31600 26340 31601 ne
rect 26340 31600 26454 31601
tri 26340 31599 26341 31600 ne
rect 26341 31599 26454 31600
tri 26341 31598 26342 31599 ne
rect 26342 31598 26454 31599
tri 26342 31597 26343 31598 ne
rect 26343 31597 26454 31598
tri 26343 31596 26344 31597 ne
rect 26344 31596 26454 31597
tri 26344 31595 26345 31596 ne
rect 26345 31595 26454 31596
tri 26345 31594 26346 31595 ne
rect 26346 31594 26454 31595
tri 26346 31593 26347 31594 ne
rect 26347 31593 26454 31594
tri 26347 31592 26348 31593 ne
rect 26348 31592 26454 31593
tri 26348 31591 26349 31592 ne
rect 26349 31591 26454 31592
tri 26349 31590 26350 31591 ne
rect 26350 31590 26454 31591
tri 26350 31589 26351 31590 ne
rect 26351 31589 26454 31590
tri 26351 31544 26396 31589 ne
rect 26396 31578 26454 31589
rect 26500 31589 26582 31624
tri 26582 31589 26627 31634 sw
rect 70802 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 26500 31578 26627 31589
rect 26396 31544 26627 31578
tri 26627 31544 26672 31589 sw
tri 26396 31499 26441 31544 ne
rect 26441 31499 26672 31544
tri 26672 31499 26717 31544 sw
rect 70802 31532 71000 31590
tri 26441 31454 26486 31499 ne
rect 26486 31492 26717 31499
rect 26486 31454 26586 31492
tri 26486 31410 26530 31454 ne
rect 26530 31446 26586 31454
rect 26632 31455 26717 31492
tri 26717 31455 26761 31499 sw
rect 70802 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31446 26761 31455
rect 26530 31410 26761 31446
tri 26761 31410 26806 31455 sw
rect 70802 31428 71000 31486
tri 26530 31409 26531 31410 ne
rect 26531 31409 26806 31410
tri 26531 31401 26539 31409 ne
rect 26539 31401 26806 31409
tri 26539 31400 26540 31401 ne
rect 26540 31400 26806 31401
tri 26540 31399 26541 31400 ne
rect 26541 31399 26806 31400
tri 26541 31398 26542 31399 ne
rect 26542 31398 26806 31399
tri 26542 31397 26543 31398 ne
rect 26543 31397 26806 31398
tri 26543 31396 26544 31397 ne
rect 26544 31396 26806 31397
tri 26544 31395 26545 31396 ne
rect 26545 31395 26806 31396
tri 26545 31394 26546 31395 ne
rect 26546 31394 26806 31395
tri 26546 31393 26547 31394 ne
rect 26547 31393 26806 31394
tri 26547 31392 26548 31393 ne
rect 26548 31392 26806 31393
tri 26548 31391 26549 31392 ne
rect 26549 31391 26806 31392
tri 26549 31390 26550 31391 ne
rect 26550 31390 26806 31391
tri 26550 31389 26551 31390 ne
rect 26551 31389 26806 31390
tri 26551 31388 26552 31389 ne
rect 26552 31388 26806 31389
tri 26552 31387 26553 31388 ne
rect 26553 31387 26806 31388
tri 26553 31386 26554 31387 ne
rect 26554 31386 26806 31387
tri 26554 31385 26555 31386 ne
rect 26555 31385 26806 31386
tri 26555 31384 26556 31385 ne
rect 26556 31384 26806 31385
tri 26556 31383 26557 31384 ne
rect 26557 31383 26806 31384
tri 26557 31382 26558 31383 ne
rect 26558 31382 26806 31383
tri 26558 31381 26559 31382 ne
rect 26559 31381 26806 31382
tri 26559 31380 26560 31381 ne
rect 26560 31380 26806 31381
tri 26560 31379 26561 31380 ne
rect 26561 31379 26806 31380
tri 26561 31378 26562 31379 ne
rect 26562 31378 26806 31379
tri 26562 31377 26563 31378 ne
rect 26563 31377 26806 31378
tri 26563 31376 26564 31377 ne
rect 26564 31376 26806 31377
tri 26564 31375 26565 31376 ne
rect 26565 31375 26806 31376
tri 26565 31374 26566 31375 ne
rect 26566 31374 26806 31375
tri 26566 31373 26567 31374 ne
rect 26567 31373 26806 31374
tri 26567 31372 26568 31373 ne
rect 26568 31372 26806 31373
tri 26568 31371 26569 31372 ne
rect 26569 31371 26806 31372
tri 26569 31370 26570 31371 ne
rect 26570 31370 26806 31371
tri 26570 31369 26571 31370 ne
rect 26571 31369 26806 31370
tri 26571 31368 26572 31369 ne
rect 26572 31368 26806 31369
tri 26572 31367 26573 31368 ne
rect 26573 31367 26806 31368
tri 26573 31366 26574 31367 ne
rect 26574 31366 26806 31367
tri 26574 31365 26575 31366 ne
rect 26575 31365 26806 31366
tri 26806 31365 26851 31410 sw
rect 70802 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
tri 26575 31364 26576 31365 ne
rect 26576 31364 26851 31365
tri 26576 31363 26577 31364 ne
rect 26577 31363 26851 31364
tri 26577 31362 26578 31363 ne
rect 26578 31362 26851 31363
tri 26578 31361 26579 31362 ne
rect 26579 31361 26851 31362
tri 26579 31360 26580 31361 ne
rect 26580 31360 26851 31361
tri 26580 31359 26581 31360 ne
rect 26581 31359 26718 31360
tri 26581 31358 26582 31359 ne
rect 26582 31358 26718 31359
tri 26582 31357 26583 31358 ne
rect 26583 31357 26718 31358
tri 26583 31356 26584 31357 ne
rect 26584 31356 26718 31357
tri 26584 31355 26585 31356 ne
rect 26585 31355 26718 31356
tri 26585 31354 26586 31355 ne
rect 26586 31354 26718 31355
tri 26586 31353 26587 31354 ne
rect 26587 31353 26718 31354
tri 26587 31352 26588 31353 ne
rect 26588 31352 26718 31353
tri 26588 31351 26589 31352 ne
rect 26589 31351 26718 31352
tri 26589 31350 26590 31351 ne
rect 26590 31350 26718 31351
tri 26590 31349 26591 31350 ne
rect 26591 31349 26718 31350
tri 26591 31348 26592 31349 ne
rect 26592 31348 26718 31349
tri 26592 31347 26593 31348 ne
rect 26593 31347 26718 31348
tri 26593 31346 26594 31347 ne
rect 26594 31346 26718 31347
tri 26594 31345 26595 31346 ne
rect 26595 31345 26718 31346
tri 26595 31344 26596 31345 ne
rect 26596 31344 26718 31345
tri 26596 31343 26597 31344 ne
rect 26597 31343 26718 31344
tri 26597 31342 26598 31343 ne
rect 26598 31342 26718 31343
tri 26598 31341 26599 31342 ne
rect 26599 31341 26718 31342
tri 26599 31340 26600 31341 ne
rect 26600 31340 26718 31341
tri 26600 31339 26601 31340 ne
rect 26601 31339 26718 31340
tri 26601 31338 26602 31339 ne
rect 26602 31338 26718 31339
tri 26602 31337 26603 31338 ne
rect 26603 31337 26718 31338
tri 26603 31336 26604 31337 ne
rect 26604 31336 26718 31337
tri 26604 31335 26605 31336 ne
rect 26605 31335 26718 31336
tri 26605 31334 26606 31335 ne
rect 26606 31334 26718 31335
tri 26606 31333 26607 31334 ne
rect 26607 31333 26718 31334
tri 26607 31332 26608 31333 ne
rect 26608 31332 26718 31333
tri 26608 31331 26609 31332 ne
rect 26609 31331 26718 31332
tri 26609 31330 26610 31331 ne
rect 26610 31330 26718 31331
tri 26610 31329 26611 31330 ne
rect 26611 31329 26718 31330
tri 26611 31328 26612 31329 ne
rect 26612 31328 26718 31329
tri 26612 31327 26613 31328 ne
rect 26613 31327 26718 31328
tri 26613 31326 26614 31327 ne
rect 26614 31326 26718 31327
tri 26614 31325 26615 31326 ne
rect 26615 31325 26718 31326
tri 26615 31324 26616 31325 ne
rect 26616 31324 26718 31325
tri 26616 31323 26617 31324 ne
rect 26617 31323 26718 31324
tri 26617 31322 26618 31323 ne
rect 26618 31322 26718 31323
tri 26618 31321 26619 31322 ne
rect 26619 31321 26718 31322
tri 26619 31320 26620 31321 ne
rect 26620 31320 26718 31321
tri 26620 31319 26621 31320 ne
rect 26621 31319 26718 31320
tri 26621 31318 26622 31319 ne
rect 26622 31318 26718 31319
tri 26622 31317 26623 31318 ne
rect 26623 31317 26718 31318
tri 26623 31316 26624 31317 ne
rect 26624 31316 26718 31317
tri 26624 31315 26625 31316 ne
rect 26625 31315 26718 31316
tri 26625 31314 26626 31315 ne
rect 26626 31314 26718 31315
rect 26764 31320 26851 31360
tri 26851 31320 26896 31365 sw
rect 70802 31324 71000 31382
rect 26764 31314 26896 31320
tri 26626 31313 26627 31314 ne
rect 26627 31313 26896 31314
tri 26896 31313 26903 31320 sw
tri 26627 31268 26672 31313 ne
rect 26672 31268 26903 31313
tri 26903 31268 26948 31313 sw
rect 70802 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
tri 26672 31243 26697 31268 ne
rect 26697 31243 26948 31268
tri 26697 31198 26742 31243 ne
rect 26742 31228 26948 31243
rect 26742 31198 26850 31228
tri 26742 31153 26787 31198 ne
rect 26787 31182 26850 31198
rect 26896 31223 26948 31228
tri 26948 31223 26993 31268 sw
rect 26896 31182 26993 31223
rect 26787 31178 26993 31182
tri 26993 31178 27038 31223 sw
rect 70802 31220 71000 31278
rect 26787 31172 27038 31178
tri 27038 31172 27044 31178 sw
rect 70802 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 26787 31153 27044 31172
tri 26787 31127 26813 31153 ne
rect 26813 31127 27044 31153
tri 27044 31127 27089 31172 sw
tri 26813 31126 26814 31127 ne
rect 26814 31126 27089 31127
tri 26814 31125 26815 31126 ne
rect 26815 31125 27089 31126
tri 26815 31124 26816 31125 ne
rect 26816 31124 27089 31125
tri 26816 31123 26817 31124 ne
rect 26817 31123 27089 31124
tri 26817 31122 26818 31123 ne
rect 26818 31122 27089 31123
tri 26818 31121 26819 31122 ne
rect 26819 31121 27089 31122
tri 26819 31120 26820 31121 ne
rect 26820 31120 27089 31121
tri 26820 31119 26821 31120 ne
rect 26821 31119 27089 31120
tri 26821 31118 26822 31119 ne
rect 26822 31118 27089 31119
tri 26822 31117 26823 31118 ne
rect 26823 31117 27089 31118
tri 26823 31116 26824 31117 ne
rect 26824 31116 27089 31117
tri 26824 31115 26825 31116 ne
rect 26825 31115 27089 31116
tri 26825 31114 26826 31115 ne
rect 26826 31114 27089 31115
tri 26826 31113 26827 31114 ne
rect 26827 31113 27089 31114
tri 26827 31112 26828 31113 ne
rect 26828 31112 27089 31113
tri 26828 31111 26829 31112 ne
rect 26829 31111 27089 31112
tri 26829 31110 26830 31111 ne
rect 26830 31110 27089 31111
tri 26830 31109 26831 31110 ne
rect 26831 31109 27089 31110
tri 26831 31108 26832 31109 ne
rect 26832 31108 27089 31109
tri 26832 31107 26833 31108 ne
rect 26833 31107 27089 31108
tri 26833 31106 26834 31107 ne
rect 26834 31106 27089 31107
tri 26834 31105 26835 31106 ne
rect 26835 31105 27089 31106
tri 26835 31104 26836 31105 ne
rect 26836 31104 27089 31105
tri 26836 31103 26837 31104 ne
rect 26837 31103 27089 31104
tri 26837 31102 26838 31103 ne
rect 26838 31102 27089 31103
tri 26838 31101 26839 31102 ne
rect 26839 31101 27089 31102
tri 26839 31100 26840 31101 ne
rect 26840 31100 27089 31101
tri 26840 31099 26841 31100 ne
rect 26841 31099 27089 31100
tri 26841 31098 26842 31099 ne
rect 26842 31098 27089 31099
tri 26842 31097 26843 31098 ne
rect 26843 31097 27089 31098
tri 26843 31096 26844 31097 ne
rect 26844 31096 27089 31097
tri 26844 31095 26845 31096 ne
rect 26845 31095 26982 31096
tri 26845 31094 26846 31095 ne
rect 26846 31094 26982 31095
tri 26846 31093 26847 31094 ne
rect 26847 31093 26982 31094
tri 26847 31092 26848 31093 ne
rect 26848 31092 26982 31093
tri 26848 31091 26849 31092 ne
rect 26849 31091 26982 31092
tri 26849 31090 26850 31091 ne
rect 26850 31090 26982 31091
tri 26850 31089 26851 31090 ne
rect 26851 31089 26982 31090
tri 26851 31088 26852 31089 ne
rect 26852 31088 26982 31089
tri 26852 31087 26853 31088 ne
rect 26853 31087 26982 31088
tri 26853 31086 26854 31087 ne
rect 26854 31086 26982 31087
tri 26854 31085 26855 31086 ne
rect 26855 31085 26982 31086
tri 26855 31084 26856 31085 ne
rect 26856 31084 26982 31085
tri 26856 31083 26857 31084 ne
rect 26857 31083 26982 31084
tri 26857 31082 26858 31083 ne
rect 26858 31082 26982 31083
tri 26858 31081 26859 31082 ne
rect 26859 31081 26982 31082
tri 26859 31080 26860 31081 ne
rect 26860 31080 26982 31081
tri 26860 31079 26861 31080 ne
rect 26861 31079 26982 31080
tri 26861 31078 26862 31079 ne
rect 26862 31078 26982 31079
tri 26862 31077 26863 31078 ne
rect 26863 31077 26982 31078
tri 26863 31076 26864 31077 ne
rect 26864 31076 26982 31077
tri 26864 31075 26865 31076 ne
rect 26865 31075 26982 31076
tri 26865 31074 26866 31075 ne
rect 26866 31074 26982 31075
tri 26866 31073 26867 31074 ne
rect 26867 31073 26982 31074
tri 26867 31072 26868 31073 ne
rect 26868 31072 26982 31073
tri 26868 31071 26869 31072 ne
rect 26869 31071 26982 31072
tri 26869 31070 26870 31071 ne
rect 26870 31070 26982 31071
tri 26870 31069 26871 31070 ne
rect 26871 31069 26982 31070
tri 26871 31068 26872 31069 ne
rect 26872 31068 26982 31069
tri 26872 31067 26873 31068 ne
rect 26873 31067 26982 31068
tri 26873 31066 26874 31067 ne
rect 26874 31066 26982 31067
tri 26874 31065 26875 31066 ne
rect 26875 31065 26982 31066
tri 26875 31064 26876 31065 ne
rect 26876 31064 26982 31065
tri 26876 31063 26877 31064 ne
rect 26877 31063 26982 31064
tri 26877 31062 26878 31063 ne
rect 26878 31062 26982 31063
tri 26878 31061 26879 31062 ne
rect 26879 31061 26982 31062
tri 26879 31060 26880 31061 ne
rect 26880 31060 26982 31061
tri 26880 31059 26881 31060 ne
rect 26881 31059 26982 31060
tri 26881 31058 26882 31059 ne
rect 26882 31058 26982 31059
tri 26882 31057 26883 31058 ne
rect 26883 31057 26982 31058
tri 26883 31056 26884 31057 ne
rect 26884 31056 26982 31057
tri 26884 31055 26885 31056 ne
rect 26885 31055 26982 31056
tri 26885 31054 26886 31055 ne
rect 26886 31054 26982 31055
tri 26886 31053 26887 31054 ne
rect 26887 31053 26982 31054
tri 26887 31052 26888 31053 ne
rect 26888 31052 26982 31053
tri 26888 31051 26889 31052 ne
rect 26889 31051 26982 31052
tri 26889 31050 26890 31051 ne
rect 26890 31050 26982 31051
rect 27028 31082 27089 31096
tri 27089 31082 27134 31127 sw
rect 70802 31116 71000 31174
rect 27028 31050 27134 31082
tri 26890 31049 26891 31050 ne
rect 26891 31049 27134 31050
tri 26891 31048 26892 31049 ne
rect 26892 31048 27134 31049
tri 26892 31047 26893 31048 ne
rect 26893 31047 27134 31048
tri 26893 31046 26894 31047 ne
rect 26894 31046 27134 31047
tri 26894 31045 26895 31046 ne
rect 26895 31045 27134 31046
tri 26895 31044 26896 31045 ne
rect 26896 31044 27134 31045
tri 26896 31043 26897 31044 ne
rect 26897 31043 27134 31044
tri 26897 31042 26898 31043 ne
rect 26898 31042 27134 31043
tri 26898 31041 26899 31042 ne
rect 26899 31041 27134 31042
tri 26899 31040 26900 31041 ne
rect 26900 31040 27134 31041
tri 26900 31039 26901 31040 ne
rect 26901 31039 27134 31040
tri 26901 31038 26902 31039 ne
rect 26902 31038 27134 31039
tri 26902 31037 26903 31038 ne
rect 26903 31037 27134 31038
tri 27134 31037 27179 31082 sw
rect 70802 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
tri 26903 30999 26941 31037 ne
rect 26941 30999 27179 31037
tri 27179 30999 27217 31037 sw
rect 70802 31012 71000 31070
tri 26941 30954 26986 30999 ne
rect 26986 30964 27217 30999
rect 26986 30954 27114 30964
tri 26986 30923 27017 30954 ne
rect 27017 30923 27114 30954
tri 27017 30878 27062 30923 ne
rect 27062 30918 27114 30923
rect 27160 30954 27217 30964
tri 27217 30954 27262 30999 sw
rect 70802 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 27160 30918 27262 30954
rect 27062 30909 27262 30918
tri 27262 30909 27307 30954 sw
rect 27062 30878 27307 30909
tri 27062 30853 27087 30878 ne
rect 27087 30864 27307 30878
tri 27307 30864 27352 30909 sw
rect 70802 30908 71000 30966
rect 27087 30853 27352 30864
tri 27087 30852 27088 30853 ne
rect 27088 30852 27352 30853
tri 27088 30851 27089 30852 ne
rect 27089 30851 27352 30852
tri 27352 30851 27365 30864 sw
rect 70802 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
tri 27089 30850 27090 30851 ne
rect 27090 30850 27365 30851
tri 27090 30849 27091 30850 ne
rect 27091 30849 27365 30850
tri 27091 30848 27092 30849 ne
rect 27092 30848 27365 30849
tri 27092 30847 27093 30848 ne
rect 27093 30847 27365 30848
tri 27093 30846 27094 30847 ne
rect 27094 30846 27365 30847
tri 27094 30845 27095 30846 ne
rect 27095 30845 27365 30846
tri 27095 30844 27096 30845 ne
rect 27096 30844 27365 30845
tri 27096 30843 27097 30844 ne
rect 27097 30843 27365 30844
tri 27097 30842 27098 30843 ne
rect 27098 30842 27365 30843
tri 27098 30841 27099 30842 ne
rect 27099 30841 27365 30842
tri 27099 30840 27100 30841 ne
rect 27100 30840 27365 30841
tri 27100 30839 27101 30840 ne
rect 27101 30839 27365 30840
tri 27101 30838 27102 30839 ne
rect 27102 30838 27365 30839
tri 27102 30837 27103 30838 ne
rect 27103 30837 27365 30838
tri 27103 30836 27104 30837 ne
rect 27104 30836 27365 30837
tri 27104 30835 27105 30836 ne
rect 27105 30835 27365 30836
tri 27105 30834 27106 30835 ne
rect 27106 30834 27365 30835
tri 27106 30833 27107 30834 ne
rect 27107 30833 27365 30834
tri 27107 30832 27108 30833 ne
rect 27108 30832 27365 30833
tri 27108 30831 27109 30832 ne
rect 27109 30831 27246 30832
tri 27109 30830 27110 30831 ne
rect 27110 30830 27246 30831
tri 27110 30829 27111 30830 ne
rect 27111 30829 27246 30830
tri 27111 30828 27112 30829 ne
rect 27112 30828 27246 30829
tri 27112 30827 27113 30828 ne
rect 27113 30827 27246 30828
tri 27113 30826 27114 30827 ne
rect 27114 30826 27246 30827
tri 27114 30825 27115 30826 ne
rect 27115 30825 27246 30826
tri 27115 30824 27116 30825 ne
rect 27116 30824 27246 30825
tri 27116 30823 27117 30824 ne
rect 27117 30823 27246 30824
tri 27117 30822 27118 30823 ne
rect 27118 30822 27246 30823
tri 27118 30821 27119 30822 ne
rect 27119 30821 27246 30822
tri 27119 30820 27120 30821 ne
rect 27120 30820 27246 30821
tri 27120 30819 27121 30820 ne
rect 27121 30819 27246 30820
tri 27121 30818 27122 30819 ne
rect 27122 30818 27246 30819
tri 27122 30817 27123 30818 ne
rect 27123 30817 27246 30818
tri 27123 30816 27124 30817 ne
rect 27124 30816 27246 30817
tri 27124 30815 27125 30816 ne
rect 27125 30815 27246 30816
tri 27125 30814 27126 30815 ne
rect 27126 30814 27246 30815
tri 27126 30813 27127 30814 ne
rect 27127 30813 27246 30814
tri 27127 30812 27128 30813 ne
rect 27128 30812 27246 30813
tri 27128 30811 27129 30812 ne
rect 27129 30811 27246 30812
tri 27129 30810 27130 30811 ne
rect 27130 30810 27246 30811
tri 27130 30809 27131 30810 ne
rect 27131 30809 27246 30810
tri 27131 30808 27132 30809 ne
rect 27132 30808 27246 30809
tri 27132 30807 27133 30808 ne
rect 27133 30807 27246 30808
tri 27133 30806 27134 30807 ne
rect 27134 30806 27246 30807
tri 27134 30805 27135 30806 ne
rect 27135 30805 27246 30806
tri 27135 30804 27136 30805 ne
rect 27136 30804 27246 30805
tri 27136 30803 27137 30804 ne
rect 27137 30803 27246 30804
tri 27137 30802 27138 30803 ne
rect 27138 30802 27246 30803
tri 27138 30801 27139 30802 ne
rect 27139 30801 27246 30802
tri 27139 30800 27140 30801 ne
rect 27140 30800 27246 30801
tri 27140 30799 27141 30800 ne
rect 27141 30799 27246 30800
tri 27141 30798 27142 30799 ne
rect 27142 30798 27246 30799
tri 27142 30797 27143 30798 ne
rect 27143 30797 27246 30798
tri 27143 30796 27144 30797 ne
rect 27144 30796 27246 30797
tri 27144 30795 27145 30796 ne
rect 27145 30795 27246 30796
tri 27145 30794 27146 30795 ne
rect 27146 30794 27246 30795
tri 27146 30793 27147 30794 ne
rect 27147 30793 27246 30794
tri 27147 30792 27148 30793 ne
rect 27148 30792 27246 30793
tri 27148 30791 27149 30792 ne
rect 27149 30791 27246 30792
tri 27149 30790 27150 30791 ne
rect 27150 30790 27246 30791
tri 27150 30789 27151 30790 ne
rect 27151 30789 27246 30790
tri 27151 30788 27152 30789 ne
rect 27152 30788 27246 30789
tri 27152 30787 27153 30788 ne
rect 27153 30787 27246 30788
tri 27153 30786 27154 30787 ne
rect 27154 30786 27246 30787
rect 27292 30806 27365 30832
tri 27365 30806 27410 30851 sw
rect 27292 30786 27410 30806
tri 27154 30785 27155 30786 ne
rect 27155 30785 27410 30786
tri 27155 30784 27156 30785 ne
rect 27156 30784 27410 30785
tri 27156 30783 27157 30784 ne
rect 27157 30783 27410 30784
tri 27157 30782 27158 30783 ne
rect 27158 30782 27410 30783
tri 27158 30781 27159 30782 ne
rect 27159 30781 27410 30782
tri 27159 30780 27160 30781 ne
rect 27160 30780 27410 30781
tri 27160 30779 27161 30780 ne
rect 27161 30779 27410 30780
tri 27161 30778 27162 30779 ne
rect 27162 30778 27410 30779
tri 27162 30777 27163 30778 ne
rect 27163 30777 27410 30778
tri 27163 30776 27164 30777 ne
rect 27164 30776 27410 30777
tri 27164 30775 27165 30776 ne
rect 27165 30775 27410 30776
tri 27165 30774 27166 30775 ne
rect 27166 30774 27410 30775
tri 27166 30773 27167 30774 ne
rect 27167 30773 27410 30774
tri 27167 30772 27168 30773 ne
rect 27168 30772 27410 30773
tri 27168 30771 27169 30772 ne
rect 27169 30771 27410 30772
tri 27169 30770 27170 30771 ne
rect 27170 30770 27410 30771
tri 27170 30769 27171 30770 ne
rect 27171 30769 27410 30770
tri 27171 30768 27172 30769 ne
rect 27172 30768 27410 30769
tri 27172 30767 27173 30768 ne
rect 27173 30767 27410 30768
tri 27173 30766 27174 30767 ne
rect 27174 30766 27410 30767
tri 27174 30765 27175 30766 ne
rect 27175 30765 27410 30766
tri 27175 30764 27176 30765 ne
rect 27176 30764 27410 30765
tri 27176 30763 27177 30764 ne
rect 27177 30763 27410 30764
tri 27177 30762 27178 30763 ne
rect 27178 30762 27410 30763
tri 27178 30761 27179 30762 ne
rect 27179 30761 27410 30762
tri 27410 30761 27455 30806 sw
rect 70802 30804 71000 30862
tri 27179 30716 27224 30761 ne
rect 27224 30716 27455 30761
tri 27455 30716 27500 30761 sw
rect 70802 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27224 30678 27262 30716 ne
rect 27262 30700 27500 30716
rect 27262 30678 27378 30700
tri 27262 30671 27269 30678 ne
rect 27269 30671 27378 30678
tri 27269 30633 27307 30671 ne
rect 27307 30654 27378 30671
rect 27424 30678 27500 30700
tri 27500 30678 27538 30716 sw
rect 70802 30700 71000 30758
rect 27424 30654 27538 30678
rect 27307 30633 27538 30654
tri 27538 30633 27583 30678 sw
rect 70802 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
tri 27307 30588 27352 30633 ne
rect 27352 30588 27583 30633
tri 27583 30588 27628 30633 sw
rect 70802 30596 71000 30654
tri 27352 30578 27362 30588 ne
rect 27362 30578 27628 30588
tri 27362 30577 27363 30578 ne
rect 27363 30577 27628 30578
tri 27363 30576 27364 30577 ne
rect 27364 30576 27628 30577
tri 27364 30575 27365 30576 ne
rect 27365 30575 27628 30576
tri 27365 30574 27366 30575 ne
rect 27366 30574 27628 30575
tri 27366 30573 27367 30574 ne
rect 27367 30573 27628 30574
tri 27367 30572 27368 30573 ne
rect 27368 30572 27628 30573
tri 27368 30571 27369 30572 ne
rect 27369 30571 27628 30572
tri 27369 30570 27370 30571 ne
rect 27370 30570 27628 30571
tri 27370 30569 27371 30570 ne
rect 27371 30569 27628 30570
tri 27371 30568 27372 30569 ne
rect 27372 30568 27628 30569
tri 27372 30567 27373 30568 ne
rect 27373 30567 27510 30568
tri 27373 30566 27374 30567 ne
rect 27374 30566 27510 30567
tri 27374 30565 27375 30566 ne
rect 27375 30565 27510 30566
tri 27375 30564 27376 30565 ne
rect 27376 30564 27510 30565
tri 27376 30563 27377 30564 ne
rect 27377 30563 27510 30564
tri 27377 30562 27378 30563 ne
rect 27378 30562 27510 30563
tri 27378 30561 27379 30562 ne
rect 27379 30561 27510 30562
tri 27379 30560 27380 30561 ne
rect 27380 30560 27510 30561
tri 27380 30559 27381 30560 ne
rect 27381 30559 27510 30560
tri 27381 30558 27382 30559 ne
rect 27382 30558 27510 30559
tri 27382 30557 27383 30558 ne
rect 27383 30557 27510 30558
tri 27383 30556 27384 30557 ne
rect 27384 30556 27510 30557
tri 27384 30555 27385 30556 ne
rect 27385 30555 27510 30556
tri 27385 30554 27386 30555 ne
rect 27386 30554 27510 30555
tri 27386 30553 27387 30554 ne
rect 27387 30553 27510 30554
tri 27387 30552 27388 30553 ne
rect 27388 30552 27510 30553
tri 27388 30551 27389 30552 ne
rect 27389 30551 27510 30552
tri 27389 30550 27390 30551 ne
rect 27390 30550 27510 30551
tri 27390 30549 27391 30550 ne
rect 27391 30549 27510 30550
tri 27391 30548 27392 30549 ne
rect 27392 30548 27510 30549
tri 27392 30547 27393 30548 ne
rect 27393 30547 27510 30548
tri 27393 30546 27394 30547 ne
rect 27394 30546 27510 30547
tri 27394 30545 27395 30546 ne
rect 27395 30545 27510 30546
tri 27395 30544 27396 30545 ne
rect 27396 30544 27510 30545
tri 27396 30543 27397 30544 ne
rect 27397 30543 27510 30544
tri 27397 30542 27398 30543 ne
rect 27398 30542 27510 30543
tri 27398 30541 27399 30542 ne
rect 27399 30541 27510 30542
tri 27399 30540 27400 30541 ne
rect 27400 30540 27510 30541
tri 27400 30539 27401 30540 ne
rect 27401 30539 27510 30540
tri 27401 30538 27402 30539 ne
rect 27402 30538 27510 30539
tri 27402 30537 27403 30538 ne
rect 27403 30537 27510 30538
tri 27403 30536 27404 30537 ne
rect 27404 30536 27510 30537
tri 27404 30535 27405 30536 ne
rect 27405 30535 27510 30536
tri 27405 30534 27406 30535 ne
rect 27406 30534 27510 30535
tri 27406 30533 27407 30534 ne
rect 27407 30533 27510 30534
tri 27407 30532 27408 30533 ne
rect 27408 30532 27510 30533
tri 27408 30531 27409 30532 ne
rect 27409 30531 27510 30532
tri 27409 30530 27410 30531 ne
rect 27410 30530 27510 30531
tri 27410 30529 27411 30530 ne
rect 27411 30529 27510 30530
tri 27411 30528 27412 30529 ne
rect 27412 30528 27510 30529
tri 27412 30527 27413 30528 ne
rect 27413 30527 27510 30528
tri 27413 30526 27414 30527 ne
rect 27414 30526 27510 30527
tri 27414 30525 27415 30526 ne
rect 27415 30525 27510 30526
tri 27415 30524 27416 30525 ne
rect 27416 30524 27510 30525
tri 27416 30523 27417 30524 ne
rect 27417 30523 27510 30524
tri 27417 30522 27418 30523 ne
rect 27418 30522 27510 30523
rect 27556 30543 27628 30568
tri 27628 30543 27673 30588 sw
rect 70802 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30530 27673 30543
tri 27673 30530 27686 30543 sw
rect 27556 30522 27686 30530
tri 27418 30521 27419 30522 ne
rect 27419 30521 27686 30522
tri 27419 30520 27420 30521 ne
rect 27420 30520 27686 30521
tri 27420 30519 27421 30520 ne
rect 27421 30519 27686 30520
tri 27421 30518 27422 30519 ne
rect 27422 30518 27686 30519
tri 27422 30517 27423 30518 ne
rect 27423 30517 27686 30518
tri 27423 30516 27424 30517 ne
rect 27424 30516 27686 30517
tri 27424 30515 27425 30516 ne
rect 27425 30515 27686 30516
tri 27425 30514 27426 30515 ne
rect 27426 30514 27686 30515
tri 27426 30513 27427 30514 ne
rect 27427 30513 27686 30514
tri 27427 30512 27428 30513 ne
rect 27428 30512 27686 30513
tri 27428 30511 27429 30512 ne
rect 27429 30511 27686 30512
tri 27429 30510 27430 30511 ne
rect 27430 30510 27686 30511
tri 27430 30509 27431 30510 ne
rect 27431 30509 27686 30510
tri 27431 30508 27432 30509 ne
rect 27432 30508 27686 30509
tri 27432 30507 27433 30508 ne
rect 27433 30507 27686 30508
tri 27433 30506 27434 30507 ne
rect 27434 30506 27686 30507
tri 27434 30505 27435 30506 ne
rect 27435 30505 27686 30506
tri 27435 30504 27436 30505 ne
rect 27436 30504 27686 30505
tri 27436 30503 27437 30504 ne
rect 27437 30503 27686 30504
tri 27437 30502 27438 30503 ne
rect 27438 30502 27686 30503
tri 27438 30501 27439 30502 ne
rect 27439 30501 27686 30502
tri 27439 30500 27440 30501 ne
rect 27440 30500 27686 30501
tri 27440 30499 27441 30500 ne
rect 27441 30499 27686 30500
tri 27441 30498 27442 30499 ne
rect 27442 30498 27686 30499
tri 27442 30497 27443 30498 ne
rect 27443 30497 27686 30498
tri 27443 30496 27444 30497 ne
rect 27444 30496 27686 30497
tri 27444 30495 27445 30496 ne
rect 27445 30495 27686 30496
tri 27445 30494 27446 30495 ne
rect 27446 30494 27686 30495
tri 27446 30493 27447 30494 ne
rect 27447 30493 27686 30494
tri 27447 30492 27448 30493 ne
rect 27448 30492 27686 30493
tri 27448 30491 27449 30492 ne
rect 27449 30491 27686 30492
tri 27449 30490 27450 30491 ne
rect 27450 30490 27686 30491
tri 27450 30489 27451 30490 ne
rect 27451 30489 27686 30490
tri 27451 30488 27452 30489 ne
rect 27452 30488 27686 30489
tri 27452 30487 27453 30488 ne
rect 27453 30487 27686 30488
tri 27453 30486 27454 30487 ne
rect 27454 30486 27686 30487
tri 27454 30485 27455 30486 ne
rect 27455 30485 27686 30486
tri 27686 30485 27731 30530 sw
rect 70802 30492 71000 30550
tri 27455 30440 27500 30485 ne
rect 27500 30440 27731 30485
tri 27731 30440 27776 30485 sw
rect 70802 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
tri 27500 30395 27545 30440 ne
rect 27545 30436 27776 30440
rect 27545 30395 27642 30436
tri 27545 30350 27590 30395 ne
rect 27590 30390 27642 30395
rect 27688 30395 27776 30436
tri 27776 30395 27821 30440 sw
rect 27688 30390 27821 30395
rect 27590 30357 27821 30390
tri 27821 30357 27859 30395 sw
rect 70802 30388 71000 30446
rect 27590 30350 27859 30357
tri 27590 30312 27628 30350 ne
rect 27628 30312 27859 30350
tri 27859 30312 27904 30357 sw
rect 70802 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27628 30305 27635 30312 ne
rect 27635 30305 27904 30312
tri 27635 30304 27636 30305 ne
rect 27636 30304 27904 30305
tri 27636 30303 27637 30304 ne
rect 27637 30303 27774 30304
tri 27637 30302 27638 30303 ne
rect 27638 30302 27774 30303
tri 27638 30301 27639 30302 ne
rect 27639 30301 27774 30302
tri 27639 30300 27640 30301 ne
rect 27640 30300 27774 30301
tri 27640 30299 27641 30300 ne
rect 27641 30299 27774 30300
tri 27641 30298 27642 30299 ne
rect 27642 30298 27774 30299
tri 27642 30297 27643 30298 ne
rect 27643 30297 27774 30298
tri 27643 30296 27644 30297 ne
rect 27644 30296 27774 30297
tri 27644 30295 27645 30296 ne
rect 27645 30295 27774 30296
tri 27645 30294 27646 30295 ne
rect 27646 30294 27774 30295
tri 27646 30293 27647 30294 ne
rect 27647 30293 27774 30294
tri 27647 30292 27648 30293 ne
rect 27648 30292 27774 30293
tri 27648 30291 27649 30292 ne
rect 27649 30291 27774 30292
tri 27649 30290 27650 30291 ne
rect 27650 30290 27774 30291
tri 27650 30289 27651 30290 ne
rect 27651 30289 27774 30290
tri 27651 30288 27652 30289 ne
rect 27652 30288 27774 30289
tri 27652 30287 27653 30288 ne
rect 27653 30287 27774 30288
tri 27653 30286 27654 30287 ne
rect 27654 30286 27774 30287
tri 27654 30285 27655 30286 ne
rect 27655 30285 27774 30286
tri 27655 30284 27656 30285 ne
rect 27656 30284 27774 30285
tri 27656 30283 27657 30284 ne
rect 27657 30283 27774 30284
tri 27657 30282 27658 30283 ne
rect 27658 30282 27774 30283
tri 27658 30281 27659 30282 ne
rect 27659 30281 27774 30282
tri 27659 30280 27660 30281 ne
rect 27660 30280 27774 30281
tri 27660 30279 27661 30280 ne
rect 27661 30279 27774 30280
tri 27661 30278 27662 30279 ne
rect 27662 30278 27774 30279
tri 27662 30277 27663 30278 ne
rect 27663 30277 27774 30278
tri 27663 30276 27664 30277 ne
rect 27664 30276 27774 30277
tri 27664 30275 27665 30276 ne
rect 27665 30275 27774 30276
tri 27665 30274 27666 30275 ne
rect 27666 30274 27774 30275
tri 27666 30273 27667 30274 ne
rect 27667 30273 27774 30274
tri 27667 30272 27668 30273 ne
rect 27668 30272 27774 30273
tri 27668 30271 27669 30272 ne
rect 27669 30271 27774 30272
tri 27669 30270 27670 30271 ne
rect 27670 30270 27774 30271
tri 27670 30269 27671 30270 ne
rect 27671 30269 27774 30270
tri 27671 30268 27672 30269 ne
rect 27672 30268 27774 30269
tri 27672 30267 27673 30268 ne
rect 27673 30267 27774 30268
tri 27673 30266 27674 30267 ne
rect 27674 30266 27774 30267
tri 27674 30265 27675 30266 ne
rect 27675 30265 27774 30266
tri 27675 30264 27676 30265 ne
rect 27676 30264 27774 30265
tri 27676 30263 27677 30264 ne
rect 27677 30263 27774 30264
tri 27677 30262 27678 30263 ne
rect 27678 30262 27774 30263
tri 27678 30261 27679 30262 ne
rect 27679 30261 27774 30262
tri 27679 30260 27680 30261 ne
rect 27680 30260 27774 30261
tri 27680 30259 27681 30260 ne
rect 27681 30259 27774 30260
tri 27681 30258 27682 30259 ne
rect 27682 30258 27774 30259
rect 27820 30267 27904 30304
tri 27904 30267 27949 30312 sw
rect 70802 30284 71000 30342
rect 27820 30258 27949 30267
tri 27682 30257 27683 30258 ne
rect 27683 30257 27949 30258
tri 27683 30256 27684 30257 ne
rect 27684 30256 27949 30257
tri 27684 30255 27685 30256 ne
rect 27685 30255 27949 30256
tri 27685 30254 27686 30255 ne
rect 27686 30254 27949 30255
tri 27686 30253 27687 30254 ne
rect 27687 30253 27949 30254
tri 27687 30252 27688 30253 ne
rect 27688 30252 27949 30253
tri 27688 30251 27689 30252 ne
rect 27689 30251 27949 30252
tri 27689 30250 27690 30251 ne
rect 27690 30250 27949 30251
tri 27690 30249 27691 30250 ne
rect 27691 30249 27949 30250
tri 27691 30248 27692 30249 ne
rect 27692 30248 27949 30249
tri 27692 30247 27693 30248 ne
rect 27693 30247 27949 30248
tri 27693 30246 27694 30247 ne
rect 27694 30246 27949 30247
tri 27694 30245 27695 30246 ne
rect 27695 30245 27949 30246
tri 27695 30244 27696 30245 ne
rect 27696 30244 27949 30245
tri 27696 30243 27697 30244 ne
rect 27697 30243 27949 30244
tri 27697 30242 27698 30243 ne
rect 27698 30242 27949 30243
tri 27698 30241 27699 30242 ne
rect 27699 30241 27949 30242
tri 27699 30240 27700 30241 ne
rect 27700 30240 27949 30241
tri 27700 30239 27701 30240 ne
rect 27701 30239 27949 30240
tri 27701 30238 27702 30239 ne
rect 27702 30238 27949 30239
tri 27702 30237 27703 30238 ne
rect 27703 30237 27949 30238
tri 27703 30236 27704 30237 ne
rect 27704 30236 27949 30237
tri 27704 30235 27705 30236 ne
rect 27705 30235 27949 30236
tri 27705 30234 27706 30235 ne
rect 27706 30234 27949 30235
tri 27706 30233 27707 30234 ne
rect 27707 30233 27949 30234
tri 27707 30232 27708 30233 ne
rect 27708 30232 27949 30233
tri 27708 30231 27709 30232 ne
rect 27709 30231 27949 30232
tri 27709 30230 27710 30231 ne
rect 27710 30230 27949 30231
tri 27710 30229 27711 30230 ne
rect 27711 30229 27949 30230
tri 27711 30228 27712 30229 ne
rect 27712 30228 27949 30229
tri 27712 30227 27713 30228 ne
rect 27713 30227 27949 30228
tri 27713 30226 27714 30227 ne
rect 27714 30226 27949 30227
tri 27714 30225 27715 30226 ne
rect 27715 30225 27949 30226
tri 27715 30224 27716 30225 ne
rect 27716 30224 27949 30225
tri 27716 30223 27717 30224 ne
rect 27717 30223 27949 30224
tri 27717 30222 27718 30223 ne
rect 27718 30222 27949 30223
tri 27949 30222 27994 30267 sw
rect 70802 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27718 30221 27719 30222 ne
rect 27719 30221 27994 30222
tri 27719 30220 27720 30221 ne
rect 27720 30220 27994 30221
tri 27720 30219 27721 30220 ne
rect 27721 30219 27994 30220
tri 27721 30218 27722 30219 ne
rect 27722 30218 27994 30219
tri 27722 30217 27723 30218 ne
rect 27723 30217 27994 30218
tri 27723 30216 27724 30217 ne
rect 27724 30216 27994 30217
tri 27724 30215 27725 30216 ne
rect 27725 30215 27994 30216
tri 27725 30214 27726 30215 ne
rect 27726 30214 27994 30215
tri 27726 30213 27727 30214 ne
rect 27727 30213 27994 30214
tri 27727 30212 27728 30213 ne
rect 27728 30212 27994 30213
tri 27728 30211 27729 30212 ne
rect 27729 30211 27994 30212
tri 27729 30210 27730 30211 ne
rect 27730 30210 27994 30211
tri 27730 30209 27731 30210 ne
rect 27731 30209 27994 30210
tri 27994 30209 28007 30222 sw
tri 27731 30164 27776 30209 ne
rect 27776 30172 28007 30209
rect 27776 30164 27906 30172
tri 27776 30149 27791 30164 ne
rect 27791 30149 27906 30164
tri 27791 30104 27836 30149 ne
rect 27836 30126 27906 30149
rect 27952 30164 28007 30172
tri 28007 30164 28052 30209 sw
rect 70802 30180 71000 30238
rect 27952 30126 28052 30164
rect 27836 30119 28052 30126
tri 28052 30119 28097 30164 sw
rect 70802 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 27836 30104 28097 30119
tri 27836 30059 27881 30104 ne
rect 27881 30074 28097 30104
tri 28097 30074 28142 30119 sw
rect 70802 30076 71000 30134
rect 27881 30068 28142 30074
tri 28142 30068 28148 30074 sw
rect 27881 30059 28148 30068
tri 27881 30029 27911 30059 ne
rect 27911 30040 28148 30059
rect 27911 30029 28038 30040
tri 27911 30028 27912 30029 ne
rect 27912 30028 28038 30029
tri 27912 30027 27913 30028 ne
rect 27913 30027 28038 30028
tri 27913 30026 27914 30027 ne
rect 27914 30026 28038 30027
tri 27914 30025 27915 30026 ne
rect 27915 30025 28038 30026
tri 27915 30024 27916 30025 ne
rect 27916 30024 28038 30025
tri 27916 30023 27917 30024 ne
rect 27917 30023 28038 30024
tri 27917 30022 27918 30023 ne
rect 27918 30022 28038 30023
tri 27918 30021 27919 30022 ne
rect 27919 30021 28038 30022
tri 27919 30020 27920 30021 ne
rect 27920 30020 28038 30021
tri 27920 30019 27921 30020 ne
rect 27921 30019 28038 30020
tri 27921 30018 27922 30019 ne
rect 27922 30018 28038 30019
tri 27922 30017 27923 30018 ne
rect 27923 30017 28038 30018
tri 27923 30016 27924 30017 ne
rect 27924 30016 28038 30017
tri 27924 30015 27925 30016 ne
rect 27925 30015 28038 30016
tri 27925 30014 27926 30015 ne
rect 27926 30014 28038 30015
tri 27926 30013 27927 30014 ne
rect 27927 30013 28038 30014
tri 27927 30012 27928 30013 ne
rect 27928 30012 28038 30013
tri 27928 30011 27929 30012 ne
rect 27929 30011 28038 30012
tri 27929 30010 27930 30011 ne
rect 27930 30010 28038 30011
tri 27930 30009 27931 30010 ne
rect 27931 30009 28038 30010
tri 27931 30008 27932 30009 ne
rect 27932 30008 28038 30009
tri 27932 30007 27933 30008 ne
rect 27933 30007 28038 30008
tri 27933 30006 27934 30007 ne
rect 27934 30006 28038 30007
tri 27934 30005 27935 30006 ne
rect 27935 30005 28038 30006
tri 27935 30004 27936 30005 ne
rect 27936 30004 28038 30005
tri 27936 30003 27937 30004 ne
rect 27937 30003 28038 30004
tri 27937 30002 27938 30003 ne
rect 27938 30002 28038 30003
tri 27938 30001 27939 30002 ne
rect 27939 30001 28038 30002
tri 27939 30000 27940 30001 ne
rect 27940 30000 28038 30001
tri 27940 29999 27941 30000 ne
rect 27941 29999 28038 30000
tri 27941 29998 27942 29999 ne
rect 27942 29998 28038 29999
tri 27942 29997 27943 29998 ne
rect 27943 29997 28038 29998
tri 27943 29996 27944 29997 ne
rect 27944 29996 28038 29997
tri 27944 29995 27945 29996 ne
rect 27945 29995 28038 29996
tri 27945 29994 27946 29995 ne
rect 27946 29994 28038 29995
rect 28084 30023 28148 30040
tri 28148 30023 28193 30068 sw
rect 70802 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 29994 28193 30023
tri 27946 29993 27947 29994 ne
rect 27947 29993 28193 29994
tri 27947 29992 27948 29993 ne
rect 27948 29992 28193 29993
tri 27948 29991 27949 29992 ne
rect 27949 29991 28193 29992
tri 27949 29990 27950 29991 ne
rect 27950 29990 28193 29991
tri 27950 29989 27951 29990 ne
rect 27951 29989 28193 29990
tri 27951 29988 27952 29989 ne
rect 27952 29988 28193 29989
tri 27952 29987 27953 29988 ne
rect 27953 29987 28193 29988
tri 27953 29986 27954 29987 ne
rect 27954 29986 28193 29987
tri 27954 29985 27955 29986 ne
rect 27955 29985 28193 29986
tri 27955 29984 27956 29985 ne
rect 27956 29984 28193 29985
tri 27956 29983 27957 29984 ne
rect 27957 29983 28193 29984
tri 27957 29982 27958 29983 ne
rect 27958 29982 28193 29983
tri 27958 29981 27959 29982 ne
rect 27959 29981 28193 29982
tri 27959 29980 27960 29981 ne
rect 27960 29980 28193 29981
tri 27960 29979 27961 29980 ne
rect 27961 29979 28193 29980
tri 27961 29978 27962 29979 ne
rect 27962 29978 28193 29979
tri 28193 29978 28238 30023 sw
tri 27962 29977 27963 29978 ne
rect 27963 29977 28238 29978
tri 27963 29976 27964 29977 ne
rect 27964 29976 28238 29977
tri 27964 29975 27965 29976 ne
rect 27965 29975 28238 29976
tri 27965 29974 27966 29975 ne
rect 27966 29974 28238 29975
tri 27966 29973 27967 29974 ne
rect 27967 29973 28238 29974
tri 27967 29972 27968 29973 ne
rect 27968 29972 28238 29973
tri 27968 29971 27969 29972 ne
rect 27969 29971 28238 29972
tri 27969 29970 27970 29971 ne
rect 27970 29970 28238 29971
tri 27970 29969 27971 29970 ne
rect 27971 29969 28238 29970
tri 27971 29968 27972 29969 ne
rect 27972 29968 28238 29969
tri 27972 29967 27973 29968 ne
rect 27973 29967 28238 29968
tri 27973 29966 27974 29967 ne
rect 27974 29966 28238 29967
tri 27974 29965 27975 29966 ne
rect 27975 29965 28238 29966
tri 27975 29964 27976 29965 ne
rect 27976 29964 28238 29965
tri 27976 29963 27977 29964 ne
rect 27977 29963 28238 29964
tri 27977 29962 27978 29963 ne
rect 27978 29962 28238 29963
tri 27978 29961 27979 29962 ne
rect 27979 29961 28238 29962
tri 27979 29960 27980 29961 ne
rect 27980 29960 28238 29961
tri 27980 29959 27981 29960 ne
rect 27981 29959 28238 29960
tri 27981 29958 27982 29959 ne
rect 27982 29958 28238 29959
tri 27982 29957 27983 29958 ne
rect 27983 29957 28238 29958
tri 27983 29956 27984 29957 ne
rect 27984 29956 28238 29957
tri 27984 29955 27985 29956 ne
rect 27985 29955 28238 29956
tri 27985 29954 27986 29955 ne
rect 27986 29954 28238 29955
tri 27986 29953 27987 29954 ne
rect 27987 29953 28238 29954
tri 27987 29952 27988 29953 ne
rect 27988 29952 28238 29953
tri 27988 29951 27989 29952 ne
rect 27989 29951 28238 29952
tri 27989 29950 27990 29951 ne
rect 27990 29950 28238 29951
tri 27990 29949 27991 29950 ne
rect 27991 29949 28238 29950
tri 27991 29948 27992 29949 ne
rect 27992 29948 28238 29949
tri 27992 29947 27993 29948 ne
rect 27993 29947 28238 29948
tri 27993 29946 27994 29947 ne
rect 27994 29946 28238 29947
tri 27994 29945 27995 29946 ne
rect 27995 29945 28238 29946
tri 27995 29944 27996 29945 ne
rect 27996 29944 28238 29945
tri 27996 29943 27997 29944 ne
rect 27997 29943 28238 29944
tri 27997 29942 27998 29943 ne
rect 27998 29942 28238 29943
tri 27998 29941 27999 29942 ne
rect 27999 29941 28238 29942
tri 27999 29940 28000 29941 ne
rect 28000 29940 28238 29941
tri 28000 29939 28001 29940 ne
rect 28001 29939 28238 29940
tri 28001 29938 28002 29939 ne
rect 28002 29938 28238 29939
tri 28002 29937 28003 29938 ne
rect 28003 29937 28238 29938
tri 28003 29936 28004 29937 ne
rect 28004 29936 28238 29937
tri 28004 29935 28005 29936 ne
rect 28005 29935 28238 29936
tri 28005 29934 28006 29935 ne
rect 28006 29934 28238 29935
tri 28006 29933 28007 29934 ne
rect 28007 29933 28238 29934
tri 28238 29933 28283 29978 sw
rect 70802 29972 71000 30030
tri 28007 29901 28039 29933 ne
rect 28039 29908 28283 29933
rect 28039 29901 28170 29908
tri 28039 29856 28084 29901 ne
rect 28084 29862 28170 29901
rect 28216 29901 28283 29908
tri 28283 29901 28315 29933 sw
rect 70802 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 28216 29862 28315 29901
rect 28084 29856 28315 29862
tri 28315 29856 28360 29901 sw
rect 70802 29868 71000 29926
tri 28084 29829 28111 29856 ne
rect 28111 29829 28360 29856
tri 28111 29784 28156 29829 ne
rect 28156 29811 28360 29829
tri 28360 29811 28405 29856 sw
rect 70802 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28156 29784 28405 29811
tri 28156 29755 28185 29784 ne
rect 28185 29776 28405 29784
rect 28185 29755 28302 29776
tri 28185 29754 28186 29755 ne
rect 28186 29754 28302 29755
tri 28186 29753 28187 29754 ne
rect 28187 29753 28302 29754
tri 28187 29752 28188 29753 ne
rect 28188 29752 28302 29753
tri 28188 29751 28189 29752 ne
rect 28189 29751 28302 29752
tri 28189 29750 28190 29751 ne
rect 28190 29750 28302 29751
tri 28190 29749 28191 29750 ne
rect 28191 29749 28302 29750
tri 28191 29748 28192 29749 ne
rect 28192 29748 28302 29749
tri 28192 29747 28193 29748 ne
rect 28193 29747 28302 29748
tri 28193 29746 28194 29747 ne
rect 28194 29746 28302 29747
tri 28194 29745 28195 29746 ne
rect 28195 29745 28302 29746
tri 28195 29744 28196 29745 ne
rect 28196 29744 28302 29745
tri 28196 29743 28197 29744 ne
rect 28197 29743 28302 29744
tri 28197 29742 28198 29743 ne
rect 28198 29742 28302 29743
tri 28198 29741 28199 29742 ne
rect 28199 29741 28302 29742
tri 28199 29740 28200 29741 ne
rect 28200 29740 28302 29741
tri 28200 29739 28201 29740 ne
rect 28201 29739 28302 29740
tri 28201 29738 28202 29739 ne
rect 28202 29738 28302 29739
tri 28202 29737 28203 29738 ne
rect 28203 29737 28302 29738
tri 28203 29736 28204 29737 ne
rect 28204 29736 28302 29737
tri 28204 29735 28205 29736 ne
rect 28205 29735 28302 29736
tri 28205 29734 28206 29735 ne
rect 28206 29734 28302 29735
tri 28206 29733 28207 29734 ne
rect 28207 29733 28302 29734
tri 28207 29732 28208 29733 ne
rect 28208 29732 28302 29733
tri 28208 29731 28209 29732 ne
rect 28209 29731 28302 29732
tri 28209 29730 28210 29731 ne
rect 28210 29730 28302 29731
rect 28348 29766 28405 29776
tri 28405 29766 28450 29811 sw
rect 28348 29747 28450 29766
tri 28450 29747 28469 29766 sw
rect 70802 29764 71000 29822
rect 28348 29730 28469 29747
tri 28210 29729 28211 29730 ne
rect 28211 29729 28469 29730
tri 28211 29728 28212 29729 ne
rect 28212 29728 28469 29729
tri 28212 29727 28213 29728 ne
rect 28213 29727 28469 29728
tri 28213 29726 28214 29727 ne
rect 28214 29726 28469 29727
tri 28214 29725 28215 29726 ne
rect 28215 29725 28469 29726
tri 28215 29724 28216 29725 ne
rect 28216 29724 28469 29725
tri 28216 29723 28217 29724 ne
rect 28217 29723 28469 29724
tri 28217 29722 28218 29723 ne
rect 28218 29722 28469 29723
tri 28218 29721 28219 29722 ne
rect 28219 29721 28469 29722
tri 28219 29720 28220 29721 ne
rect 28220 29720 28469 29721
tri 28220 29719 28221 29720 ne
rect 28221 29719 28469 29720
tri 28221 29718 28222 29719 ne
rect 28222 29718 28469 29719
tri 28222 29717 28223 29718 ne
rect 28223 29717 28469 29718
tri 28223 29716 28224 29717 ne
rect 28224 29716 28469 29717
tri 28224 29715 28225 29716 ne
rect 28225 29715 28469 29716
tri 28225 29714 28226 29715 ne
rect 28226 29714 28469 29715
tri 28226 29713 28227 29714 ne
rect 28227 29713 28469 29714
tri 28227 29712 28228 29713 ne
rect 28228 29712 28469 29713
tri 28228 29711 28229 29712 ne
rect 28229 29711 28469 29712
tri 28229 29710 28230 29711 ne
rect 28230 29710 28469 29711
tri 28230 29709 28231 29710 ne
rect 28231 29709 28469 29710
tri 28231 29708 28232 29709 ne
rect 28232 29708 28469 29709
tri 28232 29707 28233 29708 ne
rect 28233 29707 28469 29708
tri 28233 29706 28234 29707 ne
rect 28234 29706 28469 29707
tri 28234 29705 28235 29706 ne
rect 28235 29705 28469 29706
tri 28235 29704 28236 29705 ne
rect 28236 29704 28469 29705
tri 28236 29703 28237 29704 ne
rect 28237 29703 28469 29704
tri 28237 29702 28238 29703 ne
rect 28238 29702 28469 29703
tri 28469 29702 28514 29747 sw
rect 70802 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
tri 28238 29701 28239 29702 ne
rect 28239 29701 28514 29702
tri 28239 29700 28240 29701 ne
rect 28240 29700 28514 29701
tri 28240 29699 28241 29700 ne
rect 28241 29699 28514 29700
tri 28241 29698 28242 29699 ne
rect 28242 29698 28514 29699
tri 28242 29697 28243 29698 ne
rect 28243 29697 28514 29698
tri 28243 29696 28244 29697 ne
rect 28244 29696 28514 29697
tri 28244 29695 28245 29696 ne
rect 28245 29695 28514 29696
tri 28245 29694 28246 29695 ne
rect 28246 29694 28514 29695
tri 28246 29693 28247 29694 ne
rect 28247 29693 28514 29694
tri 28247 29692 28248 29693 ne
rect 28248 29692 28514 29693
tri 28248 29691 28249 29692 ne
rect 28249 29691 28514 29692
tri 28249 29690 28250 29691 ne
rect 28250 29690 28514 29691
tri 28250 29689 28251 29690 ne
rect 28251 29689 28514 29690
tri 28251 29688 28252 29689 ne
rect 28252 29688 28514 29689
tri 28252 29687 28253 29688 ne
rect 28253 29687 28514 29688
tri 28253 29686 28254 29687 ne
rect 28254 29686 28514 29687
tri 28254 29685 28255 29686 ne
rect 28255 29685 28514 29686
tri 28255 29684 28256 29685 ne
rect 28256 29684 28514 29685
tri 28256 29683 28257 29684 ne
rect 28257 29683 28514 29684
tri 28257 29682 28258 29683 ne
rect 28258 29682 28514 29683
tri 28258 29681 28259 29682 ne
rect 28259 29681 28514 29682
tri 28259 29680 28260 29681 ne
rect 28260 29680 28514 29681
tri 28260 29679 28261 29680 ne
rect 28261 29679 28514 29680
tri 28261 29678 28262 29679 ne
rect 28262 29678 28514 29679
tri 28262 29677 28263 29678 ne
rect 28263 29677 28514 29678
tri 28263 29676 28264 29677 ne
rect 28264 29676 28514 29677
tri 28264 29675 28265 29676 ne
rect 28265 29675 28514 29676
tri 28265 29674 28266 29675 ne
rect 28266 29674 28514 29675
tri 28266 29673 28267 29674 ne
rect 28267 29673 28514 29674
tri 28267 29672 28268 29673 ne
rect 28268 29672 28514 29673
tri 28268 29671 28269 29672 ne
rect 28269 29671 28514 29672
tri 28269 29670 28270 29671 ne
rect 28270 29670 28514 29671
tri 28270 29669 28271 29670 ne
rect 28271 29669 28514 29670
tri 28271 29668 28272 29669 ne
rect 28272 29668 28514 29669
tri 28272 29667 28273 29668 ne
rect 28273 29667 28514 29668
tri 28273 29666 28274 29667 ne
rect 28274 29666 28514 29667
tri 28274 29665 28275 29666 ne
rect 28275 29665 28514 29666
tri 28275 29664 28276 29665 ne
rect 28276 29664 28514 29665
tri 28276 29663 28277 29664 ne
rect 28277 29663 28514 29664
tri 28277 29662 28278 29663 ne
rect 28278 29662 28514 29663
tri 28278 29661 28279 29662 ne
rect 28279 29661 28514 29662
tri 28279 29660 28280 29661 ne
rect 28280 29660 28514 29661
tri 28280 29659 28281 29660 ne
rect 28281 29659 28514 29660
tri 28281 29658 28282 29659 ne
rect 28282 29658 28514 29659
tri 28282 29657 28283 29658 ne
rect 28283 29657 28514 29658
tri 28514 29657 28559 29702 sw
rect 70802 29660 71000 29718
tri 28283 29612 28328 29657 ne
rect 28328 29644 28559 29657
rect 28328 29612 28434 29644
tri 28328 29580 28360 29612 ne
rect 28360 29598 28434 29612
rect 28480 29612 28559 29644
tri 28559 29612 28604 29657 sw
rect 70802 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 28480 29598 28604 29612
rect 28360 29580 28604 29598
tri 28604 29580 28636 29612 sw
tri 28360 29567 28373 29580 ne
rect 28373 29567 28636 29580
tri 28373 29535 28405 29567 ne
rect 28405 29535 28636 29567
tri 28636 29535 28681 29580 sw
rect 70802 29556 71000 29614
tri 28405 29490 28450 29535 ne
rect 28450 29512 28681 29535
rect 28450 29490 28566 29512
tri 28450 29481 28459 29490 ne
rect 28459 29481 28566 29490
tri 28459 29480 28460 29481 ne
rect 28460 29480 28566 29481
tri 28460 29479 28461 29480 ne
rect 28461 29479 28566 29480
tri 28461 29478 28462 29479 ne
rect 28462 29478 28566 29479
tri 28462 29477 28463 29478 ne
rect 28463 29477 28566 29478
tri 28463 29476 28464 29477 ne
rect 28464 29476 28566 29477
tri 28464 29475 28465 29476 ne
rect 28465 29475 28566 29476
tri 28465 29474 28466 29475 ne
rect 28466 29474 28566 29475
tri 28466 29473 28467 29474 ne
rect 28467 29473 28566 29474
tri 28467 29472 28468 29473 ne
rect 28468 29472 28566 29473
tri 28468 29471 28469 29472 ne
rect 28469 29471 28566 29472
tri 28469 29470 28470 29471 ne
rect 28470 29470 28566 29471
tri 28470 29469 28471 29470 ne
rect 28471 29469 28566 29470
tri 28471 29468 28472 29469 ne
rect 28472 29468 28566 29469
tri 28472 29467 28473 29468 ne
rect 28473 29467 28566 29468
tri 28473 29466 28474 29467 ne
rect 28474 29466 28566 29467
rect 28612 29490 28681 29512
tri 28681 29490 28726 29535 sw
rect 70802 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29466 28726 29490
tri 28474 29465 28475 29466 ne
rect 28475 29465 28726 29466
tri 28475 29464 28476 29465 ne
rect 28476 29464 28726 29465
tri 28476 29463 28477 29464 ne
rect 28477 29463 28726 29464
tri 28477 29462 28478 29463 ne
rect 28478 29462 28726 29463
tri 28478 29461 28479 29462 ne
rect 28479 29461 28726 29462
tri 28479 29460 28480 29461 ne
rect 28480 29460 28726 29461
tri 28480 29459 28481 29460 ne
rect 28481 29459 28726 29460
tri 28481 29458 28482 29459 ne
rect 28482 29458 28726 29459
tri 28482 29457 28483 29458 ne
rect 28483 29457 28726 29458
tri 28483 29456 28484 29457 ne
rect 28484 29456 28726 29457
tri 28484 29455 28485 29456 ne
rect 28485 29455 28726 29456
tri 28485 29454 28486 29455 ne
rect 28486 29454 28726 29455
tri 28486 29453 28487 29454 ne
rect 28487 29453 28726 29454
tri 28487 29452 28488 29453 ne
rect 28488 29452 28726 29453
tri 28488 29451 28489 29452 ne
rect 28489 29451 28726 29452
tri 28489 29450 28490 29451 ne
rect 28490 29450 28726 29451
tri 28490 29449 28491 29450 ne
rect 28491 29449 28726 29450
tri 28491 29448 28492 29449 ne
rect 28492 29448 28726 29449
tri 28492 29447 28493 29448 ne
rect 28493 29447 28726 29448
tri 28493 29446 28494 29447 ne
rect 28494 29446 28726 29447
tri 28494 29445 28495 29446 ne
rect 28495 29445 28726 29446
tri 28726 29445 28771 29490 sw
rect 70802 29452 71000 29510
tri 28495 29444 28496 29445 ne
rect 28496 29444 28771 29445
tri 28496 29443 28497 29444 ne
rect 28497 29443 28771 29444
tri 28497 29442 28498 29443 ne
rect 28498 29442 28771 29443
tri 28498 29441 28499 29442 ne
rect 28499 29441 28771 29442
tri 28499 29440 28500 29441 ne
rect 28500 29440 28771 29441
tri 28500 29439 28501 29440 ne
rect 28501 29439 28771 29440
tri 28501 29438 28502 29439 ne
rect 28502 29438 28771 29439
tri 28502 29437 28503 29438 ne
rect 28503 29437 28771 29438
tri 28503 29436 28504 29437 ne
rect 28504 29436 28771 29437
tri 28504 29435 28505 29436 ne
rect 28505 29435 28771 29436
tri 28505 29434 28506 29435 ne
rect 28506 29434 28771 29435
tri 28506 29433 28507 29434 ne
rect 28507 29433 28771 29434
tri 28507 29432 28508 29433 ne
rect 28508 29432 28771 29433
tri 28508 29431 28509 29432 ne
rect 28509 29431 28771 29432
tri 28509 29430 28510 29431 ne
rect 28510 29430 28771 29431
tri 28510 29429 28511 29430 ne
rect 28511 29429 28771 29430
tri 28511 29428 28512 29429 ne
rect 28512 29428 28771 29429
tri 28512 29427 28513 29428 ne
rect 28513 29427 28771 29428
tri 28513 29426 28514 29427 ne
rect 28514 29426 28771 29427
tri 28771 29426 28790 29445 sw
tri 28514 29425 28515 29426 ne
rect 28515 29425 28790 29426
tri 28515 29424 28516 29425 ne
rect 28516 29424 28790 29425
tri 28516 29423 28517 29424 ne
rect 28517 29423 28790 29424
tri 28517 29422 28518 29423 ne
rect 28518 29422 28790 29423
tri 28518 29421 28519 29422 ne
rect 28519 29421 28790 29422
tri 28519 29420 28520 29421 ne
rect 28520 29420 28790 29421
tri 28520 29419 28521 29420 ne
rect 28521 29419 28790 29420
tri 28521 29418 28522 29419 ne
rect 28522 29418 28790 29419
tri 28522 29417 28523 29418 ne
rect 28523 29417 28790 29418
tri 28523 29416 28524 29417 ne
rect 28524 29416 28790 29417
tri 28524 29415 28525 29416 ne
rect 28525 29415 28790 29416
tri 28525 29414 28526 29415 ne
rect 28526 29414 28790 29415
tri 28526 29413 28527 29414 ne
rect 28527 29413 28790 29414
tri 28527 29412 28528 29413 ne
rect 28528 29412 28790 29413
tri 28528 29411 28529 29412 ne
rect 28529 29411 28790 29412
tri 28529 29410 28530 29411 ne
rect 28530 29410 28790 29411
tri 28530 29409 28531 29410 ne
rect 28531 29409 28790 29410
tri 28531 29408 28532 29409 ne
rect 28532 29408 28790 29409
tri 28532 29407 28533 29408 ne
rect 28533 29407 28790 29408
tri 28533 29406 28534 29407 ne
rect 28534 29406 28790 29407
tri 28534 29405 28535 29406 ne
rect 28535 29405 28790 29406
tri 28535 29404 28536 29405 ne
rect 28536 29404 28790 29405
tri 28536 29403 28537 29404 ne
rect 28537 29403 28790 29404
tri 28537 29402 28538 29403 ne
rect 28538 29402 28790 29403
tri 28538 29401 28539 29402 ne
rect 28539 29401 28790 29402
tri 28539 29400 28540 29401 ne
rect 28540 29400 28790 29401
tri 28540 29399 28541 29400 ne
rect 28541 29399 28790 29400
tri 28541 29398 28542 29399 ne
rect 28542 29398 28790 29399
tri 28542 29397 28543 29398 ne
rect 28543 29397 28790 29398
tri 28543 29396 28544 29397 ne
rect 28544 29396 28790 29397
tri 28544 29395 28545 29396 ne
rect 28545 29395 28790 29396
tri 28545 29394 28546 29395 ne
rect 28546 29394 28790 29395
tri 28546 29393 28547 29394 ne
rect 28547 29393 28790 29394
tri 28547 29392 28548 29393 ne
rect 28548 29392 28790 29393
tri 28548 29391 28549 29392 ne
rect 28549 29391 28790 29392
tri 28549 29390 28550 29391 ne
rect 28550 29390 28790 29391
tri 28550 29389 28551 29390 ne
rect 28551 29389 28790 29390
tri 28551 29388 28552 29389 ne
rect 28552 29388 28790 29389
tri 28552 29387 28553 29388 ne
rect 28553 29387 28790 29388
tri 28553 29386 28554 29387 ne
rect 28554 29386 28790 29387
tri 28554 29385 28555 29386 ne
rect 28555 29385 28790 29386
tri 28555 29384 28556 29385 ne
rect 28556 29384 28790 29385
tri 28556 29383 28557 29384 ne
rect 28557 29383 28790 29384
tri 28557 29382 28558 29383 ne
rect 28558 29382 28790 29383
tri 28558 29381 28559 29382 ne
rect 28559 29381 28790 29382
tri 28790 29381 28835 29426 sw
rect 70802 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28559 29336 28604 29381 ne
rect 28604 29380 28835 29381
rect 28604 29336 28698 29380
tri 28604 29291 28649 29336 ne
rect 28649 29334 28698 29336
rect 28744 29336 28835 29380
tri 28835 29336 28880 29381 sw
rect 70802 29348 71000 29406
rect 28744 29334 28880 29336
rect 28649 29291 28880 29334
tri 28880 29291 28925 29336 sw
rect 70802 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28649 29246 28694 29291 ne
rect 28694 29259 28925 29291
tri 28925 29259 28957 29291 sw
rect 28694 29248 28957 29259
rect 28694 29246 28830 29248
tri 28694 29214 28726 29246 ne
rect 28726 29214 28830 29246
tri 28726 29206 28734 29214 ne
rect 28734 29206 28830 29214
tri 28734 29205 28735 29206 ne
rect 28735 29205 28830 29206
tri 28735 29204 28736 29205 ne
rect 28736 29204 28830 29205
tri 28736 29203 28737 29204 ne
rect 28737 29203 28830 29204
tri 28737 29202 28738 29203 ne
rect 28738 29202 28830 29203
rect 28876 29214 28957 29248
tri 28957 29214 29002 29259 sw
rect 70802 29244 71000 29302
rect 28876 29202 29002 29214
tri 28738 29201 28739 29202 ne
rect 28739 29201 29002 29202
tri 28739 29200 28740 29201 ne
rect 28740 29200 29002 29201
tri 28740 29199 28741 29200 ne
rect 28741 29199 29002 29200
tri 28741 29198 28742 29199 ne
rect 28742 29198 29002 29199
tri 28742 29197 28743 29198 ne
rect 28743 29197 29002 29198
tri 28743 29196 28744 29197 ne
rect 28744 29196 29002 29197
tri 28744 29195 28745 29196 ne
rect 28745 29195 29002 29196
tri 28745 29194 28746 29195 ne
rect 28746 29194 29002 29195
tri 28746 29193 28747 29194 ne
rect 28747 29193 29002 29194
tri 28747 29192 28748 29193 ne
rect 28748 29192 29002 29193
tri 28748 29191 28749 29192 ne
rect 28749 29191 29002 29192
tri 28749 29190 28750 29191 ne
rect 28750 29190 29002 29191
tri 28750 29189 28751 29190 ne
rect 28751 29189 29002 29190
tri 28751 29188 28752 29189 ne
rect 28752 29188 29002 29189
tri 28752 29187 28753 29188 ne
rect 28753 29187 29002 29188
tri 28753 29186 28754 29187 ne
rect 28754 29186 29002 29187
tri 28754 29185 28755 29186 ne
rect 28755 29185 29002 29186
tri 28755 29184 28756 29185 ne
rect 28756 29184 29002 29185
tri 28756 29183 28757 29184 ne
rect 28757 29183 29002 29184
tri 28757 29182 28758 29183 ne
rect 28758 29182 29002 29183
tri 28758 29181 28759 29182 ne
rect 28759 29181 29002 29182
tri 28759 29180 28760 29181 ne
rect 28760 29180 29002 29181
tri 28760 29179 28761 29180 ne
rect 28761 29179 29002 29180
tri 28761 29178 28762 29179 ne
rect 28762 29178 29002 29179
tri 28762 29177 28763 29178 ne
rect 28763 29177 29002 29178
tri 28763 29176 28764 29177 ne
rect 28764 29176 29002 29177
tri 28764 29175 28765 29176 ne
rect 28765 29175 29002 29176
tri 28765 29174 28766 29175 ne
rect 28766 29174 29002 29175
tri 28766 29173 28767 29174 ne
rect 28767 29173 29002 29174
tri 28767 29172 28768 29173 ne
rect 28768 29172 29002 29173
tri 28768 29171 28769 29172 ne
rect 28769 29171 29002 29172
tri 28769 29170 28770 29171 ne
rect 28770 29170 29002 29171
tri 28770 29169 28771 29170 ne
rect 28771 29169 29002 29170
tri 29002 29169 29047 29214 sw
rect 70802 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
tri 28771 29168 28772 29169 ne
rect 28772 29168 29047 29169
tri 28772 29167 28773 29168 ne
rect 28773 29167 29047 29168
tri 28773 29166 28774 29167 ne
rect 28774 29166 29047 29167
tri 28774 29165 28775 29166 ne
rect 28775 29165 29047 29166
tri 28775 29164 28776 29165 ne
rect 28776 29164 29047 29165
tri 28776 29163 28777 29164 ne
rect 28777 29163 29047 29164
tri 28777 29162 28778 29163 ne
rect 28778 29162 29047 29163
tri 28778 29161 28779 29162 ne
rect 28779 29161 29047 29162
tri 28779 29160 28780 29161 ne
rect 28780 29160 29047 29161
tri 28780 29159 28781 29160 ne
rect 28781 29159 29047 29160
tri 28781 29158 28782 29159 ne
rect 28782 29158 29047 29159
tri 28782 29157 28783 29158 ne
rect 28783 29157 29047 29158
tri 28783 29156 28784 29157 ne
rect 28784 29156 29047 29157
tri 28784 29155 28785 29156 ne
rect 28785 29155 29047 29156
tri 28785 29154 28786 29155 ne
rect 28786 29154 29047 29155
tri 28786 29153 28787 29154 ne
rect 28787 29153 29047 29154
tri 28787 29152 28788 29153 ne
rect 28788 29152 29047 29153
tri 28788 29151 28789 29152 ne
rect 28789 29151 29047 29152
tri 28789 29150 28790 29151 ne
rect 28790 29150 29047 29151
tri 28790 29149 28791 29150 ne
rect 28791 29149 29047 29150
tri 28791 29148 28792 29149 ne
rect 28792 29148 29047 29149
tri 28792 29147 28793 29148 ne
rect 28793 29147 29047 29148
tri 28793 29146 28794 29147 ne
rect 28794 29146 29047 29147
tri 28794 29145 28795 29146 ne
rect 28795 29145 29047 29146
tri 28795 29144 28796 29145 ne
rect 28796 29144 29047 29145
tri 28796 29143 28797 29144 ne
rect 28797 29143 29047 29144
tri 28797 29142 28798 29143 ne
rect 28798 29142 29047 29143
tri 28798 29141 28799 29142 ne
rect 28799 29141 29047 29142
tri 28799 29140 28800 29141 ne
rect 28800 29140 29047 29141
tri 28800 29139 28801 29140 ne
rect 28801 29139 29047 29140
tri 28801 29138 28802 29139 ne
rect 28802 29138 29047 29139
tri 28802 29137 28803 29138 ne
rect 28803 29137 29047 29138
tri 28803 29136 28804 29137 ne
rect 28804 29136 29047 29137
tri 28804 29135 28805 29136 ne
rect 28805 29135 29047 29136
tri 28805 29134 28806 29135 ne
rect 28806 29134 29047 29135
tri 28806 29133 28807 29134 ne
rect 28807 29133 29047 29134
tri 28807 29132 28808 29133 ne
rect 28808 29132 29047 29133
tri 28808 29131 28809 29132 ne
rect 28809 29131 29047 29132
tri 28809 29130 28810 29131 ne
rect 28810 29130 29047 29131
tri 28810 29129 28811 29130 ne
rect 28811 29129 29047 29130
tri 28811 29128 28812 29129 ne
rect 28812 29128 29047 29129
tri 28812 29127 28813 29128 ne
rect 28813 29127 29047 29128
tri 28813 29126 28814 29127 ne
rect 28814 29126 29047 29127
tri 28814 29125 28815 29126 ne
rect 28815 29125 29047 29126
tri 28815 29124 28816 29125 ne
rect 28816 29124 29047 29125
tri 29047 29124 29092 29169 sw
rect 70802 29140 71000 29198
tri 28816 29123 28817 29124 ne
rect 28817 29123 29092 29124
tri 28817 29122 28818 29123 ne
rect 28818 29122 29092 29123
tri 28818 29121 28819 29122 ne
rect 28819 29121 29092 29122
tri 28819 29120 28820 29121 ne
rect 28820 29120 29092 29121
tri 28820 29119 28821 29120 ne
rect 28821 29119 29092 29120
tri 28821 29118 28822 29119 ne
rect 28822 29118 29092 29119
tri 28822 29117 28823 29118 ne
rect 28823 29117 29092 29118
tri 28823 29116 28824 29117 ne
rect 28824 29116 29092 29117
tri 28824 29115 28825 29116 ne
rect 28825 29115 28962 29116
tri 28825 29114 28826 29115 ne
rect 28826 29114 28962 29115
tri 28826 29113 28827 29114 ne
rect 28827 29113 28962 29114
tri 28827 29112 28828 29113 ne
rect 28828 29112 28962 29113
tri 28828 29111 28829 29112 ne
rect 28829 29111 28962 29112
tri 28829 29110 28830 29111 ne
rect 28830 29110 28962 29111
tri 28830 29109 28831 29110 ne
rect 28831 29109 28962 29110
tri 28831 29108 28832 29109 ne
rect 28832 29108 28962 29109
tri 28832 29107 28833 29108 ne
rect 28833 29107 28962 29108
tri 28833 29106 28834 29107 ne
rect 28834 29106 28962 29107
tri 28834 29105 28835 29106 ne
rect 28835 29105 28962 29106
tri 28835 29060 28880 29105 ne
rect 28880 29070 28962 29105
rect 29008 29105 29092 29116
tri 29092 29105 29111 29124 sw
rect 29008 29070 29111 29105
rect 28880 29060 29111 29070
tri 29111 29060 29156 29105 sw
rect 70802 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
tri 28880 29054 28886 29060 ne
rect 28886 29054 29156 29060
tri 28886 29009 28931 29054 ne
rect 28931 29015 29156 29054
tri 29156 29015 29201 29060 sw
rect 70802 29036 71000 29094
rect 28931 29009 29201 29015
tri 28931 28964 28976 29009 ne
rect 28976 28984 29201 29009
rect 28976 28964 29094 28984
tri 28976 28932 29008 28964 ne
rect 29008 28938 29094 28964
rect 29140 28970 29201 28984
tri 29201 28970 29246 29015 sw
rect 70802 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 29140 28964 29246 28970
tri 29246 28964 29252 28970 sw
rect 29140 28938 29252 28964
rect 29008 28932 29252 28938
tri 29008 28931 29009 28932 ne
rect 29009 28931 29252 28932
tri 29009 28930 29010 28931 ne
rect 29010 28930 29252 28931
tri 29010 28929 29011 28930 ne
rect 29011 28929 29252 28930
tri 29011 28928 29012 28929 ne
rect 29012 28928 29252 28929
tri 29012 28927 29013 28928 ne
rect 29013 28927 29252 28928
tri 29013 28926 29014 28927 ne
rect 29014 28926 29252 28927
tri 29014 28925 29015 28926 ne
rect 29015 28925 29252 28926
tri 29015 28924 29016 28925 ne
rect 29016 28924 29252 28925
tri 29016 28923 29017 28924 ne
rect 29017 28923 29252 28924
tri 29017 28922 29018 28923 ne
rect 29018 28922 29252 28923
tri 29018 28921 29019 28922 ne
rect 29019 28921 29252 28922
tri 29019 28920 29020 28921 ne
rect 29020 28920 29252 28921
tri 29020 28919 29021 28920 ne
rect 29021 28919 29252 28920
tri 29252 28919 29297 28964 sw
rect 70802 28932 71000 28990
tri 29021 28918 29022 28919 ne
rect 29022 28918 29297 28919
tri 29022 28917 29023 28918 ne
rect 29023 28917 29297 28918
tri 29023 28916 29024 28917 ne
rect 29024 28916 29297 28917
tri 29024 28915 29025 28916 ne
rect 29025 28915 29297 28916
tri 29025 28914 29026 28915 ne
rect 29026 28914 29297 28915
tri 29026 28913 29027 28914 ne
rect 29027 28913 29297 28914
tri 29027 28912 29028 28913 ne
rect 29028 28912 29297 28913
tri 29028 28911 29029 28912 ne
rect 29029 28911 29297 28912
tri 29029 28910 29030 28911 ne
rect 29030 28910 29297 28911
tri 29030 28909 29031 28910 ne
rect 29031 28909 29297 28910
tri 29031 28908 29032 28909 ne
rect 29032 28908 29297 28909
tri 29032 28907 29033 28908 ne
rect 29033 28907 29297 28908
tri 29033 28906 29034 28907 ne
rect 29034 28906 29297 28907
tri 29034 28905 29035 28906 ne
rect 29035 28905 29297 28906
tri 29035 28904 29036 28905 ne
rect 29036 28904 29297 28905
tri 29036 28903 29037 28904 ne
rect 29037 28903 29297 28904
tri 29037 28902 29038 28903 ne
rect 29038 28902 29297 28903
tri 29038 28901 29039 28902 ne
rect 29039 28901 29297 28902
tri 29039 28900 29040 28901 ne
rect 29040 28900 29297 28901
tri 29040 28899 29041 28900 ne
rect 29041 28899 29297 28900
tri 29041 28898 29042 28899 ne
rect 29042 28898 29297 28899
tri 29042 28897 29043 28898 ne
rect 29043 28897 29297 28898
tri 29043 28896 29044 28897 ne
rect 29044 28896 29297 28897
tri 29044 28895 29045 28896 ne
rect 29045 28895 29297 28896
tri 29045 28894 29046 28895 ne
rect 29046 28894 29297 28895
tri 29046 28893 29047 28894 ne
rect 29047 28893 29297 28894
tri 29047 28892 29048 28893 ne
rect 29048 28892 29297 28893
tri 29048 28891 29049 28892 ne
rect 29049 28891 29297 28892
tri 29049 28890 29050 28891 ne
rect 29050 28890 29297 28891
tri 29050 28889 29051 28890 ne
rect 29051 28889 29297 28890
tri 29051 28888 29052 28889 ne
rect 29052 28888 29297 28889
tri 29052 28887 29053 28888 ne
rect 29053 28887 29297 28888
tri 29053 28886 29054 28887 ne
rect 29054 28886 29297 28887
tri 29054 28885 29055 28886 ne
rect 29055 28885 29297 28886
tri 29055 28884 29056 28885 ne
rect 29056 28884 29297 28885
tri 29056 28883 29057 28884 ne
rect 29057 28883 29297 28884
tri 29057 28882 29058 28883 ne
rect 29058 28882 29297 28883
tri 29058 28881 29059 28882 ne
rect 29059 28881 29297 28882
tri 29059 28880 29060 28881 ne
rect 29060 28880 29297 28881
tri 29060 28879 29061 28880 ne
rect 29061 28879 29297 28880
tri 29061 28878 29062 28879 ne
rect 29062 28878 29297 28879
tri 29062 28877 29063 28878 ne
rect 29063 28877 29297 28878
tri 29063 28876 29064 28877 ne
rect 29064 28876 29297 28877
tri 29064 28875 29065 28876 ne
rect 29065 28875 29297 28876
tri 29065 28874 29066 28875 ne
rect 29066 28874 29297 28875
tri 29297 28874 29342 28919 sw
rect 70802 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29066 28873 29067 28874 ne
rect 29067 28873 29342 28874
tri 29067 28872 29068 28873 ne
rect 29068 28872 29342 28873
tri 29068 28871 29069 28872 ne
rect 29069 28871 29342 28872
tri 29069 28870 29070 28871 ne
rect 29070 28870 29342 28871
tri 29070 28869 29071 28870 ne
rect 29071 28869 29342 28870
tri 29071 28868 29072 28869 ne
rect 29072 28868 29342 28869
tri 29072 28867 29073 28868 ne
rect 29073 28867 29342 28868
tri 29073 28866 29074 28867 ne
rect 29074 28866 29342 28867
tri 29074 28865 29075 28866 ne
rect 29075 28865 29342 28866
tri 29075 28864 29076 28865 ne
rect 29076 28864 29342 28865
tri 29076 28863 29077 28864 ne
rect 29077 28863 29342 28864
tri 29077 28862 29078 28863 ne
rect 29078 28862 29342 28863
tri 29078 28861 29079 28862 ne
rect 29079 28861 29342 28862
tri 29079 28860 29080 28861 ne
rect 29080 28860 29342 28861
tri 29080 28859 29081 28860 ne
rect 29081 28859 29342 28860
tri 29081 28858 29082 28859 ne
rect 29082 28858 29342 28859
tri 29082 28857 29083 28858 ne
rect 29083 28857 29342 28858
tri 29083 28856 29084 28857 ne
rect 29084 28856 29342 28857
tri 29084 28855 29085 28856 ne
rect 29085 28855 29342 28856
tri 29085 28854 29086 28855 ne
rect 29086 28854 29342 28855
tri 29086 28853 29087 28854 ne
rect 29087 28853 29342 28854
tri 29087 28852 29088 28853 ne
rect 29088 28852 29342 28853
tri 29088 28851 29089 28852 ne
rect 29089 28851 29226 28852
tri 29089 28850 29090 28851 ne
rect 29090 28850 29226 28851
tri 29090 28849 29091 28850 ne
rect 29091 28849 29226 28850
tri 29091 28848 29092 28849 ne
rect 29092 28848 29226 28849
tri 29092 28847 29093 28848 ne
rect 29093 28847 29226 28848
tri 29093 28846 29094 28847 ne
rect 29094 28846 29226 28847
tri 29094 28845 29095 28846 ne
rect 29095 28845 29226 28846
tri 29095 28844 29096 28845 ne
rect 29096 28844 29226 28845
tri 29096 28843 29097 28844 ne
rect 29097 28843 29226 28844
tri 29097 28842 29098 28843 ne
rect 29098 28842 29226 28843
tri 29098 28841 29099 28842 ne
rect 29099 28841 29226 28842
tri 29099 28840 29100 28841 ne
rect 29100 28840 29226 28841
tri 29100 28839 29101 28840 ne
rect 29101 28839 29226 28840
tri 29101 28838 29102 28839 ne
rect 29102 28838 29226 28839
tri 29102 28837 29103 28838 ne
rect 29103 28837 29226 28838
tri 29103 28836 29104 28837 ne
rect 29104 28836 29226 28837
tri 29104 28835 29105 28836 ne
rect 29105 28835 29226 28836
tri 29105 28834 29106 28835 ne
rect 29106 28834 29226 28835
tri 29106 28833 29107 28834 ne
rect 29107 28833 29226 28834
tri 29107 28832 29108 28833 ne
rect 29108 28832 29226 28833
tri 29108 28831 29109 28832 ne
rect 29109 28831 29226 28832
tri 29109 28830 29110 28831 ne
rect 29110 28830 29226 28831
tri 29110 28829 29111 28830 ne
rect 29111 28829 29226 28830
tri 29111 28803 29137 28829 ne
rect 29137 28806 29226 28829
rect 29272 28829 29342 28852
tri 29342 28829 29387 28874 sw
rect 29272 28806 29387 28829
rect 29137 28803 29387 28806
tri 29387 28803 29413 28829 sw
rect 70802 28828 71000 28886
tri 29137 28758 29182 28803 ne
rect 29182 28758 29413 28803
tri 29413 28758 29458 28803 sw
rect 70802 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
tri 29182 28735 29205 28758 ne
rect 29205 28735 29458 28758
tri 29205 28690 29250 28735 ne
rect 29250 28720 29458 28735
rect 29250 28690 29358 28720
tri 29250 28657 29283 28690 ne
rect 29283 28674 29358 28690
rect 29404 28713 29458 28720
tri 29458 28713 29503 28758 sw
rect 70802 28724 71000 28782
rect 29404 28674 29503 28713
rect 29283 28668 29503 28674
tri 29503 28668 29548 28713 sw
rect 70802 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 29283 28657 29548 28668
tri 29283 28656 29284 28657 ne
rect 29284 28656 29548 28657
tri 29284 28655 29285 28656 ne
rect 29285 28655 29548 28656
tri 29285 28654 29286 28655 ne
rect 29286 28654 29548 28655
tri 29286 28653 29287 28654 ne
rect 29287 28653 29548 28654
tri 29287 28652 29288 28653 ne
rect 29288 28652 29548 28653
tri 29288 28651 29289 28652 ne
rect 29289 28651 29548 28652
tri 29289 28650 29290 28651 ne
rect 29290 28650 29548 28651
tri 29290 28649 29291 28650 ne
rect 29291 28649 29548 28650
tri 29291 28648 29292 28649 ne
rect 29292 28648 29548 28649
tri 29292 28647 29293 28648 ne
rect 29293 28647 29548 28648
tri 29293 28646 29294 28647 ne
rect 29294 28646 29548 28647
tri 29294 28645 29295 28646 ne
rect 29295 28645 29548 28646
tri 29295 28644 29296 28645 ne
rect 29296 28644 29548 28645
tri 29296 28643 29297 28644 ne
rect 29297 28643 29548 28644
tri 29548 28643 29573 28668 sw
tri 29297 28642 29298 28643 ne
rect 29298 28642 29573 28643
tri 29298 28641 29299 28642 ne
rect 29299 28641 29573 28642
tri 29299 28640 29300 28641 ne
rect 29300 28640 29573 28641
tri 29300 28639 29301 28640 ne
rect 29301 28639 29573 28640
tri 29301 28638 29302 28639 ne
rect 29302 28638 29573 28639
tri 29302 28637 29303 28638 ne
rect 29303 28637 29573 28638
tri 29303 28636 29304 28637 ne
rect 29304 28636 29573 28637
tri 29304 28635 29305 28636 ne
rect 29305 28635 29573 28636
tri 29305 28634 29306 28635 ne
rect 29306 28634 29573 28635
tri 29306 28633 29307 28634 ne
rect 29307 28633 29573 28634
tri 29307 28632 29308 28633 ne
rect 29308 28632 29573 28633
tri 29308 28631 29309 28632 ne
rect 29309 28631 29573 28632
tri 29309 28630 29310 28631 ne
rect 29310 28630 29573 28631
tri 29310 28629 29311 28630 ne
rect 29311 28629 29573 28630
tri 29311 28628 29312 28629 ne
rect 29312 28628 29573 28629
tri 29312 28627 29313 28628 ne
rect 29313 28627 29573 28628
tri 29313 28626 29314 28627 ne
rect 29314 28626 29573 28627
tri 29314 28625 29315 28626 ne
rect 29315 28625 29573 28626
tri 29315 28624 29316 28625 ne
rect 29316 28624 29573 28625
tri 29316 28623 29317 28624 ne
rect 29317 28623 29573 28624
tri 29317 28622 29318 28623 ne
rect 29318 28622 29573 28623
tri 29318 28621 29319 28622 ne
rect 29319 28621 29573 28622
tri 29319 28620 29320 28621 ne
rect 29320 28620 29573 28621
tri 29320 28619 29321 28620 ne
rect 29321 28619 29573 28620
tri 29321 28618 29322 28619 ne
rect 29322 28618 29573 28619
tri 29322 28617 29323 28618 ne
rect 29323 28617 29573 28618
tri 29323 28616 29324 28617 ne
rect 29324 28616 29573 28617
tri 29324 28615 29325 28616 ne
rect 29325 28615 29573 28616
tri 29325 28614 29326 28615 ne
rect 29326 28614 29573 28615
tri 29326 28613 29327 28614 ne
rect 29327 28613 29573 28614
tri 29327 28612 29328 28613 ne
rect 29328 28612 29573 28613
tri 29328 28611 29329 28612 ne
rect 29329 28611 29573 28612
tri 29329 28610 29330 28611 ne
rect 29330 28610 29573 28611
tri 29330 28609 29331 28610 ne
rect 29331 28609 29573 28610
tri 29331 28608 29332 28609 ne
rect 29332 28608 29573 28609
tri 29332 28607 29333 28608 ne
rect 29333 28607 29573 28608
tri 29333 28606 29334 28607 ne
rect 29334 28606 29573 28607
tri 29334 28605 29335 28606 ne
rect 29335 28605 29573 28606
tri 29335 28604 29336 28605 ne
rect 29336 28604 29573 28605
tri 29336 28603 29337 28604 ne
rect 29337 28603 29573 28604
tri 29337 28602 29338 28603 ne
rect 29338 28602 29573 28603
tri 29338 28601 29339 28602 ne
rect 29339 28601 29573 28602
tri 29339 28600 29340 28601 ne
rect 29340 28600 29573 28601
tri 29340 28599 29341 28600 ne
rect 29341 28599 29573 28600
tri 29341 28598 29342 28599 ne
rect 29342 28598 29573 28599
tri 29573 28598 29618 28643 sw
rect 70802 28620 71000 28678
tri 29342 28597 29343 28598 ne
rect 29343 28597 29618 28598
tri 29343 28596 29344 28597 ne
rect 29344 28596 29618 28597
tri 29344 28595 29345 28596 ne
rect 29345 28595 29618 28596
tri 29345 28594 29346 28595 ne
rect 29346 28594 29618 28595
tri 29346 28593 29347 28594 ne
rect 29347 28593 29618 28594
tri 29347 28592 29348 28593 ne
rect 29348 28592 29618 28593
tri 29348 28591 29349 28592 ne
rect 29349 28591 29618 28592
tri 29349 28590 29350 28591 ne
rect 29350 28590 29618 28591
tri 29350 28589 29351 28590 ne
rect 29351 28589 29618 28590
tri 29351 28588 29352 28589 ne
rect 29352 28588 29618 28589
tri 29352 28587 29353 28588 ne
rect 29353 28587 29490 28588
tri 29353 28586 29354 28587 ne
rect 29354 28586 29490 28587
tri 29354 28585 29355 28586 ne
rect 29355 28585 29490 28586
tri 29355 28584 29356 28585 ne
rect 29356 28584 29490 28585
tri 29356 28583 29357 28584 ne
rect 29357 28583 29490 28584
tri 29357 28582 29358 28583 ne
rect 29358 28582 29490 28583
tri 29358 28581 29359 28582 ne
rect 29359 28581 29490 28582
tri 29359 28580 29360 28581 ne
rect 29360 28580 29490 28581
tri 29360 28579 29361 28580 ne
rect 29361 28579 29490 28580
tri 29361 28578 29362 28579 ne
rect 29362 28578 29490 28579
tri 29362 28577 29363 28578 ne
rect 29363 28577 29490 28578
tri 29363 28576 29364 28577 ne
rect 29364 28576 29490 28577
tri 29364 28575 29365 28576 ne
rect 29365 28575 29490 28576
tri 29365 28574 29366 28575 ne
rect 29366 28574 29490 28575
tri 29366 28573 29367 28574 ne
rect 29367 28573 29490 28574
tri 29367 28572 29368 28573 ne
rect 29368 28572 29490 28573
tri 29368 28571 29369 28572 ne
rect 29369 28571 29490 28572
tri 29369 28570 29370 28571 ne
rect 29370 28570 29490 28571
tri 29370 28569 29371 28570 ne
rect 29371 28569 29490 28570
tri 29371 28568 29372 28569 ne
rect 29372 28568 29490 28569
tri 29372 28567 29373 28568 ne
rect 29373 28567 29490 28568
tri 29373 28566 29374 28567 ne
rect 29374 28566 29490 28567
tri 29374 28565 29375 28566 ne
rect 29375 28565 29490 28566
tri 29375 28564 29376 28565 ne
rect 29376 28564 29490 28565
tri 29376 28563 29377 28564 ne
rect 29377 28563 29490 28564
tri 29377 28562 29378 28563 ne
rect 29378 28562 29490 28563
tri 29378 28561 29379 28562 ne
rect 29379 28561 29490 28562
tri 29379 28560 29380 28561 ne
rect 29380 28560 29490 28561
tri 29380 28559 29381 28560 ne
rect 29381 28559 29490 28560
tri 29381 28558 29382 28559 ne
rect 29382 28558 29490 28559
tri 29382 28557 29383 28558 ne
rect 29383 28557 29490 28558
tri 29383 28556 29384 28557 ne
rect 29384 28556 29490 28557
tri 29384 28555 29385 28556 ne
rect 29385 28555 29490 28556
tri 29385 28554 29386 28555 ne
rect 29386 28554 29490 28555
tri 29386 28553 29387 28554 ne
rect 29387 28553 29490 28554
tri 29387 28508 29432 28553 ne
rect 29432 28542 29490 28553
rect 29536 28553 29618 28588
tri 29618 28553 29663 28598 sw
rect 70802 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28542 29663 28553
rect 29432 28508 29663 28542
tri 29663 28508 29708 28553 sw
rect 70802 28516 71000 28574
tri 29432 28482 29458 28508 ne
rect 29458 28482 29708 28508
tri 29708 28482 29734 28508 sw
tri 29458 28463 29477 28482 ne
rect 29477 28463 29734 28482
tri 29477 28437 29503 28463 ne
rect 29503 28456 29734 28463
rect 29503 28437 29622 28456
tri 29503 28392 29548 28437 ne
rect 29548 28410 29622 28437
rect 29668 28437 29734 28456
tri 29734 28437 29779 28482 sw
rect 70802 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29668 28410 29779 28437
rect 29548 28392 29779 28410
tri 29779 28392 29824 28437 sw
rect 70802 28412 71000 28470
tri 29548 28383 29557 28392 ne
rect 29557 28383 29824 28392
tri 29557 28382 29558 28383 ne
rect 29558 28382 29824 28383
tri 29558 28381 29559 28382 ne
rect 29559 28381 29824 28382
tri 29559 28380 29560 28381 ne
rect 29560 28380 29824 28381
tri 29560 28379 29561 28380 ne
rect 29561 28379 29824 28380
tri 29561 28378 29562 28379 ne
rect 29562 28378 29824 28379
tri 29562 28377 29563 28378 ne
rect 29563 28377 29824 28378
tri 29563 28376 29564 28377 ne
rect 29564 28376 29824 28377
tri 29564 28375 29565 28376 ne
rect 29565 28375 29824 28376
tri 29565 28374 29566 28375 ne
rect 29566 28374 29824 28375
tri 29566 28373 29567 28374 ne
rect 29567 28373 29824 28374
tri 29567 28372 29568 28373 ne
rect 29568 28372 29824 28373
tri 29568 28371 29569 28372 ne
rect 29569 28371 29824 28372
tri 29569 28370 29570 28371 ne
rect 29570 28370 29824 28371
tri 29570 28369 29571 28370 ne
rect 29571 28369 29824 28370
tri 29571 28368 29572 28369 ne
rect 29572 28368 29824 28369
tri 29572 28367 29573 28368 ne
rect 29573 28367 29824 28368
tri 29573 28366 29574 28367 ne
rect 29574 28366 29824 28367
tri 29574 28365 29575 28366 ne
rect 29575 28365 29824 28366
tri 29575 28364 29576 28365 ne
rect 29576 28364 29824 28365
tri 29576 28363 29577 28364 ne
rect 29577 28363 29824 28364
tri 29577 28362 29578 28363 ne
rect 29578 28362 29824 28363
tri 29578 28361 29579 28362 ne
rect 29579 28361 29824 28362
tri 29579 28360 29580 28361 ne
rect 29580 28360 29824 28361
tri 29580 28359 29581 28360 ne
rect 29581 28359 29824 28360
tri 29581 28358 29582 28359 ne
rect 29582 28358 29824 28359
tri 29582 28357 29583 28358 ne
rect 29583 28357 29824 28358
tri 29583 28356 29584 28357 ne
rect 29584 28356 29824 28357
tri 29584 28355 29585 28356 ne
rect 29585 28355 29824 28356
tri 29585 28354 29586 28355 ne
rect 29586 28354 29824 28355
tri 29586 28353 29587 28354 ne
rect 29587 28353 29824 28354
tri 29587 28352 29588 28353 ne
rect 29588 28352 29824 28353
tri 29588 28351 29589 28352 ne
rect 29589 28351 29824 28352
tri 29589 28350 29590 28351 ne
rect 29590 28350 29824 28351
tri 29590 28349 29591 28350 ne
rect 29591 28349 29824 28350
tri 29591 28348 29592 28349 ne
rect 29592 28348 29824 28349
tri 29592 28347 29593 28348 ne
rect 29593 28347 29824 28348
tri 29824 28347 29869 28392 sw
rect 70802 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29593 28346 29594 28347 ne
rect 29594 28346 29869 28347
tri 29594 28345 29595 28346 ne
rect 29595 28345 29869 28346
tri 29595 28344 29596 28345 ne
rect 29596 28344 29869 28345
tri 29596 28343 29597 28344 ne
rect 29597 28343 29869 28344
tri 29597 28342 29598 28343 ne
rect 29598 28342 29869 28343
tri 29598 28341 29599 28342 ne
rect 29599 28341 29869 28342
tri 29599 28340 29600 28341 ne
rect 29600 28340 29869 28341
tri 29600 28339 29601 28340 ne
rect 29601 28339 29869 28340
tri 29601 28338 29602 28339 ne
rect 29602 28338 29869 28339
tri 29602 28337 29603 28338 ne
rect 29603 28337 29869 28338
tri 29603 28336 29604 28337 ne
rect 29604 28336 29869 28337
tri 29604 28335 29605 28336 ne
rect 29605 28335 29869 28336
tri 29605 28334 29606 28335 ne
rect 29606 28334 29869 28335
tri 29606 28333 29607 28334 ne
rect 29607 28333 29869 28334
tri 29607 28332 29608 28333 ne
rect 29608 28332 29869 28333
tri 29608 28331 29609 28332 ne
rect 29609 28331 29869 28332
tri 29609 28330 29610 28331 ne
rect 29610 28330 29869 28331
tri 29610 28329 29611 28330 ne
rect 29611 28329 29869 28330
tri 29611 28328 29612 28329 ne
rect 29612 28328 29869 28329
tri 29612 28327 29613 28328 ne
rect 29613 28327 29869 28328
tri 29613 28326 29614 28327 ne
rect 29614 28326 29869 28327
tri 29614 28325 29615 28326 ne
rect 29615 28325 29869 28326
tri 29615 28324 29616 28325 ne
rect 29616 28324 29869 28325
tri 29616 28323 29617 28324 ne
rect 29617 28323 29754 28324
tri 29617 28322 29618 28323 ne
rect 29618 28322 29754 28323
tri 29618 28321 29619 28322 ne
rect 29619 28321 29754 28322
tri 29619 28320 29620 28321 ne
rect 29620 28320 29754 28321
tri 29620 28319 29621 28320 ne
rect 29621 28319 29754 28320
tri 29621 28318 29622 28319 ne
rect 29622 28318 29754 28319
tri 29622 28317 29623 28318 ne
rect 29623 28317 29754 28318
tri 29623 28316 29624 28317 ne
rect 29624 28316 29754 28317
tri 29624 28315 29625 28316 ne
rect 29625 28315 29754 28316
tri 29625 28314 29626 28315 ne
rect 29626 28314 29754 28315
tri 29626 28313 29627 28314 ne
rect 29627 28313 29754 28314
tri 29627 28312 29628 28313 ne
rect 29628 28312 29754 28313
tri 29628 28311 29629 28312 ne
rect 29629 28311 29754 28312
tri 29629 28310 29630 28311 ne
rect 29630 28310 29754 28311
tri 29630 28309 29631 28310 ne
rect 29631 28309 29754 28310
tri 29631 28308 29632 28309 ne
rect 29632 28308 29754 28309
tri 29632 28307 29633 28308 ne
rect 29633 28307 29754 28308
tri 29633 28306 29634 28307 ne
rect 29634 28306 29754 28307
tri 29634 28305 29635 28306 ne
rect 29635 28305 29754 28306
tri 29635 28304 29636 28305 ne
rect 29636 28304 29754 28305
tri 29636 28303 29637 28304 ne
rect 29637 28303 29754 28304
tri 29637 28302 29638 28303 ne
rect 29638 28302 29754 28303
tri 29638 28301 29639 28302 ne
rect 29639 28301 29754 28302
tri 29639 28300 29640 28301 ne
rect 29640 28300 29754 28301
tri 29640 28299 29641 28300 ne
rect 29641 28299 29754 28300
tri 29641 28298 29642 28299 ne
rect 29642 28298 29754 28299
tri 29642 28297 29643 28298 ne
rect 29643 28297 29754 28298
tri 29643 28296 29644 28297 ne
rect 29644 28296 29754 28297
tri 29644 28295 29645 28296 ne
rect 29645 28295 29754 28296
tri 29645 28294 29646 28295 ne
rect 29646 28294 29754 28295
tri 29646 28293 29647 28294 ne
rect 29647 28293 29754 28294
tri 29647 28292 29648 28293 ne
rect 29648 28292 29754 28293
tri 29648 28291 29649 28292 ne
rect 29649 28291 29754 28292
tri 29649 28290 29650 28291 ne
rect 29650 28290 29754 28291
tri 29650 28289 29651 28290 ne
rect 29651 28289 29754 28290
tri 29651 28288 29652 28289 ne
rect 29652 28288 29754 28289
tri 29652 28287 29653 28288 ne
rect 29653 28287 29754 28288
tri 29653 28286 29654 28287 ne
rect 29654 28286 29754 28287
tri 29654 28285 29655 28286 ne
rect 29655 28285 29754 28286
tri 29655 28284 29656 28285 ne
rect 29656 28284 29754 28285
tri 29656 28283 29657 28284 ne
rect 29657 28283 29754 28284
tri 29657 28282 29658 28283 ne
rect 29658 28282 29754 28283
tri 29658 28281 29659 28282 ne
rect 29659 28281 29754 28282
tri 29659 28280 29660 28281 ne
rect 29660 28280 29754 28281
tri 29660 28279 29661 28280 ne
rect 29661 28279 29754 28280
tri 29661 28278 29662 28279 ne
rect 29662 28278 29754 28279
rect 29800 28322 29869 28324
tri 29869 28322 29894 28347 sw
rect 29800 28278 29894 28322
tri 29662 28277 29663 28278 ne
rect 29663 28277 29894 28278
tri 29894 28277 29939 28322 sw
rect 70802 28308 71000 28366
tri 29663 28232 29708 28277 ne
rect 29708 28232 29939 28277
tri 29939 28232 29984 28277 sw
rect 70802 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
tri 29708 28187 29753 28232 ne
rect 29753 28192 29984 28232
rect 29753 28187 29886 28192
tri 29753 28142 29798 28187 ne
rect 29798 28146 29886 28187
rect 29932 28187 29984 28192
tri 29984 28187 30029 28232 sw
rect 70802 28204 71000 28262
rect 29932 28161 30029 28187
tri 30029 28161 30055 28187 sw
rect 29932 28146 30055 28161
rect 29798 28142 30055 28146
tri 29798 28116 29824 28142 ne
rect 29824 28116 30055 28142
tri 30055 28116 30100 28161 sw
rect 70802 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
tri 29824 28109 29831 28116 ne
rect 29831 28109 30100 28116
tri 29831 28108 29832 28109 ne
rect 29832 28108 30100 28109
tri 29832 28107 29833 28108 ne
rect 29833 28107 30100 28108
tri 29833 28106 29834 28107 ne
rect 29834 28106 30100 28107
tri 29834 28105 29835 28106 ne
rect 29835 28105 30100 28106
tri 29835 28104 29836 28105 ne
rect 29836 28104 30100 28105
tri 29836 28103 29837 28104 ne
rect 29837 28103 30100 28104
tri 29837 28102 29838 28103 ne
rect 29838 28102 30100 28103
tri 29838 28101 29839 28102 ne
rect 29839 28101 30100 28102
tri 29839 28100 29840 28101 ne
rect 29840 28100 30100 28101
tri 29840 28099 29841 28100 ne
rect 29841 28099 30100 28100
tri 29841 28098 29842 28099 ne
rect 29842 28098 30100 28099
tri 29842 28097 29843 28098 ne
rect 29843 28097 30100 28098
tri 29843 28096 29844 28097 ne
rect 29844 28096 30100 28097
tri 29844 28095 29845 28096 ne
rect 29845 28095 30100 28096
tri 29845 28094 29846 28095 ne
rect 29846 28094 30100 28095
tri 29846 28093 29847 28094 ne
rect 29847 28093 30100 28094
tri 29847 28092 29848 28093 ne
rect 29848 28092 30100 28093
tri 29848 28091 29849 28092 ne
rect 29849 28091 30100 28092
tri 29849 28090 29850 28091 ne
rect 29850 28090 30100 28091
tri 29850 28089 29851 28090 ne
rect 29851 28089 30100 28090
tri 29851 28088 29852 28089 ne
rect 29852 28088 30100 28089
tri 29852 28087 29853 28088 ne
rect 29853 28087 30100 28088
tri 29853 28086 29854 28087 ne
rect 29854 28086 30100 28087
tri 29854 28085 29855 28086 ne
rect 29855 28085 30100 28086
tri 29855 28084 29856 28085 ne
rect 29856 28084 30100 28085
tri 29856 28083 29857 28084 ne
rect 29857 28083 30100 28084
tri 29857 28082 29858 28083 ne
rect 29858 28082 30100 28083
tri 29858 28081 29859 28082 ne
rect 29859 28081 30100 28082
tri 29859 28080 29860 28081 ne
rect 29860 28080 30100 28081
tri 29860 28079 29861 28080 ne
rect 29861 28079 30100 28080
tri 29861 28078 29862 28079 ne
rect 29862 28078 30100 28079
tri 29862 28077 29863 28078 ne
rect 29863 28077 30100 28078
tri 29863 28076 29864 28077 ne
rect 29864 28076 30100 28077
tri 29864 28075 29865 28076 ne
rect 29865 28075 30100 28076
tri 29865 28074 29866 28075 ne
rect 29866 28074 30100 28075
tri 29866 28073 29867 28074 ne
rect 29867 28073 30100 28074
tri 29867 28072 29868 28073 ne
rect 29868 28072 30100 28073
tri 29868 28071 29869 28072 ne
rect 29869 28071 30100 28072
tri 30100 28071 30145 28116 sw
rect 70802 28100 71000 28158
tri 29869 28070 29870 28071 ne
rect 29870 28070 30145 28071
tri 29870 28069 29871 28070 ne
rect 29871 28069 30145 28070
tri 29871 28068 29872 28069 ne
rect 29872 28068 30145 28069
tri 29872 28067 29873 28068 ne
rect 29873 28067 30145 28068
tri 29873 28066 29874 28067 ne
rect 29874 28066 30145 28067
tri 29874 28065 29875 28066 ne
rect 29875 28065 30145 28066
tri 29875 28064 29876 28065 ne
rect 29876 28064 30145 28065
tri 29876 28063 29877 28064 ne
rect 29877 28063 30145 28064
tri 29877 28062 29878 28063 ne
rect 29878 28062 30145 28063
tri 29878 28061 29879 28062 ne
rect 29879 28061 30145 28062
tri 29879 28060 29880 28061 ne
rect 29880 28060 30145 28061
tri 29880 28059 29881 28060 ne
rect 29881 28059 30018 28060
tri 29881 28058 29882 28059 ne
rect 29882 28058 30018 28059
tri 29882 28057 29883 28058 ne
rect 29883 28057 30018 28058
tri 29883 28056 29884 28057 ne
rect 29884 28056 30018 28057
tri 29884 28055 29885 28056 ne
rect 29885 28055 30018 28056
tri 29885 28054 29886 28055 ne
rect 29886 28054 30018 28055
tri 29886 28053 29887 28054 ne
rect 29887 28053 30018 28054
tri 29887 28052 29888 28053 ne
rect 29888 28052 30018 28053
tri 29888 28051 29889 28052 ne
rect 29889 28051 30018 28052
tri 29889 28050 29890 28051 ne
rect 29890 28050 30018 28051
tri 29890 28049 29891 28050 ne
rect 29891 28049 30018 28050
tri 29891 28048 29892 28049 ne
rect 29892 28048 30018 28049
tri 29892 28047 29893 28048 ne
rect 29893 28047 30018 28048
tri 29893 28046 29894 28047 ne
rect 29894 28046 30018 28047
tri 29894 28045 29895 28046 ne
rect 29895 28045 30018 28046
tri 29895 28044 29896 28045 ne
rect 29896 28044 30018 28045
tri 29896 28043 29897 28044 ne
rect 29897 28043 30018 28044
tri 29897 28042 29898 28043 ne
rect 29898 28042 30018 28043
tri 29898 28041 29899 28042 ne
rect 29899 28041 30018 28042
tri 29899 28040 29900 28041 ne
rect 29900 28040 30018 28041
tri 29900 28039 29901 28040 ne
rect 29901 28039 30018 28040
tri 29901 28038 29902 28039 ne
rect 29902 28038 30018 28039
tri 29902 28037 29903 28038 ne
rect 29903 28037 30018 28038
tri 29903 28036 29904 28037 ne
rect 29904 28036 30018 28037
tri 29904 28035 29905 28036 ne
rect 29905 28035 30018 28036
tri 29905 28034 29906 28035 ne
rect 29906 28034 30018 28035
tri 29906 28033 29907 28034 ne
rect 29907 28033 30018 28034
tri 29907 28032 29908 28033 ne
rect 29908 28032 30018 28033
tri 29908 28031 29909 28032 ne
rect 29909 28031 30018 28032
tri 29909 28030 29910 28031 ne
rect 29910 28030 30018 28031
tri 29910 28029 29911 28030 ne
rect 29911 28029 30018 28030
tri 29911 28028 29912 28029 ne
rect 29912 28028 30018 28029
tri 29912 28027 29913 28028 ne
rect 29913 28027 30018 28028
tri 29913 28026 29914 28027 ne
rect 29914 28026 30018 28027
tri 29914 28025 29915 28026 ne
rect 29915 28025 30018 28026
tri 29915 28024 29916 28025 ne
rect 29916 28024 30018 28025
tri 29916 28023 29917 28024 ne
rect 29917 28023 30018 28024
tri 29917 28022 29918 28023 ne
rect 29918 28022 30018 28023
tri 29918 28021 29919 28022 ne
rect 29919 28021 30018 28022
tri 29919 28020 29920 28021 ne
rect 29920 28020 30018 28021
tri 29920 28019 29921 28020 ne
rect 29921 28019 30018 28020
tri 29921 28018 29922 28019 ne
rect 29922 28018 30018 28019
tri 29922 28017 29923 28018 ne
rect 29923 28017 30018 28018
tri 29923 28016 29924 28017 ne
rect 29924 28016 30018 28017
tri 29924 28015 29925 28016 ne
rect 29925 28015 30018 28016
tri 29925 28014 29926 28015 ne
rect 29926 28014 30018 28015
rect 30064 28026 30145 28060
tri 30145 28026 30190 28071 sw
rect 70802 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28014 30190 28026
tri 29926 28013 29927 28014 ne
rect 29927 28013 30190 28014
tri 29927 28012 29928 28013 ne
rect 29928 28012 30190 28013
tri 29928 28011 29929 28012 ne
rect 29929 28011 30190 28012
tri 29929 28010 29930 28011 ne
rect 29930 28010 30190 28011
tri 29930 28009 29931 28010 ne
rect 29931 28009 30190 28010
tri 29931 28008 29932 28009 ne
rect 29932 28008 30190 28009
tri 29932 28007 29933 28008 ne
rect 29933 28007 30190 28008
tri 29933 28006 29934 28007 ne
rect 29934 28006 30190 28007
tri 29934 28005 29935 28006 ne
rect 29935 28005 30190 28006
tri 29935 28004 29936 28005 ne
rect 29936 28004 30190 28005
tri 29936 28003 29937 28004 ne
rect 29937 28003 30190 28004
tri 29937 28002 29938 28003 ne
rect 29938 28002 30190 28003
tri 29938 28001 29939 28002 ne
rect 29939 28001 30190 28002
tri 30190 28001 30215 28026 sw
tri 29939 27960 29980 28001 ne
rect 29980 27960 30215 28001
tri 29980 27915 30025 27960 ne
rect 30025 27956 30215 27960
tri 30215 27956 30260 28001 sw
rect 70802 27996 71000 28054
rect 30025 27928 30260 27956
rect 30025 27915 30150 27928
tri 30025 27870 30070 27915 ne
rect 30070 27882 30150 27915
rect 30196 27911 30260 27928
tri 30260 27911 30305 27956 sw
rect 70802 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 30196 27882 30305 27911
rect 30070 27870 30305 27882
tri 30070 27834 30106 27870 ne
rect 30106 27866 30305 27870
tri 30305 27866 30350 27911 sw
rect 70802 27892 71000 27950
rect 30106 27860 30350 27866
tri 30350 27860 30356 27866 sw
rect 30106 27834 30356 27860
tri 30106 27833 30107 27834 ne
rect 30107 27833 30356 27834
tri 30107 27832 30108 27833 ne
rect 30108 27832 30356 27833
tri 30108 27831 30109 27832 ne
rect 30109 27831 30356 27832
tri 30109 27830 30110 27831 ne
rect 30110 27830 30356 27831
tri 30110 27829 30111 27830 ne
rect 30111 27829 30356 27830
tri 30111 27828 30112 27829 ne
rect 30112 27828 30356 27829
tri 30112 27827 30113 27828 ne
rect 30113 27827 30356 27828
tri 30113 27826 30114 27827 ne
rect 30114 27826 30356 27827
tri 30114 27825 30115 27826 ne
rect 30115 27825 30356 27826
tri 30115 27824 30116 27825 ne
rect 30116 27824 30356 27825
tri 30116 27823 30117 27824 ne
rect 30117 27823 30356 27824
tri 30117 27822 30118 27823 ne
rect 30118 27822 30356 27823
tri 30118 27821 30119 27822 ne
rect 30119 27821 30356 27822
tri 30119 27820 30120 27821 ne
rect 30120 27820 30356 27821
tri 30120 27819 30121 27820 ne
rect 30121 27819 30356 27820
tri 30121 27818 30122 27819 ne
rect 30122 27818 30356 27819
tri 30122 27817 30123 27818 ne
rect 30123 27817 30356 27818
tri 30123 27816 30124 27817 ne
rect 30124 27816 30356 27817
tri 30124 27815 30125 27816 ne
rect 30125 27815 30356 27816
tri 30356 27815 30401 27860 sw
rect 70802 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30125 27814 30126 27815 ne
rect 30126 27814 30401 27815
tri 30126 27813 30127 27814 ne
rect 30127 27813 30401 27814
tri 30127 27812 30128 27813 ne
rect 30128 27812 30401 27813
tri 30128 27811 30129 27812 ne
rect 30129 27811 30401 27812
tri 30129 27810 30130 27811 ne
rect 30130 27810 30401 27811
tri 30130 27809 30131 27810 ne
rect 30131 27809 30401 27810
tri 30131 27808 30132 27809 ne
rect 30132 27808 30401 27809
tri 30132 27807 30133 27808 ne
rect 30133 27807 30401 27808
tri 30133 27806 30134 27807 ne
rect 30134 27806 30401 27807
tri 30134 27805 30135 27806 ne
rect 30135 27805 30401 27806
tri 30135 27804 30136 27805 ne
rect 30136 27804 30401 27805
tri 30136 27803 30137 27804 ne
rect 30137 27803 30401 27804
tri 30137 27802 30138 27803 ne
rect 30138 27802 30401 27803
tri 30138 27801 30139 27802 ne
rect 30139 27801 30401 27802
tri 30139 27800 30140 27801 ne
rect 30140 27800 30401 27801
tri 30140 27799 30141 27800 ne
rect 30141 27799 30401 27800
tri 30141 27798 30142 27799 ne
rect 30142 27798 30401 27799
tri 30142 27797 30143 27798 ne
rect 30143 27797 30401 27798
tri 30143 27796 30144 27797 ne
rect 30144 27796 30401 27797
tri 30144 27795 30145 27796 ne
rect 30145 27795 30282 27796
tri 30145 27794 30146 27795 ne
rect 30146 27794 30282 27795
tri 30146 27793 30147 27794 ne
rect 30147 27793 30282 27794
tri 30147 27792 30148 27793 ne
rect 30148 27792 30282 27793
tri 30148 27791 30149 27792 ne
rect 30149 27791 30282 27792
tri 30149 27790 30150 27791 ne
rect 30150 27790 30282 27791
tri 30150 27789 30151 27790 ne
rect 30151 27789 30282 27790
tri 30151 27788 30152 27789 ne
rect 30152 27788 30282 27789
tri 30152 27787 30153 27788 ne
rect 30153 27787 30282 27788
tri 30153 27786 30154 27787 ne
rect 30154 27786 30282 27787
tri 30154 27785 30155 27786 ne
rect 30155 27785 30282 27786
tri 30155 27784 30156 27785 ne
rect 30156 27784 30282 27785
tri 30156 27783 30157 27784 ne
rect 30157 27783 30282 27784
tri 30157 27782 30158 27783 ne
rect 30158 27782 30282 27783
tri 30158 27781 30159 27782 ne
rect 30159 27781 30282 27782
tri 30159 27780 30160 27781 ne
rect 30160 27780 30282 27781
tri 30160 27779 30161 27780 ne
rect 30161 27779 30282 27780
tri 30161 27778 30162 27779 ne
rect 30162 27778 30282 27779
tri 30162 27777 30163 27778 ne
rect 30163 27777 30282 27778
tri 30163 27776 30164 27777 ne
rect 30164 27776 30282 27777
tri 30164 27775 30165 27776 ne
rect 30165 27775 30282 27776
tri 30165 27774 30166 27775 ne
rect 30166 27774 30282 27775
tri 30166 27773 30167 27774 ne
rect 30167 27773 30282 27774
tri 30167 27772 30168 27773 ne
rect 30168 27772 30282 27773
tri 30168 27771 30169 27772 ne
rect 30169 27771 30282 27772
tri 30169 27770 30170 27771 ne
rect 30170 27770 30282 27771
tri 30170 27769 30171 27770 ne
rect 30171 27769 30282 27770
tri 30171 27768 30172 27769 ne
rect 30172 27768 30282 27769
tri 30172 27767 30173 27768 ne
rect 30173 27767 30282 27768
tri 30173 27766 30174 27767 ne
rect 30174 27766 30282 27767
tri 30174 27765 30175 27766 ne
rect 30175 27765 30282 27766
tri 30175 27764 30176 27765 ne
rect 30176 27764 30282 27765
tri 30176 27763 30177 27764 ne
rect 30177 27763 30282 27764
tri 30177 27762 30178 27763 ne
rect 30178 27762 30282 27763
tri 30178 27761 30179 27762 ne
rect 30179 27761 30282 27762
tri 30179 27760 30180 27761 ne
rect 30180 27760 30282 27761
tri 30180 27759 30181 27760 ne
rect 30181 27759 30282 27760
tri 30181 27758 30182 27759 ne
rect 30182 27758 30282 27759
tri 30182 27757 30183 27758 ne
rect 30183 27757 30282 27758
tri 30183 27756 30184 27757 ne
rect 30184 27756 30282 27757
tri 30184 27755 30185 27756 ne
rect 30185 27755 30282 27756
tri 30185 27754 30186 27755 ne
rect 30186 27754 30282 27755
tri 30186 27753 30187 27754 ne
rect 30187 27753 30282 27754
tri 30187 27752 30188 27753 ne
rect 30188 27752 30282 27753
tri 30188 27751 30189 27752 ne
rect 30189 27751 30282 27752
tri 30189 27750 30190 27751 ne
rect 30190 27750 30282 27751
rect 30328 27770 30401 27796
tri 30401 27770 30446 27815 sw
rect 70802 27788 71000 27846
rect 30328 27750 30446 27770
tri 30190 27749 30191 27750 ne
rect 30191 27749 30446 27750
tri 30191 27748 30192 27749 ne
rect 30192 27748 30446 27749
tri 30192 27747 30193 27748 ne
rect 30193 27747 30446 27748
tri 30193 27746 30194 27747 ne
rect 30194 27746 30446 27747
tri 30194 27745 30195 27746 ne
rect 30195 27745 30446 27746
tri 30195 27744 30196 27745 ne
rect 30196 27744 30446 27745
tri 30196 27743 30197 27744 ne
rect 30197 27743 30446 27744
tri 30197 27742 30198 27743 ne
rect 30198 27742 30446 27743
tri 30198 27741 30199 27742 ne
rect 30199 27741 30446 27742
tri 30199 27740 30200 27741 ne
rect 30200 27740 30446 27741
tri 30200 27739 30201 27740 ne
rect 30201 27739 30446 27740
tri 30201 27738 30202 27739 ne
rect 30202 27738 30446 27739
tri 30202 27737 30203 27738 ne
rect 30203 27737 30446 27738
tri 30203 27736 30204 27737 ne
rect 30204 27736 30446 27737
tri 30204 27735 30205 27736 ne
rect 30205 27735 30446 27736
tri 30205 27734 30206 27735 ne
rect 30206 27734 30446 27735
tri 30206 27733 30207 27734 ne
rect 30207 27733 30446 27734
tri 30207 27732 30208 27733 ne
rect 30208 27732 30446 27733
tri 30208 27731 30209 27732 ne
rect 30209 27731 30446 27732
tri 30209 27730 30210 27731 ne
rect 30210 27730 30446 27731
tri 30210 27729 30211 27730 ne
rect 30211 27729 30446 27730
tri 30211 27728 30212 27729 ne
rect 30212 27728 30446 27729
tri 30212 27727 30213 27728 ne
rect 30213 27727 30446 27728
tri 30213 27726 30214 27727 ne
rect 30214 27726 30446 27727
tri 30214 27725 30215 27726 ne
rect 30215 27725 30446 27726
tri 30446 27725 30491 27770 sw
rect 70802 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
tri 30215 27705 30235 27725 ne
rect 30235 27705 30491 27725
tri 30491 27705 30511 27725 sw
tri 30235 27660 30280 27705 ne
rect 30280 27664 30511 27705
rect 30280 27660 30414 27664
tri 30280 27640 30300 27660 ne
rect 30300 27640 30414 27660
tri 30300 27595 30345 27640 ne
rect 30345 27618 30414 27640
rect 30460 27660 30511 27664
tri 30511 27660 30556 27705 sw
rect 70802 27684 71000 27742
rect 30460 27618 30556 27660
rect 30345 27615 30556 27618
tri 30556 27615 30601 27660 sw
rect 70802 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30345 27595 30601 27615
tri 30345 27560 30380 27595 ne
rect 30380 27570 30601 27595
tri 30601 27570 30646 27615 sw
rect 70802 27580 71000 27638
rect 30380 27560 30646 27570
tri 30380 27559 30381 27560 ne
rect 30381 27559 30646 27560
tri 30381 27558 30382 27559 ne
rect 30382 27558 30646 27559
tri 30382 27557 30383 27558 ne
rect 30383 27557 30646 27558
tri 30383 27556 30384 27557 ne
rect 30384 27556 30646 27557
tri 30384 27555 30385 27556 ne
rect 30385 27555 30646 27556
tri 30385 27554 30386 27555 ne
rect 30386 27554 30646 27555
tri 30386 27553 30387 27554 ne
rect 30387 27553 30646 27554
tri 30387 27552 30388 27553 ne
rect 30388 27552 30646 27553
tri 30388 27551 30389 27552 ne
rect 30389 27551 30646 27552
tri 30389 27550 30390 27551 ne
rect 30390 27550 30646 27551
tri 30390 27549 30391 27550 ne
rect 30391 27549 30646 27550
tri 30391 27548 30392 27549 ne
rect 30392 27548 30646 27549
tri 30392 27547 30393 27548 ne
rect 30393 27547 30646 27548
tri 30393 27546 30394 27547 ne
rect 30394 27546 30646 27547
tri 30394 27545 30395 27546 ne
rect 30395 27545 30646 27546
tri 30395 27544 30396 27545 ne
rect 30396 27544 30646 27545
tri 30396 27543 30397 27544 ne
rect 30397 27543 30646 27544
tri 30397 27542 30398 27543 ne
rect 30398 27542 30646 27543
tri 30398 27541 30399 27542 ne
rect 30399 27541 30646 27542
tri 30399 27540 30400 27541 ne
rect 30400 27540 30646 27541
tri 30400 27539 30401 27540 ne
rect 30401 27539 30646 27540
tri 30646 27539 30677 27570 sw
tri 30401 27538 30402 27539 ne
rect 30402 27538 30677 27539
tri 30402 27537 30403 27538 ne
rect 30403 27537 30677 27538
tri 30403 27536 30404 27537 ne
rect 30404 27536 30677 27537
tri 30404 27535 30405 27536 ne
rect 30405 27535 30677 27536
tri 30405 27534 30406 27535 ne
rect 30406 27534 30677 27535
tri 30406 27533 30407 27534 ne
rect 30407 27533 30677 27534
tri 30407 27532 30408 27533 ne
rect 30408 27532 30677 27533
tri 30408 27531 30409 27532 ne
rect 30409 27531 30546 27532
tri 30409 27530 30410 27531 ne
rect 30410 27530 30546 27531
tri 30410 27529 30411 27530 ne
rect 30411 27529 30546 27530
tri 30411 27528 30412 27529 ne
rect 30412 27528 30546 27529
tri 30412 27527 30413 27528 ne
rect 30413 27527 30546 27528
tri 30413 27526 30414 27527 ne
rect 30414 27526 30546 27527
tri 30414 27525 30415 27526 ne
rect 30415 27525 30546 27526
tri 30415 27524 30416 27525 ne
rect 30416 27524 30546 27525
tri 30416 27523 30417 27524 ne
rect 30417 27523 30546 27524
tri 30417 27522 30418 27523 ne
rect 30418 27522 30546 27523
tri 30418 27521 30419 27522 ne
rect 30419 27521 30546 27522
tri 30419 27520 30420 27521 ne
rect 30420 27520 30546 27521
tri 30420 27519 30421 27520 ne
rect 30421 27519 30546 27520
tri 30421 27518 30422 27519 ne
rect 30422 27518 30546 27519
tri 30422 27517 30423 27518 ne
rect 30423 27517 30546 27518
tri 30423 27516 30424 27517 ne
rect 30424 27516 30546 27517
tri 30424 27515 30425 27516 ne
rect 30425 27515 30546 27516
tri 30425 27514 30426 27515 ne
rect 30426 27514 30546 27515
tri 30426 27513 30427 27514 ne
rect 30427 27513 30546 27514
tri 30427 27512 30428 27513 ne
rect 30428 27512 30546 27513
tri 30428 27511 30429 27512 ne
rect 30429 27511 30546 27512
tri 30429 27510 30430 27511 ne
rect 30430 27510 30546 27511
tri 30430 27509 30431 27510 ne
rect 30431 27509 30546 27510
tri 30431 27508 30432 27509 ne
rect 30432 27508 30546 27509
tri 30432 27507 30433 27508 ne
rect 30433 27507 30546 27508
tri 30433 27506 30434 27507 ne
rect 30434 27506 30546 27507
tri 30434 27505 30435 27506 ne
rect 30435 27505 30546 27506
tri 30435 27504 30436 27505 ne
rect 30436 27504 30546 27505
tri 30436 27503 30437 27504 ne
rect 30437 27503 30546 27504
tri 30437 27502 30438 27503 ne
rect 30438 27502 30546 27503
tri 30438 27501 30439 27502 ne
rect 30439 27501 30546 27502
tri 30439 27500 30440 27501 ne
rect 30440 27500 30546 27501
tri 30440 27499 30441 27500 ne
rect 30441 27499 30546 27500
tri 30441 27498 30442 27499 ne
rect 30442 27498 30546 27499
tri 30442 27497 30443 27498 ne
rect 30443 27497 30546 27498
tri 30443 27496 30444 27497 ne
rect 30444 27496 30546 27497
tri 30444 27495 30445 27496 ne
rect 30445 27495 30546 27496
tri 30445 27494 30446 27495 ne
rect 30446 27494 30546 27495
tri 30446 27493 30447 27494 ne
rect 30447 27493 30546 27494
tri 30447 27492 30448 27493 ne
rect 30448 27492 30546 27493
tri 30448 27491 30449 27492 ne
rect 30449 27491 30546 27492
tri 30449 27490 30450 27491 ne
rect 30450 27490 30546 27491
tri 30450 27489 30451 27490 ne
rect 30451 27489 30546 27490
tri 30451 27488 30452 27489 ne
rect 30452 27488 30546 27489
tri 30452 27487 30453 27488 ne
rect 30453 27487 30546 27488
tri 30453 27486 30454 27487 ne
rect 30454 27486 30546 27487
rect 30592 27494 30677 27532
tri 30677 27494 30722 27539 sw
rect 70802 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 30592 27486 30722 27494
tri 30454 27485 30455 27486 ne
rect 30455 27485 30722 27486
tri 30455 27484 30456 27485 ne
rect 30456 27484 30722 27485
tri 30456 27483 30457 27484 ne
rect 30457 27483 30722 27484
tri 30457 27482 30458 27483 ne
rect 30458 27482 30722 27483
tri 30458 27481 30459 27482 ne
rect 30459 27481 30722 27482
tri 30459 27480 30460 27481 ne
rect 30460 27480 30722 27481
tri 30460 27479 30461 27480 ne
rect 30461 27479 30722 27480
tri 30461 27478 30462 27479 ne
rect 30462 27478 30722 27479
tri 30462 27477 30463 27478 ne
rect 30463 27477 30722 27478
tri 30463 27476 30464 27477 ne
rect 30464 27476 30722 27477
tri 30464 27475 30465 27476 ne
rect 30465 27475 30722 27476
tri 30465 27474 30466 27475 ne
rect 30466 27474 30722 27475
tri 30466 27473 30467 27474 ne
rect 30467 27473 30722 27474
tri 30467 27472 30468 27473 ne
rect 30468 27472 30722 27473
tri 30468 27471 30469 27472 ne
rect 30469 27471 30722 27472
tri 30469 27470 30470 27471 ne
rect 30470 27470 30722 27471
tri 30470 27469 30471 27470 ne
rect 30471 27469 30722 27470
tri 30471 27468 30472 27469 ne
rect 30472 27468 30722 27469
tri 30472 27467 30473 27468 ne
rect 30473 27467 30722 27468
tri 30473 27466 30474 27467 ne
rect 30474 27466 30722 27467
tri 30474 27465 30475 27466 ne
rect 30475 27465 30722 27466
tri 30475 27464 30476 27465 ne
rect 30476 27464 30722 27465
tri 30476 27463 30477 27464 ne
rect 30477 27463 30722 27464
tri 30477 27462 30478 27463 ne
rect 30478 27462 30722 27463
tri 30478 27461 30479 27462 ne
rect 30479 27461 30722 27462
tri 30479 27460 30480 27461 ne
rect 30480 27460 30722 27461
tri 30480 27459 30481 27460 ne
rect 30481 27459 30722 27460
tri 30481 27458 30482 27459 ne
rect 30482 27458 30722 27459
tri 30482 27457 30483 27458 ne
rect 30483 27457 30722 27458
tri 30483 27456 30484 27457 ne
rect 30484 27456 30722 27457
tri 30484 27455 30485 27456 ne
rect 30485 27455 30722 27456
tri 30485 27454 30486 27455 ne
rect 30486 27454 30722 27455
tri 30486 27453 30487 27454 ne
rect 30487 27453 30722 27454
tri 30487 27452 30488 27453 ne
rect 30488 27452 30722 27453
tri 30488 27451 30489 27452 ne
rect 30489 27451 30722 27452
tri 30489 27450 30490 27451 ne
rect 30490 27450 30722 27451
tri 30490 27449 30491 27450 ne
rect 30491 27449 30722 27450
tri 30722 27449 30767 27494 sw
rect 70802 27476 71000 27534
tri 30491 27404 30536 27449 ne
rect 30536 27404 30767 27449
tri 30767 27404 30812 27449 sw
rect 70802 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30536 27384 30556 27404 ne
rect 30556 27400 30812 27404
rect 30556 27384 30678 27400
tri 30556 27359 30581 27384 ne
rect 30581 27359 30678 27384
tri 30581 27339 30601 27359 ne
rect 30601 27354 30678 27359
rect 30724 27384 30812 27400
tri 30812 27384 30832 27404 sw
rect 30724 27354 30832 27384
rect 30601 27339 30832 27354
tri 30832 27339 30877 27384 sw
rect 70802 27372 71000 27430
tri 30601 27294 30646 27339 ne
rect 30646 27294 30877 27339
tri 30877 27294 30922 27339 sw
rect 70802 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
tri 30646 27285 30655 27294 ne
rect 30655 27285 30922 27294
tri 30655 27284 30656 27285 ne
rect 30656 27284 30922 27285
tri 30656 27283 30657 27284 ne
rect 30657 27283 30922 27284
tri 30657 27282 30658 27283 ne
rect 30658 27282 30922 27283
tri 30658 27281 30659 27282 ne
rect 30659 27281 30922 27282
tri 30659 27280 30660 27281 ne
rect 30660 27280 30922 27281
tri 30660 27279 30661 27280 ne
rect 30661 27279 30922 27280
tri 30661 27278 30662 27279 ne
rect 30662 27278 30922 27279
tri 30662 27277 30663 27278 ne
rect 30663 27277 30922 27278
tri 30663 27276 30664 27277 ne
rect 30664 27276 30922 27277
tri 30664 27275 30665 27276 ne
rect 30665 27275 30922 27276
tri 30665 27274 30666 27275 ne
rect 30666 27274 30922 27275
tri 30666 27273 30667 27274 ne
rect 30667 27273 30922 27274
tri 30667 27272 30668 27273 ne
rect 30668 27272 30922 27273
tri 30668 27271 30669 27272 ne
rect 30669 27271 30922 27272
tri 30669 27270 30670 27271 ne
rect 30670 27270 30922 27271
tri 30670 27269 30671 27270 ne
rect 30671 27269 30922 27270
tri 30671 27268 30672 27269 ne
rect 30672 27268 30922 27269
tri 30672 27267 30673 27268 ne
rect 30673 27267 30810 27268
tri 30673 27266 30674 27267 ne
rect 30674 27266 30810 27267
tri 30674 27265 30675 27266 ne
rect 30675 27265 30810 27266
tri 30675 27264 30676 27265 ne
rect 30676 27264 30810 27265
tri 30676 27263 30677 27264 ne
rect 30677 27263 30810 27264
tri 30677 27262 30678 27263 ne
rect 30678 27262 30810 27263
tri 30678 27261 30679 27262 ne
rect 30679 27261 30810 27262
tri 30679 27260 30680 27261 ne
rect 30680 27260 30810 27261
tri 30680 27259 30681 27260 ne
rect 30681 27259 30810 27260
tri 30681 27258 30682 27259 ne
rect 30682 27258 30810 27259
tri 30682 27257 30683 27258 ne
rect 30683 27257 30810 27258
tri 30683 27256 30684 27257 ne
rect 30684 27256 30810 27257
tri 30684 27255 30685 27256 ne
rect 30685 27255 30810 27256
tri 30685 27254 30686 27255 ne
rect 30686 27254 30810 27255
tri 30686 27253 30687 27254 ne
rect 30687 27253 30810 27254
tri 30687 27252 30688 27253 ne
rect 30688 27252 30810 27253
tri 30688 27251 30689 27252 ne
rect 30689 27251 30810 27252
tri 30689 27250 30690 27251 ne
rect 30690 27250 30810 27251
tri 30690 27249 30691 27250 ne
rect 30691 27249 30810 27250
tri 30691 27248 30692 27249 ne
rect 30692 27248 30810 27249
tri 30692 27247 30693 27248 ne
rect 30693 27247 30810 27248
tri 30693 27246 30694 27247 ne
rect 30694 27246 30810 27247
tri 30694 27245 30695 27246 ne
rect 30695 27245 30810 27246
tri 30695 27244 30696 27245 ne
rect 30696 27244 30810 27245
tri 30696 27243 30697 27244 ne
rect 30697 27243 30810 27244
tri 30697 27242 30698 27243 ne
rect 30698 27242 30810 27243
tri 30698 27241 30699 27242 ne
rect 30699 27241 30810 27242
tri 30699 27240 30700 27241 ne
rect 30700 27240 30810 27241
tri 30700 27239 30701 27240 ne
rect 30701 27239 30810 27240
tri 30701 27238 30702 27239 ne
rect 30702 27238 30810 27239
tri 30702 27237 30703 27238 ne
rect 30703 27237 30810 27238
tri 30703 27236 30704 27237 ne
rect 30704 27236 30810 27237
tri 30704 27235 30705 27236 ne
rect 30705 27235 30810 27236
tri 30705 27234 30706 27235 ne
rect 30706 27234 30810 27235
tri 30706 27233 30707 27234 ne
rect 30707 27233 30810 27234
tri 30707 27232 30708 27233 ne
rect 30708 27232 30810 27233
tri 30708 27231 30709 27232 ne
rect 30709 27231 30810 27232
tri 30709 27230 30710 27231 ne
rect 30710 27230 30810 27231
tri 30710 27229 30711 27230 ne
rect 30711 27229 30810 27230
tri 30711 27228 30712 27229 ne
rect 30712 27228 30810 27229
tri 30712 27227 30713 27228 ne
rect 30713 27227 30810 27228
tri 30713 27226 30714 27227 ne
rect 30714 27226 30810 27227
tri 30714 27225 30715 27226 ne
rect 30715 27225 30810 27226
tri 30715 27224 30716 27225 ne
rect 30716 27224 30810 27225
tri 30716 27223 30717 27224 ne
rect 30717 27223 30810 27224
tri 30717 27222 30718 27223 ne
rect 30718 27222 30810 27223
rect 30856 27249 30922 27268
tri 30922 27249 30967 27294 sw
rect 70802 27268 71000 27326
rect 30856 27222 30967 27249
tri 30718 27221 30719 27222 ne
rect 30719 27221 30967 27222
tri 30719 27220 30720 27221 ne
rect 30720 27220 30967 27221
tri 30720 27219 30721 27220 ne
rect 30721 27219 30967 27220
tri 30721 27218 30722 27219 ne
rect 30722 27218 30967 27219
tri 30967 27218 30998 27249 sw
rect 70802 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30722 27217 30723 27218 ne
rect 30723 27217 30998 27218
tri 30723 27216 30724 27217 ne
rect 30724 27216 30998 27217
tri 30724 27215 30725 27216 ne
rect 30725 27215 30998 27216
tri 30725 27214 30726 27215 ne
rect 30726 27214 30998 27215
tri 30726 27213 30727 27214 ne
rect 30727 27213 30998 27214
tri 30727 27212 30728 27213 ne
rect 30728 27212 30998 27213
tri 30728 27211 30729 27212 ne
rect 30729 27211 30998 27212
tri 30729 27210 30730 27211 ne
rect 30730 27210 30998 27211
tri 30730 27209 30731 27210 ne
rect 30731 27209 30998 27210
tri 30731 27208 30732 27209 ne
rect 30732 27208 30998 27209
tri 30732 27207 30733 27208 ne
rect 30733 27207 30998 27208
tri 30733 27206 30734 27207 ne
rect 30734 27206 30998 27207
tri 30734 27205 30735 27206 ne
rect 30735 27205 30998 27206
tri 30735 27204 30736 27205 ne
rect 30736 27204 30998 27205
tri 30736 27203 30737 27204 ne
rect 30737 27203 30998 27204
tri 30737 27202 30738 27203 ne
rect 30738 27202 30998 27203
tri 30738 27201 30739 27202 ne
rect 30739 27201 30998 27202
tri 30739 27200 30740 27201 ne
rect 30740 27200 30998 27201
tri 30740 27199 30741 27200 ne
rect 30741 27199 30998 27200
tri 30741 27198 30742 27199 ne
rect 30742 27198 30998 27199
tri 30742 27197 30743 27198 ne
rect 30743 27197 30998 27198
tri 30743 27196 30744 27197 ne
rect 30744 27196 30998 27197
tri 30744 27195 30745 27196 ne
rect 30745 27195 30998 27196
tri 30745 27194 30746 27195 ne
rect 30746 27194 30998 27195
tri 30746 27193 30747 27194 ne
rect 30747 27193 30998 27194
tri 30747 27192 30748 27193 ne
rect 30748 27192 30998 27193
tri 30748 27191 30749 27192 ne
rect 30749 27191 30998 27192
tri 30749 27190 30750 27191 ne
rect 30750 27190 30998 27191
tri 30750 27189 30751 27190 ne
rect 30751 27189 30998 27190
tri 30751 27188 30752 27189 ne
rect 30752 27188 30998 27189
tri 30752 27187 30753 27188 ne
rect 30753 27187 30998 27188
tri 30753 27186 30754 27187 ne
rect 30754 27186 30998 27187
tri 30754 27185 30755 27186 ne
rect 30755 27185 30998 27186
tri 30755 27184 30756 27185 ne
rect 30756 27184 30998 27185
tri 30756 27183 30757 27184 ne
rect 30757 27183 30998 27184
tri 30757 27182 30758 27183 ne
rect 30758 27182 30998 27183
tri 30758 27181 30759 27182 ne
rect 30759 27181 30998 27182
tri 30759 27180 30760 27181 ne
rect 30760 27180 30998 27181
tri 30760 27179 30761 27180 ne
rect 30761 27179 30998 27180
tri 30761 27178 30762 27179 ne
rect 30762 27178 30998 27179
tri 30762 27177 30763 27178 ne
rect 30763 27177 30998 27178
tri 30763 27176 30764 27177 ne
rect 30764 27176 30998 27177
tri 30764 27175 30765 27176 ne
rect 30765 27175 30998 27176
tri 30765 27174 30766 27175 ne
rect 30766 27174 30998 27175
tri 30766 27173 30767 27174 ne
rect 30767 27173 30998 27174
tri 30998 27173 31043 27218 sw
tri 30767 27128 30812 27173 ne
rect 30812 27136 31043 27173
rect 30812 27128 30942 27136
tri 30812 27083 30857 27128 ne
rect 30857 27090 30942 27128
rect 30988 27128 31043 27136
tri 31043 27128 31088 27173 sw
rect 70802 27164 71000 27222
rect 30988 27090 31088 27128
rect 30857 27083 31088 27090
tri 31088 27083 31133 27128 sw
rect 70802 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
tri 30857 27038 30902 27083 ne
rect 30902 27063 31133 27083
tri 31133 27063 31153 27083 sw
rect 30902 27038 31153 27063
tri 30902 27018 30922 27038 ne
rect 30922 27018 31153 27038
tri 31153 27018 31198 27063 sw
rect 70802 27060 71000 27118
tri 30922 27011 30929 27018 ne
rect 30929 27011 31198 27018
tri 30929 27010 30930 27011 ne
rect 30930 27010 31198 27011
tri 30930 27009 30931 27010 ne
rect 30931 27009 31198 27010
tri 30931 27008 30932 27009 ne
rect 30932 27008 31198 27009
tri 30932 27007 30933 27008 ne
rect 30933 27007 31198 27008
tri 30933 27006 30934 27007 ne
rect 30934 27006 31198 27007
tri 30934 27005 30935 27006 ne
rect 30935 27005 31198 27006
tri 30935 27004 30936 27005 ne
rect 30936 27004 31198 27005
tri 30936 27003 30937 27004 ne
rect 30937 27003 31074 27004
tri 30937 27002 30938 27003 ne
rect 30938 27002 31074 27003
tri 30938 27001 30939 27002 ne
rect 30939 27001 31074 27002
tri 30939 27000 30940 27001 ne
rect 30940 27000 31074 27001
tri 30940 26999 30941 27000 ne
rect 30941 26999 31074 27000
tri 30941 26998 30942 26999 ne
rect 30942 26998 31074 26999
tri 30942 26997 30943 26998 ne
rect 30943 26997 31074 26998
tri 30943 26996 30944 26997 ne
rect 30944 26996 31074 26997
tri 30944 26995 30945 26996 ne
rect 30945 26995 31074 26996
tri 30945 26994 30946 26995 ne
rect 30946 26994 31074 26995
tri 30946 26993 30947 26994 ne
rect 30947 26993 31074 26994
tri 30947 26992 30948 26993 ne
rect 30948 26992 31074 26993
tri 30948 26991 30949 26992 ne
rect 30949 26991 31074 26992
tri 30949 26990 30950 26991 ne
rect 30950 26990 31074 26991
tri 30950 26989 30951 26990 ne
rect 30951 26989 31074 26990
tri 30951 26988 30952 26989 ne
rect 30952 26988 31074 26989
tri 30952 26987 30953 26988 ne
rect 30953 26987 31074 26988
tri 30953 26986 30954 26987 ne
rect 30954 26986 31074 26987
tri 30954 26985 30955 26986 ne
rect 30955 26985 31074 26986
tri 30955 26984 30956 26985 ne
rect 30956 26984 31074 26985
tri 30956 26983 30957 26984 ne
rect 30957 26983 31074 26984
tri 30957 26982 30958 26983 ne
rect 30958 26982 31074 26983
tri 30958 26981 30959 26982 ne
rect 30959 26981 31074 26982
tri 30959 26980 30960 26981 ne
rect 30960 26980 31074 26981
tri 30960 26979 30961 26980 ne
rect 30961 26979 31074 26980
tri 30961 26978 30962 26979 ne
rect 30962 26978 31074 26979
tri 30962 26977 30963 26978 ne
rect 30963 26977 31074 26978
tri 30963 26976 30964 26977 ne
rect 30964 26976 31074 26977
tri 30964 26975 30965 26976 ne
rect 30965 26975 31074 26976
tri 30965 26974 30966 26975 ne
rect 30966 26974 31074 26975
tri 30966 26973 30967 26974 ne
rect 30967 26973 31074 26974
tri 30967 26972 30968 26973 ne
rect 30968 26972 31074 26973
tri 30968 26971 30969 26972 ne
rect 30969 26971 31074 26972
tri 30969 26970 30970 26971 ne
rect 30970 26970 31074 26971
tri 30970 26969 30971 26970 ne
rect 30971 26969 31074 26970
tri 30971 26968 30972 26969 ne
rect 30972 26968 31074 26969
tri 30972 26967 30973 26968 ne
rect 30973 26967 31074 26968
tri 30973 26966 30974 26967 ne
rect 30974 26966 31074 26967
tri 30974 26965 30975 26966 ne
rect 30975 26965 31074 26966
tri 30975 26964 30976 26965 ne
rect 30976 26964 31074 26965
tri 30976 26963 30977 26964 ne
rect 30977 26963 31074 26964
tri 30977 26962 30978 26963 ne
rect 30978 26962 31074 26963
tri 30978 26961 30979 26962 ne
rect 30979 26961 31074 26962
tri 30979 26960 30980 26961 ne
rect 30980 26960 31074 26961
tri 30980 26959 30981 26960 ne
rect 30981 26959 31074 26960
tri 30981 26958 30982 26959 ne
rect 30982 26958 31074 26959
rect 31120 26973 31198 27004
tri 31198 26973 31243 27018 sw
rect 70802 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 31120 26958 31243 26973
tri 30982 26957 30983 26958 ne
rect 30983 26957 31243 26958
tri 30983 26956 30984 26957 ne
rect 30984 26956 31243 26957
tri 30984 26955 30985 26956 ne
rect 30985 26955 31243 26956
tri 30985 26954 30986 26955 ne
rect 30986 26954 31243 26955
tri 30986 26953 30987 26954 ne
rect 30987 26953 31243 26954
tri 30987 26952 30988 26953 ne
rect 30988 26952 31243 26953
tri 30988 26951 30989 26952 ne
rect 30989 26951 31243 26952
tri 30989 26950 30990 26951 ne
rect 30990 26950 31243 26951
tri 30990 26949 30991 26950 ne
rect 30991 26949 31243 26950
tri 30991 26948 30992 26949 ne
rect 30992 26948 31243 26949
tri 30992 26947 30993 26948 ne
rect 30993 26947 31243 26948
tri 30993 26946 30994 26947 ne
rect 30994 26946 31243 26947
tri 30994 26945 30995 26946 ne
rect 30995 26945 31243 26946
tri 30995 26944 30996 26945 ne
rect 30996 26944 31243 26945
tri 30996 26943 30997 26944 ne
rect 30997 26943 31243 26944
tri 30997 26942 30998 26943 ne
rect 30998 26942 31243 26943
tri 30998 26941 30999 26942 ne
rect 30999 26941 31243 26942
tri 30999 26940 31000 26941 ne
rect 31000 26940 31243 26941
tri 31000 26939 31001 26940 ne
rect 31001 26939 31243 26940
tri 31001 26938 31002 26939 ne
rect 31002 26938 31243 26939
tri 31002 26937 31003 26938 ne
rect 31003 26937 31243 26938
tri 31003 26936 31004 26937 ne
rect 31004 26936 31243 26937
tri 31004 26935 31005 26936 ne
rect 31005 26935 31243 26936
tri 31005 26934 31006 26935 ne
rect 31006 26934 31243 26935
tri 31006 26933 31007 26934 ne
rect 31007 26933 31243 26934
tri 31007 26932 31008 26933 ne
rect 31008 26932 31243 26933
tri 31008 26931 31009 26932 ne
rect 31009 26931 31243 26932
tri 31009 26930 31010 26931 ne
rect 31010 26930 31243 26931
tri 31010 26929 31011 26930 ne
rect 31011 26929 31243 26930
tri 31011 26928 31012 26929 ne
rect 31012 26928 31243 26929
tri 31243 26928 31288 26973 sw
rect 70802 26956 71000 27014
tri 31012 26927 31013 26928 ne
rect 31013 26927 31288 26928
tri 31013 26926 31014 26927 ne
rect 31014 26926 31288 26927
tri 31014 26925 31015 26926 ne
rect 31015 26925 31288 26926
tri 31015 26924 31016 26925 ne
rect 31016 26924 31288 26925
tri 31016 26923 31017 26924 ne
rect 31017 26923 31288 26924
tri 31017 26922 31018 26923 ne
rect 31018 26922 31288 26923
tri 31018 26921 31019 26922 ne
rect 31019 26921 31288 26922
tri 31019 26920 31020 26921 ne
rect 31020 26920 31288 26921
tri 31020 26919 31021 26920 ne
rect 31021 26919 31288 26920
tri 31021 26918 31022 26919 ne
rect 31022 26918 31288 26919
tri 31022 26917 31023 26918 ne
rect 31023 26917 31288 26918
tri 31023 26916 31024 26917 ne
rect 31024 26916 31288 26917
tri 31024 26915 31025 26916 ne
rect 31025 26915 31288 26916
tri 31025 26914 31026 26915 ne
rect 31026 26914 31288 26915
tri 31026 26913 31027 26914 ne
rect 31027 26913 31288 26914
tri 31027 26912 31028 26913 ne
rect 31028 26912 31288 26913
tri 31028 26911 31029 26912 ne
rect 31029 26911 31288 26912
tri 31029 26910 31030 26911 ne
rect 31030 26910 31288 26911
tri 31030 26909 31031 26910 ne
rect 31031 26909 31288 26910
tri 31031 26908 31032 26909 ne
rect 31032 26908 31288 26909
tri 31032 26907 31033 26908 ne
rect 31033 26907 31288 26908
tri 31033 26906 31034 26907 ne
rect 31034 26906 31288 26907
tri 31034 26905 31035 26906 ne
rect 31035 26905 31288 26906
tri 31035 26904 31036 26905 ne
rect 31036 26904 31288 26905
tri 31036 26903 31037 26904 ne
rect 31037 26903 31288 26904
tri 31037 26902 31038 26903 ne
rect 31038 26902 31288 26903
tri 31038 26901 31039 26902 ne
rect 31039 26901 31288 26902
tri 31039 26900 31040 26901 ne
rect 31040 26900 31288 26901
tri 31040 26899 31041 26900 ne
rect 31041 26899 31288 26900
tri 31041 26898 31042 26899 ne
rect 31042 26898 31288 26899
tri 31042 26897 31043 26898 ne
rect 31043 26897 31288 26898
tri 31288 26897 31319 26928 sw
rect 70802 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31043 26866 31074 26897 ne
rect 31074 26872 31319 26897
rect 31074 26866 31206 26872
tri 31074 26821 31119 26866 ne
rect 31119 26826 31206 26866
rect 31252 26852 31319 26872
tri 31319 26852 31364 26897 sw
rect 70802 26852 71000 26910
rect 31252 26826 31364 26852
rect 31119 26821 31364 26826
tri 31119 26776 31164 26821 ne
rect 31164 26807 31364 26821
tri 31364 26807 31409 26852 sw
rect 31164 26776 31409 26807
tri 31164 26737 31203 26776 ne
rect 31203 26762 31409 26776
tri 31409 26762 31454 26807 sw
rect 70802 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 31203 26756 31454 26762
tri 31454 26756 31460 26762 sw
rect 31203 26740 31460 26756
rect 31203 26737 31338 26740
tri 31203 26736 31204 26737 ne
rect 31204 26736 31338 26737
tri 31204 26735 31205 26736 ne
rect 31205 26735 31338 26736
tri 31205 26734 31206 26735 ne
rect 31206 26734 31338 26735
tri 31206 26733 31207 26734 ne
rect 31207 26733 31338 26734
tri 31207 26732 31208 26733 ne
rect 31208 26732 31338 26733
tri 31208 26731 31209 26732 ne
rect 31209 26731 31338 26732
tri 31209 26730 31210 26731 ne
rect 31210 26730 31338 26731
tri 31210 26729 31211 26730 ne
rect 31211 26729 31338 26730
tri 31211 26728 31212 26729 ne
rect 31212 26728 31338 26729
tri 31212 26727 31213 26728 ne
rect 31213 26727 31338 26728
tri 31213 26726 31214 26727 ne
rect 31214 26726 31338 26727
tri 31214 26725 31215 26726 ne
rect 31215 26725 31338 26726
tri 31215 26724 31216 26725 ne
rect 31216 26724 31338 26725
tri 31216 26723 31217 26724 ne
rect 31217 26723 31338 26724
tri 31217 26722 31218 26723 ne
rect 31218 26722 31338 26723
tri 31218 26721 31219 26722 ne
rect 31219 26721 31338 26722
tri 31219 26720 31220 26721 ne
rect 31220 26720 31338 26721
tri 31220 26719 31221 26720 ne
rect 31221 26719 31338 26720
tri 31221 26718 31222 26719 ne
rect 31222 26718 31338 26719
tri 31222 26717 31223 26718 ne
rect 31223 26717 31338 26718
tri 31223 26716 31224 26717 ne
rect 31224 26716 31338 26717
tri 31224 26715 31225 26716 ne
rect 31225 26715 31338 26716
tri 31225 26714 31226 26715 ne
rect 31226 26714 31338 26715
tri 31226 26713 31227 26714 ne
rect 31227 26713 31338 26714
tri 31227 26712 31228 26713 ne
rect 31228 26712 31338 26713
tri 31228 26711 31229 26712 ne
rect 31229 26711 31338 26712
tri 31229 26710 31230 26711 ne
rect 31230 26710 31338 26711
tri 31230 26709 31231 26710 ne
rect 31231 26709 31338 26710
tri 31231 26708 31232 26709 ne
rect 31232 26708 31338 26709
tri 31232 26707 31233 26708 ne
rect 31233 26707 31338 26708
tri 31233 26706 31234 26707 ne
rect 31234 26706 31338 26707
tri 31234 26705 31235 26706 ne
rect 31235 26705 31338 26706
tri 31235 26704 31236 26705 ne
rect 31236 26704 31338 26705
tri 31236 26703 31237 26704 ne
rect 31237 26703 31338 26704
tri 31237 26702 31238 26703 ne
rect 31238 26702 31338 26703
tri 31238 26701 31239 26702 ne
rect 31239 26701 31338 26702
tri 31239 26700 31240 26701 ne
rect 31240 26700 31338 26701
tri 31240 26699 31241 26700 ne
rect 31241 26699 31338 26700
tri 31241 26698 31242 26699 ne
rect 31242 26698 31338 26699
tri 31242 26697 31243 26698 ne
rect 31243 26697 31338 26698
tri 31243 26696 31244 26697 ne
rect 31244 26696 31338 26697
tri 31244 26695 31245 26696 ne
rect 31245 26695 31338 26696
tri 31245 26694 31246 26695 ne
rect 31246 26694 31338 26695
rect 31384 26711 31460 26740
tri 31460 26711 31505 26756 sw
rect 70802 26748 71000 26806
rect 31384 26694 31505 26711
tri 31246 26693 31247 26694 ne
rect 31247 26693 31505 26694
tri 31247 26692 31248 26693 ne
rect 31248 26692 31505 26693
tri 31248 26691 31249 26692 ne
rect 31249 26691 31505 26692
tri 31249 26690 31250 26691 ne
rect 31250 26690 31505 26691
tri 31250 26689 31251 26690 ne
rect 31251 26689 31505 26690
tri 31251 26688 31252 26689 ne
rect 31252 26688 31505 26689
tri 31252 26687 31253 26688 ne
rect 31253 26687 31505 26688
tri 31253 26686 31254 26687 ne
rect 31254 26686 31505 26687
tri 31254 26685 31255 26686 ne
rect 31255 26685 31505 26686
tri 31255 26684 31256 26685 ne
rect 31256 26684 31505 26685
tri 31256 26683 31257 26684 ne
rect 31257 26683 31505 26684
tri 31257 26682 31258 26683 ne
rect 31258 26682 31505 26683
tri 31258 26681 31259 26682 ne
rect 31259 26681 31505 26682
tri 31259 26680 31260 26681 ne
rect 31260 26680 31505 26681
tri 31260 26679 31261 26680 ne
rect 31261 26679 31505 26680
tri 31261 26678 31262 26679 ne
rect 31262 26678 31505 26679
tri 31262 26677 31263 26678 ne
rect 31263 26677 31505 26678
tri 31263 26676 31264 26677 ne
rect 31264 26676 31505 26677
tri 31264 26675 31265 26676 ne
rect 31265 26675 31505 26676
tri 31265 26674 31266 26675 ne
rect 31266 26674 31505 26675
tri 31266 26673 31267 26674 ne
rect 31267 26673 31505 26674
tri 31267 26672 31268 26673 ne
rect 31268 26672 31505 26673
tri 31268 26671 31269 26672 ne
rect 31269 26671 31505 26672
tri 31269 26670 31270 26671 ne
rect 31270 26670 31505 26671
tri 31270 26669 31271 26670 ne
rect 31271 26669 31505 26670
tri 31271 26668 31272 26669 ne
rect 31272 26668 31505 26669
tri 31272 26667 31273 26668 ne
rect 31273 26667 31505 26668
tri 31273 26666 31274 26667 ne
rect 31274 26666 31505 26667
tri 31505 26666 31550 26711 sw
rect 70802 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
tri 31274 26665 31275 26666 ne
rect 31275 26665 31550 26666
tri 31275 26664 31276 26665 ne
rect 31276 26664 31550 26665
tri 31276 26663 31277 26664 ne
rect 31277 26663 31550 26664
tri 31277 26662 31278 26663 ne
rect 31278 26662 31550 26663
tri 31278 26661 31279 26662 ne
rect 31279 26661 31550 26662
tri 31279 26660 31280 26661 ne
rect 31280 26660 31550 26661
tri 31280 26659 31281 26660 ne
rect 31281 26659 31550 26660
tri 31281 26658 31282 26659 ne
rect 31282 26658 31550 26659
tri 31282 26657 31283 26658 ne
rect 31283 26657 31550 26658
tri 31283 26656 31284 26657 ne
rect 31284 26656 31550 26657
tri 31284 26655 31285 26656 ne
rect 31285 26655 31550 26656
tri 31285 26654 31286 26655 ne
rect 31286 26654 31550 26655
tri 31286 26653 31287 26654 ne
rect 31287 26653 31550 26654
tri 31287 26652 31288 26653 ne
rect 31288 26652 31550 26653
tri 31288 26651 31289 26652 ne
rect 31289 26651 31550 26652
tri 31289 26650 31290 26651 ne
rect 31290 26650 31550 26651
tri 31290 26649 31291 26650 ne
rect 31291 26649 31550 26650
tri 31291 26648 31292 26649 ne
rect 31292 26648 31550 26649
tri 31292 26647 31293 26648 ne
rect 31293 26647 31550 26648
tri 31293 26646 31294 26647 ne
rect 31294 26646 31550 26647
tri 31294 26645 31295 26646 ne
rect 31295 26645 31550 26646
tri 31295 26644 31296 26645 ne
rect 31296 26644 31550 26645
tri 31296 26643 31297 26644 ne
rect 31297 26643 31550 26644
tri 31297 26642 31298 26643 ne
rect 31298 26642 31550 26643
tri 31298 26641 31299 26642 ne
rect 31299 26641 31550 26642
tri 31299 26640 31300 26641 ne
rect 31300 26640 31550 26641
tri 31300 26639 31301 26640 ne
rect 31301 26639 31550 26640
tri 31301 26638 31302 26639 ne
rect 31302 26638 31550 26639
tri 31302 26637 31303 26638 ne
rect 31303 26637 31550 26638
tri 31303 26636 31304 26637 ne
rect 31304 26636 31550 26637
tri 31304 26635 31305 26636 ne
rect 31305 26635 31550 26636
tri 31305 26634 31306 26635 ne
rect 31306 26634 31550 26635
tri 31306 26633 31307 26634 ne
rect 31307 26633 31550 26634
tri 31307 26632 31308 26633 ne
rect 31308 26632 31550 26633
tri 31308 26631 31309 26632 ne
rect 31309 26631 31550 26632
tri 31309 26630 31310 26631 ne
rect 31310 26630 31550 26631
tri 31310 26629 31311 26630 ne
rect 31311 26629 31550 26630
tri 31311 26628 31312 26629 ne
rect 31312 26628 31550 26629
tri 31312 26627 31313 26628 ne
rect 31313 26627 31550 26628
tri 31313 26626 31314 26627 ne
rect 31314 26626 31550 26627
tri 31314 26625 31315 26626 ne
rect 31315 26625 31550 26626
tri 31315 26624 31316 26625 ne
rect 31316 26624 31550 26625
tri 31316 26623 31317 26624 ne
rect 31317 26623 31550 26624
tri 31317 26622 31318 26623 ne
rect 31318 26622 31550 26623
tri 31318 26621 31319 26622 ne
rect 31319 26621 31550 26622
tri 31550 26621 31595 26666 sw
rect 70802 26644 71000 26702
tri 31319 26607 31333 26621 ne
rect 31333 26608 31595 26621
rect 31333 26607 31470 26608
tri 31333 26562 31378 26607 ne
rect 31378 26562 31470 26607
rect 31516 26607 31595 26608
tri 31595 26607 31609 26621 sw
rect 31516 26562 31609 26607
tri 31609 26562 31654 26607 sw
rect 70802 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
tri 31378 26546 31394 26562 ne
rect 31394 26546 31654 26562
tri 31394 26501 31439 26546 ne
rect 31439 26517 31654 26546
tri 31654 26517 31699 26562 sw
rect 70802 26540 71000 26598
rect 31439 26501 31699 26517
tri 31439 26462 31478 26501 ne
rect 31478 26476 31699 26501
rect 31478 26462 31602 26476
tri 31478 26461 31479 26462 ne
rect 31479 26461 31602 26462
tri 31479 26460 31480 26461 ne
rect 31480 26460 31602 26461
tri 31480 26459 31481 26460 ne
rect 31481 26459 31602 26460
tri 31481 26458 31482 26459 ne
rect 31482 26458 31602 26459
tri 31482 26457 31483 26458 ne
rect 31483 26457 31602 26458
tri 31483 26456 31484 26457 ne
rect 31484 26456 31602 26457
tri 31484 26455 31485 26456 ne
rect 31485 26455 31602 26456
tri 31485 26454 31486 26455 ne
rect 31486 26454 31602 26455
tri 31486 26453 31487 26454 ne
rect 31487 26453 31602 26454
tri 31487 26452 31488 26453 ne
rect 31488 26452 31602 26453
tri 31488 26451 31489 26452 ne
rect 31489 26451 31602 26452
tri 31489 26450 31490 26451 ne
rect 31490 26450 31602 26451
tri 31490 26449 31491 26450 ne
rect 31491 26449 31602 26450
tri 31491 26448 31492 26449 ne
rect 31492 26448 31602 26449
tri 31492 26447 31493 26448 ne
rect 31493 26447 31602 26448
tri 31493 26446 31494 26447 ne
rect 31494 26446 31602 26447
tri 31494 26445 31495 26446 ne
rect 31495 26445 31602 26446
tri 31495 26444 31496 26445 ne
rect 31496 26444 31602 26445
tri 31496 26443 31497 26444 ne
rect 31497 26443 31602 26444
tri 31497 26442 31498 26443 ne
rect 31498 26442 31602 26443
tri 31498 26441 31499 26442 ne
rect 31499 26441 31602 26442
tri 31499 26440 31500 26441 ne
rect 31500 26440 31602 26441
tri 31500 26439 31501 26440 ne
rect 31501 26439 31602 26440
tri 31501 26438 31502 26439 ne
rect 31502 26438 31602 26439
tri 31502 26437 31503 26438 ne
rect 31503 26437 31602 26438
tri 31503 26436 31504 26437 ne
rect 31504 26436 31602 26437
tri 31504 26435 31505 26436 ne
rect 31505 26435 31602 26436
tri 31505 26434 31506 26435 ne
rect 31506 26434 31602 26435
tri 31506 26433 31507 26434 ne
rect 31507 26433 31602 26434
tri 31507 26432 31508 26433 ne
rect 31508 26432 31602 26433
tri 31508 26431 31509 26432 ne
rect 31509 26431 31602 26432
tri 31509 26430 31510 26431 ne
rect 31510 26430 31602 26431
rect 31648 26472 31699 26476
tri 31699 26472 31744 26517 sw
rect 70802 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 31648 26435 31744 26472
tri 31744 26435 31781 26472 sw
rect 70802 26436 71000 26494
rect 31648 26430 31781 26435
tri 31510 26429 31511 26430 ne
rect 31511 26429 31781 26430
tri 31511 26428 31512 26429 ne
rect 31512 26428 31781 26429
tri 31512 26427 31513 26428 ne
rect 31513 26427 31781 26428
tri 31513 26426 31514 26427 ne
rect 31514 26426 31781 26427
tri 31514 26425 31515 26426 ne
rect 31515 26425 31781 26426
tri 31515 26424 31516 26425 ne
rect 31516 26424 31781 26425
tri 31516 26423 31517 26424 ne
rect 31517 26423 31781 26424
tri 31517 26422 31518 26423 ne
rect 31518 26422 31781 26423
tri 31518 26421 31519 26422 ne
rect 31519 26421 31781 26422
tri 31519 26420 31520 26421 ne
rect 31520 26420 31781 26421
tri 31520 26419 31521 26420 ne
rect 31521 26419 31781 26420
tri 31521 26418 31522 26419 ne
rect 31522 26418 31781 26419
tri 31522 26417 31523 26418 ne
rect 31523 26417 31781 26418
tri 31523 26416 31524 26417 ne
rect 31524 26416 31781 26417
tri 31524 26415 31525 26416 ne
rect 31525 26415 31781 26416
tri 31525 26414 31526 26415 ne
rect 31526 26414 31781 26415
tri 31526 26413 31527 26414 ne
rect 31527 26413 31781 26414
tri 31527 26412 31528 26413 ne
rect 31528 26412 31781 26413
tri 31528 26411 31529 26412 ne
rect 31529 26411 31781 26412
tri 31529 26410 31530 26411 ne
rect 31530 26410 31781 26411
tri 31530 26409 31531 26410 ne
rect 31531 26409 31781 26410
tri 31531 26408 31532 26409 ne
rect 31532 26408 31781 26409
tri 31532 26407 31533 26408 ne
rect 31533 26407 31781 26408
tri 31533 26406 31534 26407 ne
rect 31534 26406 31781 26407
tri 31534 26405 31535 26406 ne
rect 31535 26405 31781 26406
tri 31535 26404 31536 26405 ne
rect 31536 26404 31781 26405
tri 31536 26403 31537 26404 ne
rect 31537 26403 31781 26404
tri 31537 26402 31538 26403 ne
rect 31538 26402 31781 26403
tri 31538 26401 31539 26402 ne
rect 31539 26401 31781 26402
tri 31539 26400 31540 26401 ne
rect 31540 26400 31781 26401
tri 31540 26399 31541 26400 ne
rect 31541 26399 31781 26400
tri 31541 26398 31542 26399 ne
rect 31542 26398 31781 26399
tri 31542 26397 31543 26398 ne
rect 31543 26397 31781 26398
tri 31543 26396 31544 26397 ne
rect 31544 26396 31781 26397
tri 31544 26395 31545 26396 ne
rect 31545 26395 31781 26396
tri 31545 26394 31546 26395 ne
rect 31546 26394 31781 26395
tri 31546 26393 31547 26394 ne
rect 31547 26393 31781 26394
tri 31547 26392 31548 26393 ne
rect 31548 26392 31781 26393
tri 31548 26391 31549 26392 ne
rect 31549 26391 31781 26392
tri 31549 26390 31550 26391 ne
rect 31550 26390 31781 26391
tri 31781 26390 31826 26435 sw
rect 70802 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31550 26389 31551 26390 ne
rect 31551 26389 31826 26390
tri 31551 26388 31552 26389 ne
rect 31552 26388 31826 26389
tri 31552 26387 31553 26388 ne
rect 31553 26387 31826 26388
tri 31553 26386 31554 26387 ne
rect 31554 26386 31826 26387
tri 31554 26385 31555 26386 ne
rect 31555 26385 31826 26386
tri 31555 26384 31556 26385 ne
rect 31556 26384 31826 26385
tri 31556 26383 31557 26384 ne
rect 31557 26383 31826 26384
tri 31557 26382 31558 26383 ne
rect 31558 26382 31826 26383
tri 31558 26381 31559 26382 ne
rect 31559 26381 31826 26382
tri 31559 26380 31560 26381 ne
rect 31560 26380 31826 26381
tri 31560 26379 31561 26380 ne
rect 31561 26379 31826 26380
tri 31561 26378 31562 26379 ne
rect 31562 26378 31826 26379
tri 31562 26377 31563 26378 ne
rect 31563 26377 31826 26378
tri 31563 26376 31564 26377 ne
rect 31564 26376 31826 26377
tri 31564 26375 31565 26376 ne
rect 31565 26375 31826 26376
tri 31565 26374 31566 26375 ne
rect 31566 26374 31826 26375
tri 31566 26373 31567 26374 ne
rect 31567 26373 31826 26374
tri 31567 26372 31568 26373 ne
rect 31568 26372 31826 26373
tri 31568 26371 31569 26372 ne
rect 31569 26371 31826 26372
tri 31569 26370 31570 26371 ne
rect 31570 26370 31826 26371
tri 31570 26369 31571 26370 ne
rect 31571 26369 31826 26370
tri 31571 26368 31572 26369 ne
rect 31572 26368 31826 26369
tri 31572 26367 31573 26368 ne
rect 31573 26367 31826 26368
tri 31573 26366 31574 26367 ne
rect 31574 26366 31826 26367
tri 31574 26365 31575 26366 ne
rect 31575 26365 31826 26366
tri 31575 26364 31576 26365 ne
rect 31576 26364 31826 26365
tri 31576 26363 31577 26364 ne
rect 31577 26363 31826 26364
tri 31577 26362 31578 26363 ne
rect 31578 26362 31826 26363
tri 31578 26361 31579 26362 ne
rect 31579 26361 31826 26362
tri 31579 26360 31580 26361 ne
rect 31580 26360 31826 26361
tri 31580 26359 31581 26360 ne
rect 31581 26359 31826 26360
tri 31581 26358 31582 26359 ne
rect 31582 26358 31826 26359
tri 31582 26357 31583 26358 ne
rect 31583 26357 31826 26358
tri 31583 26356 31584 26357 ne
rect 31584 26356 31826 26357
tri 31584 26355 31585 26356 ne
rect 31585 26355 31826 26356
tri 31585 26354 31586 26355 ne
rect 31586 26354 31826 26355
tri 31586 26353 31587 26354 ne
rect 31587 26353 31826 26354
tri 31587 26352 31588 26353 ne
rect 31588 26352 31826 26353
tri 31588 26351 31589 26352 ne
rect 31589 26351 31826 26352
tri 31589 26350 31590 26351 ne
rect 31590 26350 31826 26351
tri 31590 26349 31591 26350 ne
rect 31591 26349 31826 26350
tri 31591 26348 31592 26349 ne
rect 31592 26348 31826 26349
tri 31592 26347 31593 26348 ne
rect 31593 26347 31826 26348
tri 31593 26346 31594 26347 ne
rect 31594 26346 31826 26347
tri 31594 26345 31595 26346 ne
rect 31595 26345 31826 26346
tri 31826 26345 31871 26390 sw
tri 31595 26300 31640 26345 ne
rect 31640 26344 31871 26345
rect 31640 26300 31734 26344
tri 31640 26286 31654 26300 ne
rect 31654 26298 31734 26300
rect 31780 26300 31871 26344
tri 31871 26300 31916 26345 sw
rect 70802 26332 71000 26390
rect 31780 26298 31916 26300
rect 31654 26286 31916 26298
tri 31916 26286 31930 26300 sw
rect 70802 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31654 26255 31685 26286 ne
rect 31685 26255 31930 26286
tri 31685 26241 31699 26255 ne
rect 31699 26241 31930 26255
tri 31930 26241 31975 26286 sw
tri 31699 26196 31744 26241 ne
rect 31744 26212 31975 26241
rect 31744 26196 31866 26212
tri 31744 26188 31752 26196 ne
rect 31752 26188 31866 26196
tri 31752 26187 31753 26188 ne
rect 31753 26187 31866 26188
tri 31753 26186 31754 26187 ne
rect 31754 26186 31866 26187
tri 31754 26185 31755 26186 ne
rect 31755 26185 31866 26186
tri 31755 26184 31756 26185 ne
rect 31756 26184 31866 26185
tri 31756 26183 31757 26184 ne
rect 31757 26183 31866 26184
tri 31757 26182 31758 26183 ne
rect 31758 26182 31866 26183
tri 31758 26181 31759 26182 ne
rect 31759 26181 31866 26182
tri 31759 26180 31760 26181 ne
rect 31760 26180 31866 26181
tri 31760 26179 31761 26180 ne
rect 31761 26179 31866 26180
tri 31761 26178 31762 26179 ne
rect 31762 26178 31866 26179
tri 31762 26177 31763 26178 ne
rect 31763 26177 31866 26178
tri 31763 26176 31764 26177 ne
rect 31764 26176 31866 26177
tri 31764 26175 31765 26176 ne
rect 31765 26175 31866 26176
tri 31765 26174 31766 26175 ne
rect 31766 26174 31866 26175
tri 31766 26173 31767 26174 ne
rect 31767 26173 31866 26174
tri 31767 26172 31768 26173 ne
rect 31768 26172 31866 26173
tri 31768 26171 31769 26172 ne
rect 31769 26171 31866 26172
tri 31769 26170 31770 26171 ne
rect 31770 26170 31866 26171
tri 31770 26169 31771 26170 ne
rect 31771 26169 31866 26170
tri 31771 26168 31772 26169 ne
rect 31772 26168 31866 26169
tri 31772 26167 31773 26168 ne
rect 31773 26167 31866 26168
tri 31773 26166 31774 26167 ne
rect 31774 26166 31866 26167
rect 31912 26196 31975 26212
tri 31975 26196 32020 26241 sw
rect 70802 26228 71000 26286
rect 31912 26166 32020 26196
tri 31774 26165 31775 26166 ne
rect 31775 26165 32020 26166
tri 31775 26164 31776 26165 ne
rect 31776 26164 32020 26165
tri 31776 26163 31777 26164 ne
rect 31777 26163 32020 26164
tri 31777 26162 31778 26163 ne
rect 31778 26162 32020 26163
tri 31778 26161 31779 26162 ne
rect 31779 26161 32020 26162
tri 31779 26160 31780 26161 ne
rect 31780 26160 32020 26161
tri 31780 26159 31781 26160 ne
rect 31781 26159 32020 26160
tri 31781 26158 31782 26159 ne
rect 31782 26158 32020 26159
tri 31782 26157 31783 26158 ne
rect 31783 26157 32020 26158
tri 31783 26156 31784 26157 ne
rect 31784 26156 32020 26157
tri 31784 26155 31785 26156 ne
rect 31785 26155 32020 26156
tri 31785 26154 31786 26155 ne
rect 31786 26154 32020 26155
tri 31786 26153 31787 26154 ne
rect 31787 26153 32020 26154
tri 31787 26152 31788 26153 ne
rect 31788 26152 32020 26153
tri 31788 26151 31789 26152 ne
rect 31789 26151 32020 26152
tri 32020 26151 32065 26196 sw
rect 70802 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
tri 31789 26150 31790 26151 ne
rect 31790 26150 32065 26151
tri 31790 26149 31791 26150 ne
rect 31791 26149 32065 26150
tri 31791 26148 31792 26149 ne
rect 31792 26148 32065 26149
tri 31792 26147 31793 26148 ne
rect 31793 26147 32065 26148
tri 31793 26146 31794 26147 ne
rect 31794 26146 32065 26147
tri 31794 26145 31795 26146 ne
rect 31795 26145 32065 26146
tri 31795 26144 31796 26145 ne
rect 31796 26144 32065 26145
tri 31796 26143 31797 26144 ne
rect 31797 26143 32065 26144
tri 31797 26142 31798 26143 ne
rect 31798 26142 32065 26143
tri 31798 26141 31799 26142 ne
rect 31799 26141 32065 26142
tri 31799 26140 31800 26141 ne
rect 31800 26140 32065 26141
tri 31800 26139 31801 26140 ne
rect 31801 26139 32065 26140
tri 31801 26138 31802 26139 ne
rect 31802 26138 32065 26139
tri 31802 26137 31803 26138 ne
rect 31803 26137 32065 26138
tri 31803 26136 31804 26137 ne
rect 31804 26136 32065 26137
tri 31804 26135 31805 26136 ne
rect 31805 26135 32065 26136
tri 31805 26134 31806 26135 ne
rect 31806 26134 32065 26135
tri 31806 26133 31807 26134 ne
rect 31807 26133 32065 26134
tri 31807 26132 31808 26133 ne
rect 31808 26132 32065 26133
tri 31808 26131 31809 26132 ne
rect 31809 26131 32065 26132
tri 31809 26130 31810 26131 ne
rect 31810 26130 32065 26131
tri 31810 26129 31811 26130 ne
rect 31811 26129 32065 26130
tri 31811 26128 31812 26129 ne
rect 31812 26128 32065 26129
tri 31812 26127 31813 26128 ne
rect 31813 26127 32065 26128
tri 31813 26126 31814 26127 ne
rect 31814 26126 32065 26127
tri 31814 26125 31815 26126 ne
rect 31815 26125 32065 26126
tri 31815 26124 31816 26125 ne
rect 31816 26124 32065 26125
tri 31816 26123 31817 26124 ne
rect 31817 26123 32065 26124
tri 31817 26122 31818 26123 ne
rect 31818 26122 32065 26123
tri 31818 26121 31819 26122 ne
rect 31819 26121 32065 26122
tri 31819 26120 31820 26121 ne
rect 31820 26120 32065 26121
tri 31820 26119 31821 26120 ne
rect 31821 26119 32065 26120
tri 31821 26118 31822 26119 ne
rect 31822 26118 32065 26119
tri 31822 26117 31823 26118 ne
rect 31823 26117 32065 26118
tri 31823 26116 31824 26117 ne
rect 31824 26116 32065 26117
tri 31824 26115 31825 26116 ne
rect 31825 26115 32065 26116
tri 31825 26114 31826 26115 ne
rect 31826 26114 32065 26115
tri 32065 26114 32102 26151 sw
rect 70802 26124 71000 26182
tri 31826 26113 31827 26114 ne
rect 31827 26113 32102 26114
tri 31827 26112 31828 26113 ne
rect 31828 26112 32102 26113
tri 31828 26111 31829 26112 ne
rect 31829 26111 32102 26112
tri 31829 26110 31830 26111 ne
rect 31830 26110 32102 26111
tri 31830 26109 31831 26110 ne
rect 31831 26109 32102 26110
tri 31831 26108 31832 26109 ne
rect 31832 26108 32102 26109
tri 31832 26107 31833 26108 ne
rect 31833 26107 32102 26108
tri 31833 26106 31834 26107 ne
rect 31834 26106 32102 26107
tri 31834 26105 31835 26106 ne
rect 31835 26105 32102 26106
tri 31835 26104 31836 26105 ne
rect 31836 26104 32102 26105
tri 31836 26103 31837 26104 ne
rect 31837 26103 32102 26104
tri 31837 26102 31838 26103 ne
rect 31838 26102 32102 26103
tri 31838 26101 31839 26102 ne
rect 31839 26101 32102 26102
tri 31839 26100 31840 26101 ne
rect 31840 26100 32102 26101
tri 31840 26099 31841 26100 ne
rect 31841 26099 32102 26100
tri 31841 26098 31842 26099 ne
rect 31842 26098 32102 26099
tri 31842 26097 31843 26098 ne
rect 31843 26097 32102 26098
tri 31843 26096 31844 26097 ne
rect 31844 26096 32102 26097
tri 31844 26095 31845 26096 ne
rect 31845 26095 32102 26096
tri 31845 26094 31846 26095 ne
rect 31846 26094 32102 26095
tri 31846 26093 31847 26094 ne
rect 31847 26093 32102 26094
tri 31847 26092 31848 26093 ne
rect 31848 26092 32102 26093
tri 31848 26091 31849 26092 ne
rect 31849 26091 32102 26092
tri 31849 26090 31850 26091 ne
rect 31850 26090 32102 26091
tri 31850 26089 31851 26090 ne
rect 31851 26089 32102 26090
tri 31851 26088 31852 26089 ne
rect 31852 26088 32102 26089
tri 31852 26087 31853 26088 ne
rect 31853 26087 32102 26088
tri 31853 26086 31854 26087 ne
rect 31854 26086 32102 26087
tri 31854 26085 31855 26086 ne
rect 31855 26085 32102 26086
tri 31855 26084 31856 26085 ne
rect 31856 26084 32102 26085
tri 31856 26083 31857 26084 ne
rect 31857 26083 32102 26084
tri 31857 26082 31858 26083 ne
rect 31858 26082 32102 26083
tri 31858 26081 31859 26082 ne
rect 31859 26081 32102 26082
tri 31859 26080 31860 26081 ne
rect 31860 26080 32102 26081
tri 31860 26079 31861 26080 ne
rect 31861 26079 31998 26080
tri 31861 26078 31862 26079 ne
rect 31862 26078 31998 26079
tri 31862 26077 31863 26078 ne
rect 31863 26077 31998 26078
tri 31863 26076 31864 26077 ne
rect 31864 26076 31998 26077
tri 31864 26075 31865 26076 ne
rect 31865 26075 31998 26076
tri 31865 26074 31866 26075 ne
rect 31866 26074 31998 26075
tri 31866 26073 31867 26074 ne
rect 31867 26073 31998 26074
tri 31867 26072 31868 26073 ne
rect 31868 26072 31998 26073
tri 31868 26071 31869 26072 ne
rect 31869 26071 31998 26072
tri 31869 26070 31870 26071 ne
rect 31870 26070 31998 26071
tri 31870 26069 31871 26070 ne
rect 31871 26069 31998 26070
tri 31871 26024 31916 26069 ne
rect 31916 26034 31998 26069
rect 32044 26069 32102 26080
tri 32102 26069 32147 26114 sw
rect 70802 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26034 32147 26069
rect 31916 26024 32147 26034
tri 32147 26024 32192 26069 sw
tri 31916 25979 31961 26024 ne
rect 31961 25979 32192 26024
tri 32192 25979 32237 26024 sw
rect 70802 26020 71000 26078
tri 31961 25934 32006 25979 ne
rect 32006 25965 32237 25979
tri 32237 25965 32251 25979 sw
rect 70802 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 32006 25948 32251 25965
rect 32006 25934 32130 25948
tri 32006 25920 32020 25934 ne
rect 32020 25920 32130 25934
tri 32020 25913 32027 25920 ne
rect 32027 25913 32130 25920
tri 32027 25912 32028 25913 ne
rect 32028 25912 32130 25913
tri 32028 25911 32029 25912 ne
rect 32029 25911 32130 25912
tri 32029 25910 32030 25911 ne
rect 32030 25910 32130 25911
tri 32030 25909 32031 25910 ne
rect 32031 25909 32130 25910
tri 32031 25908 32032 25909 ne
rect 32032 25908 32130 25909
tri 32032 25907 32033 25908 ne
rect 32033 25907 32130 25908
tri 32033 25906 32034 25907 ne
rect 32034 25906 32130 25907
tri 32034 25905 32035 25906 ne
rect 32035 25905 32130 25906
tri 32035 25904 32036 25905 ne
rect 32036 25904 32130 25905
tri 32036 25903 32037 25904 ne
rect 32037 25903 32130 25904
tri 32037 25902 32038 25903 ne
rect 32038 25902 32130 25903
rect 32176 25920 32251 25948
tri 32251 25920 32296 25965 sw
rect 32176 25902 32296 25920
tri 32038 25901 32039 25902 ne
rect 32039 25901 32296 25902
tri 32039 25900 32040 25901 ne
rect 32040 25900 32296 25901
tri 32040 25899 32041 25900 ne
rect 32041 25899 32296 25900
tri 32041 25898 32042 25899 ne
rect 32042 25898 32296 25899
tri 32042 25897 32043 25898 ne
rect 32043 25897 32296 25898
tri 32043 25896 32044 25897 ne
rect 32044 25896 32296 25897
tri 32044 25895 32045 25896 ne
rect 32045 25895 32296 25896
tri 32045 25894 32046 25895 ne
rect 32046 25894 32296 25895
tri 32046 25893 32047 25894 ne
rect 32047 25893 32296 25894
tri 32047 25892 32048 25893 ne
rect 32048 25892 32296 25893
tri 32048 25891 32049 25892 ne
rect 32049 25891 32296 25892
tri 32049 25890 32050 25891 ne
rect 32050 25890 32296 25891
tri 32050 25889 32051 25890 ne
rect 32051 25889 32296 25890
tri 32051 25888 32052 25889 ne
rect 32052 25888 32296 25889
tri 32052 25887 32053 25888 ne
rect 32053 25887 32296 25888
tri 32053 25886 32054 25887 ne
rect 32054 25886 32296 25887
tri 32054 25885 32055 25886 ne
rect 32055 25885 32296 25886
tri 32055 25884 32056 25885 ne
rect 32056 25884 32296 25885
tri 32056 25883 32057 25884 ne
rect 32057 25883 32296 25884
tri 32057 25882 32058 25883 ne
rect 32058 25882 32296 25883
tri 32058 25881 32059 25882 ne
rect 32059 25881 32296 25882
tri 32059 25880 32060 25881 ne
rect 32060 25880 32296 25881
tri 32060 25879 32061 25880 ne
rect 32061 25879 32296 25880
tri 32061 25878 32062 25879 ne
rect 32062 25878 32296 25879
tri 32062 25877 32063 25878 ne
rect 32063 25877 32296 25878
tri 32063 25876 32064 25877 ne
rect 32064 25876 32296 25877
tri 32064 25875 32065 25876 ne
rect 32065 25875 32296 25876
tri 32296 25875 32341 25920 sw
rect 70802 25916 71000 25974
tri 32065 25874 32066 25875 ne
rect 32066 25874 32341 25875
tri 32066 25873 32067 25874 ne
rect 32067 25873 32341 25874
tri 32067 25872 32068 25873 ne
rect 32068 25872 32341 25873
tri 32068 25871 32069 25872 ne
rect 32069 25871 32341 25872
tri 32069 25870 32070 25871 ne
rect 32070 25870 32341 25871
tri 32070 25869 32071 25870 ne
rect 32071 25869 32341 25870
tri 32071 25868 32072 25869 ne
rect 32072 25868 32341 25869
tri 32072 25867 32073 25868 ne
rect 32073 25867 32341 25868
tri 32073 25866 32074 25867 ne
rect 32074 25866 32341 25867
tri 32074 25865 32075 25866 ne
rect 32075 25865 32341 25866
tri 32075 25864 32076 25865 ne
rect 32076 25864 32341 25865
tri 32076 25863 32077 25864 ne
rect 32077 25863 32341 25864
tri 32077 25862 32078 25863 ne
rect 32078 25862 32341 25863
tri 32078 25861 32079 25862 ne
rect 32079 25861 32341 25862
tri 32079 25860 32080 25861 ne
rect 32080 25860 32341 25861
tri 32080 25859 32081 25860 ne
rect 32081 25859 32341 25860
tri 32081 25858 32082 25859 ne
rect 32082 25858 32341 25859
tri 32082 25857 32083 25858 ne
rect 32083 25857 32341 25858
tri 32083 25856 32084 25857 ne
rect 32084 25856 32341 25857
tri 32084 25855 32085 25856 ne
rect 32085 25855 32341 25856
tri 32085 25854 32086 25855 ne
rect 32086 25854 32341 25855
tri 32086 25853 32087 25854 ne
rect 32087 25853 32341 25854
tri 32087 25852 32088 25853 ne
rect 32088 25852 32341 25853
tri 32088 25851 32089 25852 ne
rect 32089 25851 32341 25852
tri 32089 25850 32090 25851 ne
rect 32090 25850 32341 25851
tri 32090 25849 32091 25850 ne
rect 32091 25849 32341 25850
tri 32091 25848 32092 25849 ne
rect 32092 25848 32341 25849
tri 32092 25847 32093 25848 ne
rect 32093 25847 32341 25848
tri 32093 25846 32094 25847 ne
rect 32094 25846 32341 25847
tri 32094 25845 32095 25846 ne
rect 32095 25845 32341 25846
tri 32095 25844 32096 25845 ne
rect 32096 25844 32341 25845
tri 32096 25843 32097 25844 ne
rect 32097 25843 32341 25844
tri 32097 25842 32098 25843 ne
rect 32098 25842 32341 25843
tri 32098 25841 32099 25842 ne
rect 32099 25841 32341 25842
tri 32099 25840 32100 25841 ne
rect 32100 25840 32341 25841
tri 32100 25839 32101 25840 ne
rect 32101 25839 32341 25840
tri 32101 25838 32102 25839 ne
rect 32102 25838 32341 25839
tri 32102 25837 32103 25838 ne
rect 32103 25837 32341 25838
tri 32103 25836 32104 25837 ne
rect 32104 25836 32341 25837
tri 32104 25835 32105 25836 ne
rect 32105 25835 32341 25836
tri 32105 25834 32106 25835 ne
rect 32106 25834 32341 25835
tri 32106 25833 32107 25834 ne
rect 32107 25833 32341 25834
tri 32107 25832 32108 25833 ne
rect 32108 25832 32341 25833
tri 32108 25831 32109 25832 ne
rect 32109 25831 32341 25832
tri 32109 25830 32110 25831 ne
rect 32110 25830 32341 25831
tri 32341 25830 32386 25875 sw
rect 70802 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32110 25829 32111 25830 ne
rect 32111 25829 32386 25830
tri 32111 25828 32112 25829 ne
rect 32112 25828 32386 25829
tri 32112 25827 32113 25828 ne
rect 32113 25827 32386 25828
tri 32113 25826 32114 25827 ne
rect 32114 25826 32386 25827
tri 32114 25825 32115 25826 ne
rect 32115 25825 32386 25826
tri 32115 25824 32116 25825 ne
rect 32116 25824 32386 25825
tri 32116 25823 32117 25824 ne
rect 32117 25823 32386 25824
tri 32117 25822 32118 25823 ne
rect 32118 25822 32386 25823
tri 32118 25821 32119 25822 ne
rect 32119 25821 32386 25822
tri 32119 25820 32120 25821 ne
rect 32120 25820 32386 25821
tri 32120 25819 32121 25820 ne
rect 32121 25819 32386 25820
tri 32121 25818 32122 25819 ne
rect 32122 25818 32386 25819
tri 32122 25817 32123 25818 ne
rect 32123 25817 32386 25818
tri 32123 25816 32124 25817 ne
rect 32124 25816 32386 25817
tri 32124 25815 32125 25816 ne
rect 32125 25815 32262 25816
tri 32125 25814 32126 25815 ne
rect 32126 25814 32262 25815
tri 32126 25813 32127 25814 ne
rect 32127 25813 32262 25814
tri 32127 25812 32128 25813 ne
rect 32128 25812 32262 25813
tri 32128 25811 32129 25812 ne
rect 32129 25811 32262 25812
tri 32129 25810 32130 25811 ne
rect 32130 25810 32262 25811
tri 32130 25809 32131 25810 ne
rect 32131 25809 32262 25810
tri 32131 25808 32132 25809 ne
rect 32132 25808 32262 25809
tri 32132 25807 32133 25808 ne
rect 32133 25807 32262 25808
tri 32133 25806 32134 25807 ne
rect 32134 25806 32262 25807
tri 32134 25805 32135 25806 ne
rect 32135 25805 32262 25806
tri 32135 25804 32136 25805 ne
rect 32136 25804 32262 25805
tri 32136 25803 32137 25804 ne
rect 32137 25803 32262 25804
tri 32137 25802 32138 25803 ne
rect 32138 25802 32262 25803
tri 32138 25801 32139 25802 ne
rect 32139 25801 32262 25802
tri 32139 25800 32140 25801 ne
rect 32140 25800 32262 25801
tri 32140 25799 32141 25800 ne
rect 32141 25799 32262 25800
tri 32141 25798 32142 25799 ne
rect 32142 25798 32262 25799
tri 32142 25797 32143 25798 ne
rect 32143 25797 32262 25798
tri 32143 25796 32144 25797 ne
rect 32144 25796 32262 25797
tri 32144 25795 32145 25796 ne
rect 32145 25795 32262 25796
tri 32145 25794 32146 25795 ne
rect 32146 25794 32262 25795
tri 32146 25793 32147 25794 ne
rect 32147 25793 32262 25794
tri 32147 25771 32169 25793 ne
rect 32169 25771 32262 25793
tri 32169 25726 32214 25771 ne
rect 32214 25770 32262 25771
rect 32308 25793 32386 25816
tri 32386 25793 32423 25830 sw
rect 70802 25812 71000 25870
rect 32308 25770 32423 25793
rect 32214 25748 32423 25770
tri 32423 25748 32468 25793 sw
rect 70802 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 32214 25726 32468 25748
tri 32214 25681 32259 25726 ne
rect 32259 25703 32468 25726
tri 32468 25703 32513 25748 sw
rect 70802 25708 71000 25766
rect 32259 25684 32513 25703
rect 32259 25681 32394 25684
tri 32259 25639 32301 25681 ne
rect 32301 25639 32394 25681
tri 32301 25638 32302 25639 ne
rect 32302 25638 32394 25639
rect 32440 25658 32513 25684
tri 32513 25658 32558 25703 sw
rect 70802 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25652 32558 25658
tri 32558 25652 32564 25658 sw
rect 32440 25638 32564 25652
tri 32302 25637 32303 25638 ne
rect 32303 25637 32564 25638
tri 32303 25636 32304 25637 ne
rect 32304 25636 32564 25637
tri 32304 25635 32305 25636 ne
rect 32305 25635 32564 25636
tri 32305 25634 32306 25635 ne
rect 32306 25634 32564 25635
tri 32306 25633 32307 25634 ne
rect 32307 25633 32564 25634
tri 32307 25632 32308 25633 ne
rect 32308 25632 32564 25633
tri 32308 25631 32309 25632 ne
rect 32309 25631 32564 25632
tri 32309 25630 32310 25631 ne
rect 32310 25630 32564 25631
tri 32310 25629 32311 25630 ne
rect 32311 25629 32564 25630
tri 32311 25628 32312 25629 ne
rect 32312 25628 32564 25629
tri 32312 25627 32313 25628 ne
rect 32313 25627 32564 25628
tri 32313 25626 32314 25627 ne
rect 32314 25626 32564 25627
tri 32314 25625 32315 25626 ne
rect 32315 25625 32564 25626
tri 32315 25624 32316 25625 ne
rect 32316 25624 32564 25625
tri 32316 25623 32317 25624 ne
rect 32317 25623 32564 25624
tri 32317 25622 32318 25623 ne
rect 32318 25622 32564 25623
tri 32318 25621 32319 25622 ne
rect 32319 25621 32564 25622
tri 32319 25620 32320 25621 ne
rect 32320 25620 32564 25621
tri 32320 25619 32321 25620 ne
rect 32321 25619 32564 25620
tri 32321 25618 32322 25619 ne
rect 32322 25618 32564 25619
tri 32322 25617 32323 25618 ne
rect 32323 25617 32564 25618
tri 32323 25616 32324 25617 ne
rect 32324 25616 32564 25617
tri 32324 25615 32325 25616 ne
rect 32325 25615 32564 25616
tri 32325 25614 32326 25615 ne
rect 32326 25614 32564 25615
tri 32326 25613 32327 25614 ne
rect 32327 25613 32564 25614
tri 32327 25612 32328 25613 ne
rect 32328 25612 32564 25613
tri 32328 25611 32329 25612 ne
rect 32329 25611 32564 25612
tri 32329 25610 32330 25611 ne
rect 32330 25610 32564 25611
tri 32330 25609 32331 25610 ne
rect 32331 25609 32564 25610
tri 32331 25608 32332 25609 ne
rect 32332 25608 32564 25609
tri 32332 25607 32333 25608 ne
rect 32333 25607 32564 25608
tri 32564 25607 32609 25652 sw
tri 32333 25606 32334 25607 ne
rect 32334 25606 32609 25607
tri 32334 25605 32335 25606 ne
rect 32335 25605 32609 25606
tri 32335 25604 32336 25605 ne
rect 32336 25604 32609 25605
tri 32336 25603 32337 25604 ne
rect 32337 25603 32609 25604
tri 32337 25602 32338 25603 ne
rect 32338 25602 32609 25603
tri 32338 25601 32339 25602 ne
rect 32339 25601 32609 25602
tri 32339 25600 32340 25601 ne
rect 32340 25600 32609 25601
tri 32340 25599 32341 25600 ne
rect 32341 25599 32609 25600
tri 32341 25598 32342 25599 ne
rect 32342 25598 32609 25599
tri 32342 25597 32343 25598 ne
rect 32343 25597 32609 25598
tri 32343 25596 32344 25597 ne
rect 32344 25596 32609 25597
tri 32344 25595 32345 25596 ne
rect 32345 25595 32609 25596
tri 32345 25594 32346 25595 ne
rect 32346 25594 32609 25595
tri 32346 25593 32347 25594 ne
rect 32347 25593 32609 25594
tri 32347 25592 32348 25593 ne
rect 32348 25592 32609 25593
tri 32348 25591 32349 25592 ne
rect 32349 25591 32609 25592
tri 32349 25590 32350 25591 ne
rect 32350 25590 32609 25591
tri 32350 25589 32351 25590 ne
rect 32351 25589 32609 25590
tri 32351 25588 32352 25589 ne
rect 32352 25588 32609 25589
tri 32352 25587 32353 25588 ne
rect 32353 25587 32609 25588
tri 32353 25586 32354 25587 ne
rect 32354 25586 32609 25587
tri 32354 25585 32355 25586 ne
rect 32355 25585 32609 25586
tri 32355 25584 32356 25585 ne
rect 32356 25584 32609 25585
tri 32356 25583 32357 25584 ne
rect 32357 25583 32609 25584
tri 32357 25582 32358 25583 ne
rect 32358 25582 32609 25583
tri 32358 25581 32359 25582 ne
rect 32359 25581 32609 25582
tri 32359 25580 32360 25581 ne
rect 32360 25580 32609 25581
tri 32360 25579 32361 25580 ne
rect 32361 25579 32609 25580
tri 32361 25578 32362 25579 ne
rect 32362 25578 32609 25579
tri 32362 25577 32363 25578 ne
rect 32363 25577 32609 25578
tri 32363 25576 32364 25577 ne
rect 32364 25576 32609 25577
tri 32364 25575 32365 25576 ne
rect 32365 25575 32609 25576
tri 32365 25574 32366 25575 ne
rect 32366 25574 32609 25575
tri 32366 25573 32367 25574 ne
rect 32367 25573 32609 25574
tri 32367 25572 32368 25573 ne
rect 32368 25572 32609 25573
tri 32368 25571 32369 25572 ne
rect 32369 25571 32609 25572
tri 32369 25570 32370 25571 ne
rect 32370 25570 32609 25571
tri 32370 25569 32371 25570 ne
rect 32371 25569 32609 25570
tri 32371 25568 32372 25569 ne
rect 32372 25568 32609 25569
tri 32372 25567 32373 25568 ne
rect 32373 25567 32609 25568
tri 32373 25566 32374 25567 ne
rect 32374 25566 32609 25567
tri 32374 25565 32375 25566 ne
rect 32375 25565 32609 25566
tri 32375 25564 32376 25565 ne
rect 32376 25564 32609 25565
tri 32376 25563 32377 25564 ne
rect 32377 25563 32609 25564
tri 32377 25562 32378 25563 ne
rect 32378 25562 32609 25563
tri 32609 25562 32654 25607 sw
rect 70802 25604 71000 25662
tri 32378 25561 32379 25562 ne
rect 32379 25561 32654 25562
tri 32379 25560 32380 25561 ne
rect 32380 25560 32654 25561
tri 32380 25559 32381 25560 ne
rect 32381 25559 32654 25560
tri 32381 25558 32382 25559 ne
rect 32382 25558 32654 25559
tri 32382 25557 32383 25558 ne
rect 32383 25557 32654 25558
tri 32383 25556 32384 25557 ne
rect 32384 25556 32654 25557
tri 32384 25555 32385 25556 ne
rect 32385 25555 32654 25556
tri 32385 25554 32386 25555 ne
rect 32386 25554 32654 25555
tri 32386 25553 32387 25554 ne
rect 32387 25553 32654 25554
tri 32387 25552 32388 25553 ne
rect 32388 25552 32654 25553
tri 32388 25551 32389 25552 ne
rect 32389 25551 32526 25552
tri 32389 25550 32390 25551 ne
rect 32390 25550 32526 25551
tri 32390 25549 32391 25550 ne
rect 32391 25549 32526 25550
tri 32391 25548 32392 25549 ne
rect 32392 25548 32526 25549
tri 32392 25547 32393 25548 ne
rect 32393 25547 32526 25548
tri 32393 25546 32394 25547 ne
rect 32394 25546 32526 25547
tri 32394 25545 32395 25546 ne
rect 32395 25545 32526 25546
tri 32395 25544 32396 25545 ne
rect 32396 25544 32526 25545
tri 32396 25543 32397 25544 ne
rect 32397 25543 32526 25544
tri 32397 25542 32398 25543 ne
rect 32398 25542 32526 25543
tri 32398 25541 32399 25542 ne
rect 32399 25541 32526 25542
tri 32399 25540 32400 25541 ne
rect 32400 25540 32526 25541
tri 32400 25539 32401 25540 ne
rect 32401 25539 32526 25540
tri 32401 25538 32402 25539 ne
rect 32402 25538 32526 25539
tri 32402 25537 32403 25538 ne
rect 32403 25537 32526 25538
tri 32403 25536 32404 25537 ne
rect 32404 25536 32526 25537
tri 32404 25535 32405 25536 ne
rect 32405 25535 32526 25536
tri 32405 25534 32406 25535 ne
rect 32406 25534 32526 25535
tri 32406 25533 32407 25534 ne
rect 32407 25533 32526 25534
tri 32407 25532 32408 25533 ne
rect 32408 25532 32526 25533
tri 32408 25531 32409 25532 ne
rect 32409 25531 32526 25532
tri 32409 25530 32410 25531 ne
rect 32410 25530 32526 25531
tri 32410 25529 32411 25530 ne
rect 32411 25529 32526 25530
tri 32411 25528 32412 25529 ne
rect 32412 25528 32526 25529
tri 32412 25527 32413 25528 ne
rect 32413 25527 32526 25528
tri 32413 25526 32414 25527 ne
rect 32414 25526 32526 25527
tri 32414 25525 32415 25526 ne
rect 32415 25525 32526 25526
tri 32415 25524 32416 25525 ne
rect 32416 25524 32526 25525
tri 32416 25523 32417 25524 ne
rect 32417 25523 32526 25524
tri 32417 25522 32418 25523 ne
rect 32418 25522 32526 25523
tri 32418 25521 32419 25522 ne
rect 32419 25521 32526 25522
tri 32419 25520 32420 25521 ne
rect 32420 25520 32526 25521
tri 32420 25519 32421 25520 ne
rect 32421 25519 32526 25520
tri 32421 25518 32422 25519 ne
rect 32422 25518 32526 25519
tri 32422 25517 32423 25518 ne
rect 32423 25517 32526 25518
tri 32423 25509 32431 25517 ne
rect 32431 25509 32526 25517
tri 32431 25464 32476 25509 ne
rect 32476 25506 32526 25509
rect 32572 25517 32654 25552
tri 32654 25517 32699 25562 sw
rect 70802 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32572 25509 32699 25517
tri 32699 25509 32707 25517 sw
rect 32572 25506 32707 25509
rect 32476 25464 32707 25506
tri 32707 25464 32752 25509 sw
rect 70802 25500 71000 25558
tri 32476 25451 32489 25464 ne
rect 32489 25451 32752 25464
tri 32489 25406 32534 25451 ne
rect 32534 25420 32752 25451
rect 32534 25406 32658 25420
tri 32534 25365 32575 25406 ne
rect 32575 25374 32658 25406
rect 32704 25419 32752 25420
tri 32752 25419 32797 25464 sw
rect 70802 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32704 25374 32797 25419
tri 32797 25374 32842 25419 sw
rect 70802 25396 71000 25454
rect 32575 25365 32842 25374
tri 32575 25364 32576 25365 ne
rect 32576 25364 32842 25365
tri 32576 25363 32577 25364 ne
rect 32577 25363 32842 25364
tri 32577 25362 32578 25363 ne
rect 32578 25362 32842 25363
tri 32578 25361 32579 25362 ne
rect 32579 25361 32842 25362
tri 32579 25360 32580 25361 ne
rect 32580 25360 32842 25361
tri 32580 25359 32581 25360 ne
rect 32581 25359 32842 25360
tri 32581 25358 32582 25359 ne
rect 32582 25358 32842 25359
tri 32582 25357 32583 25358 ne
rect 32583 25357 32842 25358
tri 32583 25356 32584 25357 ne
rect 32584 25356 32842 25357
tri 32584 25355 32585 25356 ne
rect 32585 25355 32842 25356
tri 32585 25354 32586 25355 ne
rect 32586 25354 32842 25355
tri 32586 25353 32587 25354 ne
rect 32587 25353 32842 25354
tri 32587 25352 32588 25353 ne
rect 32588 25352 32842 25353
tri 32588 25351 32589 25352 ne
rect 32589 25351 32842 25352
tri 32589 25350 32590 25351 ne
rect 32590 25350 32842 25351
tri 32590 25349 32591 25350 ne
rect 32591 25349 32842 25350
tri 32591 25348 32592 25349 ne
rect 32592 25348 32842 25349
tri 32592 25347 32593 25348 ne
rect 32593 25347 32842 25348
tri 32593 25346 32594 25347 ne
rect 32594 25346 32842 25347
tri 32594 25345 32595 25346 ne
rect 32595 25345 32842 25346
tri 32595 25344 32596 25345 ne
rect 32596 25344 32842 25345
tri 32596 25343 32597 25344 ne
rect 32597 25343 32842 25344
tri 32597 25342 32598 25343 ne
rect 32598 25342 32842 25343
tri 32598 25341 32599 25342 ne
rect 32599 25341 32842 25342
tri 32599 25340 32600 25341 ne
rect 32600 25340 32842 25341
tri 32600 25339 32601 25340 ne
rect 32601 25339 32842 25340
tri 32601 25338 32602 25339 ne
rect 32602 25338 32842 25339
tri 32602 25337 32603 25338 ne
rect 32603 25337 32842 25338
tri 32603 25336 32604 25337 ne
rect 32604 25336 32842 25337
tri 32604 25335 32605 25336 ne
rect 32605 25335 32842 25336
tri 32605 25334 32606 25335 ne
rect 32606 25334 32842 25335
tri 32606 25333 32607 25334 ne
rect 32607 25333 32842 25334
tri 32607 25332 32608 25333 ne
rect 32608 25332 32842 25333
tri 32608 25331 32609 25332 ne
rect 32609 25331 32842 25332
tri 32842 25331 32885 25374 sw
rect 70802 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
tri 32609 25330 32610 25331 ne
rect 32610 25330 32885 25331
tri 32610 25329 32611 25330 ne
rect 32611 25329 32885 25330
tri 32611 25328 32612 25329 ne
rect 32612 25328 32885 25329
tri 32612 25327 32613 25328 ne
rect 32613 25327 32885 25328
tri 32613 25326 32614 25327 ne
rect 32614 25326 32885 25327
tri 32614 25325 32615 25326 ne
rect 32615 25325 32885 25326
tri 32615 25324 32616 25325 ne
rect 32616 25324 32885 25325
tri 32616 25323 32617 25324 ne
rect 32617 25323 32885 25324
tri 32617 25322 32618 25323 ne
rect 32618 25322 32885 25323
tri 32618 25321 32619 25322 ne
rect 32619 25321 32885 25322
tri 32619 25320 32620 25321 ne
rect 32620 25320 32885 25321
tri 32620 25319 32621 25320 ne
rect 32621 25319 32885 25320
tri 32621 25318 32622 25319 ne
rect 32622 25318 32885 25319
tri 32622 25317 32623 25318 ne
rect 32623 25317 32885 25318
tri 32623 25316 32624 25317 ne
rect 32624 25316 32885 25317
tri 32624 25315 32625 25316 ne
rect 32625 25315 32885 25316
tri 32625 25314 32626 25315 ne
rect 32626 25314 32885 25315
tri 32626 25313 32627 25314 ne
rect 32627 25313 32885 25314
tri 32627 25312 32628 25313 ne
rect 32628 25312 32885 25313
tri 32628 25311 32629 25312 ne
rect 32629 25311 32885 25312
tri 32629 25310 32630 25311 ne
rect 32630 25310 32885 25311
tri 32630 25309 32631 25310 ne
rect 32631 25309 32885 25310
tri 32631 25308 32632 25309 ne
rect 32632 25308 32885 25309
tri 32632 25307 32633 25308 ne
rect 32633 25307 32885 25308
tri 32633 25306 32634 25307 ne
rect 32634 25306 32885 25307
tri 32634 25305 32635 25306 ne
rect 32635 25305 32885 25306
tri 32635 25304 32636 25305 ne
rect 32636 25304 32885 25305
tri 32636 25303 32637 25304 ne
rect 32637 25303 32885 25304
tri 32637 25302 32638 25303 ne
rect 32638 25302 32885 25303
tri 32638 25301 32639 25302 ne
rect 32639 25301 32885 25302
tri 32639 25300 32640 25301 ne
rect 32640 25300 32885 25301
tri 32640 25299 32641 25300 ne
rect 32641 25299 32885 25300
tri 32641 25298 32642 25299 ne
rect 32642 25298 32885 25299
tri 32642 25297 32643 25298 ne
rect 32643 25297 32885 25298
tri 32643 25296 32644 25297 ne
rect 32644 25296 32885 25297
tri 32644 25295 32645 25296 ne
rect 32645 25295 32885 25296
tri 32645 25294 32646 25295 ne
rect 32646 25294 32885 25295
tri 32646 25293 32647 25294 ne
rect 32647 25293 32885 25294
tri 32647 25292 32648 25293 ne
rect 32648 25292 32885 25293
tri 32648 25291 32649 25292 ne
rect 32649 25291 32885 25292
tri 32649 25290 32650 25291 ne
rect 32650 25290 32885 25291
tri 32650 25289 32651 25290 ne
rect 32651 25289 32885 25290
tri 32651 25288 32652 25289 ne
rect 32652 25288 32885 25289
tri 32652 25287 32653 25288 ne
rect 32653 25287 32790 25288
tri 32653 25286 32654 25287 ne
rect 32654 25286 32790 25287
tri 32654 25285 32655 25286 ne
rect 32655 25285 32790 25286
tri 32655 25284 32656 25285 ne
rect 32656 25284 32790 25285
tri 32656 25283 32657 25284 ne
rect 32657 25283 32790 25284
tri 32657 25282 32658 25283 ne
rect 32658 25282 32790 25283
tri 32658 25281 32659 25282 ne
rect 32659 25281 32790 25282
tri 32659 25280 32660 25281 ne
rect 32660 25280 32790 25281
tri 32660 25279 32661 25280 ne
rect 32661 25279 32790 25280
tri 32661 25278 32662 25279 ne
rect 32662 25278 32790 25279
tri 32662 25277 32663 25278 ne
rect 32663 25277 32790 25278
tri 32663 25276 32664 25277 ne
rect 32664 25276 32790 25277
tri 32664 25275 32665 25276 ne
rect 32665 25275 32790 25276
tri 32665 25274 32666 25275 ne
rect 32666 25274 32790 25275
tri 32666 25273 32667 25274 ne
rect 32667 25273 32790 25274
tri 32667 25272 32668 25273 ne
rect 32668 25272 32790 25273
tri 32668 25271 32669 25272 ne
rect 32669 25271 32790 25272
tri 32669 25270 32670 25271 ne
rect 32670 25270 32790 25271
tri 32670 25269 32671 25270 ne
rect 32671 25269 32790 25270
tri 32671 25268 32672 25269 ne
rect 32672 25268 32790 25269
tri 32672 25267 32673 25268 ne
rect 32673 25267 32790 25268
tri 32673 25266 32674 25267 ne
rect 32674 25266 32790 25267
tri 32674 25265 32675 25266 ne
rect 32675 25265 32790 25266
tri 32675 25264 32676 25265 ne
rect 32676 25264 32790 25265
tri 32676 25263 32677 25264 ne
rect 32677 25263 32790 25264
tri 32677 25262 32678 25263 ne
rect 32678 25262 32790 25263
tri 32678 25261 32679 25262 ne
rect 32679 25261 32790 25262
tri 32679 25260 32680 25261 ne
rect 32680 25260 32790 25261
tri 32680 25259 32681 25260 ne
rect 32681 25259 32790 25260
tri 32681 25258 32682 25259 ne
rect 32682 25258 32790 25259
tri 32682 25257 32683 25258 ne
rect 32683 25257 32790 25258
tri 32683 25256 32684 25257 ne
rect 32684 25256 32790 25257
tri 32684 25255 32685 25256 ne
rect 32685 25255 32790 25256
tri 32685 25254 32686 25255 ne
rect 32686 25254 32790 25255
tri 32686 25253 32687 25254 ne
rect 32687 25253 32790 25254
tri 32687 25252 32688 25253 ne
rect 32688 25252 32790 25253
tri 32688 25251 32689 25252 ne
rect 32689 25251 32790 25252
tri 32689 25250 32690 25251 ne
rect 32690 25250 32790 25251
tri 32690 25249 32691 25250 ne
rect 32691 25249 32790 25250
tri 32691 25248 32692 25249 ne
rect 32692 25248 32790 25249
tri 32692 25247 32693 25248 ne
rect 32693 25247 32790 25248
tri 32693 25246 32694 25247 ne
rect 32694 25246 32790 25247
tri 32694 25245 32695 25246 ne
rect 32695 25245 32790 25246
tri 32695 25244 32696 25245 ne
rect 32696 25244 32790 25245
tri 32696 25243 32697 25244 ne
rect 32697 25243 32790 25244
tri 32697 25242 32698 25243 ne
rect 32698 25242 32790 25243
rect 32836 25286 32885 25288
tri 32885 25286 32930 25331 sw
rect 70802 25292 71000 25350
rect 32836 25242 32930 25286
tri 32698 25241 32699 25242 ne
rect 32699 25241 32930 25242
tri 32930 25241 32975 25286 sw
rect 70802 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
tri 32699 25196 32744 25241 ne
rect 32744 25196 32975 25241
tri 32975 25196 33020 25241 sw
tri 32744 25188 32752 25196 ne
rect 32752 25188 33020 25196
tri 33020 25188 33028 25196 sw
rect 70802 25188 71000 25246
tri 32752 25151 32789 25188 ne
rect 32789 25156 33028 25188
rect 32789 25151 32922 25156
tri 32789 25143 32797 25151 ne
rect 32797 25143 32922 25151
tri 32797 25098 32842 25143 ne
rect 32842 25110 32922 25143
rect 32968 25143 33028 25156
tri 33028 25143 33073 25188 sw
rect 32968 25110 33073 25143
rect 32842 25098 33073 25110
tri 33073 25098 33118 25143 sw
rect 70802 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
tri 32842 25090 32850 25098 ne
rect 32850 25090 33118 25098
tri 32850 25089 32851 25090 ne
rect 32851 25089 33118 25090
tri 32851 25088 32852 25089 ne
rect 32852 25088 33118 25089
tri 32852 25087 32853 25088 ne
rect 32853 25087 33118 25088
tri 32853 25086 32854 25087 ne
rect 32854 25086 33118 25087
tri 32854 25085 32855 25086 ne
rect 32855 25085 33118 25086
tri 32855 25084 32856 25085 ne
rect 32856 25084 33118 25085
tri 32856 25083 32857 25084 ne
rect 32857 25083 33118 25084
tri 32857 25082 32858 25083 ne
rect 32858 25082 33118 25083
tri 32858 25081 32859 25082 ne
rect 32859 25081 33118 25082
tri 32859 25080 32860 25081 ne
rect 32860 25080 33118 25081
tri 32860 25079 32861 25080 ne
rect 32861 25079 33118 25080
tri 32861 25078 32862 25079 ne
rect 32862 25078 33118 25079
tri 32862 25077 32863 25078 ne
rect 32863 25077 33118 25078
tri 32863 25076 32864 25077 ne
rect 32864 25076 33118 25077
tri 32864 25075 32865 25076 ne
rect 32865 25075 33118 25076
tri 32865 25074 32866 25075 ne
rect 32866 25074 33118 25075
tri 32866 25073 32867 25074 ne
rect 32867 25073 33118 25074
tri 32867 25072 32868 25073 ne
rect 32868 25072 33118 25073
tri 32868 25071 32869 25072 ne
rect 32869 25071 33118 25072
tri 32869 25070 32870 25071 ne
rect 32870 25070 33118 25071
tri 32870 25069 32871 25070 ne
rect 32871 25069 33118 25070
tri 32871 25068 32872 25069 ne
rect 32872 25068 33118 25069
tri 32872 25067 32873 25068 ne
rect 32873 25067 33118 25068
tri 32873 25066 32874 25067 ne
rect 32874 25066 33118 25067
tri 32874 25065 32875 25066 ne
rect 32875 25065 33118 25066
tri 32875 25064 32876 25065 ne
rect 32876 25064 33118 25065
tri 32876 25063 32877 25064 ne
rect 32877 25063 33118 25064
tri 32877 25062 32878 25063 ne
rect 32878 25062 33118 25063
tri 32878 25061 32879 25062 ne
rect 32879 25061 33118 25062
tri 32879 25060 32880 25061 ne
rect 32880 25060 33118 25061
tri 32880 25059 32881 25060 ne
rect 32881 25059 33118 25060
tri 32881 25058 32882 25059 ne
rect 32882 25058 33118 25059
tri 32882 25057 32883 25058 ne
rect 32883 25057 33118 25058
tri 32883 25056 32884 25057 ne
rect 32884 25056 33118 25057
tri 32884 25055 32885 25056 ne
rect 32885 25055 33118 25056
tri 32885 25054 32886 25055 ne
rect 32886 25054 33118 25055
tri 32886 25053 32887 25054 ne
rect 32887 25053 33118 25054
tri 33118 25053 33163 25098 sw
rect 70802 25084 71000 25142
tri 32887 25052 32888 25053 ne
rect 32888 25052 33163 25053
tri 32888 25051 32889 25052 ne
rect 32889 25051 33163 25052
tri 32889 25050 32890 25051 ne
rect 32890 25050 33163 25051
tri 32890 25049 32891 25050 ne
rect 32891 25049 33163 25050
tri 32891 25048 32892 25049 ne
rect 32892 25048 33163 25049
tri 32892 25047 32893 25048 ne
rect 32893 25047 33163 25048
tri 32893 25046 32894 25047 ne
rect 32894 25046 33163 25047
tri 32894 25045 32895 25046 ne
rect 32895 25045 33163 25046
tri 32895 25044 32896 25045 ne
rect 32896 25044 33163 25045
tri 32896 25043 32897 25044 ne
rect 32897 25043 33163 25044
tri 32897 25042 32898 25043 ne
rect 32898 25042 33163 25043
tri 32898 25041 32899 25042 ne
rect 32899 25041 33163 25042
tri 32899 25040 32900 25041 ne
rect 32900 25040 33163 25041
tri 32900 25039 32901 25040 ne
rect 32901 25039 33163 25040
tri 32901 25038 32902 25039 ne
rect 32902 25038 33163 25039
tri 32902 25037 32903 25038 ne
rect 32903 25037 33163 25038
tri 32903 25036 32904 25037 ne
rect 32904 25036 33163 25037
tri 32904 25035 32905 25036 ne
rect 32905 25035 33163 25036
tri 32905 25034 32906 25035 ne
rect 32906 25034 33163 25035
tri 32906 25033 32907 25034 ne
rect 32907 25033 33163 25034
tri 32907 25032 32908 25033 ne
rect 32908 25032 33163 25033
tri 32908 25031 32909 25032 ne
rect 32909 25031 33163 25032
tri 32909 25030 32910 25031 ne
rect 32910 25030 33163 25031
tri 32910 25029 32911 25030 ne
rect 32911 25029 33163 25030
tri 32911 25028 32912 25029 ne
rect 32912 25028 33163 25029
tri 32912 25027 32913 25028 ne
rect 32913 25027 33163 25028
tri 32913 25026 32914 25027 ne
rect 32914 25026 33163 25027
tri 32914 25025 32915 25026 ne
rect 32915 25025 33163 25026
tri 32915 25024 32916 25025 ne
rect 32916 25024 33163 25025
tri 32916 25023 32917 25024 ne
rect 32917 25023 33054 25024
tri 32917 25022 32918 25023 ne
rect 32918 25022 33054 25023
tri 32918 25021 32919 25022 ne
rect 32919 25021 33054 25022
tri 32919 25020 32920 25021 ne
rect 32920 25020 33054 25021
tri 32920 25019 32921 25020 ne
rect 32921 25019 33054 25020
tri 32921 25018 32922 25019 ne
rect 32922 25018 33054 25019
tri 32922 25017 32923 25018 ne
rect 32923 25017 33054 25018
tri 32923 25016 32924 25017 ne
rect 32924 25016 33054 25017
tri 32924 25015 32925 25016 ne
rect 32925 25015 33054 25016
tri 32925 25014 32926 25015 ne
rect 32926 25014 33054 25015
tri 32926 25013 32927 25014 ne
rect 32927 25013 33054 25014
tri 32927 25012 32928 25013 ne
rect 32928 25012 33054 25013
tri 32928 25011 32929 25012 ne
rect 32929 25011 33054 25012
tri 32929 25010 32930 25011 ne
rect 32930 25010 33054 25011
tri 32930 25009 32931 25010 ne
rect 32931 25009 33054 25010
tri 32931 25008 32932 25009 ne
rect 32932 25008 33054 25009
tri 32932 25007 32933 25008 ne
rect 32933 25007 33054 25008
tri 32933 25006 32934 25007 ne
rect 32934 25006 33054 25007
tri 32934 25005 32935 25006 ne
rect 32935 25005 33054 25006
tri 32935 25004 32936 25005 ne
rect 32936 25004 33054 25005
tri 32936 25003 32937 25004 ne
rect 32937 25003 33054 25004
tri 32937 25002 32938 25003 ne
rect 32938 25002 33054 25003
tri 32938 25001 32939 25002 ne
rect 32939 25001 33054 25002
tri 32939 25000 32940 25001 ne
rect 32940 25000 33054 25001
tri 32940 24999 32941 25000 ne
rect 32941 24999 33054 25000
tri 32941 24998 32942 24999 ne
rect 32942 24998 33054 24999
tri 32942 24997 32943 24998 ne
rect 32943 24997 33054 24998
tri 32943 24996 32944 24997 ne
rect 32944 24996 33054 24997
tri 32944 24995 32945 24996 ne
rect 32945 24995 33054 24996
tri 32945 24994 32946 24995 ne
rect 32946 24994 33054 24995
tri 32946 24993 32947 24994 ne
rect 32947 24993 33054 24994
tri 32947 24992 32948 24993 ne
rect 32948 24992 33054 24993
tri 32948 24991 32949 24992 ne
rect 32949 24991 33054 24992
tri 32949 24990 32950 24991 ne
rect 32950 24990 33054 24991
tri 32950 24989 32951 24990 ne
rect 32951 24989 33054 24990
tri 32951 24988 32952 24989 ne
rect 32952 24988 33054 24989
tri 32952 24987 32953 24988 ne
rect 32953 24987 33054 24988
tri 32953 24986 32954 24987 ne
rect 32954 24986 33054 24987
tri 32954 24985 32955 24986 ne
rect 32955 24985 33054 24986
tri 32955 24984 32956 24985 ne
rect 32956 24984 33054 24985
tri 32956 24983 32957 24984 ne
rect 32957 24983 33054 24984
tri 32957 24982 32958 24983 ne
rect 32958 24982 33054 24983
tri 32958 24981 32959 24982 ne
rect 32959 24981 33054 24982
tri 32959 24980 32960 24981 ne
rect 32960 24980 33054 24981
tri 32960 24979 32961 24980 ne
rect 32961 24979 33054 24980
tri 32961 24978 32962 24979 ne
rect 32962 24978 33054 24979
rect 33100 25010 33163 25024
tri 33163 25010 33206 25053 sw
rect 70802 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 33100 24978 33206 25010
tri 32962 24977 32963 24978 ne
rect 32963 24977 33206 24978
tri 32963 24976 32964 24977 ne
rect 32964 24976 33206 24977
tri 32964 24975 32965 24976 ne
rect 32965 24975 33206 24976
tri 32965 24974 32966 24975 ne
rect 32966 24974 33206 24975
tri 32966 24973 32967 24974 ne
rect 32967 24973 33206 24974
tri 32967 24972 32968 24973 ne
rect 32968 24972 33206 24973
tri 32968 24971 32969 24972 ne
rect 32969 24971 33206 24972
tri 32969 24970 32970 24971 ne
rect 32970 24970 33206 24971
tri 32970 24969 32971 24970 ne
rect 32971 24969 33206 24970
tri 32971 24968 32972 24969 ne
rect 32972 24968 33206 24969
tri 32972 24967 32973 24968 ne
rect 32973 24967 33206 24968
tri 32973 24966 32974 24967 ne
rect 32974 24966 33206 24967
tri 32974 24965 32975 24966 ne
rect 32975 24965 33206 24966
tri 33206 24965 33251 25010 sw
rect 70802 24980 71000 25038
tri 32975 24920 33020 24965 ne
rect 33020 24920 33251 24965
tri 33251 24920 33296 24965 sw
rect 70802 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33020 24875 33065 24920 ne
rect 33065 24892 33296 24920
rect 33065 24875 33186 24892
tri 33065 24830 33110 24875 ne
rect 33110 24846 33186 24875
rect 33232 24875 33296 24892
tri 33296 24875 33341 24920 sw
rect 70802 24876 71000 24934
rect 33232 24867 33341 24875
tri 33341 24867 33349 24875 sw
rect 33232 24846 33349 24867
rect 33110 24830 33349 24846
tri 33110 24822 33118 24830 ne
rect 33118 24822 33349 24830
tri 33349 24822 33394 24867 sw
rect 70802 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
tri 33118 24816 33124 24822 ne
rect 33124 24816 33394 24822
tri 33124 24815 33125 24816 ne
rect 33125 24815 33394 24816
tri 33125 24814 33126 24815 ne
rect 33126 24814 33394 24815
tri 33126 24813 33127 24814 ne
rect 33127 24813 33394 24814
tri 33127 24812 33128 24813 ne
rect 33128 24812 33394 24813
tri 33128 24811 33129 24812 ne
rect 33129 24811 33394 24812
tri 33129 24810 33130 24811 ne
rect 33130 24810 33394 24811
tri 33130 24809 33131 24810 ne
rect 33131 24809 33394 24810
tri 33131 24808 33132 24809 ne
rect 33132 24808 33394 24809
tri 33132 24807 33133 24808 ne
rect 33133 24807 33394 24808
tri 33133 24806 33134 24807 ne
rect 33134 24806 33394 24807
tri 33134 24805 33135 24806 ne
rect 33135 24805 33394 24806
tri 33135 24804 33136 24805 ne
rect 33136 24804 33394 24805
tri 33136 24803 33137 24804 ne
rect 33137 24803 33394 24804
tri 33137 24802 33138 24803 ne
rect 33138 24802 33394 24803
tri 33138 24801 33139 24802 ne
rect 33139 24801 33394 24802
tri 33139 24800 33140 24801 ne
rect 33140 24800 33394 24801
tri 33140 24799 33141 24800 ne
rect 33141 24799 33394 24800
tri 33141 24798 33142 24799 ne
rect 33142 24798 33394 24799
tri 33142 24797 33143 24798 ne
rect 33143 24797 33394 24798
tri 33143 24796 33144 24797 ne
rect 33144 24796 33394 24797
tri 33144 24795 33145 24796 ne
rect 33145 24795 33394 24796
tri 33145 24794 33146 24795 ne
rect 33146 24794 33394 24795
tri 33146 24793 33147 24794 ne
rect 33147 24793 33394 24794
tri 33147 24792 33148 24793 ne
rect 33148 24792 33394 24793
tri 33148 24791 33149 24792 ne
rect 33149 24791 33394 24792
tri 33149 24790 33150 24791 ne
rect 33150 24790 33394 24791
tri 33150 24789 33151 24790 ne
rect 33151 24789 33394 24790
tri 33151 24788 33152 24789 ne
rect 33152 24788 33394 24789
tri 33152 24787 33153 24788 ne
rect 33153 24787 33394 24788
tri 33153 24786 33154 24787 ne
rect 33154 24786 33394 24787
tri 33154 24785 33155 24786 ne
rect 33155 24785 33394 24786
tri 33155 24784 33156 24785 ne
rect 33156 24784 33394 24785
tri 33156 24783 33157 24784 ne
rect 33157 24783 33394 24784
tri 33157 24782 33158 24783 ne
rect 33158 24782 33394 24783
tri 33158 24781 33159 24782 ne
rect 33159 24781 33394 24782
tri 33159 24780 33160 24781 ne
rect 33160 24780 33394 24781
tri 33160 24779 33161 24780 ne
rect 33161 24779 33394 24780
tri 33161 24778 33162 24779 ne
rect 33162 24778 33394 24779
tri 33162 24777 33163 24778 ne
rect 33163 24777 33394 24778
tri 33394 24777 33439 24822 sw
tri 33163 24776 33164 24777 ne
rect 33164 24776 33439 24777
tri 33164 24775 33165 24776 ne
rect 33165 24775 33439 24776
tri 33165 24774 33166 24775 ne
rect 33166 24774 33439 24775
tri 33166 24773 33167 24774 ne
rect 33167 24773 33439 24774
tri 33167 24772 33168 24773 ne
rect 33168 24772 33439 24773
tri 33168 24771 33169 24772 ne
rect 33169 24771 33439 24772
tri 33169 24770 33170 24771 ne
rect 33170 24770 33439 24771
tri 33170 24769 33171 24770 ne
rect 33171 24769 33439 24770
tri 33171 24768 33172 24769 ne
rect 33172 24768 33439 24769
tri 33172 24767 33173 24768 ne
rect 33173 24767 33439 24768
tri 33173 24766 33174 24767 ne
rect 33174 24766 33439 24767
tri 33174 24765 33175 24766 ne
rect 33175 24765 33439 24766
tri 33175 24764 33176 24765 ne
rect 33176 24764 33439 24765
tri 33176 24763 33177 24764 ne
rect 33177 24763 33439 24764
tri 33177 24762 33178 24763 ne
rect 33178 24762 33439 24763
tri 33178 24761 33179 24762 ne
rect 33179 24761 33439 24762
tri 33179 24760 33180 24761 ne
rect 33180 24760 33439 24761
tri 33180 24759 33181 24760 ne
rect 33181 24759 33318 24760
tri 33181 24758 33182 24759 ne
rect 33182 24758 33318 24759
tri 33182 24757 33183 24758 ne
rect 33183 24757 33318 24758
tri 33183 24756 33184 24757 ne
rect 33184 24756 33318 24757
tri 33184 24755 33185 24756 ne
rect 33185 24755 33318 24756
tri 33185 24754 33186 24755 ne
rect 33186 24754 33318 24755
tri 33186 24753 33187 24754 ne
rect 33187 24753 33318 24754
tri 33187 24752 33188 24753 ne
rect 33188 24752 33318 24753
tri 33188 24751 33189 24752 ne
rect 33189 24751 33318 24752
tri 33189 24750 33190 24751 ne
rect 33190 24750 33318 24751
tri 33190 24749 33191 24750 ne
rect 33191 24749 33318 24750
tri 33191 24748 33192 24749 ne
rect 33192 24748 33318 24749
tri 33192 24747 33193 24748 ne
rect 33193 24747 33318 24748
tri 33193 24746 33194 24747 ne
rect 33194 24746 33318 24747
tri 33194 24745 33195 24746 ne
rect 33195 24745 33318 24746
tri 33195 24744 33196 24745 ne
rect 33196 24744 33318 24745
tri 33196 24743 33197 24744 ne
rect 33197 24743 33318 24744
tri 33197 24742 33198 24743 ne
rect 33198 24742 33318 24743
tri 33198 24741 33199 24742 ne
rect 33199 24741 33318 24742
tri 33199 24740 33200 24741 ne
rect 33200 24740 33318 24741
tri 33200 24739 33201 24740 ne
rect 33201 24739 33318 24740
tri 33201 24738 33202 24739 ne
rect 33202 24738 33318 24739
tri 33202 24737 33203 24738 ne
rect 33203 24737 33318 24738
tri 33203 24736 33204 24737 ne
rect 33204 24736 33318 24737
tri 33204 24735 33205 24736 ne
rect 33205 24735 33318 24736
tri 33205 24734 33206 24735 ne
rect 33206 24734 33318 24735
tri 33206 24733 33207 24734 ne
rect 33207 24733 33318 24734
tri 33207 24732 33208 24733 ne
rect 33208 24732 33318 24733
tri 33208 24731 33209 24732 ne
rect 33209 24731 33318 24732
tri 33209 24730 33210 24731 ne
rect 33210 24730 33318 24731
tri 33210 24729 33211 24730 ne
rect 33211 24729 33318 24730
tri 33211 24728 33212 24729 ne
rect 33212 24728 33318 24729
tri 33212 24727 33213 24728 ne
rect 33213 24727 33318 24728
tri 33213 24726 33214 24727 ne
rect 33214 24726 33318 24727
tri 33214 24725 33215 24726 ne
rect 33215 24725 33318 24726
tri 33215 24724 33216 24725 ne
rect 33216 24724 33318 24725
tri 33216 24723 33217 24724 ne
rect 33217 24723 33318 24724
tri 33217 24722 33218 24723 ne
rect 33218 24722 33318 24723
tri 33218 24721 33219 24722 ne
rect 33219 24721 33318 24722
tri 33219 24720 33220 24721 ne
rect 33220 24720 33318 24721
tri 33220 24719 33221 24720 ne
rect 33221 24719 33318 24720
tri 33221 24718 33222 24719 ne
rect 33222 24718 33318 24719
tri 33222 24717 33223 24718 ne
rect 33223 24717 33318 24718
tri 33223 24716 33224 24717 ne
rect 33224 24716 33318 24717
tri 33224 24715 33225 24716 ne
rect 33225 24715 33318 24716
tri 33225 24714 33226 24715 ne
rect 33226 24714 33318 24715
rect 33364 24732 33439 24760
tri 33439 24732 33484 24777 sw
rect 70802 24772 71000 24830
rect 33364 24714 33484 24732
tri 33226 24713 33227 24714 ne
rect 33227 24713 33484 24714
tri 33227 24712 33228 24713 ne
rect 33228 24712 33484 24713
tri 33228 24711 33229 24712 ne
rect 33229 24711 33484 24712
tri 33229 24710 33230 24711 ne
rect 33230 24710 33484 24711
tri 33230 24709 33231 24710 ne
rect 33231 24709 33484 24710
tri 33231 24708 33232 24709 ne
rect 33232 24708 33484 24709
tri 33232 24707 33233 24708 ne
rect 33233 24707 33484 24708
tri 33233 24706 33234 24707 ne
rect 33234 24706 33484 24707
tri 33234 24705 33235 24706 ne
rect 33235 24705 33484 24706
tri 33235 24704 33236 24705 ne
rect 33236 24704 33484 24705
tri 33236 24703 33237 24704 ne
rect 33237 24703 33484 24704
tri 33237 24702 33238 24703 ne
rect 33238 24702 33484 24703
tri 33238 24701 33239 24702 ne
rect 33239 24701 33484 24702
tri 33239 24700 33240 24701 ne
rect 33240 24700 33484 24701
tri 33240 24699 33241 24700 ne
rect 33241 24699 33484 24700
tri 33241 24698 33242 24699 ne
rect 33242 24698 33484 24699
tri 33242 24697 33243 24698 ne
rect 33243 24697 33484 24698
tri 33243 24696 33244 24697 ne
rect 33244 24696 33484 24697
tri 33244 24695 33245 24696 ne
rect 33245 24695 33484 24696
tri 33245 24694 33246 24695 ne
rect 33246 24694 33484 24695
tri 33246 24693 33247 24694 ne
rect 33247 24693 33484 24694
tri 33247 24692 33248 24693 ne
rect 33248 24692 33484 24693
tri 33248 24691 33249 24692 ne
rect 33249 24691 33484 24692
tri 33249 24690 33250 24691 ne
rect 33250 24690 33484 24691
tri 33250 24689 33251 24690 ne
rect 33251 24689 33484 24690
tri 33484 24689 33527 24732 sw
rect 70802 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
tri 33251 24677 33263 24689 ne
rect 33263 24677 33527 24689
tri 33263 24632 33308 24677 ne
rect 33308 24644 33527 24677
tri 33527 24644 33572 24689 sw
rect 70802 24668 71000 24726
rect 33308 24632 33572 24644
tri 33308 24587 33353 24632 ne
rect 33353 24628 33572 24632
rect 33353 24587 33450 24628
tri 33353 24542 33398 24587 ne
rect 33398 24582 33450 24587
rect 33496 24599 33572 24628
tri 33572 24599 33617 24644 sw
rect 70802 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24582 33617 24599
rect 33398 24554 33617 24582
tri 33617 24554 33662 24599 sw
rect 70802 24564 71000 24622
rect 33398 24548 33662 24554
tri 33662 24548 33668 24554 sw
rect 33398 24542 33668 24548
tri 33398 24541 33399 24542 ne
rect 33399 24541 33668 24542
tri 33399 24540 33400 24541 ne
rect 33400 24540 33668 24541
tri 33400 24539 33401 24540 ne
rect 33401 24539 33668 24540
tri 33401 24538 33402 24539 ne
rect 33402 24538 33668 24539
tri 33402 24537 33403 24538 ne
rect 33403 24537 33668 24538
tri 33403 24536 33404 24537 ne
rect 33404 24536 33668 24537
tri 33404 24535 33405 24536 ne
rect 33405 24535 33668 24536
tri 33405 24534 33406 24535 ne
rect 33406 24534 33668 24535
tri 33406 24533 33407 24534 ne
rect 33407 24533 33668 24534
tri 33407 24532 33408 24533 ne
rect 33408 24532 33668 24533
tri 33408 24531 33409 24532 ne
rect 33409 24531 33668 24532
tri 33409 24530 33410 24531 ne
rect 33410 24530 33668 24531
tri 33410 24529 33411 24530 ne
rect 33411 24529 33668 24530
tri 33411 24528 33412 24529 ne
rect 33412 24528 33668 24529
tri 33412 24527 33413 24528 ne
rect 33413 24527 33668 24528
tri 33413 24526 33414 24527 ne
rect 33414 24526 33668 24527
tri 33414 24525 33415 24526 ne
rect 33415 24525 33668 24526
tri 33415 24524 33416 24525 ne
rect 33416 24524 33668 24525
tri 33416 24523 33417 24524 ne
rect 33417 24523 33668 24524
tri 33417 24522 33418 24523 ne
rect 33418 24522 33668 24523
tri 33418 24521 33419 24522 ne
rect 33419 24521 33668 24522
tri 33419 24520 33420 24521 ne
rect 33420 24520 33668 24521
tri 33420 24519 33421 24520 ne
rect 33421 24519 33668 24520
tri 33421 24518 33422 24519 ne
rect 33422 24518 33668 24519
tri 33422 24517 33423 24518 ne
rect 33423 24517 33668 24518
tri 33423 24516 33424 24517 ne
rect 33424 24516 33668 24517
tri 33424 24515 33425 24516 ne
rect 33425 24515 33668 24516
tri 33425 24514 33426 24515 ne
rect 33426 24514 33668 24515
tri 33426 24513 33427 24514 ne
rect 33427 24513 33668 24514
tri 33427 24512 33428 24513 ne
rect 33428 24512 33668 24513
tri 33428 24511 33429 24512 ne
rect 33429 24511 33668 24512
tri 33429 24510 33430 24511 ne
rect 33430 24510 33668 24511
tri 33430 24509 33431 24510 ne
rect 33431 24509 33668 24510
tri 33431 24508 33432 24509 ne
rect 33432 24508 33668 24509
tri 33432 24507 33433 24508 ne
rect 33433 24507 33668 24508
tri 33433 24506 33434 24507 ne
rect 33434 24506 33668 24507
tri 33434 24505 33435 24506 ne
rect 33435 24505 33668 24506
tri 33435 24504 33436 24505 ne
rect 33436 24504 33668 24505
tri 33436 24503 33437 24504 ne
rect 33437 24503 33668 24504
tri 33668 24503 33713 24548 sw
rect 70802 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33437 24502 33438 24503 ne
rect 33438 24502 33713 24503
tri 33438 24501 33439 24502 ne
rect 33439 24501 33713 24502
tri 33439 24500 33440 24501 ne
rect 33440 24500 33713 24501
tri 33440 24499 33441 24500 ne
rect 33441 24499 33713 24500
tri 33441 24498 33442 24499 ne
rect 33442 24498 33713 24499
tri 33442 24497 33443 24498 ne
rect 33443 24497 33713 24498
tri 33443 24496 33444 24497 ne
rect 33444 24496 33713 24497
tri 33444 24495 33445 24496 ne
rect 33445 24495 33582 24496
tri 33445 24494 33446 24495 ne
rect 33446 24494 33582 24495
tri 33446 24493 33447 24494 ne
rect 33447 24493 33582 24494
tri 33447 24492 33448 24493 ne
rect 33448 24492 33582 24493
tri 33448 24491 33449 24492 ne
rect 33449 24491 33582 24492
tri 33449 24490 33450 24491 ne
rect 33450 24490 33582 24491
tri 33450 24489 33451 24490 ne
rect 33451 24489 33582 24490
tri 33451 24488 33452 24489 ne
rect 33452 24488 33582 24489
tri 33452 24487 33453 24488 ne
rect 33453 24487 33582 24488
tri 33453 24486 33454 24487 ne
rect 33454 24486 33582 24487
tri 33454 24485 33455 24486 ne
rect 33455 24485 33582 24486
tri 33455 24484 33456 24485 ne
rect 33456 24484 33582 24485
tri 33456 24483 33457 24484 ne
rect 33457 24483 33582 24484
tri 33457 24482 33458 24483 ne
rect 33458 24482 33582 24483
tri 33458 24481 33459 24482 ne
rect 33459 24481 33582 24482
tri 33459 24480 33460 24481 ne
rect 33460 24480 33582 24481
tri 33460 24479 33461 24480 ne
rect 33461 24479 33582 24480
tri 33461 24478 33462 24479 ne
rect 33462 24478 33582 24479
tri 33462 24477 33463 24478 ne
rect 33463 24477 33582 24478
tri 33463 24476 33464 24477 ne
rect 33464 24476 33582 24477
tri 33464 24475 33465 24476 ne
rect 33465 24475 33582 24476
tri 33465 24474 33466 24475 ne
rect 33466 24474 33582 24475
tri 33466 24473 33467 24474 ne
rect 33467 24473 33582 24474
tri 33467 24472 33468 24473 ne
rect 33468 24472 33582 24473
tri 33468 24471 33469 24472 ne
rect 33469 24471 33582 24472
tri 33469 24470 33470 24471 ne
rect 33470 24470 33582 24471
tri 33470 24469 33471 24470 ne
rect 33471 24469 33582 24470
tri 33471 24468 33472 24469 ne
rect 33472 24468 33582 24469
tri 33472 24467 33473 24468 ne
rect 33473 24467 33582 24468
tri 33473 24466 33474 24467 ne
rect 33474 24466 33582 24467
tri 33474 24465 33475 24466 ne
rect 33475 24465 33582 24466
tri 33475 24464 33476 24465 ne
rect 33476 24464 33582 24465
tri 33476 24463 33477 24464 ne
rect 33477 24463 33582 24464
tri 33477 24462 33478 24463 ne
rect 33478 24462 33582 24463
tri 33478 24461 33479 24462 ne
rect 33479 24461 33582 24462
tri 33479 24460 33480 24461 ne
rect 33480 24460 33582 24461
tri 33480 24459 33481 24460 ne
rect 33481 24459 33582 24460
tri 33481 24458 33482 24459 ne
rect 33482 24458 33582 24459
tri 33482 24457 33483 24458 ne
rect 33483 24457 33582 24458
tri 33483 24456 33484 24457 ne
rect 33484 24456 33582 24457
tri 33484 24455 33485 24456 ne
rect 33485 24455 33582 24456
tri 33485 24454 33486 24455 ne
rect 33486 24454 33582 24455
tri 33486 24453 33487 24454 ne
rect 33487 24453 33582 24454
tri 33487 24452 33488 24453 ne
rect 33488 24452 33582 24453
tri 33488 24451 33489 24452 ne
rect 33489 24451 33582 24452
tri 33489 24450 33490 24451 ne
rect 33490 24450 33582 24451
rect 33628 24458 33713 24496
tri 33713 24458 33758 24503 sw
rect 70802 24460 71000 24518
rect 33628 24450 33758 24458
tri 33490 24449 33491 24450 ne
rect 33491 24449 33758 24450
tri 33491 24448 33492 24449 ne
rect 33492 24448 33758 24449
tri 33492 24447 33493 24448 ne
rect 33493 24447 33758 24448
tri 33493 24446 33494 24447 ne
rect 33494 24446 33758 24447
tri 33494 24445 33495 24446 ne
rect 33495 24445 33758 24446
tri 33495 24444 33496 24445 ne
rect 33496 24444 33758 24445
tri 33496 24443 33497 24444 ne
rect 33497 24443 33758 24444
tri 33497 24442 33498 24443 ne
rect 33498 24442 33758 24443
tri 33498 24441 33499 24442 ne
rect 33499 24441 33758 24442
tri 33499 24440 33500 24441 ne
rect 33500 24440 33758 24441
tri 33500 24439 33501 24440 ne
rect 33501 24439 33758 24440
tri 33501 24438 33502 24439 ne
rect 33502 24438 33758 24439
tri 33502 24437 33503 24438 ne
rect 33503 24437 33758 24438
tri 33503 24436 33504 24437 ne
rect 33504 24436 33758 24437
tri 33504 24435 33505 24436 ne
rect 33505 24435 33758 24436
tri 33505 24434 33506 24435 ne
rect 33506 24434 33758 24435
tri 33506 24433 33507 24434 ne
rect 33507 24433 33758 24434
tri 33507 24432 33508 24433 ne
rect 33508 24432 33758 24433
tri 33508 24431 33509 24432 ne
rect 33509 24431 33758 24432
tri 33509 24430 33510 24431 ne
rect 33510 24430 33758 24431
tri 33510 24429 33511 24430 ne
rect 33511 24429 33758 24430
tri 33511 24428 33512 24429 ne
rect 33512 24428 33758 24429
tri 33512 24427 33513 24428 ne
rect 33513 24427 33758 24428
tri 33513 24426 33514 24427 ne
rect 33514 24426 33758 24427
tri 33514 24425 33515 24426 ne
rect 33515 24425 33758 24426
tri 33515 24424 33516 24425 ne
rect 33516 24424 33758 24425
tri 33516 24423 33517 24424 ne
rect 33517 24423 33758 24424
tri 33517 24422 33518 24423 ne
rect 33518 24422 33758 24423
tri 33518 24421 33519 24422 ne
rect 33519 24421 33758 24422
tri 33519 24420 33520 24421 ne
rect 33520 24420 33758 24421
tri 33520 24419 33521 24420 ne
rect 33521 24419 33758 24420
tri 33521 24418 33522 24419 ne
rect 33522 24418 33758 24419
tri 33522 24417 33523 24418 ne
rect 33523 24417 33758 24418
tri 33523 24416 33524 24417 ne
rect 33524 24416 33758 24417
tri 33524 24415 33525 24416 ne
rect 33525 24415 33758 24416
tri 33525 24414 33526 24415 ne
rect 33526 24414 33758 24415
tri 33526 24413 33527 24414 ne
rect 33527 24413 33758 24414
tri 33758 24413 33803 24458 sw
rect 70802 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33527 24411 33529 24413 ne
rect 33529 24411 33803 24413
tri 33803 24411 33805 24413 sw
tri 33529 24366 33574 24411 ne
rect 33574 24366 33805 24411
tri 33805 24366 33850 24411 sw
tri 33574 24357 33583 24366 ne
rect 33583 24364 33850 24366
rect 33583 24357 33714 24364
tri 33583 24312 33628 24357 ne
rect 33628 24318 33714 24357
rect 33760 24321 33850 24364
tri 33850 24321 33895 24366 sw
rect 70802 24356 71000 24414
rect 33760 24318 33895 24321
rect 33628 24312 33895 24318
tri 33628 24267 33673 24312 ne
rect 33673 24276 33895 24312
tri 33895 24276 33940 24321 sw
rect 70802 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 33673 24272 33940 24276
tri 33940 24272 33944 24276 sw
rect 33673 24267 33944 24272
tri 33673 24266 33674 24267 ne
rect 33674 24266 33944 24267
tri 33674 24265 33675 24266 ne
rect 33675 24265 33944 24266
tri 33675 24264 33676 24265 ne
rect 33676 24264 33944 24265
tri 33676 24263 33677 24264 ne
rect 33677 24263 33944 24264
tri 33677 24262 33678 24263 ne
rect 33678 24262 33944 24263
tri 33678 24261 33679 24262 ne
rect 33679 24261 33944 24262
tri 33679 24260 33680 24261 ne
rect 33680 24260 33944 24261
tri 33680 24259 33681 24260 ne
rect 33681 24259 33944 24260
tri 33681 24258 33682 24259 ne
rect 33682 24258 33944 24259
tri 33682 24257 33683 24258 ne
rect 33683 24257 33944 24258
tri 33683 24256 33684 24257 ne
rect 33684 24256 33944 24257
tri 33684 24255 33685 24256 ne
rect 33685 24255 33944 24256
tri 33685 24254 33686 24255 ne
rect 33686 24254 33944 24255
tri 33686 24253 33687 24254 ne
rect 33687 24253 33944 24254
tri 33687 24252 33688 24253 ne
rect 33688 24252 33944 24253
tri 33688 24251 33689 24252 ne
rect 33689 24251 33944 24252
tri 33689 24250 33690 24251 ne
rect 33690 24250 33944 24251
tri 33690 24249 33691 24250 ne
rect 33691 24249 33944 24250
tri 33691 24248 33692 24249 ne
rect 33692 24248 33944 24249
tri 33692 24247 33693 24248 ne
rect 33693 24247 33944 24248
tri 33693 24246 33694 24247 ne
rect 33694 24246 33944 24247
tri 33694 24245 33695 24246 ne
rect 33695 24245 33944 24246
tri 33695 24244 33696 24245 ne
rect 33696 24244 33944 24245
tri 33696 24243 33697 24244 ne
rect 33697 24243 33944 24244
tri 33697 24242 33698 24243 ne
rect 33698 24242 33944 24243
tri 33698 24241 33699 24242 ne
rect 33699 24241 33944 24242
tri 33699 24240 33700 24241 ne
rect 33700 24240 33944 24241
tri 33700 24239 33701 24240 ne
rect 33701 24239 33944 24240
tri 33701 24238 33702 24239 ne
rect 33702 24238 33944 24239
tri 33702 24237 33703 24238 ne
rect 33703 24237 33944 24238
tri 33703 24236 33704 24237 ne
rect 33704 24236 33944 24237
tri 33704 24235 33705 24236 ne
rect 33705 24235 33944 24236
tri 33705 24234 33706 24235 ne
rect 33706 24234 33944 24235
tri 33706 24233 33707 24234 ne
rect 33707 24233 33944 24234
tri 33707 24232 33708 24233 ne
rect 33708 24232 33944 24233
tri 33708 24231 33709 24232 ne
rect 33709 24231 33846 24232
tri 33709 24230 33710 24231 ne
rect 33710 24230 33846 24231
tri 33710 24229 33711 24230 ne
rect 33711 24229 33846 24230
tri 33711 24228 33712 24229 ne
rect 33712 24228 33846 24229
tri 33712 24227 33713 24228 ne
rect 33713 24227 33846 24228
tri 33713 24226 33714 24227 ne
rect 33714 24226 33846 24227
tri 33714 24225 33715 24226 ne
rect 33715 24225 33846 24226
tri 33715 24224 33716 24225 ne
rect 33716 24224 33846 24225
tri 33716 24223 33717 24224 ne
rect 33717 24223 33846 24224
tri 33717 24222 33718 24223 ne
rect 33718 24222 33846 24223
tri 33718 24221 33719 24222 ne
rect 33719 24221 33846 24222
tri 33719 24220 33720 24221 ne
rect 33720 24220 33846 24221
tri 33720 24219 33721 24220 ne
rect 33721 24219 33846 24220
tri 33721 24218 33722 24219 ne
rect 33722 24218 33846 24219
tri 33722 24217 33723 24218 ne
rect 33723 24217 33846 24218
tri 33723 24216 33724 24217 ne
rect 33724 24216 33846 24217
tri 33724 24215 33725 24216 ne
rect 33725 24215 33846 24216
tri 33725 24214 33726 24215 ne
rect 33726 24214 33846 24215
tri 33726 24213 33727 24214 ne
rect 33727 24213 33846 24214
tri 33727 24212 33728 24213 ne
rect 33728 24212 33846 24213
tri 33728 24211 33729 24212 ne
rect 33729 24211 33846 24212
tri 33729 24210 33730 24211 ne
rect 33730 24210 33846 24211
tri 33730 24209 33731 24210 ne
rect 33731 24209 33846 24210
tri 33731 24208 33732 24209 ne
rect 33732 24208 33846 24209
tri 33732 24207 33733 24208 ne
rect 33733 24207 33846 24208
tri 33733 24206 33734 24207 ne
rect 33734 24206 33846 24207
tri 33734 24205 33735 24206 ne
rect 33735 24205 33846 24206
tri 33735 24204 33736 24205 ne
rect 33736 24204 33846 24205
tri 33736 24203 33737 24204 ne
rect 33737 24203 33846 24204
tri 33737 24202 33738 24203 ne
rect 33738 24202 33846 24203
tri 33738 24201 33739 24202 ne
rect 33739 24201 33846 24202
tri 33739 24200 33740 24201 ne
rect 33740 24200 33846 24201
tri 33740 24199 33741 24200 ne
rect 33741 24199 33846 24200
tri 33741 24198 33742 24199 ne
rect 33742 24198 33846 24199
tri 33742 24197 33743 24198 ne
rect 33743 24197 33846 24198
tri 33743 24196 33744 24197 ne
rect 33744 24196 33846 24197
tri 33744 24195 33745 24196 ne
rect 33745 24195 33846 24196
tri 33745 24194 33746 24195 ne
rect 33746 24194 33846 24195
tri 33746 24193 33747 24194 ne
rect 33747 24193 33846 24194
tri 33747 24192 33748 24193 ne
rect 33748 24192 33846 24193
tri 33748 24191 33749 24192 ne
rect 33749 24191 33846 24192
tri 33749 24190 33750 24191 ne
rect 33750 24190 33846 24191
tri 33750 24189 33751 24190 ne
rect 33751 24189 33846 24190
tri 33751 24188 33752 24189 ne
rect 33752 24188 33846 24189
tri 33752 24187 33753 24188 ne
rect 33753 24187 33846 24188
tri 33753 24186 33754 24187 ne
rect 33754 24186 33846 24187
rect 33892 24227 33944 24232
tri 33944 24227 33989 24272 sw
rect 70802 24252 71000 24310
rect 33892 24186 33989 24227
tri 33754 24185 33755 24186 ne
rect 33755 24185 33989 24186
tri 33755 24184 33756 24185 ne
rect 33756 24184 33989 24185
tri 33756 24183 33757 24184 ne
rect 33757 24183 33989 24184
tri 33757 24182 33758 24183 ne
rect 33758 24182 33989 24183
tri 33989 24182 34034 24227 sw
rect 70802 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
tri 33758 24181 33759 24182 ne
rect 33759 24181 34034 24182
tri 33759 24180 33760 24181 ne
rect 33760 24180 34034 24181
tri 33760 24179 33761 24180 ne
rect 33761 24179 34034 24180
tri 33761 24178 33762 24179 ne
rect 33762 24178 34034 24179
tri 33762 24177 33763 24178 ne
rect 33763 24177 34034 24178
tri 33763 24176 33764 24177 ne
rect 33764 24176 34034 24177
tri 33764 24175 33765 24176 ne
rect 33765 24175 34034 24176
tri 33765 24174 33766 24175 ne
rect 33766 24174 34034 24175
tri 33766 24173 33767 24174 ne
rect 33767 24173 34034 24174
tri 33767 24172 33768 24173 ne
rect 33768 24172 34034 24173
tri 33768 24171 33769 24172 ne
rect 33769 24171 34034 24172
tri 33769 24170 33770 24171 ne
rect 33770 24170 34034 24171
tri 33770 24169 33771 24170 ne
rect 33771 24169 34034 24170
tri 33771 24168 33772 24169 ne
rect 33772 24168 34034 24169
tri 33772 24167 33773 24168 ne
rect 33773 24167 34034 24168
tri 33773 24166 33774 24167 ne
rect 33774 24166 34034 24167
tri 33774 24165 33775 24166 ne
rect 33775 24165 34034 24166
tri 33775 24164 33776 24165 ne
rect 33776 24164 34034 24165
tri 33776 24163 33777 24164 ne
rect 33777 24163 34034 24164
tri 33777 24162 33778 24163 ne
rect 33778 24162 34034 24163
tri 33778 24161 33779 24162 ne
rect 33779 24161 34034 24162
tri 33779 24160 33780 24161 ne
rect 33780 24160 34034 24161
tri 33780 24159 33781 24160 ne
rect 33781 24159 34034 24160
tri 33781 24158 33782 24159 ne
rect 33782 24158 34034 24159
tri 33782 24157 33783 24158 ne
rect 33783 24157 34034 24158
tri 33783 24156 33784 24157 ne
rect 33784 24156 34034 24157
tri 33784 24155 33785 24156 ne
rect 33785 24155 34034 24156
tri 33785 24154 33786 24155 ne
rect 33786 24154 34034 24155
tri 33786 24153 33787 24154 ne
rect 33787 24153 34034 24154
tri 33787 24152 33788 24153 ne
rect 33788 24152 34034 24153
tri 33788 24151 33789 24152 ne
rect 33789 24151 34034 24152
tri 33789 24150 33790 24151 ne
rect 33790 24150 34034 24151
tri 33790 24149 33791 24150 ne
rect 33791 24149 34034 24150
tri 33791 24148 33792 24149 ne
rect 33792 24148 34034 24149
tri 33792 24147 33793 24148 ne
rect 33793 24147 34034 24148
tri 33793 24146 33794 24147 ne
rect 33794 24146 34034 24147
tri 33794 24145 33795 24146 ne
rect 33795 24145 34034 24146
tri 33795 24144 33796 24145 ne
rect 33796 24144 34034 24145
tri 33796 24143 33797 24144 ne
rect 33797 24143 34034 24144
tri 33797 24142 33798 24143 ne
rect 33798 24142 34034 24143
tri 33798 24141 33799 24142 ne
rect 33799 24141 34034 24142
tri 33799 24140 33800 24141 ne
rect 33800 24140 34034 24141
tri 33800 24139 33801 24140 ne
rect 33801 24139 34034 24140
tri 33801 24138 33802 24139 ne
rect 33802 24138 34034 24139
tri 33802 24137 33803 24138 ne
rect 33803 24137 34034 24138
tri 34034 24137 34079 24182 sw
rect 70802 24148 71000 24206
tri 33803 24092 33848 24137 ne
rect 33848 24100 34079 24137
rect 33848 24092 33978 24100
tri 33848 24090 33850 24092 ne
rect 33850 24090 33978 24092
tri 33850 24047 33893 24090 ne
rect 33893 24054 33978 24090
rect 34024 24092 34079 24100
tri 34079 24092 34124 24137 sw
rect 70802 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 34024 24090 34124 24092
tri 34124 24090 34126 24092 sw
rect 34024 24054 34126 24090
rect 33893 24047 34126 24054
tri 33893 24045 33895 24047 ne
rect 33895 24045 34126 24047
tri 34126 24045 34171 24090 sw
tri 33895 24000 33940 24045 ne
rect 33940 24000 34171 24045
tri 34171 24000 34216 24045 sw
rect 70802 24044 71000 24102
tri 33940 23993 33947 24000 ne
rect 33947 23993 34216 24000
tri 33947 23992 33948 23993 ne
rect 33948 23992 34216 23993
tri 33948 23991 33949 23992 ne
rect 33949 23991 34216 23992
tri 33949 23990 33950 23991 ne
rect 33950 23990 34216 23991
tri 33950 23989 33951 23990 ne
rect 33951 23989 34216 23990
tri 33951 23988 33952 23989 ne
rect 33952 23988 34216 23989
tri 33952 23987 33953 23988 ne
rect 33953 23987 34216 23988
tri 33953 23986 33954 23987 ne
rect 33954 23986 34216 23987
tri 33954 23985 33955 23986 ne
rect 33955 23985 34216 23986
tri 33955 23984 33956 23985 ne
rect 33956 23984 34216 23985
tri 33956 23983 33957 23984 ne
rect 33957 23983 34216 23984
tri 33957 23982 33958 23983 ne
rect 33958 23982 34216 23983
tri 33958 23981 33959 23982 ne
rect 33959 23981 34216 23982
tri 33959 23980 33960 23981 ne
rect 33960 23980 34216 23981
tri 33960 23979 33961 23980 ne
rect 33961 23979 34216 23980
tri 33961 23978 33962 23979 ne
rect 33962 23978 34216 23979
tri 33962 23977 33963 23978 ne
rect 33963 23977 34216 23978
tri 33963 23976 33964 23977 ne
rect 33964 23976 34216 23977
tri 33964 23975 33965 23976 ne
rect 33965 23975 34216 23976
tri 33965 23974 33966 23975 ne
rect 33966 23974 34216 23975
tri 33966 23973 33967 23974 ne
rect 33967 23973 34216 23974
tri 33967 23972 33968 23973 ne
rect 33968 23972 34216 23973
tri 33968 23971 33969 23972 ne
rect 33969 23971 34216 23972
tri 33969 23970 33970 23971 ne
rect 33970 23970 34216 23971
tri 33970 23969 33971 23970 ne
rect 33971 23969 34216 23970
tri 33971 23968 33972 23969 ne
rect 33972 23968 34216 23969
tri 33972 23967 33973 23968 ne
rect 33973 23967 34110 23968
tri 33973 23966 33974 23967 ne
rect 33974 23966 34110 23967
tri 33974 23965 33975 23966 ne
rect 33975 23965 34110 23966
tri 33975 23964 33976 23965 ne
rect 33976 23964 34110 23965
tri 33976 23963 33977 23964 ne
rect 33977 23963 34110 23964
tri 33977 23962 33978 23963 ne
rect 33978 23962 34110 23963
tri 33978 23961 33979 23962 ne
rect 33979 23961 34110 23962
tri 33979 23960 33980 23961 ne
rect 33980 23960 34110 23961
tri 33980 23959 33981 23960 ne
rect 33981 23959 34110 23960
tri 33981 23958 33982 23959 ne
rect 33982 23958 34110 23959
tri 33982 23957 33983 23958 ne
rect 33983 23957 34110 23958
tri 33983 23956 33984 23957 ne
rect 33984 23956 34110 23957
tri 33984 23955 33985 23956 ne
rect 33985 23955 34110 23956
tri 33985 23954 33986 23955 ne
rect 33986 23954 34110 23955
tri 33986 23953 33987 23954 ne
rect 33987 23953 34110 23954
tri 33987 23952 33988 23953 ne
rect 33988 23952 34110 23953
tri 33988 23951 33989 23952 ne
rect 33989 23951 34110 23952
tri 33989 23950 33990 23951 ne
rect 33990 23950 34110 23951
tri 33990 23949 33991 23950 ne
rect 33991 23949 34110 23950
tri 33991 23948 33992 23949 ne
rect 33992 23948 34110 23949
tri 33992 23947 33993 23948 ne
rect 33993 23947 34110 23948
tri 33993 23946 33994 23947 ne
rect 33994 23946 34110 23947
tri 33994 23945 33995 23946 ne
rect 33995 23945 34110 23946
tri 33995 23944 33996 23945 ne
rect 33996 23944 34110 23945
tri 33996 23943 33997 23944 ne
rect 33997 23943 34110 23944
tri 33997 23942 33998 23943 ne
rect 33998 23942 34110 23943
tri 33998 23941 33999 23942 ne
rect 33999 23941 34110 23942
tri 33999 23940 34000 23941 ne
rect 34000 23940 34110 23941
tri 34000 23939 34001 23940 ne
rect 34001 23939 34110 23940
tri 34001 23938 34002 23939 ne
rect 34002 23938 34110 23939
tri 34002 23937 34003 23938 ne
rect 34003 23937 34110 23938
tri 34003 23936 34004 23937 ne
rect 34004 23936 34110 23937
tri 34004 23935 34005 23936 ne
rect 34005 23935 34110 23936
tri 34005 23934 34006 23935 ne
rect 34006 23934 34110 23935
tri 34006 23933 34007 23934 ne
rect 34007 23933 34110 23934
tri 34007 23932 34008 23933 ne
rect 34008 23932 34110 23933
tri 34008 23931 34009 23932 ne
rect 34009 23931 34110 23932
tri 34009 23930 34010 23931 ne
rect 34010 23930 34110 23931
tri 34010 23929 34011 23930 ne
rect 34011 23929 34110 23930
tri 34011 23928 34012 23929 ne
rect 34012 23928 34110 23929
tri 34012 23927 34013 23928 ne
rect 34013 23927 34110 23928
tri 34013 23926 34014 23927 ne
rect 34014 23926 34110 23927
tri 34014 23925 34015 23926 ne
rect 34015 23925 34110 23926
tri 34015 23924 34016 23925 ne
rect 34016 23924 34110 23925
tri 34016 23923 34017 23924 ne
rect 34017 23923 34110 23924
tri 34017 23922 34018 23923 ne
rect 34018 23922 34110 23923
rect 34156 23955 34216 23968
tri 34216 23955 34261 24000 sw
rect 70802 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
rect 34156 23951 34261 23955
tri 34261 23951 34265 23955 sw
rect 34156 23922 34265 23951
tri 34018 23921 34019 23922 ne
rect 34019 23921 34265 23922
tri 34019 23920 34020 23921 ne
rect 34020 23920 34265 23921
tri 34020 23919 34021 23920 ne
rect 34021 23919 34265 23920
tri 34021 23918 34022 23919 ne
rect 34022 23918 34265 23919
tri 34022 23917 34023 23918 ne
rect 34023 23917 34265 23918
tri 34023 23916 34024 23917 ne
rect 34024 23916 34265 23917
tri 34024 23915 34025 23916 ne
rect 34025 23915 34265 23916
tri 34025 23914 34026 23915 ne
rect 34026 23914 34265 23915
tri 34026 23913 34027 23914 ne
rect 34027 23913 34265 23914
tri 34027 23912 34028 23913 ne
rect 34028 23912 34265 23913
tri 34028 23911 34029 23912 ne
rect 34029 23911 34265 23912
tri 34029 23910 34030 23911 ne
rect 34030 23910 34265 23911
tri 34030 23909 34031 23910 ne
rect 34031 23909 34265 23910
tri 34031 23908 34032 23909 ne
rect 34032 23908 34265 23909
tri 34032 23907 34033 23908 ne
rect 34033 23907 34265 23908
tri 34033 23906 34034 23907 ne
rect 34034 23906 34265 23907
tri 34265 23906 34310 23951 sw
rect 70802 23940 71000 23998
tri 34034 23905 34035 23906 ne
rect 34035 23905 34310 23906
tri 34035 23904 34036 23905 ne
rect 34036 23904 34310 23905
tri 34036 23903 34037 23904 ne
rect 34037 23903 34310 23904
tri 34037 23902 34038 23903 ne
rect 34038 23902 34310 23903
tri 34038 23901 34039 23902 ne
rect 34039 23901 34310 23902
tri 34039 23900 34040 23901 ne
rect 34040 23900 34310 23901
tri 34040 23899 34041 23900 ne
rect 34041 23899 34310 23900
tri 34041 23898 34042 23899 ne
rect 34042 23898 34310 23899
tri 34042 23897 34043 23898 ne
rect 34043 23897 34310 23898
tri 34043 23896 34044 23897 ne
rect 34044 23896 34310 23897
tri 34044 23895 34045 23896 ne
rect 34045 23895 34310 23896
tri 34045 23894 34046 23895 ne
rect 34046 23894 34310 23895
tri 34046 23893 34047 23894 ne
rect 34047 23893 34310 23894
tri 34047 23892 34048 23893 ne
rect 34048 23892 34310 23893
tri 34048 23891 34049 23892 ne
rect 34049 23891 34310 23892
tri 34049 23890 34050 23891 ne
rect 34050 23890 34310 23891
tri 34050 23889 34051 23890 ne
rect 34051 23889 34310 23890
tri 34051 23888 34052 23889 ne
rect 34052 23888 34310 23889
tri 34052 23887 34053 23888 ne
rect 34053 23887 34310 23888
tri 34053 23886 34054 23887 ne
rect 34054 23886 34310 23887
tri 34054 23885 34055 23886 ne
rect 34055 23885 34310 23886
tri 34055 23884 34056 23885 ne
rect 34056 23884 34310 23885
tri 34056 23883 34057 23884 ne
rect 34057 23883 34310 23884
tri 34057 23882 34058 23883 ne
rect 34058 23882 34310 23883
tri 34058 23881 34059 23882 ne
rect 34059 23881 34310 23882
tri 34059 23880 34060 23881 ne
rect 34060 23880 34310 23881
tri 34060 23879 34061 23880 ne
rect 34061 23879 34310 23880
tri 34061 23878 34062 23879 ne
rect 34062 23878 34310 23879
tri 34062 23877 34063 23878 ne
rect 34063 23877 34310 23878
tri 34063 23876 34064 23877 ne
rect 34064 23876 34310 23877
tri 34064 23875 34065 23876 ne
rect 34065 23875 34310 23876
tri 34065 23874 34066 23875 ne
rect 34066 23874 34310 23875
tri 34066 23873 34067 23874 ne
rect 34067 23873 34310 23874
tri 34067 23872 34068 23873 ne
rect 34068 23872 34310 23873
tri 34068 23871 34069 23872 ne
rect 34069 23871 34310 23872
tri 34069 23870 34070 23871 ne
rect 34070 23870 34310 23871
tri 34070 23869 34071 23870 ne
rect 34071 23869 34310 23870
tri 34071 23868 34072 23869 ne
rect 34072 23868 34310 23869
tri 34072 23867 34073 23868 ne
rect 34073 23867 34310 23868
tri 34073 23866 34074 23867 ne
rect 34074 23866 34310 23867
tri 34074 23865 34075 23866 ne
rect 34075 23865 34310 23866
tri 34075 23864 34076 23865 ne
rect 34076 23864 34310 23865
tri 34076 23863 34077 23864 ne
rect 34077 23863 34310 23864
tri 34077 23862 34078 23863 ne
rect 34078 23862 34310 23863
tri 34078 23861 34079 23862 ne
rect 34079 23861 34310 23862
tri 34310 23861 34355 23906 sw
rect 70802 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34079 23816 34124 23861 ne
rect 34124 23836 34355 23861
rect 34124 23816 34242 23836
tri 34124 23771 34169 23816 ne
rect 34169 23790 34242 23816
rect 34288 23816 34355 23836
tri 34355 23816 34400 23861 sw
rect 70802 23836 71000 23894
rect 34288 23790 34400 23816
rect 34169 23771 34400 23790
tri 34400 23771 34445 23816 sw
rect 70802 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
tri 34169 23726 34214 23771 ne
rect 34214 23769 34445 23771
tri 34445 23769 34447 23771 sw
rect 34214 23726 34447 23769
tri 34214 23724 34216 23726 ne
rect 34216 23724 34447 23726
tri 34447 23724 34492 23769 sw
rect 70802 23732 71000 23790
tri 34216 23718 34222 23724 ne
rect 34222 23718 34492 23724
tri 34222 23717 34223 23718 ne
rect 34223 23717 34492 23718
tri 34223 23716 34224 23717 ne
rect 34224 23716 34492 23717
tri 34224 23715 34225 23716 ne
rect 34225 23715 34492 23716
tri 34225 23714 34226 23715 ne
rect 34226 23714 34492 23715
tri 34226 23713 34227 23714 ne
rect 34227 23713 34492 23714
tri 34227 23712 34228 23713 ne
rect 34228 23712 34492 23713
tri 34228 23711 34229 23712 ne
rect 34229 23711 34492 23712
tri 34229 23710 34230 23711 ne
rect 34230 23710 34492 23711
tri 34230 23709 34231 23710 ne
rect 34231 23709 34492 23710
tri 34231 23708 34232 23709 ne
rect 34232 23708 34492 23709
tri 34232 23707 34233 23708 ne
rect 34233 23707 34492 23708
tri 34233 23706 34234 23707 ne
rect 34234 23706 34492 23707
tri 34234 23705 34235 23706 ne
rect 34235 23705 34492 23706
tri 34235 23704 34236 23705 ne
rect 34236 23704 34492 23705
tri 34236 23703 34237 23704 ne
rect 34237 23703 34374 23704
tri 34237 23702 34238 23703 ne
rect 34238 23702 34374 23703
tri 34238 23701 34239 23702 ne
rect 34239 23701 34374 23702
tri 34239 23700 34240 23701 ne
rect 34240 23700 34374 23701
tri 34240 23699 34241 23700 ne
rect 34241 23699 34374 23700
tri 34241 23698 34242 23699 ne
rect 34242 23698 34374 23699
tri 34242 23697 34243 23698 ne
rect 34243 23697 34374 23698
tri 34243 23696 34244 23697 ne
rect 34244 23696 34374 23697
tri 34244 23695 34245 23696 ne
rect 34245 23695 34374 23696
tri 34245 23694 34246 23695 ne
rect 34246 23694 34374 23695
tri 34246 23693 34247 23694 ne
rect 34247 23693 34374 23694
tri 34247 23692 34248 23693 ne
rect 34248 23692 34374 23693
tri 34248 23691 34249 23692 ne
rect 34249 23691 34374 23692
tri 34249 23690 34250 23691 ne
rect 34250 23690 34374 23691
tri 34250 23689 34251 23690 ne
rect 34251 23689 34374 23690
tri 34251 23688 34252 23689 ne
rect 34252 23688 34374 23689
tri 34252 23687 34253 23688 ne
rect 34253 23687 34374 23688
tri 34253 23686 34254 23687 ne
rect 34254 23686 34374 23687
tri 34254 23685 34255 23686 ne
rect 34255 23685 34374 23686
tri 34255 23684 34256 23685 ne
rect 34256 23684 34374 23685
tri 34256 23683 34257 23684 ne
rect 34257 23683 34374 23684
tri 34257 23682 34258 23683 ne
rect 34258 23682 34374 23683
tri 34258 23681 34259 23682 ne
rect 34259 23681 34374 23682
tri 34259 23680 34260 23681 ne
rect 34260 23680 34374 23681
tri 34260 23679 34261 23680 ne
rect 34261 23679 34374 23680
tri 34261 23678 34262 23679 ne
rect 34262 23678 34374 23679
tri 34262 23677 34263 23678 ne
rect 34263 23677 34374 23678
tri 34263 23676 34264 23677 ne
rect 34264 23676 34374 23677
tri 34264 23675 34265 23676 ne
rect 34265 23675 34374 23676
tri 34265 23674 34266 23675 ne
rect 34266 23674 34374 23675
tri 34266 23673 34267 23674 ne
rect 34267 23673 34374 23674
tri 34267 23672 34268 23673 ne
rect 34268 23672 34374 23673
tri 34268 23671 34269 23672 ne
rect 34269 23671 34374 23672
tri 34269 23670 34270 23671 ne
rect 34270 23670 34374 23671
tri 34270 23669 34271 23670 ne
rect 34271 23669 34374 23670
tri 34271 23668 34272 23669 ne
rect 34272 23668 34374 23669
tri 34272 23667 34273 23668 ne
rect 34273 23667 34374 23668
tri 34273 23666 34274 23667 ne
rect 34274 23666 34374 23667
tri 34274 23665 34275 23666 ne
rect 34275 23665 34374 23666
tri 34275 23664 34276 23665 ne
rect 34276 23664 34374 23665
tri 34276 23663 34277 23664 ne
rect 34277 23663 34374 23664
tri 34277 23662 34278 23663 ne
rect 34278 23662 34374 23663
tri 34278 23661 34279 23662 ne
rect 34279 23661 34374 23662
tri 34279 23660 34280 23661 ne
rect 34280 23660 34374 23661
tri 34280 23659 34281 23660 ne
rect 34281 23659 34374 23660
tri 34281 23658 34282 23659 ne
rect 34282 23658 34374 23659
rect 34420 23679 34492 23704
tri 34492 23679 34537 23724 sw
rect 70802 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23658 34537 23679
tri 34282 23657 34283 23658 ne
rect 34283 23657 34537 23658
tri 34283 23656 34284 23657 ne
rect 34284 23656 34537 23657
tri 34284 23655 34285 23656 ne
rect 34285 23655 34537 23656
tri 34285 23654 34286 23655 ne
rect 34286 23654 34537 23655
tri 34286 23653 34287 23654 ne
rect 34287 23653 34537 23654
tri 34287 23652 34288 23653 ne
rect 34288 23652 34537 23653
tri 34288 23651 34289 23652 ne
rect 34289 23651 34537 23652
tri 34289 23650 34290 23651 ne
rect 34290 23650 34537 23651
tri 34290 23649 34291 23650 ne
rect 34291 23649 34537 23650
tri 34291 23648 34292 23649 ne
rect 34292 23648 34537 23649
tri 34292 23647 34293 23648 ne
rect 34293 23647 34537 23648
tri 34293 23646 34294 23647 ne
rect 34294 23646 34537 23647
tri 34294 23645 34295 23646 ne
rect 34295 23645 34537 23646
tri 34295 23644 34296 23645 ne
rect 34296 23644 34537 23645
tri 34296 23643 34297 23644 ne
rect 34297 23643 34537 23644
tri 34297 23642 34298 23643 ne
rect 34298 23642 34537 23643
tri 34298 23641 34299 23642 ne
rect 34299 23641 34537 23642
tri 34299 23640 34300 23641 ne
rect 34300 23640 34537 23641
tri 34300 23639 34301 23640 ne
rect 34301 23639 34537 23640
tri 34301 23638 34302 23639 ne
rect 34302 23638 34537 23639
tri 34302 23637 34303 23638 ne
rect 34303 23637 34537 23638
tri 34303 23636 34304 23637 ne
rect 34304 23636 34537 23637
tri 34304 23635 34305 23636 ne
rect 34305 23635 34537 23636
tri 34305 23634 34306 23635 ne
rect 34306 23634 34537 23635
tri 34537 23634 34582 23679 sw
tri 34306 23633 34307 23634 ne
rect 34307 23633 34582 23634
tri 34307 23632 34308 23633 ne
rect 34308 23632 34582 23633
tri 34308 23631 34309 23632 ne
rect 34309 23631 34582 23632
tri 34309 23630 34310 23631 ne
rect 34310 23630 34582 23631
tri 34582 23630 34586 23634 sw
tri 34310 23629 34311 23630 ne
rect 34311 23629 34586 23630
tri 34311 23628 34312 23629 ne
rect 34312 23628 34586 23629
tri 34312 23627 34313 23628 ne
rect 34313 23627 34586 23628
tri 34313 23626 34314 23627 ne
rect 34314 23626 34586 23627
tri 34314 23625 34315 23626 ne
rect 34315 23625 34586 23626
tri 34315 23624 34316 23625 ne
rect 34316 23624 34586 23625
tri 34316 23623 34317 23624 ne
rect 34317 23623 34586 23624
tri 34317 23622 34318 23623 ne
rect 34318 23622 34586 23623
tri 34318 23621 34319 23622 ne
rect 34319 23621 34586 23622
tri 34319 23620 34320 23621 ne
rect 34320 23620 34586 23621
tri 34320 23619 34321 23620 ne
rect 34321 23619 34586 23620
tri 34321 23618 34322 23619 ne
rect 34322 23618 34586 23619
tri 34322 23617 34323 23618 ne
rect 34323 23617 34586 23618
tri 34323 23616 34324 23617 ne
rect 34324 23616 34586 23617
tri 34324 23615 34325 23616 ne
rect 34325 23615 34586 23616
tri 34325 23614 34326 23615 ne
rect 34326 23614 34586 23615
tri 34326 23613 34327 23614 ne
rect 34327 23613 34586 23614
tri 34327 23612 34328 23613 ne
rect 34328 23612 34586 23613
tri 34328 23611 34329 23612 ne
rect 34329 23611 34586 23612
tri 34329 23610 34330 23611 ne
rect 34330 23610 34586 23611
tri 34330 23609 34331 23610 ne
rect 34331 23609 34586 23610
tri 34331 23608 34332 23609 ne
rect 34332 23608 34586 23609
tri 34332 23607 34333 23608 ne
rect 34333 23607 34586 23608
tri 34333 23606 34334 23607 ne
rect 34334 23606 34586 23607
tri 34334 23605 34335 23606 ne
rect 34335 23605 34586 23606
tri 34335 23604 34336 23605 ne
rect 34336 23604 34586 23605
tri 34336 23603 34337 23604 ne
rect 34337 23603 34586 23604
tri 34337 23602 34338 23603 ne
rect 34338 23602 34586 23603
tri 34338 23601 34339 23602 ne
rect 34339 23601 34586 23602
tri 34339 23600 34340 23601 ne
rect 34340 23600 34586 23601
tri 34340 23599 34341 23600 ne
rect 34341 23599 34586 23600
tri 34341 23598 34342 23599 ne
rect 34342 23598 34586 23599
tri 34342 23597 34343 23598 ne
rect 34343 23597 34586 23598
tri 34343 23596 34344 23597 ne
rect 34344 23596 34586 23597
tri 34344 23595 34345 23596 ne
rect 34345 23595 34586 23596
tri 34345 23594 34346 23595 ne
rect 34346 23594 34586 23595
tri 34346 23593 34347 23594 ne
rect 34347 23593 34586 23594
tri 34347 23592 34348 23593 ne
rect 34348 23592 34586 23593
tri 34348 23591 34349 23592 ne
rect 34349 23591 34586 23592
tri 34349 23590 34350 23591 ne
rect 34350 23590 34586 23591
tri 34350 23589 34351 23590 ne
rect 34351 23589 34586 23590
tri 34351 23588 34352 23589 ne
rect 34352 23588 34586 23589
tri 34352 23587 34353 23588 ne
rect 34353 23587 34586 23588
tri 34353 23586 34354 23587 ne
rect 34354 23586 34586 23587
tri 34354 23585 34355 23586 ne
rect 34355 23585 34586 23586
tri 34586 23585 34631 23630 sw
rect 70802 23628 71000 23686
tri 34355 23582 34358 23585 ne
rect 34358 23582 34631 23585
tri 34358 23537 34403 23582 ne
rect 34403 23572 34631 23582
rect 34403 23537 34506 23572
tri 34403 23492 34448 23537 ne
rect 34448 23526 34506 23537
rect 34552 23540 34631 23572
tri 34631 23540 34676 23585 sw
rect 70802 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 34552 23526 34676 23540
rect 34448 23495 34676 23526
tri 34676 23495 34721 23540 sw
rect 70802 23524 71000 23582
rect 34448 23492 34721 23495
tri 34448 23447 34493 23492 ne
rect 34493 23450 34721 23492
tri 34721 23450 34766 23495 sw
rect 70802 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
rect 34493 23448 34766 23450
tri 34766 23448 34768 23450 sw
rect 34493 23447 34768 23448
tri 34493 23444 34496 23447 ne
rect 34496 23444 34768 23447
tri 34496 23443 34497 23444 ne
rect 34497 23443 34768 23444
tri 34497 23442 34498 23443 ne
rect 34498 23442 34768 23443
tri 34498 23441 34499 23442 ne
rect 34499 23441 34768 23442
tri 34499 23440 34500 23441 ne
rect 34500 23440 34768 23441
tri 34500 23439 34501 23440 ne
rect 34501 23439 34638 23440
tri 34501 23438 34502 23439 ne
rect 34502 23438 34638 23439
tri 34502 23437 34503 23438 ne
rect 34503 23437 34638 23438
tri 34503 23436 34504 23437 ne
rect 34504 23436 34638 23437
tri 34504 23435 34505 23436 ne
rect 34505 23435 34638 23436
tri 34505 23434 34506 23435 ne
rect 34506 23434 34638 23435
tri 34506 23433 34507 23434 ne
rect 34507 23433 34638 23434
tri 34507 23432 34508 23433 ne
rect 34508 23432 34638 23433
tri 34508 23431 34509 23432 ne
rect 34509 23431 34638 23432
tri 34509 23430 34510 23431 ne
rect 34510 23430 34638 23431
tri 34510 23429 34511 23430 ne
rect 34511 23429 34638 23430
tri 34511 23428 34512 23429 ne
rect 34512 23428 34638 23429
tri 34512 23427 34513 23428 ne
rect 34513 23427 34638 23428
tri 34513 23426 34514 23427 ne
rect 34514 23426 34638 23427
tri 34514 23425 34515 23426 ne
rect 34515 23425 34638 23426
tri 34515 23424 34516 23425 ne
rect 34516 23424 34638 23425
tri 34516 23423 34517 23424 ne
rect 34517 23423 34638 23424
tri 34517 23422 34518 23423 ne
rect 34518 23422 34638 23423
tri 34518 23421 34519 23422 ne
rect 34519 23421 34638 23422
tri 34519 23420 34520 23421 ne
rect 34520 23420 34638 23421
tri 34520 23419 34521 23420 ne
rect 34521 23419 34638 23420
tri 34521 23418 34522 23419 ne
rect 34522 23418 34638 23419
tri 34522 23417 34523 23418 ne
rect 34523 23417 34638 23418
tri 34523 23416 34524 23417 ne
rect 34524 23416 34638 23417
tri 34524 23415 34525 23416 ne
rect 34525 23415 34638 23416
tri 34525 23414 34526 23415 ne
rect 34526 23414 34638 23415
tri 34526 23413 34527 23414 ne
rect 34527 23413 34638 23414
tri 34527 23412 34528 23413 ne
rect 34528 23412 34638 23413
tri 34528 23411 34529 23412 ne
rect 34529 23411 34638 23412
tri 34529 23410 34530 23411 ne
rect 34530 23410 34638 23411
tri 34530 23409 34531 23410 ne
rect 34531 23409 34638 23410
tri 34531 23408 34532 23409 ne
rect 34532 23408 34638 23409
tri 34532 23407 34533 23408 ne
rect 34533 23407 34638 23408
tri 34533 23406 34534 23407 ne
rect 34534 23406 34638 23407
tri 34534 23405 34535 23406 ne
rect 34535 23405 34638 23406
tri 34535 23404 34536 23405 ne
rect 34536 23404 34638 23405
tri 34536 23403 34537 23404 ne
rect 34537 23403 34638 23404
tri 34537 23402 34538 23403 ne
rect 34538 23402 34638 23403
tri 34538 23401 34539 23402 ne
rect 34539 23401 34638 23402
tri 34539 23400 34540 23401 ne
rect 34540 23400 34638 23401
tri 34540 23399 34541 23400 ne
rect 34541 23399 34638 23400
tri 34541 23398 34542 23399 ne
rect 34542 23398 34638 23399
tri 34542 23397 34543 23398 ne
rect 34543 23397 34638 23398
tri 34543 23396 34544 23397 ne
rect 34544 23396 34638 23397
tri 34544 23395 34545 23396 ne
rect 34545 23395 34638 23396
tri 34545 23394 34546 23395 ne
rect 34546 23394 34638 23395
rect 34684 23403 34768 23440
tri 34768 23403 34813 23448 sw
rect 70802 23420 71000 23478
rect 34684 23394 34813 23403
tri 34546 23393 34547 23394 ne
rect 34547 23393 34813 23394
tri 34547 23392 34548 23393 ne
rect 34548 23392 34813 23393
tri 34548 23391 34549 23392 ne
rect 34549 23391 34813 23392
tri 34549 23390 34550 23391 ne
rect 34550 23390 34813 23391
tri 34550 23389 34551 23390 ne
rect 34551 23389 34813 23390
tri 34551 23388 34552 23389 ne
rect 34552 23388 34813 23389
tri 34552 23387 34553 23388 ne
rect 34553 23387 34813 23388
tri 34553 23386 34554 23387 ne
rect 34554 23386 34813 23387
tri 34554 23385 34555 23386 ne
rect 34555 23385 34813 23386
tri 34555 23384 34556 23385 ne
rect 34556 23384 34813 23385
tri 34556 23383 34557 23384 ne
rect 34557 23383 34813 23384
tri 34557 23382 34558 23383 ne
rect 34558 23382 34813 23383
tri 34558 23381 34559 23382 ne
rect 34559 23381 34813 23382
tri 34559 23380 34560 23381 ne
rect 34560 23380 34813 23381
tri 34560 23379 34561 23380 ne
rect 34561 23379 34813 23380
tri 34561 23378 34562 23379 ne
rect 34562 23378 34813 23379
tri 34562 23377 34563 23378 ne
rect 34563 23377 34813 23378
tri 34563 23376 34564 23377 ne
rect 34564 23376 34813 23377
tri 34564 23375 34565 23376 ne
rect 34565 23375 34813 23376
tri 34565 23374 34566 23375 ne
rect 34566 23374 34813 23375
tri 34566 23373 34567 23374 ne
rect 34567 23373 34813 23374
tri 34567 23372 34568 23373 ne
rect 34568 23372 34813 23373
tri 34568 23371 34569 23372 ne
rect 34569 23371 34813 23372
tri 34569 23370 34570 23371 ne
rect 34570 23370 34813 23371
tri 34570 23369 34571 23370 ne
rect 34571 23369 34813 23370
tri 34571 23368 34572 23369 ne
rect 34572 23368 34813 23369
tri 34572 23367 34573 23368 ne
rect 34573 23367 34813 23368
tri 34573 23366 34574 23367 ne
rect 34574 23366 34813 23367
tri 34574 23365 34575 23366 ne
rect 34575 23365 34813 23366
tri 34575 23364 34576 23365 ne
rect 34576 23364 34813 23365
tri 34576 23363 34577 23364 ne
rect 34577 23363 34813 23364
tri 34577 23362 34578 23363 ne
rect 34578 23362 34813 23363
tri 34578 23361 34579 23362 ne
rect 34579 23361 34813 23362
tri 34579 23360 34580 23361 ne
rect 34580 23360 34813 23361
tri 34580 23359 34581 23360 ne
rect 34581 23359 34813 23360
tri 34581 23358 34582 23359 ne
rect 34582 23358 34813 23359
tri 34813 23358 34858 23403 sw
rect 70802 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34582 23357 34583 23358 ne
rect 34583 23357 34858 23358
tri 34583 23356 34584 23357 ne
rect 34584 23356 34858 23357
tri 34584 23355 34585 23356 ne
rect 34585 23355 34858 23356
tri 34585 23354 34586 23355 ne
rect 34586 23354 34858 23355
tri 34586 23353 34587 23354 ne
rect 34587 23353 34858 23354
tri 34587 23352 34588 23353 ne
rect 34588 23352 34858 23353
tri 34588 23351 34589 23352 ne
rect 34589 23351 34858 23352
tri 34589 23350 34590 23351 ne
rect 34590 23350 34858 23351
tri 34590 23349 34591 23350 ne
rect 34591 23349 34858 23350
tri 34591 23348 34592 23349 ne
rect 34592 23348 34858 23349
tri 34592 23347 34593 23348 ne
rect 34593 23347 34858 23348
tri 34593 23346 34594 23347 ne
rect 34594 23346 34858 23347
tri 34594 23345 34595 23346 ne
rect 34595 23345 34858 23346
tri 34595 23344 34596 23345 ne
rect 34596 23344 34858 23345
tri 34596 23343 34597 23344 ne
rect 34597 23343 34858 23344
tri 34597 23342 34598 23343 ne
rect 34598 23342 34858 23343
tri 34598 23341 34599 23342 ne
rect 34599 23341 34858 23342
tri 34599 23340 34600 23341 ne
rect 34600 23340 34858 23341
tri 34600 23339 34601 23340 ne
rect 34601 23339 34858 23340
tri 34601 23338 34602 23339 ne
rect 34602 23338 34858 23339
tri 34602 23337 34603 23338 ne
rect 34603 23337 34858 23338
tri 34603 23336 34604 23337 ne
rect 34604 23336 34858 23337
tri 34604 23335 34605 23336 ne
rect 34605 23335 34858 23336
tri 34605 23334 34606 23335 ne
rect 34606 23334 34858 23335
tri 34606 23333 34607 23334 ne
rect 34607 23333 34858 23334
tri 34607 23332 34608 23333 ne
rect 34608 23332 34858 23333
tri 34608 23331 34609 23332 ne
rect 34609 23331 34858 23332
tri 34609 23330 34610 23331 ne
rect 34610 23330 34858 23331
tri 34610 23329 34611 23330 ne
rect 34611 23329 34858 23330
tri 34611 23328 34612 23329 ne
rect 34612 23328 34858 23329
tri 34612 23327 34613 23328 ne
rect 34613 23327 34858 23328
tri 34613 23326 34614 23327 ne
rect 34614 23326 34858 23327
tri 34614 23325 34615 23326 ne
rect 34615 23325 34858 23326
tri 34615 23324 34616 23325 ne
rect 34616 23324 34858 23325
tri 34616 23323 34617 23324 ne
rect 34617 23323 34858 23324
tri 34617 23322 34618 23323 ne
rect 34618 23322 34858 23323
tri 34618 23321 34619 23322 ne
rect 34619 23321 34858 23322
tri 34619 23320 34620 23321 ne
rect 34620 23320 34858 23321
tri 34620 23319 34621 23320 ne
rect 34621 23319 34858 23320
tri 34621 23318 34622 23319 ne
rect 34622 23318 34858 23319
tri 34622 23317 34623 23318 ne
rect 34623 23317 34858 23318
tri 34623 23316 34624 23317 ne
rect 34624 23316 34858 23317
tri 34624 23315 34625 23316 ne
rect 34625 23315 34858 23316
tri 34625 23314 34626 23315 ne
rect 34626 23314 34858 23315
tri 34626 23313 34627 23314 ne
rect 34627 23313 34858 23314
tri 34858 23313 34903 23358 sw
rect 70802 23316 71000 23374
tri 34627 23312 34628 23313 ne
rect 34628 23312 34903 23313
tri 34628 23311 34629 23312 ne
rect 34629 23311 34903 23312
tri 34629 23310 34630 23311 ne
rect 34630 23310 34903 23311
tri 34630 23309 34631 23310 ne
rect 34631 23309 34903 23310
tri 34903 23309 34907 23313 sw
tri 34631 23264 34676 23309 ne
rect 34676 23308 34907 23309
rect 34676 23264 34770 23308
tri 34676 23263 34677 23264 ne
rect 34677 23263 34770 23264
tri 34677 23218 34722 23263 ne
rect 34722 23262 34770 23263
rect 34816 23268 34907 23308
tri 34907 23268 34948 23309 sw
rect 70802 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 34816 23262 34948 23268
rect 34722 23223 34948 23262
tri 34948 23223 34993 23268 sw
rect 34722 23218 34993 23223
tri 34722 23173 34767 23218 ne
rect 34767 23178 34993 23218
tri 34993 23178 35038 23223 sw
rect 70802 23212 71000 23270
rect 34767 23176 35038 23178
rect 34767 23173 34902 23176
tri 34767 23169 34771 23173 ne
rect 34771 23169 34902 23173
tri 34771 23168 34772 23169 ne
rect 34772 23168 34902 23169
tri 34772 23167 34773 23168 ne
rect 34773 23167 34902 23168
tri 34773 23166 34774 23167 ne
rect 34774 23166 34902 23167
tri 34774 23165 34775 23166 ne
rect 34775 23165 34902 23166
tri 34775 23164 34776 23165 ne
rect 34776 23164 34902 23165
tri 34776 23163 34777 23164 ne
rect 34777 23163 34902 23164
tri 34777 23162 34778 23163 ne
rect 34778 23162 34902 23163
tri 34778 23161 34779 23162 ne
rect 34779 23161 34902 23162
tri 34779 23160 34780 23161 ne
rect 34780 23160 34902 23161
tri 34780 23159 34781 23160 ne
rect 34781 23159 34902 23160
tri 34781 23158 34782 23159 ne
rect 34782 23158 34902 23159
tri 34782 23157 34783 23158 ne
rect 34783 23157 34902 23158
tri 34783 23156 34784 23157 ne
rect 34784 23156 34902 23157
tri 34784 23155 34785 23156 ne
rect 34785 23155 34902 23156
tri 34785 23154 34786 23155 ne
rect 34786 23154 34902 23155
tri 34786 23153 34787 23154 ne
rect 34787 23153 34902 23154
tri 34787 23152 34788 23153 ne
rect 34788 23152 34902 23153
tri 34788 23151 34789 23152 ne
rect 34789 23151 34902 23152
tri 34789 23150 34790 23151 ne
rect 34790 23150 34902 23151
tri 34790 23149 34791 23150 ne
rect 34791 23149 34902 23150
tri 34791 23148 34792 23149 ne
rect 34792 23148 34902 23149
tri 34792 23147 34793 23148 ne
rect 34793 23147 34902 23148
tri 34793 23146 34794 23147 ne
rect 34794 23146 34902 23147
tri 34794 23145 34795 23146 ne
rect 34795 23145 34902 23146
tri 34795 23144 34796 23145 ne
rect 34796 23144 34902 23145
tri 34796 23143 34797 23144 ne
rect 34797 23143 34902 23144
tri 34797 23142 34798 23143 ne
rect 34798 23142 34902 23143
tri 34798 23141 34799 23142 ne
rect 34799 23141 34902 23142
tri 34799 23140 34800 23141 ne
rect 34800 23140 34902 23141
tri 34800 23139 34801 23140 ne
rect 34801 23139 34902 23140
tri 34801 23138 34802 23139 ne
rect 34802 23138 34902 23139
tri 34802 23137 34803 23138 ne
rect 34803 23137 34902 23138
tri 34803 23136 34804 23137 ne
rect 34804 23136 34902 23137
tri 34804 23135 34805 23136 ne
rect 34805 23135 34902 23136
tri 34805 23134 34806 23135 ne
rect 34806 23134 34902 23135
tri 34806 23133 34807 23134 ne
rect 34807 23133 34902 23134
tri 34807 23132 34808 23133 ne
rect 34808 23132 34902 23133
tri 34808 23131 34809 23132 ne
rect 34809 23131 34902 23132
tri 34809 23130 34810 23131 ne
rect 34810 23130 34902 23131
rect 34948 23168 35038 23176
tri 35038 23168 35048 23178 sw
rect 34948 23130 35048 23168
tri 34810 23129 34811 23130 ne
rect 34811 23129 35048 23130
tri 34811 23128 34812 23129 ne
rect 34812 23128 35048 23129
tri 34812 23127 34813 23128 ne
rect 34813 23127 35048 23128
tri 34813 23126 34814 23127 ne
rect 34814 23126 35048 23127
tri 34814 23125 34815 23126 ne
rect 34815 23125 35048 23126
tri 34815 23124 34816 23125 ne
rect 34816 23124 35048 23125
tri 34816 23123 34817 23124 ne
rect 34817 23123 35048 23124
tri 35048 23123 35093 23168 sw
rect 70802 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
tri 34817 23122 34818 23123 ne
rect 34818 23122 35093 23123
tri 34818 23121 34819 23122 ne
rect 34819 23121 35093 23122
tri 34819 23120 34820 23121 ne
rect 34820 23120 35093 23121
tri 34820 23119 34821 23120 ne
rect 34821 23119 35093 23120
tri 34821 23118 34822 23119 ne
rect 34822 23118 35093 23119
tri 34822 23117 34823 23118 ne
rect 34823 23117 35093 23118
tri 34823 23116 34824 23117 ne
rect 34824 23116 35093 23117
tri 34824 23115 34825 23116 ne
rect 34825 23115 35093 23116
tri 34825 23114 34826 23115 ne
rect 34826 23114 35093 23115
tri 34826 23113 34827 23114 ne
rect 34827 23113 35093 23114
tri 34827 23112 34828 23113 ne
rect 34828 23112 35093 23113
tri 34828 23111 34829 23112 ne
rect 34829 23111 35093 23112
tri 34829 23110 34830 23111 ne
rect 34830 23110 35093 23111
tri 34830 23109 34831 23110 ne
rect 34831 23109 35093 23110
tri 34831 23108 34832 23109 ne
rect 34832 23108 35093 23109
tri 34832 23107 34833 23108 ne
rect 34833 23107 35093 23108
tri 34833 23106 34834 23107 ne
rect 34834 23106 35093 23107
tri 34834 23105 34835 23106 ne
rect 34835 23105 35093 23106
tri 34835 23104 34836 23105 ne
rect 34836 23104 35093 23105
tri 34836 23103 34837 23104 ne
rect 34837 23103 35093 23104
tri 34837 23102 34838 23103 ne
rect 34838 23102 35093 23103
tri 34838 23101 34839 23102 ne
rect 34839 23101 35093 23102
tri 34839 23100 34840 23101 ne
rect 34840 23100 35093 23101
tri 34840 23099 34841 23100 ne
rect 34841 23099 35093 23100
tri 34841 23098 34842 23099 ne
rect 34842 23098 35093 23099
tri 34842 23097 34843 23098 ne
rect 34843 23097 35093 23098
tri 34843 23096 34844 23097 ne
rect 34844 23096 35093 23097
tri 34844 23095 34845 23096 ne
rect 34845 23095 35093 23096
tri 34845 23094 34846 23095 ne
rect 34846 23094 35093 23095
tri 34846 23093 34847 23094 ne
rect 34847 23093 35093 23094
tri 34847 23092 34848 23093 ne
rect 34848 23092 35093 23093
tri 34848 23091 34849 23092 ne
rect 34849 23091 35093 23092
tri 34849 23090 34850 23091 ne
rect 34850 23090 35093 23091
tri 34850 23089 34851 23090 ne
rect 34851 23089 35093 23090
tri 34851 23088 34852 23089 ne
rect 34852 23088 35093 23089
tri 34852 23087 34853 23088 ne
rect 34853 23087 35093 23088
tri 34853 23086 34854 23087 ne
rect 34854 23086 35093 23087
tri 34854 23085 34855 23086 ne
rect 34855 23085 35093 23086
tri 34855 23084 34856 23085 ne
rect 34856 23084 35093 23085
tri 34856 23083 34857 23084 ne
rect 34857 23083 35093 23084
tri 34857 23082 34858 23083 ne
rect 34858 23082 35093 23083
tri 34858 23081 34859 23082 ne
rect 34859 23081 35093 23082
tri 34859 23080 34860 23081 ne
rect 34860 23080 35093 23081
tri 34860 23079 34861 23080 ne
rect 34861 23079 35093 23080
tri 34861 23078 34862 23079 ne
rect 34862 23078 35093 23079
tri 35093 23078 35138 23123 sw
rect 70802 23108 71000 23166
tri 34862 23077 34863 23078 ne
rect 34863 23077 35138 23078
tri 34863 23076 34864 23077 ne
rect 34864 23076 35138 23077
tri 34864 23075 34865 23076 ne
rect 34865 23075 35138 23076
tri 34865 23074 34866 23075 ne
rect 34866 23074 35138 23075
tri 34866 23073 34867 23074 ne
rect 34867 23073 35138 23074
tri 34867 23072 34868 23073 ne
rect 34868 23072 35138 23073
tri 34868 23071 34869 23072 ne
rect 34869 23071 35138 23072
tri 34869 23070 34870 23071 ne
rect 34870 23070 35138 23071
tri 34870 23069 34871 23070 ne
rect 34871 23069 35138 23070
tri 34871 23068 34872 23069 ne
rect 34872 23068 35138 23069
tri 34872 23067 34873 23068 ne
rect 34873 23067 35138 23068
tri 34873 23066 34874 23067 ne
rect 34874 23066 35138 23067
tri 34874 23065 34875 23066 ne
rect 34875 23065 35138 23066
tri 34875 23064 34876 23065 ne
rect 34876 23064 35138 23065
tri 34876 23063 34877 23064 ne
rect 34877 23063 35138 23064
tri 34877 23062 34878 23063 ne
rect 34878 23062 35138 23063
tri 34878 23061 34879 23062 ne
rect 34879 23061 35138 23062
tri 34879 23060 34880 23061 ne
rect 34880 23060 35138 23061
tri 34880 23059 34881 23060 ne
rect 34881 23059 35138 23060
tri 34881 23058 34882 23059 ne
rect 34882 23058 35138 23059
tri 34882 23057 34883 23058 ne
rect 34883 23057 35138 23058
tri 34883 23056 34884 23057 ne
rect 34884 23056 35138 23057
tri 34884 23055 34885 23056 ne
rect 34885 23055 35138 23056
tri 34885 23054 34886 23055 ne
rect 34886 23054 35138 23055
tri 34886 23053 34887 23054 ne
rect 34887 23053 35138 23054
tri 34887 23052 34888 23053 ne
rect 34888 23052 35138 23053
tri 34888 23051 34889 23052 ne
rect 34889 23051 35138 23052
tri 34889 23050 34890 23051 ne
rect 34890 23050 35138 23051
tri 34890 23049 34891 23050 ne
rect 34891 23049 35138 23050
tri 34891 23048 34892 23049 ne
rect 34892 23048 35138 23049
tri 34892 23047 34893 23048 ne
rect 34893 23047 35138 23048
tri 34893 23046 34894 23047 ne
rect 34894 23046 35138 23047
tri 34894 23045 34895 23046 ne
rect 34895 23045 35138 23046
tri 34895 23044 34896 23045 ne
rect 34896 23044 35138 23045
tri 34896 23043 34897 23044 ne
rect 34897 23043 35034 23044
tri 34897 23042 34898 23043 ne
rect 34898 23042 35034 23043
tri 34898 23041 34899 23042 ne
rect 34899 23041 35034 23042
tri 34899 23040 34900 23041 ne
rect 34900 23040 35034 23041
tri 34900 23039 34901 23040 ne
rect 34901 23039 35034 23040
tri 34901 23038 34902 23039 ne
rect 34902 23038 35034 23039
tri 34902 23037 34903 23038 ne
rect 34903 23037 35034 23038
tri 34903 23036 34904 23037 ne
rect 34904 23036 35034 23037
tri 34904 23035 34905 23036 ne
rect 34905 23035 35034 23036
tri 34905 23034 34906 23035 ne
rect 34906 23034 35034 23035
tri 34906 23033 34907 23034 ne
rect 34907 23033 35034 23034
tri 34907 22992 34948 23033 ne
rect 34948 22998 35034 23033
rect 35080 23033 35138 23044
tri 35138 23033 35183 23078 sw
rect 70802 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 35080 22998 35183 23033
rect 34948 22992 35183 22998
tri 35183 22992 35224 23033 sw
rect 70802 23004 71000 23062
tri 34948 22988 34952 22992 ne
rect 34952 22988 35224 22992
tri 34952 22947 34993 22988 ne
rect 34993 22947 35224 22988
tri 35224 22947 35269 22992 sw
rect 70802 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 34993 22902 35038 22947 ne
rect 35038 22912 35269 22947
rect 35038 22902 35166 22912
tri 35038 22895 35045 22902 ne
rect 35045 22895 35166 22902
tri 35045 22894 35046 22895 ne
rect 35046 22894 35166 22895
tri 35046 22893 35047 22894 ne
rect 35047 22893 35166 22894
tri 35047 22892 35048 22893 ne
rect 35048 22892 35166 22893
tri 35048 22891 35049 22892 ne
rect 35049 22891 35166 22892
tri 35049 22890 35050 22891 ne
rect 35050 22890 35166 22891
tri 35050 22889 35051 22890 ne
rect 35051 22889 35166 22890
tri 35051 22888 35052 22889 ne
rect 35052 22888 35166 22889
tri 35052 22887 35053 22888 ne
rect 35053 22887 35166 22888
tri 35053 22886 35054 22887 ne
rect 35054 22886 35166 22887
tri 35054 22885 35055 22886 ne
rect 35055 22885 35166 22886
tri 35055 22884 35056 22885 ne
rect 35056 22884 35166 22885
tri 35056 22883 35057 22884 ne
rect 35057 22883 35166 22884
tri 35057 22882 35058 22883 ne
rect 35058 22882 35166 22883
tri 35058 22881 35059 22882 ne
rect 35059 22881 35166 22882
tri 35059 22880 35060 22881 ne
rect 35060 22880 35166 22881
tri 35060 22879 35061 22880 ne
rect 35061 22879 35166 22880
tri 35061 22878 35062 22879 ne
rect 35062 22878 35166 22879
tri 35062 22877 35063 22878 ne
rect 35063 22877 35166 22878
tri 35063 22876 35064 22877 ne
rect 35064 22876 35166 22877
tri 35064 22875 35065 22876 ne
rect 35065 22875 35166 22876
tri 35065 22874 35066 22875 ne
rect 35066 22874 35166 22875
tri 35066 22873 35067 22874 ne
rect 35067 22873 35166 22874
tri 35067 22872 35068 22873 ne
rect 35068 22872 35166 22873
tri 35068 22871 35069 22872 ne
rect 35069 22871 35166 22872
tri 35069 22870 35070 22871 ne
rect 35070 22870 35166 22871
tri 35070 22869 35071 22870 ne
rect 35071 22869 35166 22870
tri 35071 22868 35072 22869 ne
rect 35072 22868 35166 22869
tri 35072 22867 35073 22868 ne
rect 35073 22867 35166 22868
tri 35073 22866 35074 22867 ne
rect 35074 22866 35166 22867
rect 35212 22902 35269 22912
tri 35269 22902 35314 22947 sw
rect 35212 22866 35314 22902
tri 35074 22865 35075 22866 ne
rect 35075 22865 35314 22866
tri 35075 22864 35076 22865 ne
rect 35076 22864 35314 22865
tri 35076 22863 35077 22864 ne
rect 35077 22863 35314 22864
tri 35077 22862 35078 22863 ne
rect 35078 22862 35314 22863
tri 35078 22861 35079 22862 ne
rect 35079 22861 35314 22862
tri 35079 22860 35080 22861 ne
rect 35080 22860 35314 22861
tri 35080 22859 35081 22860 ne
rect 35081 22859 35314 22860
tri 35081 22858 35082 22859 ne
rect 35082 22858 35314 22859
tri 35082 22857 35083 22858 ne
rect 35083 22857 35314 22858
tri 35314 22857 35359 22902 sw
rect 70802 22900 71000 22958
tri 35083 22856 35084 22857 ne
rect 35084 22856 35359 22857
tri 35084 22855 35085 22856 ne
rect 35085 22855 35359 22856
tri 35085 22854 35086 22855 ne
rect 35086 22854 35359 22855
tri 35086 22853 35087 22854 ne
rect 35087 22853 35359 22854
tri 35087 22852 35088 22853 ne
rect 35088 22852 35359 22853
tri 35088 22851 35089 22852 ne
rect 35089 22851 35359 22852
tri 35089 22850 35090 22851 ne
rect 35090 22850 35359 22851
tri 35090 22849 35091 22850 ne
rect 35091 22849 35359 22850
tri 35091 22848 35092 22849 ne
rect 35092 22848 35359 22849
tri 35092 22847 35093 22848 ne
rect 35093 22847 35359 22848
tri 35359 22847 35369 22857 sw
rect 70802 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
tri 35093 22846 35094 22847 ne
rect 35094 22846 35369 22847
tri 35094 22845 35095 22846 ne
rect 35095 22845 35369 22846
tri 35095 22844 35096 22845 ne
rect 35096 22844 35369 22845
tri 35096 22843 35097 22844 ne
rect 35097 22843 35369 22844
tri 35097 22842 35098 22843 ne
rect 35098 22842 35369 22843
tri 35098 22841 35099 22842 ne
rect 35099 22841 35369 22842
tri 35099 22840 35100 22841 ne
rect 35100 22840 35369 22841
tri 35100 22839 35101 22840 ne
rect 35101 22839 35369 22840
tri 35101 22838 35102 22839 ne
rect 35102 22838 35369 22839
tri 35102 22837 35103 22838 ne
rect 35103 22837 35369 22838
tri 35103 22836 35104 22837 ne
rect 35104 22836 35369 22837
tri 35104 22835 35105 22836 ne
rect 35105 22835 35369 22836
tri 35105 22834 35106 22835 ne
rect 35106 22834 35369 22835
tri 35106 22833 35107 22834 ne
rect 35107 22833 35369 22834
tri 35107 22832 35108 22833 ne
rect 35108 22832 35369 22833
tri 35108 22831 35109 22832 ne
rect 35109 22831 35369 22832
tri 35109 22830 35110 22831 ne
rect 35110 22830 35369 22831
tri 35110 22829 35111 22830 ne
rect 35111 22829 35369 22830
tri 35111 22828 35112 22829 ne
rect 35112 22828 35369 22829
tri 35112 22827 35113 22828 ne
rect 35113 22827 35369 22828
tri 35113 22826 35114 22827 ne
rect 35114 22826 35369 22827
tri 35114 22825 35115 22826 ne
rect 35115 22825 35369 22826
tri 35115 22824 35116 22825 ne
rect 35116 22824 35369 22825
tri 35116 22823 35117 22824 ne
rect 35117 22823 35369 22824
tri 35117 22822 35118 22823 ne
rect 35118 22822 35369 22823
tri 35118 22821 35119 22822 ne
rect 35119 22821 35369 22822
tri 35119 22820 35120 22821 ne
rect 35120 22820 35369 22821
tri 35120 22819 35121 22820 ne
rect 35121 22819 35369 22820
tri 35121 22818 35122 22819 ne
rect 35122 22818 35369 22819
tri 35122 22817 35123 22818 ne
rect 35123 22817 35369 22818
tri 35123 22816 35124 22817 ne
rect 35124 22816 35369 22817
tri 35124 22815 35125 22816 ne
rect 35125 22815 35369 22816
tri 35125 22814 35126 22815 ne
rect 35126 22814 35369 22815
tri 35126 22813 35127 22814 ne
rect 35127 22813 35369 22814
tri 35127 22812 35128 22813 ne
rect 35128 22812 35369 22813
tri 35128 22811 35129 22812 ne
rect 35129 22811 35369 22812
tri 35129 22810 35130 22811 ne
rect 35130 22810 35369 22811
tri 35130 22809 35131 22810 ne
rect 35131 22809 35369 22810
tri 35131 22808 35132 22809 ne
rect 35132 22808 35369 22809
tri 35132 22807 35133 22808 ne
rect 35133 22807 35369 22808
tri 35133 22806 35134 22807 ne
rect 35134 22806 35369 22807
tri 35134 22805 35135 22806 ne
rect 35135 22805 35369 22806
tri 35135 22804 35136 22805 ne
rect 35136 22804 35369 22805
tri 35136 22803 35137 22804 ne
rect 35137 22803 35369 22804
tri 35137 22802 35138 22803 ne
rect 35138 22802 35369 22803
tri 35369 22802 35414 22847 sw
tri 35138 22801 35139 22802 ne
rect 35139 22801 35414 22802
tri 35139 22800 35140 22801 ne
rect 35140 22800 35414 22801
tri 35140 22799 35141 22800 ne
rect 35141 22799 35414 22800
tri 35141 22798 35142 22799 ne
rect 35142 22798 35414 22799
tri 35142 22797 35143 22798 ne
rect 35143 22797 35414 22798
tri 35143 22796 35144 22797 ne
rect 35144 22796 35414 22797
tri 35144 22795 35145 22796 ne
rect 35145 22795 35414 22796
tri 35145 22794 35146 22795 ne
rect 35146 22794 35414 22795
tri 35146 22793 35147 22794 ne
rect 35147 22793 35414 22794
tri 35147 22792 35148 22793 ne
rect 35148 22792 35414 22793
tri 35148 22791 35149 22792 ne
rect 35149 22791 35414 22792
tri 35149 22790 35150 22791 ne
rect 35150 22790 35414 22791
tri 35150 22789 35151 22790 ne
rect 35151 22789 35414 22790
tri 35151 22788 35152 22789 ne
rect 35152 22788 35414 22789
tri 35152 22787 35153 22788 ne
rect 35153 22787 35414 22788
tri 35153 22786 35154 22787 ne
rect 35154 22786 35414 22787
tri 35154 22785 35155 22786 ne
rect 35155 22785 35414 22786
tri 35155 22784 35156 22785 ne
rect 35156 22784 35414 22785
tri 35156 22783 35157 22784 ne
rect 35157 22783 35414 22784
tri 35157 22782 35158 22783 ne
rect 35158 22782 35414 22783
tri 35158 22781 35159 22782 ne
rect 35159 22781 35414 22782
tri 35159 22780 35160 22781 ne
rect 35160 22780 35414 22781
tri 35160 22779 35161 22780 ne
rect 35161 22779 35298 22780
tri 35161 22778 35162 22779 ne
rect 35162 22778 35298 22779
tri 35162 22777 35163 22778 ne
rect 35163 22777 35298 22778
tri 35163 22776 35164 22777 ne
rect 35164 22776 35298 22777
tri 35164 22775 35165 22776 ne
rect 35165 22775 35298 22776
tri 35165 22774 35166 22775 ne
rect 35166 22774 35298 22775
tri 35166 22773 35167 22774 ne
rect 35167 22773 35298 22774
tri 35167 22772 35168 22773 ne
rect 35168 22772 35298 22773
tri 35168 22771 35169 22772 ne
rect 35169 22771 35298 22772
tri 35169 22770 35170 22771 ne
rect 35170 22770 35298 22771
tri 35170 22769 35171 22770 ne
rect 35171 22769 35298 22770
tri 35171 22768 35172 22769 ne
rect 35172 22768 35298 22769
tri 35172 22767 35173 22768 ne
rect 35173 22767 35298 22768
tri 35173 22766 35174 22767 ne
rect 35174 22766 35298 22767
tri 35174 22765 35175 22766 ne
rect 35175 22765 35298 22766
tri 35175 22764 35176 22765 ne
rect 35176 22764 35298 22765
tri 35176 22763 35177 22764 ne
rect 35177 22763 35298 22764
tri 35177 22762 35178 22763 ne
rect 35178 22762 35298 22763
tri 35178 22761 35179 22762 ne
rect 35179 22761 35298 22762
tri 35179 22760 35180 22761 ne
rect 35180 22760 35298 22761
tri 35180 22759 35181 22760 ne
rect 35181 22759 35298 22760
tri 35181 22758 35182 22759 ne
rect 35182 22758 35298 22759
tri 35182 22757 35183 22758 ne
rect 35183 22757 35298 22758
tri 35183 22712 35228 22757 ne
rect 35228 22734 35298 22757
rect 35344 22757 35414 22780
tri 35414 22757 35459 22802 sw
rect 70802 22796 71000 22854
rect 35344 22734 35459 22757
rect 35228 22712 35459 22734
tri 35459 22712 35504 22757 sw
rect 70802 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
tri 35228 22667 35273 22712 ne
rect 35273 22671 35504 22712
tri 35504 22671 35545 22712 sw
rect 70802 22692 71000 22750
rect 35273 22667 35545 22671
tri 35273 22626 35314 22667 ne
rect 35314 22648 35545 22667
rect 35314 22626 35430 22648
tri 35314 22622 35318 22626 ne
rect 35318 22622 35430 22626
tri 35318 22621 35319 22622 ne
rect 35319 22621 35430 22622
tri 35319 22620 35320 22621 ne
rect 35320 22620 35430 22621
tri 35320 22619 35321 22620 ne
rect 35321 22619 35430 22620
tri 35321 22618 35322 22619 ne
rect 35322 22618 35430 22619
tri 35322 22617 35323 22618 ne
rect 35323 22617 35430 22618
tri 35323 22616 35324 22617 ne
rect 35324 22616 35430 22617
tri 35324 22615 35325 22616 ne
rect 35325 22615 35430 22616
tri 35325 22614 35326 22615 ne
rect 35326 22614 35430 22615
tri 35326 22613 35327 22614 ne
rect 35327 22613 35430 22614
tri 35327 22612 35328 22613 ne
rect 35328 22612 35430 22613
tri 35328 22611 35329 22612 ne
rect 35329 22611 35430 22612
tri 35329 22610 35330 22611 ne
rect 35330 22610 35430 22611
tri 35330 22609 35331 22610 ne
rect 35331 22609 35430 22610
tri 35331 22608 35332 22609 ne
rect 35332 22608 35430 22609
tri 35332 22607 35333 22608 ne
rect 35333 22607 35430 22608
tri 35333 22606 35334 22607 ne
rect 35334 22606 35430 22607
tri 35334 22605 35335 22606 ne
rect 35335 22605 35430 22606
tri 35335 22604 35336 22605 ne
rect 35336 22604 35430 22605
tri 35336 22603 35337 22604 ne
rect 35337 22603 35430 22604
tri 35337 22602 35338 22603 ne
rect 35338 22602 35430 22603
rect 35476 22626 35545 22648
tri 35545 22626 35590 22671 sw
rect 70802 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22602 35590 22626
tri 35338 22601 35339 22602 ne
rect 35339 22601 35590 22602
tri 35339 22600 35340 22601 ne
rect 35340 22600 35590 22601
tri 35340 22599 35341 22600 ne
rect 35341 22599 35590 22600
tri 35341 22598 35342 22599 ne
rect 35342 22598 35590 22599
tri 35342 22597 35343 22598 ne
rect 35343 22597 35590 22598
tri 35343 22596 35344 22597 ne
rect 35344 22596 35590 22597
tri 35344 22595 35345 22596 ne
rect 35345 22595 35590 22596
tri 35345 22594 35346 22595 ne
rect 35346 22594 35590 22595
tri 35346 22593 35347 22594 ne
rect 35347 22593 35590 22594
tri 35347 22592 35348 22593 ne
rect 35348 22592 35590 22593
tri 35348 22591 35349 22592 ne
rect 35349 22591 35590 22592
tri 35349 22590 35350 22591 ne
rect 35350 22590 35590 22591
tri 35350 22589 35351 22590 ne
rect 35351 22589 35590 22590
tri 35351 22588 35352 22589 ne
rect 35352 22588 35590 22589
tri 35352 22587 35353 22588 ne
rect 35353 22587 35590 22588
tri 35353 22586 35354 22587 ne
rect 35354 22586 35590 22587
tri 35354 22585 35355 22586 ne
rect 35355 22585 35590 22586
tri 35355 22584 35356 22585 ne
rect 35356 22584 35590 22585
tri 35356 22583 35357 22584 ne
rect 35357 22583 35590 22584
tri 35357 22582 35358 22583 ne
rect 35358 22582 35590 22583
tri 35358 22581 35359 22582 ne
rect 35359 22581 35590 22582
tri 35590 22581 35635 22626 sw
rect 70802 22588 71000 22646
tri 35359 22580 35360 22581 ne
rect 35360 22580 35635 22581
tri 35360 22579 35361 22580 ne
rect 35361 22579 35635 22580
tri 35361 22578 35362 22579 ne
rect 35362 22578 35635 22579
tri 35362 22577 35363 22578 ne
rect 35363 22577 35635 22578
tri 35363 22576 35364 22577 ne
rect 35364 22576 35635 22577
tri 35364 22575 35365 22576 ne
rect 35365 22575 35635 22576
tri 35365 22574 35366 22575 ne
rect 35366 22574 35635 22575
tri 35366 22573 35367 22574 ne
rect 35367 22573 35635 22574
tri 35367 22572 35368 22573 ne
rect 35368 22572 35635 22573
tri 35368 22571 35369 22572 ne
rect 35369 22571 35635 22572
tri 35369 22570 35370 22571 ne
rect 35370 22570 35635 22571
tri 35370 22569 35371 22570 ne
rect 35371 22569 35635 22570
tri 35371 22568 35372 22569 ne
rect 35372 22568 35635 22569
tri 35372 22567 35373 22568 ne
rect 35373 22567 35635 22568
tri 35373 22566 35374 22567 ne
rect 35374 22566 35635 22567
tri 35374 22565 35375 22566 ne
rect 35375 22565 35635 22566
tri 35375 22564 35376 22565 ne
rect 35376 22564 35635 22565
tri 35376 22563 35377 22564 ne
rect 35377 22563 35635 22564
tri 35377 22562 35378 22563 ne
rect 35378 22562 35635 22563
tri 35378 22561 35379 22562 ne
rect 35379 22561 35635 22562
tri 35379 22560 35380 22561 ne
rect 35380 22560 35635 22561
tri 35380 22559 35381 22560 ne
rect 35381 22559 35635 22560
tri 35381 22558 35382 22559 ne
rect 35382 22558 35635 22559
tri 35382 22557 35383 22558 ne
rect 35383 22557 35635 22558
tri 35383 22556 35384 22557 ne
rect 35384 22556 35635 22557
tri 35384 22555 35385 22556 ne
rect 35385 22555 35635 22556
tri 35385 22554 35386 22555 ne
rect 35386 22554 35635 22555
tri 35386 22553 35387 22554 ne
rect 35387 22553 35635 22554
tri 35387 22552 35388 22553 ne
rect 35388 22552 35635 22553
tri 35388 22551 35389 22552 ne
rect 35389 22551 35635 22552
tri 35389 22550 35390 22551 ne
rect 35390 22550 35635 22551
tri 35390 22549 35391 22550 ne
rect 35391 22549 35635 22550
tri 35391 22548 35392 22549 ne
rect 35392 22548 35635 22549
tri 35392 22547 35393 22548 ne
rect 35393 22547 35635 22548
tri 35393 22546 35394 22547 ne
rect 35394 22546 35635 22547
tri 35394 22545 35395 22546 ne
rect 35395 22545 35635 22546
tri 35395 22544 35396 22545 ne
rect 35396 22544 35635 22545
tri 35396 22543 35397 22544 ne
rect 35397 22543 35635 22544
tri 35397 22542 35398 22543 ne
rect 35398 22542 35635 22543
tri 35398 22541 35399 22542 ne
rect 35399 22541 35635 22542
tri 35399 22540 35400 22541 ne
rect 35400 22540 35635 22541
tri 35400 22539 35401 22540 ne
rect 35401 22539 35635 22540
tri 35401 22538 35402 22539 ne
rect 35402 22538 35635 22539
tri 35402 22537 35403 22538 ne
rect 35403 22537 35635 22538
tri 35403 22536 35404 22537 ne
rect 35404 22536 35635 22537
tri 35635 22536 35680 22581 sw
rect 70802 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35404 22535 35405 22536 ne
rect 35405 22535 35680 22536
tri 35405 22534 35406 22535 ne
rect 35406 22534 35680 22535
tri 35406 22533 35407 22534 ne
rect 35407 22533 35680 22534
tri 35407 22532 35408 22533 ne
rect 35408 22532 35680 22533
tri 35408 22531 35409 22532 ne
rect 35409 22531 35680 22532
tri 35409 22530 35410 22531 ne
rect 35410 22530 35680 22531
tri 35410 22529 35411 22530 ne
rect 35411 22529 35680 22530
tri 35411 22528 35412 22529 ne
rect 35412 22528 35680 22529
tri 35412 22527 35413 22528 ne
rect 35413 22527 35680 22528
tri 35413 22526 35414 22527 ne
rect 35414 22526 35680 22527
tri 35680 22526 35690 22536 sw
tri 35414 22525 35415 22526 ne
rect 35415 22525 35690 22526
tri 35415 22524 35416 22525 ne
rect 35416 22524 35690 22525
tri 35416 22523 35417 22524 ne
rect 35417 22523 35690 22524
tri 35417 22522 35418 22523 ne
rect 35418 22522 35690 22523
tri 35418 22521 35419 22522 ne
rect 35419 22521 35690 22522
tri 35419 22520 35420 22521 ne
rect 35420 22520 35690 22521
tri 35420 22519 35421 22520 ne
rect 35421 22519 35690 22520
tri 35421 22518 35422 22519 ne
rect 35422 22518 35690 22519
tri 35422 22517 35423 22518 ne
rect 35423 22517 35690 22518
tri 35423 22516 35424 22517 ne
rect 35424 22516 35690 22517
tri 35424 22515 35425 22516 ne
rect 35425 22515 35562 22516
tri 35425 22514 35426 22515 ne
rect 35426 22514 35562 22515
tri 35426 22513 35427 22514 ne
rect 35427 22513 35562 22514
tri 35427 22512 35428 22513 ne
rect 35428 22512 35562 22513
tri 35428 22511 35429 22512 ne
rect 35429 22511 35562 22512
tri 35429 22510 35430 22511 ne
rect 35430 22510 35562 22511
tri 35430 22509 35431 22510 ne
rect 35431 22509 35562 22510
tri 35431 22508 35432 22509 ne
rect 35432 22508 35562 22509
tri 35432 22507 35433 22508 ne
rect 35433 22507 35562 22508
tri 35433 22506 35434 22507 ne
rect 35434 22506 35562 22507
tri 35434 22505 35435 22506 ne
rect 35435 22505 35562 22506
tri 35435 22504 35436 22505 ne
rect 35436 22504 35562 22505
tri 35436 22503 35437 22504 ne
rect 35437 22503 35562 22504
tri 35437 22502 35438 22503 ne
rect 35438 22502 35562 22503
tri 35438 22501 35439 22502 ne
rect 35439 22501 35562 22502
tri 35439 22500 35440 22501 ne
rect 35440 22500 35562 22501
tri 35440 22499 35441 22500 ne
rect 35441 22499 35562 22500
tri 35441 22498 35442 22499 ne
rect 35442 22498 35562 22499
tri 35442 22497 35443 22498 ne
rect 35443 22497 35562 22498
tri 35443 22496 35444 22497 ne
rect 35444 22496 35562 22497
tri 35444 22495 35445 22496 ne
rect 35445 22495 35562 22496
tri 35445 22494 35446 22495 ne
rect 35446 22494 35562 22495
tri 35446 22493 35447 22494 ne
rect 35447 22493 35562 22494
tri 35447 22492 35448 22493 ne
rect 35448 22492 35562 22493
tri 35448 22491 35449 22492 ne
rect 35449 22491 35562 22492
tri 35449 22490 35450 22491 ne
rect 35450 22490 35562 22491
tri 35450 22489 35451 22490 ne
rect 35451 22489 35562 22490
tri 35451 22488 35452 22489 ne
rect 35452 22488 35562 22489
tri 35452 22487 35453 22488 ne
rect 35453 22487 35562 22488
tri 35453 22486 35454 22487 ne
rect 35454 22486 35562 22487
tri 35454 22485 35455 22486 ne
rect 35455 22485 35562 22486
tri 35455 22484 35456 22485 ne
rect 35456 22484 35562 22485
tri 35456 22483 35457 22484 ne
rect 35457 22483 35562 22484
tri 35457 22482 35458 22483 ne
rect 35458 22482 35562 22483
tri 35458 22481 35459 22482 ne
rect 35459 22481 35562 22482
tri 35459 22436 35504 22481 ne
rect 35504 22470 35562 22481
rect 35608 22481 35690 22516
tri 35690 22481 35735 22526 sw
rect 70802 22484 71000 22542
rect 35608 22470 35735 22481
rect 35504 22436 35735 22470
tri 35735 22436 35780 22481 sw
rect 70802 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35504 22391 35549 22436 ne
rect 35549 22391 35780 22436
tri 35780 22391 35825 22436 sw
tri 35549 22346 35594 22391 ne
rect 35594 22384 35825 22391
rect 35594 22346 35694 22384
tri 35594 22345 35595 22346 ne
rect 35595 22345 35694 22346
tri 35595 22344 35596 22345 ne
rect 35596 22344 35694 22345
tri 35596 22343 35597 22344 ne
rect 35597 22343 35694 22344
tri 35597 22342 35598 22343 ne
rect 35598 22342 35694 22343
tri 35598 22341 35599 22342 ne
rect 35599 22341 35694 22342
tri 35599 22340 35600 22341 ne
rect 35600 22340 35694 22341
tri 35600 22339 35601 22340 ne
rect 35601 22339 35694 22340
tri 35601 22338 35602 22339 ne
rect 35602 22338 35694 22339
rect 35740 22350 35825 22384
tri 35825 22350 35866 22391 sw
rect 70802 22380 71000 22438
rect 35740 22338 35866 22350
tri 35602 22337 35603 22338 ne
rect 35603 22337 35866 22338
tri 35603 22336 35604 22337 ne
rect 35604 22336 35866 22337
tri 35604 22335 35605 22336 ne
rect 35605 22335 35866 22336
tri 35605 22334 35606 22335 ne
rect 35606 22334 35866 22335
tri 35606 22333 35607 22334 ne
rect 35607 22333 35866 22334
tri 35607 22332 35608 22333 ne
rect 35608 22332 35866 22333
tri 35608 22331 35609 22332 ne
rect 35609 22331 35866 22332
tri 35609 22330 35610 22331 ne
rect 35610 22330 35866 22331
tri 35610 22329 35611 22330 ne
rect 35611 22329 35866 22330
tri 35611 22328 35612 22329 ne
rect 35612 22328 35866 22329
tri 35612 22327 35613 22328 ne
rect 35613 22327 35866 22328
tri 35613 22326 35614 22327 ne
rect 35614 22326 35866 22327
tri 35614 22325 35615 22326 ne
rect 35615 22325 35866 22326
tri 35615 22324 35616 22325 ne
rect 35616 22324 35866 22325
tri 35616 22323 35617 22324 ne
rect 35617 22323 35866 22324
tri 35617 22322 35618 22323 ne
rect 35618 22322 35866 22323
tri 35618 22321 35619 22322 ne
rect 35619 22321 35866 22322
tri 35619 22320 35620 22321 ne
rect 35620 22320 35866 22321
tri 35620 22319 35621 22320 ne
rect 35621 22319 35866 22320
tri 35621 22318 35622 22319 ne
rect 35622 22318 35866 22319
tri 35622 22317 35623 22318 ne
rect 35623 22317 35866 22318
tri 35623 22316 35624 22317 ne
rect 35624 22316 35866 22317
tri 35624 22315 35625 22316 ne
rect 35625 22315 35866 22316
tri 35625 22314 35626 22315 ne
rect 35626 22314 35866 22315
tri 35626 22313 35627 22314 ne
rect 35627 22313 35866 22314
tri 35627 22312 35628 22313 ne
rect 35628 22312 35866 22313
tri 35628 22311 35629 22312 ne
rect 35629 22311 35866 22312
tri 35629 22310 35630 22311 ne
rect 35630 22310 35866 22311
tri 35630 22309 35631 22310 ne
rect 35631 22309 35866 22310
tri 35631 22308 35632 22309 ne
rect 35632 22308 35866 22309
tri 35632 22307 35633 22308 ne
rect 35633 22307 35866 22308
tri 35633 22306 35634 22307 ne
rect 35634 22306 35866 22307
tri 35634 22305 35635 22306 ne
rect 35635 22305 35866 22306
tri 35866 22305 35911 22350 sw
rect 70802 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35635 22304 35636 22305 ne
rect 35636 22304 35911 22305
tri 35636 22303 35637 22304 ne
rect 35637 22303 35911 22304
tri 35637 22302 35638 22303 ne
rect 35638 22302 35911 22303
tri 35638 22301 35639 22302 ne
rect 35639 22301 35911 22302
tri 35639 22300 35640 22301 ne
rect 35640 22300 35911 22301
tri 35640 22299 35641 22300 ne
rect 35641 22299 35911 22300
tri 35641 22298 35642 22299 ne
rect 35642 22298 35911 22299
tri 35642 22297 35643 22298 ne
rect 35643 22297 35911 22298
tri 35643 22296 35644 22297 ne
rect 35644 22296 35911 22297
tri 35644 22295 35645 22296 ne
rect 35645 22295 35911 22296
tri 35645 22294 35646 22295 ne
rect 35646 22294 35911 22295
tri 35646 22293 35647 22294 ne
rect 35647 22293 35911 22294
tri 35647 22292 35648 22293 ne
rect 35648 22292 35911 22293
tri 35648 22291 35649 22292 ne
rect 35649 22291 35911 22292
tri 35649 22290 35650 22291 ne
rect 35650 22290 35911 22291
tri 35650 22289 35651 22290 ne
rect 35651 22289 35911 22290
tri 35651 22288 35652 22289 ne
rect 35652 22288 35911 22289
tri 35652 22287 35653 22288 ne
rect 35653 22287 35911 22288
tri 35653 22286 35654 22287 ne
rect 35654 22286 35911 22287
tri 35654 22285 35655 22286 ne
rect 35655 22285 35911 22286
tri 35655 22284 35656 22285 ne
rect 35656 22284 35911 22285
tri 35656 22283 35657 22284 ne
rect 35657 22283 35911 22284
tri 35657 22282 35658 22283 ne
rect 35658 22282 35911 22283
tri 35658 22281 35659 22282 ne
rect 35659 22281 35911 22282
tri 35659 22280 35660 22281 ne
rect 35660 22280 35911 22281
tri 35660 22279 35661 22280 ne
rect 35661 22279 35911 22280
tri 35661 22278 35662 22279 ne
rect 35662 22278 35911 22279
tri 35662 22277 35663 22278 ne
rect 35663 22277 35911 22278
tri 35663 22276 35664 22277 ne
rect 35664 22276 35911 22277
tri 35664 22275 35665 22276 ne
rect 35665 22275 35911 22276
tri 35665 22274 35666 22275 ne
rect 35666 22274 35911 22275
tri 35666 22273 35667 22274 ne
rect 35667 22273 35911 22274
tri 35667 22272 35668 22273 ne
rect 35668 22272 35911 22273
tri 35668 22271 35669 22272 ne
rect 35669 22271 35911 22272
tri 35669 22270 35670 22271 ne
rect 35670 22270 35911 22271
tri 35670 22269 35671 22270 ne
rect 35671 22269 35911 22270
tri 35671 22268 35672 22269 ne
rect 35672 22268 35911 22269
tri 35672 22267 35673 22268 ne
rect 35673 22267 35911 22268
tri 35673 22266 35674 22267 ne
rect 35674 22266 35911 22267
tri 35674 22265 35675 22266 ne
rect 35675 22265 35911 22266
tri 35675 22264 35676 22265 ne
rect 35676 22264 35911 22265
tri 35676 22263 35677 22264 ne
rect 35677 22263 35911 22264
tri 35677 22262 35678 22263 ne
rect 35678 22262 35911 22263
tri 35678 22261 35679 22262 ne
rect 35679 22261 35911 22262
tri 35679 22260 35680 22261 ne
rect 35680 22260 35911 22261
tri 35911 22260 35956 22305 sw
rect 70802 22276 71000 22334
tri 35680 22259 35681 22260 ne
rect 35681 22259 35956 22260
tri 35681 22258 35682 22259 ne
rect 35682 22258 35956 22259
tri 35682 22257 35683 22258 ne
rect 35683 22257 35956 22258
tri 35683 22256 35684 22257 ne
rect 35684 22256 35956 22257
tri 35684 22255 35685 22256 ne
rect 35685 22255 35956 22256
tri 35685 22254 35686 22255 ne
rect 35686 22254 35956 22255
tri 35686 22253 35687 22254 ne
rect 35687 22253 35956 22254
tri 35687 22252 35688 22253 ne
rect 35688 22252 35956 22253
tri 35688 22251 35689 22252 ne
rect 35689 22251 35826 22252
tri 35689 22250 35690 22251 ne
rect 35690 22250 35826 22251
tri 35690 22249 35691 22250 ne
rect 35691 22249 35826 22250
tri 35691 22248 35692 22249 ne
rect 35692 22248 35826 22249
tri 35692 22247 35693 22248 ne
rect 35693 22247 35826 22248
tri 35693 22246 35694 22247 ne
rect 35694 22246 35826 22247
tri 35694 22245 35695 22246 ne
rect 35695 22245 35826 22246
tri 35695 22244 35696 22245 ne
rect 35696 22244 35826 22245
tri 35696 22243 35697 22244 ne
rect 35697 22243 35826 22244
tri 35697 22242 35698 22243 ne
rect 35698 22242 35826 22243
tri 35698 22241 35699 22242 ne
rect 35699 22241 35826 22242
tri 35699 22240 35700 22241 ne
rect 35700 22240 35826 22241
tri 35700 22239 35701 22240 ne
rect 35701 22239 35826 22240
tri 35701 22238 35702 22239 ne
rect 35702 22238 35826 22239
tri 35702 22237 35703 22238 ne
rect 35703 22237 35826 22238
tri 35703 22236 35704 22237 ne
rect 35704 22236 35826 22237
tri 35704 22235 35705 22236 ne
rect 35705 22235 35826 22236
tri 35705 22234 35706 22235 ne
rect 35706 22234 35826 22235
tri 35706 22233 35707 22234 ne
rect 35707 22233 35826 22234
tri 35707 22232 35708 22233 ne
rect 35708 22232 35826 22233
tri 35708 22231 35709 22232 ne
rect 35709 22231 35826 22232
tri 35709 22230 35710 22231 ne
rect 35710 22230 35826 22231
tri 35710 22229 35711 22230 ne
rect 35711 22229 35826 22230
tri 35711 22228 35712 22229 ne
rect 35712 22228 35826 22229
tri 35712 22227 35713 22228 ne
rect 35713 22227 35826 22228
tri 35713 22226 35714 22227 ne
rect 35714 22226 35826 22227
tri 35714 22225 35715 22226 ne
rect 35715 22225 35826 22226
tri 35715 22224 35716 22225 ne
rect 35716 22224 35826 22225
tri 35716 22223 35717 22224 ne
rect 35717 22223 35826 22224
tri 35717 22222 35718 22223 ne
rect 35718 22222 35826 22223
tri 35718 22221 35719 22222 ne
rect 35719 22221 35826 22222
tri 35719 22220 35720 22221 ne
rect 35720 22220 35826 22221
tri 35720 22219 35721 22220 ne
rect 35721 22219 35826 22220
tri 35721 22218 35722 22219 ne
rect 35722 22218 35826 22219
tri 35722 22217 35723 22218 ne
rect 35723 22217 35826 22218
tri 35723 22216 35724 22217 ne
rect 35724 22216 35826 22217
tri 35724 22215 35725 22216 ne
rect 35725 22215 35826 22216
tri 35725 22214 35726 22215 ne
rect 35726 22214 35826 22215
tri 35726 22213 35727 22214 ne
rect 35727 22213 35826 22214
tri 35727 22212 35728 22213 ne
rect 35728 22212 35826 22213
tri 35728 22211 35729 22212 ne
rect 35729 22211 35826 22212
tri 35729 22210 35730 22211 ne
rect 35730 22210 35826 22211
tri 35730 22209 35731 22210 ne
rect 35731 22209 35826 22210
tri 35731 22208 35732 22209 ne
rect 35732 22208 35826 22209
tri 35732 22207 35733 22208 ne
rect 35733 22207 35826 22208
tri 35733 22206 35734 22207 ne
rect 35734 22206 35826 22207
rect 35872 22215 35956 22252
tri 35956 22215 36001 22260 sw
rect 70802 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22206 36001 22215
tri 35734 22205 35735 22206 ne
rect 35735 22205 36001 22206
tri 36001 22205 36011 22215 sw
tri 35735 22160 35780 22205 ne
rect 35780 22170 36011 22205
tri 36011 22170 36046 22205 sw
rect 70802 22172 71000 22230
rect 35780 22160 36046 22170
tri 35780 22123 35817 22160 ne
rect 35817 22125 36046 22160
tri 36046 22125 36091 22170 sw
rect 70802 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 35817 22123 36091 22125
tri 35817 22078 35862 22123 ne
rect 35862 22120 36091 22123
rect 35862 22078 35958 22120
tri 35862 22072 35868 22078 ne
rect 35868 22074 35958 22078
rect 36004 22080 36091 22120
tri 36091 22080 36136 22125 sw
rect 36004 22074 36136 22080
rect 35868 22072 36136 22074
tri 35868 22071 35869 22072 ne
rect 35869 22071 36136 22072
tri 35869 22070 35870 22071 ne
rect 35870 22070 36136 22071
tri 35870 22069 35871 22070 ne
rect 35871 22069 36136 22070
tri 35871 22068 35872 22069 ne
rect 35872 22068 36136 22069
tri 35872 22067 35873 22068 ne
rect 35873 22067 36136 22068
tri 35873 22066 35874 22067 ne
rect 35874 22066 36136 22067
tri 35874 22065 35875 22066 ne
rect 35875 22065 36136 22066
tri 35875 22064 35876 22065 ne
rect 35876 22064 36136 22065
tri 36136 22064 36152 22080 sw
rect 70802 22068 71000 22126
tri 35876 22063 35877 22064 ne
rect 35877 22063 36152 22064
tri 35877 22062 35878 22063 ne
rect 35878 22062 36152 22063
tri 35878 22061 35879 22062 ne
rect 35879 22061 36152 22062
tri 35879 22060 35880 22061 ne
rect 35880 22060 36152 22061
tri 35880 22059 35881 22060 ne
rect 35881 22059 36152 22060
tri 35881 22058 35882 22059 ne
rect 35882 22058 36152 22059
tri 35882 22057 35883 22058 ne
rect 35883 22057 36152 22058
tri 35883 22056 35884 22057 ne
rect 35884 22056 36152 22057
tri 35884 22055 35885 22056 ne
rect 35885 22055 36152 22056
tri 35885 22054 35886 22055 ne
rect 35886 22054 36152 22055
tri 35886 22053 35887 22054 ne
rect 35887 22053 36152 22054
tri 35887 22052 35888 22053 ne
rect 35888 22052 36152 22053
tri 35888 22051 35889 22052 ne
rect 35889 22051 36152 22052
tri 35889 22050 35890 22051 ne
rect 35890 22050 36152 22051
tri 35890 22049 35891 22050 ne
rect 35891 22049 36152 22050
tri 35891 22048 35892 22049 ne
rect 35892 22048 36152 22049
tri 35892 22047 35893 22048 ne
rect 35893 22047 36152 22048
tri 35893 22046 35894 22047 ne
rect 35894 22046 36152 22047
tri 35894 22045 35895 22046 ne
rect 35895 22045 36152 22046
tri 35895 22044 35896 22045 ne
rect 35896 22044 36152 22045
tri 35896 22043 35897 22044 ne
rect 35897 22043 36152 22044
tri 35897 22042 35898 22043 ne
rect 35898 22042 36152 22043
tri 35898 22041 35899 22042 ne
rect 35899 22041 36152 22042
tri 35899 22040 35900 22041 ne
rect 35900 22040 36152 22041
tri 35900 22039 35901 22040 ne
rect 35901 22039 36152 22040
tri 35901 22038 35902 22039 ne
rect 35902 22038 36152 22039
tri 35902 22037 35903 22038 ne
rect 35903 22037 36152 22038
tri 35903 22036 35904 22037 ne
rect 35904 22036 36152 22037
tri 35904 22035 35905 22036 ne
rect 35905 22035 36152 22036
tri 35905 22034 35906 22035 ne
rect 35906 22034 36152 22035
tri 35906 22033 35907 22034 ne
rect 35907 22033 36152 22034
tri 35907 22032 35908 22033 ne
rect 35908 22032 36152 22033
tri 35908 22031 35909 22032 ne
rect 35909 22031 36152 22032
tri 35909 22030 35910 22031 ne
rect 35910 22030 36152 22031
tri 35910 22029 35911 22030 ne
rect 35911 22029 36152 22030
tri 35911 22028 35912 22029 ne
rect 35912 22028 36152 22029
tri 35912 22027 35913 22028 ne
rect 35913 22027 36152 22028
tri 35913 22026 35914 22027 ne
rect 35914 22026 36152 22027
tri 35914 22025 35915 22026 ne
rect 35915 22025 36152 22026
tri 35915 22024 35916 22025 ne
rect 35916 22024 36152 22025
tri 35916 22023 35917 22024 ne
rect 35917 22023 36152 22024
tri 35917 22022 35918 22023 ne
rect 35918 22022 36152 22023
tri 35918 22021 35919 22022 ne
rect 35919 22021 36152 22022
tri 35919 22020 35920 22021 ne
rect 35920 22020 36152 22021
tri 35920 22019 35921 22020 ne
rect 35921 22019 36152 22020
tri 36152 22019 36197 22064 sw
rect 70802 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35921 22018 35922 22019 ne
rect 35922 22018 36197 22019
tri 35922 22017 35923 22018 ne
rect 35923 22017 36197 22018
tri 35923 22016 35924 22017 ne
rect 35924 22016 36197 22017
tri 35924 22015 35925 22016 ne
rect 35925 22015 36197 22016
tri 35925 22014 35926 22015 ne
rect 35926 22014 36197 22015
tri 35926 22013 35927 22014 ne
rect 35927 22013 36197 22014
tri 35927 22012 35928 22013 ne
rect 35928 22012 36197 22013
tri 35928 22011 35929 22012 ne
rect 35929 22011 36197 22012
tri 35929 22010 35930 22011 ne
rect 35930 22010 36197 22011
tri 35930 22009 35931 22010 ne
rect 35931 22009 36197 22010
tri 35931 22008 35932 22009 ne
rect 35932 22008 36197 22009
tri 35932 22007 35933 22008 ne
rect 35933 22007 36197 22008
tri 35933 22006 35934 22007 ne
rect 35934 22006 36197 22007
tri 35934 22005 35935 22006 ne
rect 35935 22005 36197 22006
tri 35935 22004 35936 22005 ne
rect 35936 22004 36197 22005
tri 35936 22003 35937 22004 ne
rect 35937 22003 36197 22004
tri 35937 22002 35938 22003 ne
rect 35938 22002 36197 22003
tri 35938 22001 35939 22002 ne
rect 35939 22001 36197 22002
tri 35939 22000 35940 22001 ne
rect 35940 22000 36197 22001
tri 35940 21999 35941 22000 ne
rect 35941 21999 36197 22000
tri 35941 21998 35942 21999 ne
rect 35942 21998 36197 21999
tri 35942 21997 35943 21998 ne
rect 35943 21997 36197 21998
tri 35943 21996 35944 21997 ne
rect 35944 21996 36197 21997
tri 35944 21995 35945 21996 ne
rect 35945 21995 36197 21996
tri 35945 21994 35946 21995 ne
rect 35946 21994 36197 21995
tri 35946 21993 35947 21994 ne
rect 35947 21993 36197 21994
tri 35947 21992 35948 21993 ne
rect 35948 21992 36197 21993
tri 35948 21991 35949 21992 ne
rect 35949 21991 36197 21992
tri 35949 21990 35950 21991 ne
rect 35950 21990 36197 21991
tri 35950 21989 35951 21990 ne
rect 35951 21989 36197 21990
tri 35951 21988 35952 21989 ne
rect 35952 21988 36197 21989
tri 35952 21987 35953 21988 ne
rect 35953 21987 36090 21988
tri 35953 21986 35954 21987 ne
rect 35954 21986 36090 21987
tri 35954 21985 35955 21986 ne
rect 35955 21985 36090 21986
tri 35955 21984 35956 21985 ne
rect 35956 21984 36090 21985
tri 35956 21983 35957 21984 ne
rect 35957 21983 36090 21984
tri 35957 21982 35958 21983 ne
rect 35958 21982 36090 21983
tri 35958 21981 35959 21982 ne
rect 35959 21981 36090 21982
tri 35959 21980 35960 21981 ne
rect 35960 21980 36090 21981
tri 35960 21979 35961 21980 ne
rect 35961 21979 36090 21980
tri 35961 21978 35962 21979 ne
rect 35962 21978 36090 21979
tri 35962 21977 35963 21978 ne
rect 35963 21977 36090 21978
tri 35963 21976 35964 21977 ne
rect 35964 21976 36090 21977
tri 35964 21975 35965 21976 ne
rect 35965 21975 36090 21976
tri 35965 21974 35966 21975 ne
rect 35966 21974 36090 21975
tri 35966 21973 35967 21974 ne
rect 35967 21973 36090 21974
tri 35967 21972 35968 21973 ne
rect 35968 21972 36090 21973
tri 35968 21971 35969 21972 ne
rect 35969 21971 36090 21972
tri 35969 21970 35970 21971 ne
rect 35970 21970 36090 21971
tri 35970 21969 35971 21970 ne
rect 35971 21969 36090 21970
tri 35971 21968 35972 21969 ne
rect 35972 21968 36090 21969
tri 35972 21967 35973 21968 ne
rect 35973 21967 36090 21968
tri 35973 21966 35974 21967 ne
rect 35974 21966 36090 21967
tri 35974 21965 35975 21966 ne
rect 35975 21965 36090 21966
tri 35975 21964 35976 21965 ne
rect 35976 21964 36090 21965
tri 35976 21963 35977 21964 ne
rect 35977 21963 36090 21964
tri 35977 21962 35978 21963 ne
rect 35978 21962 36090 21963
tri 35978 21961 35979 21962 ne
rect 35979 21961 36090 21962
tri 35979 21960 35980 21961 ne
rect 35980 21960 36090 21961
tri 35980 21959 35981 21960 ne
rect 35981 21959 36090 21960
tri 35981 21958 35982 21959 ne
rect 35982 21958 36090 21959
tri 35982 21957 35983 21958 ne
rect 35983 21957 36090 21958
tri 35983 21956 35984 21957 ne
rect 35984 21956 36090 21957
tri 35984 21955 35985 21956 ne
rect 35985 21955 36090 21956
tri 35985 21954 35986 21955 ne
rect 35986 21954 36090 21955
tri 35986 21953 35987 21954 ne
rect 35987 21953 36090 21954
tri 35987 21952 35988 21953 ne
rect 35988 21952 36090 21953
tri 35988 21951 35989 21952 ne
rect 35989 21951 36090 21952
tri 35989 21950 35990 21951 ne
rect 35990 21950 36090 21951
tri 35990 21949 35991 21950 ne
rect 35991 21949 36090 21950
tri 35991 21948 35992 21949 ne
rect 35992 21948 36090 21949
tri 35992 21947 35993 21948 ne
rect 35993 21947 36090 21948
tri 35993 21946 35994 21947 ne
rect 35994 21946 36090 21947
tri 35994 21945 35995 21946 ne
rect 35995 21945 36090 21946
tri 35995 21944 35996 21945 ne
rect 35996 21944 36090 21945
tri 35996 21943 35997 21944 ne
rect 35997 21943 36090 21944
tri 35997 21942 35998 21943 ne
rect 35998 21942 36090 21943
rect 36136 21974 36197 21988
tri 36197 21974 36242 22019 sw
rect 36136 21942 36242 21974
tri 35998 21941 35999 21942 ne
rect 35999 21941 36242 21942
tri 35999 21940 36000 21941 ne
rect 36000 21940 36242 21941
tri 36000 21939 36001 21940 ne
rect 36001 21939 36242 21940
tri 36001 21938 36002 21939 ne
rect 36002 21938 36242 21939
tri 36002 21937 36003 21938 ne
rect 36003 21937 36242 21938
tri 36003 21936 36004 21937 ne
rect 36004 21936 36242 21937
tri 36004 21935 36005 21936 ne
rect 36005 21935 36242 21936
tri 36005 21934 36006 21935 ne
rect 36006 21934 36242 21935
tri 36006 21933 36007 21934 ne
rect 36007 21933 36242 21934
tri 36007 21932 36008 21933 ne
rect 36008 21932 36242 21933
tri 36008 21931 36009 21932 ne
rect 36009 21931 36242 21932
tri 36009 21930 36010 21931 ne
rect 36010 21930 36242 21931
tri 36010 21929 36011 21930 ne
rect 36011 21929 36242 21930
tri 36242 21929 36287 21974 sw
rect 70802 21964 71000 22022
tri 36011 21894 36046 21929 ne
rect 36046 21894 36287 21929
tri 36287 21894 36322 21929 sw
rect 70802 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
tri 36046 21884 36056 21894 ne
rect 36056 21884 36322 21894
tri 36056 21849 36091 21884 ne
rect 36091 21856 36322 21884
rect 36091 21849 36222 21856
tri 36091 21804 36136 21849 ne
rect 36136 21810 36222 21849
rect 36268 21849 36322 21856
tri 36322 21849 36367 21894 sw
rect 70802 21860 71000 21918
rect 36268 21810 36367 21849
rect 36136 21804 36367 21810
tri 36367 21804 36412 21849 sw
rect 70802 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
tri 36136 21797 36143 21804 ne
rect 36143 21797 36412 21804
tri 36143 21796 36144 21797 ne
rect 36144 21796 36412 21797
tri 36144 21795 36145 21796 ne
rect 36145 21795 36412 21796
tri 36145 21794 36146 21795 ne
rect 36146 21794 36412 21795
tri 36146 21793 36147 21794 ne
rect 36147 21793 36412 21794
tri 36147 21792 36148 21793 ne
rect 36148 21792 36412 21793
tri 36148 21791 36149 21792 ne
rect 36149 21791 36412 21792
tri 36149 21790 36150 21791 ne
rect 36150 21790 36412 21791
tri 36150 21789 36151 21790 ne
rect 36151 21789 36412 21790
tri 36151 21788 36152 21789 ne
rect 36152 21788 36412 21789
tri 36152 21787 36153 21788 ne
rect 36153 21787 36412 21788
tri 36153 21786 36154 21787 ne
rect 36154 21786 36412 21787
tri 36154 21785 36155 21786 ne
rect 36155 21785 36412 21786
tri 36155 21784 36156 21785 ne
rect 36156 21784 36412 21785
tri 36156 21783 36157 21784 ne
rect 36157 21783 36412 21784
tri 36157 21782 36158 21783 ne
rect 36158 21782 36412 21783
tri 36158 21781 36159 21782 ne
rect 36159 21781 36412 21782
tri 36159 21780 36160 21781 ne
rect 36160 21780 36412 21781
tri 36160 21779 36161 21780 ne
rect 36161 21779 36412 21780
tri 36161 21778 36162 21779 ne
rect 36162 21778 36412 21779
tri 36162 21777 36163 21778 ne
rect 36163 21777 36412 21778
tri 36163 21776 36164 21777 ne
rect 36164 21776 36412 21777
tri 36164 21775 36165 21776 ne
rect 36165 21775 36412 21776
tri 36165 21774 36166 21775 ne
rect 36166 21774 36412 21775
tri 36166 21773 36167 21774 ne
rect 36167 21773 36412 21774
tri 36167 21772 36168 21773 ne
rect 36168 21772 36412 21773
tri 36168 21771 36169 21772 ne
rect 36169 21771 36412 21772
tri 36169 21770 36170 21771 ne
rect 36170 21770 36412 21771
tri 36170 21769 36171 21770 ne
rect 36171 21769 36412 21770
tri 36171 21768 36172 21769 ne
rect 36172 21768 36412 21769
tri 36172 21767 36173 21768 ne
rect 36173 21767 36412 21768
tri 36173 21766 36174 21767 ne
rect 36174 21766 36412 21767
tri 36174 21765 36175 21766 ne
rect 36175 21765 36412 21766
tri 36175 21764 36176 21765 ne
rect 36176 21764 36412 21765
tri 36176 21763 36177 21764 ne
rect 36177 21763 36412 21764
tri 36177 21762 36178 21763 ne
rect 36178 21762 36412 21763
tri 36178 21761 36179 21762 ne
rect 36179 21761 36412 21762
tri 36179 21760 36180 21761 ne
rect 36180 21760 36412 21761
tri 36180 21759 36181 21760 ne
rect 36181 21759 36412 21760
tri 36412 21759 36457 21804 sw
tri 36181 21758 36182 21759 ne
rect 36182 21758 36457 21759
tri 36182 21757 36183 21758 ne
rect 36183 21757 36457 21758
tri 36183 21756 36184 21757 ne
rect 36184 21756 36457 21757
tri 36184 21755 36185 21756 ne
rect 36185 21755 36457 21756
tri 36185 21754 36186 21755 ne
rect 36186 21754 36457 21755
tri 36186 21753 36187 21754 ne
rect 36187 21753 36457 21754
tri 36187 21752 36188 21753 ne
rect 36188 21752 36457 21753
tri 36188 21751 36189 21752 ne
rect 36189 21751 36457 21752
tri 36189 21750 36190 21751 ne
rect 36190 21750 36457 21751
tri 36190 21749 36191 21750 ne
rect 36191 21749 36457 21750
tri 36191 21748 36192 21749 ne
rect 36192 21748 36457 21749
tri 36192 21747 36193 21748 ne
rect 36193 21747 36457 21748
tri 36193 21746 36194 21747 ne
rect 36194 21746 36457 21747
tri 36194 21745 36195 21746 ne
rect 36195 21745 36457 21746
tri 36195 21744 36196 21745 ne
rect 36196 21744 36457 21745
tri 36196 21743 36197 21744 ne
rect 36197 21743 36457 21744
tri 36457 21743 36473 21759 sw
rect 70802 21756 71000 21814
tri 36197 21742 36198 21743 ne
rect 36198 21742 36473 21743
tri 36198 21741 36199 21742 ne
rect 36199 21741 36473 21742
tri 36199 21740 36200 21741 ne
rect 36200 21740 36473 21741
tri 36200 21739 36201 21740 ne
rect 36201 21739 36473 21740
tri 36201 21738 36202 21739 ne
rect 36202 21738 36473 21739
tri 36202 21737 36203 21738 ne
rect 36203 21737 36473 21738
tri 36203 21736 36204 21737 ne
rect 36204 21736 36473 21737
tri 36204 21735 36205 21736 ne
rect 36205 21735 36473 21736
tri 36205 21734 36206 21735 ne
rect 36206 21734 36473 21735
tri 36206 21733 36207 21734 ne
rect 36207 21733 36473 21734
tri 36207 21732 36208 21733 ne
rect 36208 21732 36473 21733
tri 36208 21731 36209 21732 ne
rect 36209 21731 36473 21732
tri 36209 21730 36210 21731 ne
rect 36210 21730 36473 21731
tri 36210 21729 36211 21730 ne
rect 36211 21729 36473 21730
tri 36211 21728 36212 21729 ne
rect 36212 21728 36473 21729
tri 36212 21727 36213 21728 ne
rect 36213 21727 36473 21728
tri 36213 21726 36214 21727 ne
rect 36214 21726 36473 21727
tri 36214 21725 36215 21726 ne
rect 36215 21725 36473 21726
tri 36215 21724 36216 21725 ne
rect 36216 21724 36473 21725
tri 36216 21723 36217 21724 ne
rect 36217 21723 36354 21724
tri 36217 21722 36218 21723 ne
rect 36218 21722 36354 21723
tri 36218 21721 36219 21722 ne
rect 36219 21721 36354 21722
tri 36219 21720 36220 21721 ne
rect 36220 21720 36354 21721
tri 36220 21719 36221 21720 ne
rect 36221 21719 36354 21720
tri 36221 21718 36222 21719 ne
rect 36222 21718 36354 21719
tri 36222 21717 36223 21718 ne
rect 36223 21717 36354 21718
tri 36223 21716 36224 21717 ne
rect 36224 21716 36354 21717
tri 36224 21715 36225 21716 ne
rect 36225 21715 36354 21716
tri 36225 21714 36226 21715 ne
rect 36226 21714 36354 21715
tri 36226 21713 36227 21714 ne
rect 36227 21713 36354 21714
tri 36227 21712 36228 21713 ne
rect 36228 21712 36354 21713
tri 36228 21711 36229 21712 ne
rect 36229 21711 36354 21712
tri 36229 21710 36230 21711 ne
rect 36230 21710 36354 21711
tri 36230 21709 36231 21710 ne
rect 36231 21709 36354 21710
tri 36231 21708 36232 21709 ne
rect 36232 21708 36354 21709
tri 36232 21707 36233 21708 ne
rect 36233 21707 36354 21708
tri 36233 21706 36234 21707 ne
rect 36234 21706 36354 21707
tri 36234 21705 36235 21706 ne
rect 36235 21705 36354 21706
tri 36235 21704 36236 21705 ne
rect 36236 21704 36354 21705
tri 36236 21703 36237 21704 ne
rect 36237 21703 36354 21704
tri 36237 21702 36238 21703 ne
rect 36238 21702 36354 21703
tri 36238 21701 36239 21702 ne
rect 36239 21701 36354 21702
tri 36239 21700 36240 21701 ne
rect 36240 21700 36354 21701
tri 36240 21699 36241 21700 ne
rect 36241 21699 36354 21700
tri 36241 21698 36242 21699 ne
rect 36242 21698 36354 21699
tri 36242 21697 36243 21698 ne
rect 36243 21697 36354 21698
tri 36243 21696 36244 21697 ne
rect 36244 21696 36354 21697
tri 36244 21695 36245 21696 ne
rect 36245 21695 36354 21696
tri 36245 21694 36246 21695 ne
rect 36246 21694 36354 21695
tri 36246 21693 36247 21694 ne
rect 36247 21693 36354 21694
tri 36247 21692 36248 21693 ne
rect 36248 21692 36354 21693
tri 36248 21691 36249 21692 ne
rect 36249 21691 36354 21692
tri 36249 21690 36250 21691 ne
rect 36250 21690 36354 21691
tri 36250 21689 36251 21690 ne
rect 36251 21689 36354 21690
tri 36251 21688 36252 21689 ne
rect 36252 21688 36354 21689
tri 36252 21687 36253 21688 ne
rect 36253 21687 36354 21688
tri 36253 21686 36254 21687 ne
rect 36254 21686 36354 21687
tri 36254 21685 36255 21686 ne
rect 36255 21685 36354 21686
tri 36255 21684 36256 21685 ne
rect 36256 21684 36354 21685
tri 36256 21683 36257 21684 ne
rect 36257 21683 36354 21684
tri 36257 21682 36258 21683 ne
rect 36258 21682 36354 21683
tri 36258 21681 36259 21682 ne
rect 36259 21681 36354 21682
tri 36259 21680 36260 21681 ne
rect 36260 21680 36354 21681
tri 36260 21679 36261 21680 ne
rect 36261 21679 36354 21680
tri 36261 21678 36262 21679 ne
rect 36262 21678 36354 21679
rect 36400 21698 36473 21724
tri 36473 21698 36518 21743 sw
rect 70802 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 36400 21678 36518 21698
tri 36262 21677 36263 21678 ne
rect 36263 21677 36518 21678
tri 36263 21676 36264 21677 ne
rect 36264 21676 36518 21677
tri 36264 21675 36265 21676 ne
rect 36265 21675 36518 21676
tri 36265 21674 36266 21675 ne
rect 36266 21674 36518 21675
tri 36266 21673 36267 21674 ne
rect 36267 21673 36518 21674
tri 36267 21672 36268 21673 ne
rect 36268 21672 36518 21673
tri 36268 21671 36269 21672 ne
rect 36269 21671 36518 21672
tri 36269 21670 36270 21671 ne
rect 36270 21670 36518 21671
tri 36270 21669 36271 21670 ne
rect 36271 21669 36518 21670
tri 36271 21668 36272 21669 ne
rect 36272 21668 36518 21669
tri 36272 21667 36273 21668 ne
rect 36273 21667 36518 21668
tri 36273 21666 36274 21667 ne
rect 36274 21666 36518 21667
tri 36274 21665 36275 21666 ne
rect 36275 21665 36518 21666
tri 36275 21664 36276 21665 ne
rect 36276 21664 36518 21665
tri 36276 21663 36277 21664 ne
rect 36277 21663 36518 21664
tri 36277 21662 36278 21663 ne
rect 36278 21662 36518 21663
tri 36278 21661 36279 21662 ne
rect 36279 21661 36518 21662
tri 36279 21660 36280 21661 ne
rect 36280 21660 36518 21661
tri 36280 21659 36281 21660 ne
rect 36281 21659 36518 21660
tri 36281 21658 36282 21659 ne
rect 36282 21658 36518 21659
tri 36282 21657 36283 21658 ne
rect 36283 21657 36518 21658
tri 36283 21656 36284 21657 ne
rect 36284 21656 36518 21657
tri 36284 21655 36285 21656 ne
rect 36285 21655 36518 21656
tri 36285 21654 36286 21655 ne
rect 36286 21654 36518 21655
tri 36286 21653 36287 21654 ne
rect 36287 21653 36518 21654
tri 36518 21653 36563 21698 sw
tri 36287 21608 36332 21653 ne
rect 36332 21608 36563 21653
tri 36563 21608 36608 21653 sw
rect 70802 21652 71000 21710
tri 36332 21563 36377 21608 ne
rect 36377 21592 36608 21608
rect 36377 21563 36486 21592
tri 36377 21528 36412 21563 ne
rect 36412 21546 36486 21563
rect 36532 21573 36608 21592
tri 36608 21573 36643 21608 sw
rect 70802 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 36532 21546 36643 21573
rect 36412 21528 36643 21546
tri 36643 21528 36688 21573 sw
rect 70802 21548 71000 21606
tri 36412 21523 36417 21528 ne
rect 36417 21523 36688 21528
tri 36417 21522 36418 21523 ne
rect 36418 21522 36688 21523
tri 36418 21521 36419 21522 ne
rect 36419 21521 36688 21522
tri 36419 21520 36420 21521 ne
rect 36420 21520 36688 21521
tri 36420 21519 36421 21520 ne
rect 36421 21519 36688 21520
tri 36421 21518 36422 21519 ne
rect 36422 21518 36688 21519
tri 36422 21517 36423 21518 ne
rect 36423 21517 36688 21518
tri 36423 21516 36424 21517 ne
rect 36424 21516 36688 21517
tri 36424 21515 36425 21516 ne
rect 36425 21515 36688 21516
tri 36425 21514 36426 21515 ne
rect 36426 21514 36688 21515
tri 36426 21513 36427 21514 ne
rect 36427 21513 36688 21514
tri 36427 21512 36428 21513 ne
rect 36428 21512 36688 21513
tri 36428 21511 36429 21512 ne
rect 36429 21511 36688 21512
tri 36429 21510 36430 21511 ne
rect 36430 21510 36688 21511
tri 36430 21509 36431 21510 ne
rect 36431 21509 36688 21510
tri 36431 21508 36432 21509 ne
rect 36432 21508 36688 21509
tri 36432 21507 36433 21508 ne
rect 36433 21507 36688 21508
tri 36433 21506 36434 21507 ne
rect 36434 21506 36688 21507
tri 36434 21505 36435 21506 ne
rect 36435 21505 36688 21506
tri 36435 21504 36436 21505 ne
rect 36436 21504 36688 21505
tri 36436 21503 36437 21504 ne
rect 36437 21503 36688 21504
tri 36437 21502 36438 21503 ne
rect 36438 21502 36688 21503
tri 36438 21501 36439 21502 ne
rect 36439 21501 36688 21502
tri 36439 21500 36440 21501 ne
rect 36440 21500 36688 21501
tri 36440 21499 36441 21500 ne
rect 36441 21499 36688 21500
tri 36441 21498 36442 21499 ne
rect 36442 21498 36688 21499
tri 36442 21497 36443 21498 ne
rect 36443 21497 36688 21498
tri 36443 21496 36444 21497 ne
rect 36444 21496 36688 21497
tri 36444 21495 36445 21496 ne
rect 36445 21495 36688 21496
tri 36445 21494 36446 21495 ne
rect 36446 21494 36688 21495
tri 36446 21493 36447 21494 ne
rect 36447 21493 36688 21494
tri 36447 21492 36448 21493 ne
rect 36448 21492 36688 21493
tri 36448 21491 36449 21492 ne
rect 36449 21491 36688 21492
tri 36449 21490 36450 21491 ne
rect 36450 21490 36688 21491
tri 36450 21489 36451 21490 ne
rect 36451 21489 36688 21490
tri 36451 21488 36452 21489 ne
rect 36452 21488 36688 21489
tri 36452 21487 36453 21488 ne
rect 36453 21487 36688 21488
tri 36453 21486 36454 21487 ne
rect 36454 21486 36688 21487
tri 36454 21485 36455 21486 ne
rect 36455 21485 36688 21486
tri 36455 21484 36456 21485 ne
rect 36456 21484 36688 21485
tri 36456 21483 36457 21484 ne
rect 36457 21483 36688 21484
tri 36688 21483 36733 21528 sw
rect 70802 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36457 21482 36458 21483 ne
rect 36458 21482 36733 21483
tri 36458 21481 36459 21482 ne
rect 36459 21481 36733 21482
tri 36459 21480 36460 21481 ne
rect 36460 21480 36733 21481
tri 36460 21479 36461 21480 ne
rect 36461 21479 36733 21480
tri 36461 21478 36462 21479 ne
rect 36462 21478 36733 21479
tri 36462 21477 36463 21478 ne
rect 36463 21477 36733 21478
tri 36463 21476 36464 21477 ne
rect 36464 21476 36733 21477
tri 36464 21475 36465 21476 ne
rect 36465 21475 36733 21476
tri 36465 21474 36466 21475 ne
rect 36466 21474 36733 21475
tri 36466 21473 36467 21474 ne
rect 36467 21473 36733 21474
tri 36467 21472 36468 21473 ne
rect 36468 21472 36733 21473
tri 36468 21471 36469 21472 ne
rect 36469 21471 36733 21472
tri 36469 21470 36470 21471 ne
rect 36470 21470 36733 21471
tri 36470 21469 36471 21470 ne
rect 36471 21469 36733 21470
tri 36471 21468 36472 21469 ne
rect 36472 21468 36733 21469
tri 36472 21467 36473 21468 ne
rect 36473 21467 36733 21468
tri 36473 21466 36474 21467 ne
rect 36474 21466 36733 21467
tri 36474 21465 36475 21466 ne
rect 36475 21465 36733 21466
tri 36475 21464 36476 21465 ne
rect 36476 21464 36733 21465
tri 36476 21463 36477 21464 ne
rect 36477 21463 36733 21464
tri 36477 21462 36478 21463 ne
rect 36478 21462 36733 21463
tri 36478 21461 36479 21462 ne
rect 36479 21461 36733 21462
tri 36479 21460 36480 21461 ne
rect 36480 21460 36733 21461
tri 36480 21459 36481 21460 ne
rect 36481 21459 36618 21460
tri 36481 21458 36482 21459 ne
rect 36482 21458 36618 21459
tri 36482 21457 36483 21458 ne
rect 36483 21457 36618 21458
tri 36483 21456 36484 21457 ne
rect 36484 21456 36618 21457
tri 36484 21455 36485 21456 ne
rect 36485 21455 36618 21456
tri 36485 21454 36486 21455 ne
rect 36486 21454 36618 21455
tri 36486 21453 36487 21454 ne
rect 36487 21453 36618 21454
tri 36487 21452 36488 21453 ne
rect 36488 21452 36618 21453
tri 36488 21451 36489 21452 ne
rect 36489 21451 36618 21452
tri 36489 21450 36490 21451 ne
rect 36490 21450 36618 21451
tri 36490 21449 36491 21450 ne
rect 36491 21449 36618 21450
tri 36491 21448 36492 21449 ne
rect 36492 21448 36618 21449
tri 36492 21447 36493 21448 ne
rect 36493 21447 36618 21448
tri 36493 21446 36494 21447 ne
rect 36494 21446 36618 21447
tri 36494 21445 36495 21446 ne
rect 36495 21445 36618 21446
tri 36495 21444 36496 21445 ne
rect 36496 21444 36618 21445
tri 36496 21443 36497 21444 ne
rect 36497 21443 36618 21444
tri 36497 21442 36498 21443 ne
rect 36498 21442 36618 21443
tri 36498 21441 36499 21442 ne
rect 36499 21441 36618 21442
tri 36499 21440 36500 21441 ne
rect 36500 21440 36618 21441
tri 36500 21439 36501 21440 ne
rect 36501 21439 36618 21440
tri 36501 21438 36502 21439 ne
rect 36502 21438 36618 21439
tri 36502 21437 36503 21438 ne
rect 36503 21437 36618 21438
tri 36503 21436 36504 21437 ne
rect 36504 21436 36618 21437
tri 36504 21435 36505 21436 ne
rect 36505 21435 36618 21436
tri 36505 21434 36506 21435 ne
rect 36506 21434 36618 21435
tri 36506 21433 36507 21434 ne
rect 36507 21433 36618 21434
tri 36507 21432 36508 21433 ne
rect 36508 21432 36618 21433
tri 36508 21431 36509 21432 ne
rect 36509 21431 36618 21432
tri 36509 21430 36510 21431 ne
rect 36510 21430 36618 21431
tri 36510 21429 36511 21430 ne
rect 36511 21429 36618 21430
tri 36511 21428 36512 21429 ne
rect 36512 21428 36618 21429
tri 36512 21427 36513 21428 ne
rect 36513 21427 36618 21428
tri 36513 21426 36514 21427 ne
rect 36514 21426 36618 21427
tri 36514 21425 36515 21426 ne
rect 36515 21425 36618 21426
tri 36515 21424 36516 21425 ne
rect 36516 21424 36618 21425
tri 36516 21423 36517 21424 ne
rect 36517 21423 36618 21424
tri 36517 21422 36518 21423 ne
rect 36518 21422 36618 21423
tri 36518 21421 36519 21422 ne
rect 36519 21421 36618 21422
tri 36519 21420 36520 21421 ne
rect 36520 21420 36618 21421
tri 36520 21419 36521 21420 ne
rect 36521 21419 36618 21420
tri 36521 21418 36522 21419 ne
rect 36522 21418 36618 21419
tri 36522 21417 36523 21418 ne
rect 36523 21417 36618 21418
tri 36523 21416 36524 21417 ne
rect 36524 21416 36618 21417
tri 36524 21415 36525 21416 ne
rect 36525 21415 36618 21416
tri 36525 21414 36526 21415 ne
rect 36526 21414 36618 21415
rect 36664 21438 36733 21460
tri 36733 21438 36778 21483 sw
rect 70802 21444 71000 21502
rect 36664 21422 36778 21438
tri 36778 21422 36794 21438 sw
rect 36664 21414 36794 21422
tri 36526 21413 36527 21414 ne
rect 36527 21413 36794 21414
tri 36527 21412 36528 21413 ne
rect 36528 21412 36794 21413
tri 36528 21411 36529 21412 ne
rect 36529 21411 36794 21412
tri 36529 21410 36530 21411 ne
rect 36530 21410 36794 21411
tri 36530 21409 36531 21410 ne
rect 36531 21409 36794 21410
tri 36531 21408 36532 21409 ne
rect 36532 21408 36794 21409
tri 36532 21407 36533 21408 ne
rect 36533 21407 36794 21408
tri 36533 21406 36534 21407 ne
rect 36534 21406 36794 21407
tri 36534 21405 36535 21406 ne
rect 36535 21405 36794 21406
tri 36535 21404 36536 21405 ne
rect 36536 21404 36794 21405
tri 36536 21403 36537 21404 ne
rect 36537 21403 36794 21404
tri 36537 21402 36538 21403 ne
rect 36538 21402 36794 21403
tri 36538 21401 36539 21402 ne
rect 36539 21401 36794 21402
tri 36539 21400 36540 21401 ne
rect 36540 21400 36794 21401
tri 36540 21399 36541 21400 ne
rect 36541 21399 36794 21400
tri 36541 21398 36542 21399 ne
rect 36542 21398 36794 21399
tri 36542 21397 36543 21398 ne
rect 36543 21397 36794 21398
tri 36543 21396 36544 21397 ne
rect 36544 21396 36794 21397
tri 36544 21395 36545 21396 ne
rect 36545 21395 36794 21396
tri 36545 21394 36546 21395 ne
rect 36546 21394 36794 21395
tri 36546 21393 36547 21394 ne
rect 36547 21393 36794 21394
tri 36547 21392 36548 21393 ne
rect 36548 21392 36794 21393
tri 36548 21391 36549 21392 ne
rect 36549 21391 36794 21392
tri 36549 21390 36550 21391 ne
rect 36550 21390 36794 21391
tri 36550 21389 36551 21390 ne
rect 36551 21389 36794 21390
tri 36551 21388 36552 21389 ne
rect 36552 21388 36794 21389
tri 36552 21387 36553 21388 ne
rect 36553 21387 36794 21388
tri 36553 21386 36554 21387 ne
rect 36554 21386 36794 21387
tri 36554 21385 36555 21386 ne
rect 36555 21385 36794 21386
tri 36555 21384 36556 21385 ne
rect 36556 21384 36794 21385
tri 36556 21383 36557 21384 ne
rect 36557 21383 36794 21384
tri 36557 21382 36558 21383 ne
rect 36558 21382 36794 21383
tri 36558 21381 36559 21382 ne
rect 36559 21381 36794 21382
tri 36559 21380 36560 21381 ne
rect 36560 21380 36794 21381
tri 36560 21379 36561 21380 ne
rect 36561 21379 36794 21380
tri 36561 21378 36562 21379 ne
rect 36562 21378 36794 21379
tri 36562 21377 36563 21378 ne
rect 36563 21377 36794 21378
tri 36794 21377 36839 21422 sw
rect 70802 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36563 21332 36608 21377 ne
rect 36608 21332 36839 21377
tri 36839 21332 36884 21377 sw
rect 70802 21340 71000 21398
tri 36608 21287 36653 21332 ne
rect 36653 21328 36884 21332
rect 36653 21287 36750 21328
tri 36653 21249 36691 21287 ne
rect 36691 21282 36750 21287
rect 36796 21287 36884 21328
tri 36884 21287 36929 21332 sw
rect 70802 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36796 21282 36929 21287
rect 36691 21252 36929 21282
tri 36929 21252 36964 21287 sw
rect 36691 21249 36964 21252
tri 36691 21248 36692 21249 ne
rect 36692 21248 36964 21249
tri 36692 21247 36693 21248 ne
rect 36693 21247 36964 21248
tri 36693 21246 36694 21247 ne
rect 36694 21246 36964 21247
tri 36694 21245 36695 21246 ne
rect 36695 21245 36964 21246
tri 36695 21244 36696 21245 ne
rect 36696 21244 36964 21245
tri 36696 21243 36697 21244 ne
rect 36697 21243 36964 21244
tri 36697 21242 36698 21243 ne
rect 36698 21242 36964 21243
tri 36698 21241 36699 21242 ne
rect 36699 21241 36964 21242
tri 36699 21240 36700 21241 ne
rect 36700 21240 36964 21241
tri 36700 21239 36701 21240 ne
rect 36701 21239 36964 21240
tri 36701 21238 36702 21239 ne
rect 36702 21238 36964 21239
tri 36702 21237 36703 21238 ne
rect 36703 21237 36964 21238
tri 36703 21236 36704 21237 ne
rect 36704 21236 36964 21237
tri 36704 21235 36705 21236 ne
rect 36705 21235 36964 21236
tri 36705 21234 36706 21235 ne
rect 36706 21234 36964 21235
tri 36706 21233 36707 21234 ne
rect 36707 21233 36964 21234
tri 36707 21232 36708 21233 ne
rect 36708 21232 36964 21233
tri 36708 21231 36709 21232 ne
rect 36709 21231 36964 21232
tri 36709 21230 36710 21231 ne
rect 36710 21230 36964 21231
tri 36710 21229 36711 21230 ne
rect 36711 21229 36964 21230
tri 36711 21228 36712 21229 ne
rect 36712 21228 36964 21229
tri 36712 21227 36713 21228 ne
rect 36713 21227 36964 21228
tri 36713 21226 36714 21227 ne
rect 36714 21226 36964 21227
tri 36714 21225 36715 21226 ne
rect 36715 21225 36964 21226
tri 36715 21224 36716 21225 ne
rect 36716 21224 36964 21225
tri 36716 21223 36717 21224 ne
rect 36717 21223 36964 21224
tri 36717 21222 36718 21223 ne
rect 36718 21222 36964 21223
tri 36718 21221 36719 21222 ne
rect 36719 21221 36964 21222
tri 36719 21220 36720 21221 ne
rect 36720 21220 36964 21221
tri 36720 21219 36721 21220 ne
rect 36721 21219 36964 21220
tri 36721 21218 36722 21219 ne
rect 36722 21218 36964 21219
tri 36722 21217 36723 21218 ne
rect 36723 21217 36964 21218
tri 36723 21216 36724 21217 ne
rect 36724 21216 36964 21217
tri 36724 21215 36725 21216 ne
rect 36725 21215 36964 21216
tri 36725 21214 36726 21215 ne
rect 36726 21214 36964 21215
tri 36726 21213 36727 21214 ne
rect 36727 21213 36964 21214
tri 36727 21212 36728 21213 ne
rect 36728 21212 36964 21213
tri 36728 21211 36729 21212 ne
rect 36729 21211 36964 21212
tri 36729 21210 36730 21211 ne
rect 36730 21210 36964 21211
tri 36730 21209 36731 21210 ne
rect 36731 21209 36964 21210
tri 36731 21208 36732 21209 ne
rect 36732 21208 36964 21209
tri 36732 21207 36733 21208 ne
rect 36733 21207 36964 21208
tri 36964 21207 37009 21252 sw
rect 70802 21236 71000 21294
tri 36733 21206 36734 21207 ne
rect 36734 21206 37009 21207
tri 36734 21205 36735 21206 ne
rect 36735 21205 37009 21206
tri 36735 21204 36736 21205 ne
rect 36736 21204 37009 21205
tri 36736 21203 36737 21204 ne
rect 36737 21203 37009 21204
tri 36737 21202 36738 21203 ne
rect 36738 21202 37009 21203
tri 36738 21201 36739 21202 ne
rect 36739 21201 37009 21202
tri 36739 21200 36740 21201 ne
rect 36740 21200 37009 21201
tri 36740 21199 36741 21200 ne
rect 36741 21199 37009 21200
tri 36741 21198 36742 21199 ne
rect 36742 21198 37009 21199
tri 36742 21197 36743 21198 ne
rect 36743 21197 37009 21198
tri 36743 21196 36744 21197 ne
rect 36744 21196 37009 21197
tri 36744 21195 36745 21196 ne
rect 36745 21195 36882 21196
tri 36745 21194 36746 21195 ne
rect 36746 21194 36882 21195
tri 36746 21193 36747 21194 ne
rect 36747 21193 36882 21194
tri 36747 21192 36748 21193 ne
rect 36748 21192 36882 21193
tri 36748 21191 36749 21192 ne
rect 36749 21191 36882 21192
tri 36749 21190 36750 21191 ne
rect 36750 21190 36882 21191
tri 36750 21189 36751 21190 ne
rect 36751 21189 36882 21190
tri 36751 21188 36752 21189 ne
rect 36752 21188 36882 21189
tri 36752 21187 36753 21188 ne
rect 36753 21187 36882 21188
tri 36753 21186 36754 21187 ne
rect 36754 21186 36882 21187
tri 36754 21185 36755 21186 ne
rect 36755 21185 36882 21186
tri 36755 21184 36756 21185 ne
rect 36756 21184 36882 21185
tri 36756 21183 36757 21184 ne
rect 36757 21183 36882 21184
tri 36757 21182 36758 21183 ne
rect 36758 21182 36882 21183
tri 36758 21181 36759 21182 ne
rect 36759 21181 36882 21182
tri 36759 21180 36760 21181 ne
rect 36760 21180 36882 21181
tri 36760 21179 36761 21180 ne
rect 36761 21179 36882 21180
tri 36761 21178 36762 21179 ne
rect 36762 21178 36882 21179
tri 36762 21177 36763 21178 ne
rect 36763 21177 36882 21178
tri 36763 21176 36764 21177 ne
rect 36764 21176 36882 21177
tri 36764 21175 36765 21176 ne
rect 36765 21175 36882 21176
tri 36765 21174 36766 21175 ne
rect 36766 21174 36882 21175
tri 36766 21173 36767 21174 ne
rect 36767 21173 36882 21174
tri 36767 21172 36768 21173 ne
rect 36768 21172 36882 21173
tri 36768 21171 36769 21172 ne
rect 36769 21171 36882 21172
tri 36769 21170 36770 21171 ne
rect 36770 21170 36882 21171
tri 36770 21169 36771 21170 ne
rect 36771 21169 36882 21170
tri 36771 21168 36772 21169 ne
rect 36772 21168 36882 21169
tri 36772 21167 36773 21168 ne
rect 36773 21167 36882 21168
tri 36773 21166 36774 21167 ne
rect 36774 21166 36882 21167
tri 36774 21165 36775 21166 ne
rect 36775 21165 36882 21166
tri 36775 21164 36776 21165 ne
rect 36776 21164 36882 21165
tri 36776 21163 36777 21164 ne
rect 36777 21163 36882 21164
tri 36777 21162 36778 21163 ne
rect 36778 21162 36882 21163
tri 36778 21161 36779 21162 ne
rect 36779 21161 36882 21162
tri 36779 21160 36780 21161 ne
rect 36780 21160 36882 21161
tri 36780 21159 36781 21160 ne
rect 36781 21159 36882 21160
tri 36781 21158 36782 21159 ne
rect 36782 21158 36882 21159
tri 36782 21157 36783 21158 ne
rect 36783 21157 36882 21158
tri 36783 21156 36784 21157 ne
rect 36784 21156 36882 21157
tri 36784 21155 36785 21156 ne
rect 36785 21155 36882 21156
tri 36785 21154 36786 21155 ne
rect 36786 21154 36882 21155
tri 36786 21153 36787 21154 ne
rect 36787 21153 36882 21154
tri 36787 21152 36788 21153 ne
rect 36788 21152 36882 21153
tri 36788 21151 36789 21152 ne
rect 36789 21151 36882 21152
tri 36789 21150 36790 21151 ne
rect 36790 21150 36882 21151
rect 36928 21162 37009 21196
tri 37009 21162 37054 21207 sw
rect 70802 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21150 37054 21162
tri 36790 21149 36791 21150 ne
rect 36791 21149 37054 21150
tri 36791 21148 36792 21149 ne
rect 36792 21148 37054 21149
tri 36792 21147 36793 21148 ne
rect 36793 21147 37054 21148
tri 36793 21146 36794 21147 ne
rect 36794 21146 37054 21147
tri 36794 21145 36795 21146 ne
rect 36795 21145 37054 21146
tri 36795 21144 36796 21145 ne
rect 36796 21144 37054 21145
tri 36796 21143 36797 21144 ne
rect 36797 21143 37054 21144
tri 36797 21142 36798 21143 ne
rect 36798 21142 37054 21143
tri 36798 21141 36799 21142 ne
rect 36799 21141 37054 21142
tri 36799 21140 36800 21141 ne
rect 36800 21140 37054 21141
tri 36800 21139 36801 21140 ne
rect 36801 21139 37054 21140
tri 36801 21138 36802 21139 ne
rect 36802 21138 37054 21139
tri 36802 21137 36803 21138 ne
rect 36803 21137 37054 21138
tri 36803 21136 36804 21137 ne
rect 36804 21136 37054 21137
tri 36804 21135 36805 21136 ne
rect 36805 21135 37054 21136
tri 36805 21134 36806 21135 ne
rect 36806 21134 37054 21135
tri 36806 21133 36807 21134 ne
rect 36807 21133 37054 21134
tri 36807 21132 36808 21133 ne
rect 36808 21132 37054 21133
tri 36808 21131 36809 21132 ne
rect 36809 21131 37054 21132
tri 36809 21130 36810 21131 ne
rect 36810 21130 37054 21131
tri 36810 21129 36811 21130 ne
rect 36811 21129 37054 21130
tri 36811 21128 36812 21129 ne
rect 36812 21128 37054 21129
tri 36812 21127 36813 21128 ne
rect 36813 21127 37054 21128
tri 36813 21126 36814 21127 ne
rect 36814 21126 37054 21127
tri 36814 21125 36815 21126 ne
rect 36815 21125 37054 21126
tri 36815 21124 36816 21125 ne
rect 36816 21124 37054 21125
tri 36816 21123 36817 21124 ne
rect 36817 21123 37054 21124
tri 36817 21122 36818 21123 ne
rect 36818 21122 37054 21123
tri 36818 21121 36819 21122 ne
rect 36819 21121 37054 21122
tri 36819 21120 36820 21121 ne
rect 36820 21120 37054 21121
tri 36820 21119 36821 21120 ne
rect 36821 21119 37054 21120
tri 36821 21118 36822 21119 ne
rect 36822 21118 37054 21119
tri 36822 21117 36823 21118 ne
rect 36823 21117 37054 21118
tri 37054 21117 37099 21162 sw
rect 70802 21132 71000 21190
tri 36823 21116 36824 21117 ne
rect 36824 21116 37099 21117
tri 36824 21115 36825 21116 ne
rect 36825 21115 37099 21116
tri 36825 21114 36826 21115 ne
rect 36826 21114 37099 21115
tri 36826 21113 36827 21114 ne
rect 36827 21113 37099 21114
tri 36827 21112 36828 21113 ne
rect 36828 21112 37099 21113
tri 36828 21111 36829 21112 ne
rect 36829 21111 37099 21112
tri 36829 21110 36830 21111 ne
rect 36830 21110 37099 21111
tri 36830 21109 36831 21110 ne
rect 36831 21109 37099 21110
tri 36831 21108 36832 21109 ne
rect 36832 21108 37099 21109
tri 36832 21107 36833 21108 ne
rect 36833 21107 37099 21108
tri 36833 21106 36834 21107 ne
rect 36834 21106 37099 21107
tri 36834 21105 36835 21106 ne
rect 36835 21105 37099 21106
tri 36835 21104 36836 21105 ne
rect 36836 21104 37099 21105
tri 36836 21103 36837 21104 ne
rect 36837 21103 37099 21104
tri 36837 21102 36838 21103 ne
rect 36838 21102 37099 21103
tri 36838 21101 36839 21102 ne
rect 36839 21101 37099 21102
tri 37099 21101 37115 21117 sw
tri 36839 21056 36884 21101 ne
rect 36884 21072 37115 21101
tri 37115 21072 37144 21101 sw
rect 70802 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 36884 21064 37144 21072
rect 36884 21056 37014 21064
tri 36884 21029 36911 21056 ne
rect 36911 21029 37014 21056
tri 36911 20984 36956 21029 ne
rect 36956 21018 37014 21029
rect 37060 21027 37144 21064
tri 37144 21027 37189 21072 sw
rect 70802 21028 71000 21086
rect 37060 21018 37189 21027
rect 36956 20984 37189 21018
tri 36956 20974 36966 20984 ne
rect 36966 20982 37189 20984
tri 37189 20982 37234 21027 sw
rect 70802 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
rect 36966 20974 37234 20982
tri 36966 20973 36967 20974 ne
rect 36967 20973 37234 20974
tri 36967 20972 36968 20973 ne
rect 36968 20972 37234 20973
tri 36968 20971 36969 20972 ne
rect 36969 20971 37234 20972
tri 36969 20970 36970 20971 ne
rect 36970 20970 37234 20971
tri 36970 20969 36971 20970 ne
rect 36971 20969 37234 20970
tri 36971 20968 36972 20969 ne
rect 36972 20968 37234 20969
tri 36972 20967 36973 20968 ne
rect 36973 20967 37234 20968
tri 36973 20966 36974 20967 ne
rect 36974 20966 37234 20967
tri 36974 20965 36975 20966 ne
rect 36975 20965 37234 20966
tri 36975 20964 36976 20965 ne
rect 36976 20964 37234 20965
tri 36976 20963 36977 20964 ne
rect 36977 20963 37234 20964
tri 36977 20962 36978 20963 ne
rect 36978 20962 37234 20963
tri 36978 20961 36979 20962 ne
rect 36979 20961 37234 20962
tri 36979 20960 36980 20961 ne
rect 36980 20960 37234 20961
tri 37234 20960 37256 20982 sw
tri 36980 20959 36981 20960 ne
rect 36981 20959 37256 20960
tri 36981 20958 36982 20959 ne
rect 36982 20958 37256 20959
tri 36982 20957 36983 20958 ne
rect 36983 20957 37256 20958
tri 36983 20956 36984 20957 ne
rect 36984 20956 37256 20957
tri 36984 20955 36985 20956 ne
rect 36985 20955 37256 20956
tri 36985 20954 36986 20955 ne
rect 36986 20954 37256 20955
tri 36986 20953 36987 20954 ne
rect 36987 20953 37256 20954
tri 36987 20952 36988 20953 ne
rect 36988 20952 37256 20953
tri 36988 20951 36989 20952 ne
rect 36989 20951 37256 20952
tri 36989 20950 36990 20951 ne
rect 36990 20950 37256 20951
tri 36990 20949 36991 20950 ne
rect 36991 20949 37256 20950
tri 36991 20948 36992 20949 ne
rect 36992 20948 37256 20949
tri 36992 20947 36993 20948 ne
rect 36993 20947 37256 20948
tri 36993 20946 36994 20947 ne
rect 36994 20946 37256 20947
tri 36994 20945 36995 20946 ne
rect 36995 20945 37256 20946
tri 36995 20944 36996 20945 ne
rect 36996 20944 37256 20945
tri 36996 20943 36997 20944 ne
rect 36997 20943 37256 20944
tri 36997 20942 36998 20943 ne
rect 36998 20942 37256 20943
tri 36998 20941 36999 20942 ne
rect 36999 20941 37256 20942
tri 36999 20940 37000 20941 ne
rect 37000 20940 37256 20941
tri 37000 20939 37001 20940 ne
rect 37001 20939 37256 20940
tri 37001 20938 37002 20939 ne
rect 37002 20938 37256 20939
tri 37002 20937 37003 20938 ne
rect 37003 20937 37256 20938
tri 37003 20936 37004 20937 ne
rect 37004 20936 37256 20937
tri 37004 20935 37005 20936 ne
rect 37005 20935 37256 20936
tri 37005 20934 37006 20935 ne
rect 37006 20934 37256 20935
tri 37006 20933 37007 20934 ne
rect 37007 20933 37256 20934
tri 37007 20932 37008 20933 ne
rect 37008 20932 37256 20933
tri 37008 20931 37009 20932 ne
rect 37009 20931 37146 20932
tri 37009 20930 37010 20931 ne
rect 37010 20930 37146 20931
tri 37010 20929 37011 20930 ne
rect 37011 20929 37146 20930
tri 37011 20928 37012 20929 ne
rect 37012 20928 37146 20929
tri 37012 20927 37013 20928 ne
rect 37013 20927 37146 20928
tri 37013 20926 37014 20927 ne
rect 37014 20926 37146 20927
tri 37014 20925 37015 20926 ne
rect 37015 20925 37146 20926
tri 37015 20924 37016 20925 ne
rect 37016 20924 37146 20925
tri 37016 20923 37017 20924 ne
rect 37017 20923 37146 20924
tri 37017 20922 37018 20923 ne
rect 37018 20922 37146 20923
tri 37018 20921 37019 20922 ne
rect 37019 20921 37146 20922
tri 37019 20920 37020 20921 ne
rect 37020 20920 37146 20921
tri 37020 20919 37021 20920 ne
rect 37021 20919 37146 20920
tri 37021 20918 37022 20919 ne
rect 37022 20918 37146 20919
tri 37022 20917 37023 20918 ne
rect 37023 20917 37146 20918
tri 37023 20916 37024 20917 ne
rect 37024 20916 37146 20917
tri 37024 20915 37025 20916 ne
rect 37025 20915 37146 20916
tri 37025 20914 37026 20915 ne
rect 37026 20914 37146 20915
tri 37026 20913 37027 20914 ne
rect 37027 20913 37146 20914
tri 37027 20912 37028 20913 ne
rect 37028 20912 37146 20913
tri 37028 20911 37029 20912 ne
rect 37029 20911 37146 20912
tri 37029 20910 37030 20911 ne
rect 37030 20910 37146 20911
tri 37030 20909 37031 20910 ne
rect 37031 20909 37146 20910
tri 37031 20908 37032 20909 ne
rect 37032 20908 37146 20909
tri 37032 20907 37033 20908 ne
rect 37033 20907 37146 20908
tri 37033 20906 37034 20907 ne
rect 37034 20906 37146 20907
tri 37034 20905 37035 20906 ne
rect 37035 20905 37146 20906
tri 37035 20904 37036 20905 ne
rect 37036 20904 37146 20905
tri 37036 20903 37037 20904 ne
rect 37037 20903 37146 20904
tri 37037 20902 37038 20903 ne
rect 37038 20902 37146 20903
tri 37038 20901 37039 20902 ne
rect 37039 20901 37146 20902
tri 37039 20900 37040 20901 ne
rect 37040 20900 37146 20901
tri 37040 20899 37041 20900 ne
rect 37041 20899 37146 20900
tri 37041 20898 37042 20899 ne
rect 37042 20898 37146 20899
tri 37042 20897 37043 20898 ne
rect 37043 20897 37146 20898
tri 37043 20896 37044 20897 ne
rect 37044 20896 37146 20897
tri 37044 20895 37045 20896 ne
rect 37045 20895 37146 20896
tri 37045 20894 37046 20895 ne
rect 37046 20894 37146 20895
tri 37046 20893 37047 20894 ne
rect 37047 20893 37146 20894
tri 37047 20892 37048 20893 ne
rect 37048 20892 37146 20893
tri 37048 20891 37049 20892 ne
rect 37049 20891 37146 20892
tri 37049 20890 37050 20891 ne
rect 37050 20890 37146 20891
tri 37050 20889 37051 20890 ne
rect 37051 20889 37146 20890
tri 37051 20888 37052 20889 ne
rect 37052 20888 37146 20889
tri 37052 20887 37053 20888 ne
rect 37053 20887 37146 20888
tri 37053 20886 37054 20887 ne
rect 37054 20886 37146 20887
rect 37192 20915 37256 20932
tri 37256 20915 37301 20960 sw
rect 70802 20924 71000 20982
rect 37192 20886 37301 20915
tri 37054 20885 37055 20886 ne
rect 37055 20885 37301 20886
tri 37055 20884 37056 20885 ne
rect 37056 20884 37301 20885
tri 37056 20883 37057 20884 ne
rect 37057 20883 37301 20884
tri 37057 20882 37058 20883 ne
rect 37058 20882 37301 20883
tri 37058 20881 37059 20882 ne
rect 37059 20881 37301 20882
tri 37059 20880 37060 20881 ne
rect 37060 20880 37301 20881
tri 37060 20879 37061 20880 ne
rect 37061 20879 37301 20880
tri 37061 20878 37062 20879 ne
rect 37062 20878 37301 20879
tri 37062 20877 37063 20878 ne
rect 37063 20877 37301 20878
tri 37063 20876 37064 20877 ne
rect 37064 20876 37301 20877
tri 37064 20875 37065 20876 ne
rect 37065 20875 37301 20876
tri 37065 20874 37066 20875 ne
rect 37066 20874 37301 20875
tri 37066 20873 37067 20874 ne
rect 37067 20873 37301 20874
tri 37067 20872 37068 20873 ne
rect 37068 20872 37301 20873
tri 37068 20871 37069 20872 ne
rect 37069 20871 37301 20872
tri 37069 20870 37070 20871 ne
rect 37070 20870 37301 20871
tri 37301 20870 37346 20915 sw
rect 70802 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
tri 37070 20869 37071 20870 ne
rect 37071 20869 37346 20870
tri 37071 20868 37072 20869 ne
rect 37072 20868 37346 20869
tri 37072 20867 37073 20868 ne
rect 37073 20867 37346 20868
tri 37073 20866 37074 20867 ne
rect 37074 20866 37346 20867
tri 37074 20865 37075 20866 ne
rect 37075 20865 37346 20866
tri 37075 20864 37076 20865 ne
rect 37076 20864 37346 20865
tri 37076 20863 37077 20864 ne
rect 37077 20863 37346 20864
tri 37077 20862 37078 20863 ne
rect 37078 20862 37346 20863
tri 37078 20861 37079 20862 ne
rect 37079 20861 37346 20862
tri 37079 20860 37080 20861 ne
rect 37080 20860 37346 20861
tri 37080 20859 37081 20860 ne
rect 37081 20859 37346 20860
tri 37081 20858 37082 20859 ne
rect 37082 20858 37346 20859
tri 37082 20857 37083 20858 ne
rect 37083 20857 37346 20858
tri 37083 20856 37084 20857 ne
rect 37084 20856 37346 20857
tri 37084 20855 37085 20856 ne
rect 37085 20855 37346 20856
tri 37085 20854 37086 20855 ne
rect 37086 20854 37346 20855
tri 37086 20853 37087 20854 ne
rect 37087 20853 37346 20854
tri 37087 20852 37088 20853 ne
rect 37088 20852 37346 20853
tri 37088 20851 37089 20852 ne
rect 37089 20851 37346 20852
tri 37089 20850 37090 20851 ne
rect 37090 20850 37346 20851
tri 37090 20849 37091 20850 ne
rect 37091 20849 37346 20850
tri 37091 20848 37092 20849 ne
rect 37092 20848 37346 20849
tri 37092 20847 37093 20848 ne
rect 37093 20847 37346 20848
tri 37093 20846 37094 20847 ne
rect 37094 20846 37346 20847
tri 37094 20845 37095 20846 ne
rect 37095 20845 37346 20846
tri 37095 20844 37096 20845 ne
rect 37096 20844 37346 20845
tri 37096 20843 37097 20844 ne
rect 37097 20843 37346 20844
tri 37097 20842 37098 20843 ne
rect 37098 20842 37346 20843
tri 37098 20841 37099 20842 ne
rect 37099 20841 37346 20842
tri 37099 20840 37100 20841 ne
rect 37100 20840 37346 20841
tri 37100 20839 37101 20840 ne
rect 37101 20839 37346 20840
tri 37101 20838 37102 20839 ne
rect 37102 20838 37346 20839
tri 37102 20837 37103 20838 ne
rect 37103 20837 37346 20838
tri 37103 20836 37104 20837 ne
rect 37104 20836 37346 20837
tri 37104 20835 37105 20836 ne
rect 37105 20835 37346 20836
tri 37105 20834 37106 20835 ne
rect 37106 20834 37346 20835
tri 37106 20833 37107 20834 ne
rect 37107 20833 37346 20834
tri 37107 20832 37108 20833 ne
rect 37108 20832 37346 20833
tri 37108 20831 37109 20832 ne
rect 37109 20831 37346 20832
tri 37109 20830 37110 20831 ne
rect 37110 20830 37346 20831
tri 37110 20829 37111 20830 ne
rect 37111 20829 37346 20830
tri 37111 20828 37112 20829 ne
rect 37112 20828 37346 20829
tri 37112 20827 37113 20828 ne
rect 37113 20827 37346 20828
tri 37113 20826 37114 20827 ne
rect 37114 20826 37346 20827
tri 37114 20825 37115 20826 ne
rect 37115 20825 37346 20826
tri 37346 20825 37391 20870 sw
tri 37115 20796 37144 20825 ne
rect 37144 20800 37391 20825
rect 37144 20796 37278 20800
tri 37144 20780 37160 20796 ne
rect 37160 20780 37278 20796
tri 37160 20751 37189 20780 ne
rect 37189 20754 37278 20780
rect 37324 20796 37391 20800
tri 37391 20796 37420 20825 sw
rect 70802 20820 71000 20878
rect 37324 20754 37420 20796
rect 37189 20751 37420 20754
tri 37420 20751 37465 20796 sw
rect 70802 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
tri 37189 20706 37234 20751 ne
rect 37234 20706 37465 20751
tri 37465 20706 37510 20751 sw
rect 70802 20716 71000 20774
tri 37234 20700 37240 20706 ne
rect 37240 20700 37510 20706
tri 37240 20699 37241 20700 ne
rect 37241 20699 37510 20700
tri 37241 20698 37242 20699 ne
rect 37242 20698 37510 20699
tri 37242 20697 37243 20698 ne
rect 37243 20697 37510 20698
tri 37243 20696 37244 20697 ne
rect 37244 20696 37510 20697
tri 37244 20695 37245 20696 ne
rect 37245 20695 37510 20696
tri 37245 20694 37246 20695 ne
rect 37246 20694 37510 20695
tri 37246 20693 37247 20694 ne
rect 37247 20693 37510 20694
tri 37247 20692 37248 20693 ne
rect 37248 20692 37510 20693
tri 37248 20691 37249 20692 ne
rect 37249 20691 37510 20692
tri 37249 20690 37250 20691 ne
rect 37250 20690 37510 20691
tri 37250 20689 37251 20690 ne
rect 37251 20689 37510 20690
tri 37251 20688 37252 20689 ne
rect 37252 20688 37510 20689
tri 37252 20687 37253 20688 ne
rect 37253 20687 37510 20688
tri 37253 20686 37254 20687 ne
rect 37254 20686 37510 20687
tri 37254 20685 37255 20686 ne
rect 37255 20685 37510 20686
tri 37255 20684 37256 20685 ne
rect 37256 20684 37510 20685
tri 37256 20683 37257 20684 ne
rect 37257 20683 37510 20684
tri 37257 20682 37258 20683 ne
rect 37258 20682 37510 20683
tri 37258 20681 37259 20682 ne
rect 37259 20681 37510 20682
tri 37259 20680 37260 20681 ne
rect 37260 20680 37510 20681
tri 37260 20679 37261 20680 ne
rect 37261 20679 37510 20680
tri 37261 20678 37262 20679 ne
rect 37262 20678 37510 20679
tri 37262 20677 37263 20678 ne
rect 37263 20677 37510 20678
tri 37263 20676 37264 20677 ne
rect 37264 20676 37510 20677
tri 37264 20675 37265 20676 ne
rect 37265 20675 37510 20676
tri 37265 20674 37266 20675 ne
rect 37266 20674 37510 20675
tri 37266 20673 37267 20674 ne
rect 37267 20673 37510 20674
tri 37267 20672 37268 20673 ne
rect 37268 20672 37510 20673
tri 37268 20671 37269 20672 ne
rect 37269 20671 37510 20672
tri 37269 20670 37270 20671 ne
rect 37270 20670 37510 20671
tri 37270 20669 37271 20670 ne
rect 37271 20669 37510 20670
tri 37271 20668 37272 20669 ne
rect 37272 20668 37510 20669
tri 37272 20667 37273 20668 ne
rect 37273 20667 37410 20668
tri 37273 20666 37274 20667 ne
rect 37274 20666 37410 20667
tri 37274 20665 37275 20666 ne
rect 37275 20665 37410 20666
tri 37275 20664 37276 20665 ne
rect 37276 20664 37410 20665
tri 37276 20663 37277 20664 ne
rect 37277 20663 37410 20664
tri 37277 20662 37278 20663 ne
rect 37278 20662 37410 20663
tri 37278 20661 37279 20662 ne
rect 37279 20661 37410 20662
tri 37279 20660 37280 20661 ne
rect 37280 20660 37410 20661
tri 37280 20659 37281 20660 ne
rect 37281 20659 37410 20660
tri 37281 20658 37282 20659 ne
rect 37282 20658 37410 20659
tri 37282 20657 37283 20658 ne
rect 37283 20657 37410 20658
tri 37283 20656 37284 20657 ne
rect 37284 20656 37410 20657
tri 37284 20655 37285 20656 ne
rect 37285 20655 37410 20656
tri 37285 20654 37286 20655 ne
rect 37286 20654 37410 20655
tri 37286 20653 37287 20654 ne
rect 37287 20653 37410 20654
tri 37287 20652 37288 20653 ne
rect 37288 20652 37410 20653
tri 37288 20651 37289 20652 ne
rect 37289 20651 37410 20652
tri 37289 20650 37290 20651 ne
rect 37290 20650 37410 20651
tri 37290 20649 37291 20650 ne
rect 37291 20649 37410 20650
tri 37291 20648 37292 20649 ne
rect 37292 20648 37410 20649
tri 37292 20647 37293 20648 ne
rect 37293 20647 37410 20648
tri 37293 20646 37294 20647 ne
rect 37294 20646 37410 20647
tri 37294 20645 37295 20646 ne
rect 37295 20645 37410 20646
tri 37295 20644 37296 20645 ne
rect 37296 20644 37410 20645
tri 37296 20643 37297 20644 ne
rect 37297 20643 37410 20644
tri 37297 20642 37298 20643 ne
rect 37298 20642 37410 20643
tri 37298 20641 37299 20642 ne
rect 37299 20641 37410 20642
tri 37299 20640 37300 20641 ne
rect 37300 20640 37410 20641
tri 37300 20639 37301 20640 ne
rect 37301 20639 37410 20640
tri 37301 20638 37302 20639 ne
rect 37302 20638 37410 20639
tri 37302 20637 37303 20638 ne
rect 37303 20637 37410 20638
tri 37303 20636 37304 20637 ne
rect 37304 20636 37410 20637
tri 37304 20635 37305 20636 ne
rect 37305 20635 37410 20636
tri 37305 20634 37306 20635 ne
rect 37306 20634 37410 20635
tri 37306 20633 37307 20634 ne
rect 37307 20633 37410 20634
tri 37307 20632 37308 20633 ne
rect 37308 20632 37410 20633
tri 37308 20631 37309 20632 ne
rect 37309 20631 37410 20632
tri 37309 20630 37310 20631 ne
rect 37310 20630 37410 20631
tri 37310 20629 37311 20630 ne
rect 37311 20629 37410 20630
tri 37311 20628 37312 20629 ne
rect 37312 20628 37410 20629
tri 37312 20627 37313 20628 ne
rect 37313 20627 37410 20628
tri 37313 20626 37314 20627 ne
rect 37314 20626 37410 20627
tri 37314 20625 37315 20626 ne
rect 37315 20625 37410 20626
tri 37315 20624 37316 20625 ne
rect 37316 20624 37410 20625
tri 37316 20623 37317 20624 ne
rect 37317 20623 37410 20624
tri 37317 20622 37318 20623 ne
rect 37318 20622 37410 20623
rect 37456 20661 37510 20668
tri 37510 20661 37555 20706 sw
rect 70802 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 37456 20639 37555 20661
tri 37555 20639 37577 20661 sw
rect 37456 20622 37577 20639
tri 37318 20621 37319 20622 ne
rect 37319 20621 37577 20622
tri 37319 20620 37320 20621 ne
rect 37320 20620 37577 20621
tri 37320 20619 37321 20620 ne
rect 37321 20619 37577 20620
tri 37321 20618 37322 20619 ne
rect 37322 20618 37577 20619
tri 37322 20617 37323 20618 ne
rect 37323 20617 37577 20618
tri 37323 20616 37324 20617 ne
rect 37324 20616 37577 20617
tri 37324 20615 37325 20616 ne
rect 37325 20615 37577 20616
tri 37325 20614 37326 20615 ne
rect 37326 20614 37577 20615
tri 37326 20613 37327 20614 ne
rect 37327 20613 37577 20614
tri 37327 20612 37328 20613 ne
rect 37328 20612 37577 20613
tri 37328 20611 37329 20612 ne
rect 37329 20611 37577 20612
tri 37329 20610 37330 20611 ne
rect 37330 20610 37577 20611
tri 37330 20609 37331 20610 ne
rect 37331 20609 37577 20610
tri 37331 20608 37332 20609 ne
rect 37332 20608 37577 20609
tri 37332 20607 37333 20608 ne
rect 37333 20607 37577 20608
tri 37333 20606 37334 20607 ne
rect 37334 20606 37577 20607
tri 37334 20605 37335 20606 ne
rect 37335 20605 37577 20606
tri 37335 20604 37336 20605 ne
rect 37336 20604 37577 20605
tri 37336 20603 37337 20604 ne
rect 37337 20603 37577 20604
tri 37337 20602 37338 20603 ne
rect 37338 20602 37577 20603
tri 37338 20601 37339 20602 ne
rect 37339 20601 37577 20602
tri 37339 20600 37340 20601 ne
rect 37340 20600 37577 20601
tri 37340 20599 37341 20600 ne
rect 37341 20599 37577 20600
tri 37341 20598 37342 20599 ne
rect 37342 20598 37577 20599
tri 37342 20597 37343 20598 ne
rect 37343 20597 37577 20598
tri 37343 20596 37344 20597 ne
rect 37344 20596 37577 20597
tri 37344 20595 37345 20596 ne
rect 37345 20595 37577 20596
tri 37345 20594 37346 20595 ne
rect 37346 20594 37577 20595
tri 37577 20594 37622 20639 sw
rect 70802 20612 71000 20670
tri 37346 20593 37347 20594 ne
rect 37347 20593 37622 20594
tri 37347 20592 37348 20593 ne
rect 37348 20592 37622 20593
tri 37348 20591 37349 20592 ne
rect 37349 20591 37622 20592
tri 37349 20590 37350 20591 ne
rect 37350 20590 37622 20591
tri 37350 20589 37351 20590 ne
rect 37351 20589 37622 20590
tri 37351 20588 37352 20589 ne
rect 37352 20588 37622 20589
tri 37352 20587 37353 20588 ne
rect 37353 20587 37622 20588
tri 37353 20586 37354 20587 ne
rect 37354 20586 37622 20587
tri 37354 20585 37355 20586 ne
rect 37355 20585 37622 20586
tri 37355 20584 37356 20585 ne
rect 37356 20584 37622 20585
tri 37356 20583 37357 20584 ne
rect 37357 20583 37622 20584
tri 37357 20582 37358 20583 ne
rect 37358 20582 37622 20583
tri 37358 20581 37359 20582 ne
rect 37359 20581 37622 20582
tri 37359 20580 37360 20581 ne
rect 37360 20580 37622 20581
tri 37360 20579 37361 20580 ne
rect 37361 20579 37622 20580
tri 37361 20578 37362 20579 ne
rect 37362 20578 37622 20579
tri 37362 20577 37363 20578 ne
rect 37363 20577 37622 20578
tri 37363 20576 37364 20577 ne
rect 37364 20576 37622 20577
tri 37364 20575 37365 20576 ne
rect 37365 20575 37622 20576
tri 37365 20574 37366 20575 ne
rect 37366 20574 37622 20575
tri 37366 20573 37367 20574 ne
rect 37367 20573 37622 20574
tri 37367 20572 37368 20573 ne
rect 37368 20572 37622 20573
tri 37368 20571 37369 20572 ne
rect 37369 20571 37622 20572
tri 37369 20570 37370 20571 ne
rect 37370 20570 37622 20571
tri 37370 20569 37371 20570 ne
rect 37371 20569 37622 20570
tri 37371 20568 37372 20569 ne
rect 37372 20568 37622 20569
tri 37372 20567 37373 20568 ne
rect 37373 20567 37622 20568
tri 37373 20566 37374 20567 ne
rect 37374 20566 37622 20567
tri 37374 20565 37375 20566 ne
rect 37375 20565 37622 20566
tri 37375 20564 37376 20565 ne
rect 37376 20564 37622 20565
tri 37376 20563 37377 20564 ne
rect 37377 20563 37622 20564
tri 37377 20562 37378 20563 ne
rect 37378 20562 37622 20563
tri 37378 20561 37379 20562 ne
rect 37379 20561 37622 20562
tri 37379 20560 37380 20561 ne
rect 37380 20560 37622 20561
tri 37380 20559 37381 20560 ne
rect 37381 20559 37622 20560
tri 37381 20558 37382 20559 ne
rect 37382 20558 37622 20559
tri 37382 20557 37383 20558 ne
rect 37383 20557 37622 20558
tri 37383 20556 37384 20557 ne
rect 37384 20556 37622 20557
tri 37384 20555 37385 20556 ne
rect 37385 20555 37622 20556
tri 37385 20554 37386 20555 ne
rect 37386 20554 37622 20555
tri 37386 20553 37387 20554 ne
rect 37387 20553 37622 20554
tri 37387 20552 37388 20553 ne
rect 37388 20552 37622 20553
tri 37388 20551 37389 20552 ne
rect 37389 20551 37622 20552
tri 37389 20550 37390 20551 ne
rect 37390 20550 37622 20551
tri 37390 20549 37391 20550 ne
rect 37391 20549 37622 20550
tri 37622 20549 37667 20594 sw
rect 70802 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
tri 37391 20504 37436 20549 ne
rect 37436 20536 37667 20549
rect 37436 20504 37542 20536
tri 37436 20459 37481 20504 ne
rect 37481 20490 37542 20504
rect 37588 20504 37667 20536
tri 37667 20504 37712 20549 sw
rect 70802 20508 71000 20566
rect 37588 20490 37712 20504
rect 37481 20475 37712 20490
tri 37712 20475 37741 20504 sw
rect 37481 20459 37741 20475
tri 37481 20430 37510 20459 ne
rect 37510 20430 37741 20459
tri 37741 20430 37786 20475 sw
rect 70802 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
tri 37510 20425 37515 20430 ne
rect 37515 20425 37786 20430
tri 37515 20424 37516 20425 ne
rect 37516 20424 37786 20425
tri 37516 20423 37517 20424 ne
rect 37517 20423 37786 20424
tri 37517 20422 37518 20423 ne
rect 37518 20422 37786 20423
tri 37518 20421 37519 20422 ne
rect 37519 20421 37786 20422
tri 37519 20420 37520 20421 ne
rect 37520 20420 37786 20421
tri 37520 20419 37521 20420 ne
rect 37521 20419 37786 20420
tri 37521 20418 37522 20419 ne
rect 37522 20418 37786 20419
tri 37522 20417 37523 20418 ne
rect 37523 20417 37786 20418
tri 37523 20416 37524 20417 ne
rect 37524 20416 37786 20417
tri 37524 20415 37525 20416 ne
rect 37525 20415 37786 20416
tri 37525 20414 37526 20415 ne
rect 37526 20414 37786 20415
tri 37526 20413 37527 20414 ne
rect 37527 20413 37786 20414
tri 37527 20412 37528 20413 ne
rect 37528 20412 37786 20413
tri 37528 20411 37529 20412 ne
rect 37529 20411 37786 20412
tri 37529 20410 37530 20411 ne
rect 37530 20410 37786 20411
tri 37530 20409 37531 20410 ne
rect 37531 20409 37786 20410
tri 37531 20408 37532 20409 ne
rect 37532 20408 37786 20409
tri 37532 20407 37533 20408 ne
rect 37533 20407 37786 20408
tri 37533 20406 37534 20407 ne
rect 37534 20406 37786 20407
tri 37534 20405 37535 20406 ne
rect 37535 20405 37786 20406
tri 37535 20404 37536 20405 ne
rect 37536 20404 37786 20405
tri 37536 20403 37537 20404 ne
rect 37537 20403 37674 20404
tri 37537 20402 37538 20403 ne
rect 37538 20402 37674 20403
tri 37538 20401 37539 20402 ne
rect 37539 20401 37674 20402
tri 37539 20400 37540 20401 ne
rect 37540 20400 37674 20401
tri 37540 20399 37541 20400 ne
rect 37541 20399 37674 20400
tri 37541 20398 37542 20399 ne
rect 37542 20398 37674 20399
tri 37542 20397 37543 20398 ne
rect 37543 20397 37674 20398
tri 37543 20396 37544 20397 ne
rect 37544 20396 37674 20397
tri 37544 20395 37545 20396 ne
rect 37545 20395 37674 20396
tri 37545 20394 37546 20395 ne
rect 37546 20394 37674 20395
tri 37546 20393 37547 20394 ne
rect 37547 20393 37674 20394
tri 37547 20392 37548 20393 ne
rect 37548 20392 37674 20393
tri 37548 20391 37549 20392 ne
rect 37549 20391 37674 20392
tri 37549 20390 37550 20391 ne
rect 37550 20390 37674 20391
tri 37550 20389 37551 20390 ne
rect 37551 20389 37674 20390
tri 37551 20388 37552 20389 ne
rect 37552 20388 37674 20389
tri 37552 20387 37553 20388 ne
rect 37553 20387 37674 20388
tri 37553 20386 37554 20387 ne
rect 37554 20386 37674 20387
tri 37554 20385 37555 20386 ne
rect 37555 20385 37674 20386
tri 37555 20384 37556 20385 ne
rect 37556 20384 37674 20385
tri 37556 20383 37557 20384 ne
rect 37557 20383 37674 20384
tri 37557 20382 37558 20383 ne
rect 37558 20382 37674 20383
tri 37558 20381 37559 20382 ne
rect 37559 20381 37674 20382
tri 37559 20380 37560 20381 ne
rect 37560 20380 37674 20381
tri 37560 20379 37561 20380 ne
rect 37561 20379 37674 20380
tri 37561 20378 37562 20379 ne
rect 37562 20378 37674 20379
tri 37562 20377 37563 20378 ne
rect 37563 20377 37674 20378
tri 37563 20376 37564 20377 ne
rect 37564 20376 37674 20377
tri 37564 20375 37565 20376 ne
rect 37565 20375 37674 20376
tri 37565 20374 37566 20375 ne
rect 37566 20374 37674 20375
tri 37566 20373 37567 20374 ne
rect 37567 20373 37674 20374
tri 37567 20372 37568 20373 ne
rect 37568 20372 37674 20373
tri 37568 20371 37569 20372 ne
rect 37569 20371 37674 20372
tri 37569 20370 37570 20371 ne
rect 37570 20370 37674 20371
tri 37570 20369 37571 20370 ne
rect 37571 20369 37674 20370
tri 37571 20368 37572 20369 ne
rect 37572 20368 37674 20369
tri 37572 20367 37573 20368 ne
rect 37573 20367 37674 20368
tri 37573 20366 37574 20367 ne
rect 37574 20366 37674 20367
tri 37574 20365 37575 20366 ne
rect 37575 20365 37674 20366
tri 37575 20364 37576 20365 ne
rect 37576 20364 37674 20365
tri 37576 20363 37577 20364 ne
rect 37577 20363 37674 20364
tri 37577 20362 37578 20363 ne
rect 37578 20362 37674 20363
tri 37578 20361 37579 20362 ne
rect 37579 20361 37674 20362
tri 37579 20360 37580 20361 ne
rect 37580 20360 37674 20361
tri 37580 20359 37581 20360 ne
rect 37581 20359 37674 20360
tri 37581 20358 37582 20359 ne
rect 37582 20358 37674 20359
rect 37720 20385 37786 20404
tri 37786 20385 37831 20430 sw
rect 70802 20404 71000 20462
rect 37720 20358 37831 20385
tri 37582 20357 37583 20358 ne
rect 37583 20357 37831 20358
tri 37583 20356 37584 20357 ne
rect 37584 20356 37831 20357
tri 37584 20355 37585 20356 ne
rect 37585 20355 37831 20356
tri 37585 20354 37586 20355 ne
rect 37586 20354 37831 20355
tri 37586 20353 37587 20354 ne
rect 37587 20353 37831 20354
tri 37587 20352 37588 20353 ne
rect 37588 20352 37831 20353
tri 37588 20351 37589 20352 ne
rect 37589 20351 37831 20352
tri 37589 20350 37590 20351 ne
rect 37590 20350 37831 20351
tri 37590 20349 37591 20350 ne
rect 37591 20349 37831 20350
tri 37591 20348 37592 20349 ne
rect 37592 20348 37831 20349
tri 37592 20347 37593 20348 ne
rect 37593 20347 37831 20348
tri 37593 20346 37594 20347 ne
rect 37594 20346 37831 20347
tri 37594 20345 37595 20346 ne
rect 37595 20345 37831 20346
tri 37595 20344 37596 20345 ne
rect 37596 20344 37831 20345
tri 37596 20343 37597 20344 ne
rect 37597 20343 37831 20344
tri 37597 20342 37598 20343 ne
rect 37598 20342 37831 20343
tri 37598 20341 37599 20342 ne
rect 37599 20341 37831 20342
tri 37599 20340 37600 20341 ne
rect 37600 20340 37831 20341
tri 37831 20340 37876 20385 sw
rect 70802 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37600 20339 37601 20340 ne
rect 37601 20339 37876 20340
tri 37601 20338 37602 20339 ne
rect 37602 20338 37876 20339
tri 37602 20337 37603 20338 ne
rect 37603 20337 37876 20338
tri 37603 20336 37604 20337 ne
rect 37604 20336 37876 20337
tri 37604 20335 37605 20336 ne
rect 37605 20335 37876 20336
tri 37605 20334 37606 20335 ne
rect 37606 20334 37876 20335
tri 37606 20333 37607 20334 ne
rect 37607 20333 37876 20334
tri 37607 20332 37608 20333 ne
rect 37608 20332 37876 20333
tri 37608 20331 37609 20332 ne
rect 37609 20331 37876 20332
tri 37609 20330 37610 20331 ne
rect 37610 20330 37876 20331
tri 37610 20329 37611 20330 ne
rect 37611 20329 37876 20330
tri 37611 20328 37612 20329 ne
rect 37612 20328 37876 20329
tri 37612 20327 37613 20328 ne
rect 37613 20327 37876 20328
tri 37613 20326 37614 20327 ne
rect 37614 20326 37876 20327
tri 37614 20325 37615 20326 ne
rect 37615 20325 37876 20326
tri 37615 20324 37616 20325 ne
rect 37616 20324 37876 20325
tri 37616 20323 37617 20324 ne
rect 37617 20323 37876 20324
tri 37617 20322 37618 20323 ne
rect 37618 20322 37876 20323
tri 37618 20321 37619 20322 ne
rect 37619 20321 37876 20322
tri 37619 20320 37620 20321 ne
rect 37620 20320 37876 20321
tri 37620 20319 37621 20320 ne
rect 37621 20319 37876 20320
tri 37621 20318 37622 20319 ne
rect 37622 20318 37876 20319
tri 37876 20318 37898 20340 sw
tri 37622 20317 37623 20318 ne
rect 37623 20317 37898 20318
tri 37623 20316 37624 20317 ne
rect 37624 20316 37898 20317
tri 37624 20315 37625 20316 ne
rect 37625 20315 37898 20316
tri 37625 20314 37626 20315 ne
rect 37626 20314 37898 20315
tri 37626 20313 37627 20314 ne
rect 37627 20313 37898 20314
tri 37627 20312 37628 20313 ne
rect 37628 20312 37898 20313
tri 37628 20311 37629 20312 ne
rect 37629 20311 37898 20312
tri 37629 20310 37630 20311 ne
rect 37630 20310 37898 20311
tri 37630 20309 37631 20310 ne
rect 37631 20309 37898 20310
tri 37631 20308 37632 20309 ne
rect 37632 20308 37898 20309
tri 37632 20307 37633 20308 ne
rect 37633 20307 37898 20308
tri 37633 20306 37634 20307 ne
rect 37634 20306 37898 20307
tri 37634 20305 37635 20306 ne
rect 37635 20305 37898 20306
tri 37635 20304 37636 20305 ne
rect 37636 20304 37898 20305
tri 37636 20303 37637 20304 ne
rect 37637 20303 37898 20304
tri 37637 20302 37638 20303 ne
rect 37638 20302 37898 20303
tri 37638 20301 37639 20302 ne
rect 37639 20301 37898 20302
tri 37639 20300 37640 20301 ne
rect 37640 20300 37898 20301
tri 37640 20299 37641 20300 ne
rect 37641 20299 37898 20300
tri 37641 20298 37642 20299 ne
rect 37642 20298 37898 20299
tri 37642 20297 37643 20298 ne
rect 37643 20297 37898 20298
tri 37643 20296 37644 20297 ne
rect 37644 20296 37898 20297
tri 37644 20295 37645 20296 ne
rect 37645 20295 37898 20296
tri 37645 20294 37646 20295 ne
rect 37646 20294 37898 20295
tri 37646 20293 37647 20294 ne
rect 37647 20293 37898 20294
tri 37647 20292 37648 20293 ne
rect 37648 20292 37898 20293
tri 37648 20291 37649 20292 ne
rect 37649 20291 37898 20292
tri 37649 20290 37650 20291 ne
rect 37650 20290 37898 20291
tri 37650 20289 37651 20290 ne
rect 37651 20289 37898 20290
tri 37651 20288 37652 20289 ne
rect 37652 20288 37898 20289
tri 37652 20287 37653 20288 ne
rect 37653 20287 37898 20288
tri 37653 20286 37654 20287 ne
rect 37654 20286 37898 20287
tri 37654 20285 37655 20286 ne
rect 37655 20285 37898 20286
tri 37655 20284 37656 20285 ne
rect 37656 20284 37898 20285
tri 37656 20283 37657 20284 ne
rect 37657 20283 37898 20284
tri 37657 20282 37658 20283 ne
rect 37658 20282 37898 20283
tri 37658 20281 37659 20282 ne
rect 37659 20281 37898 20282
tri 37659 20280 37660 20281 ne
rect 37660 20280 37898 20281
tri 37660 20279 37661 20280 ne
rect 37661 20279 37898 20280
tri 37661 20278 37662 20279 ne
rect 37662 20278 37898 20279
tri 37662 20277 37663 20278 ne
rect 37663 20277 37898 20278
tri 37663 20276 37664 20277 ne
rect 37664 20276 37898 20277
tri 37664 20275 37665 20276 ne
rect 37665 20275 37898 20276
tri 37665 20274 37666 20275 ne
rect 37666 20274 37898 20275
tri 37666 20273 37667 20274 ne
rect 37667 20273 37898 20274
tri 37898 20273 37943 20318 sw
rect 70802 20300 71000 20358
tri 37667 20228 37712 20273 ne
rect 37712 20272 37943 20273
rect 37712 20228 37806 20272
tri 37712 20183 37757 20228 ne
rect 37757 20226 37806 20228
rect 37852 20228 37943 20272
tri 37943 20228 37988 20273 sw
rect 70802 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20226 37988 20228
rect 37757 20183 37988 20226
tri 37988 20183 38033 20228 sw
rect 70802 20196 71000 20254
tri 37757 20151 37789 20183 ne
rect 37789 20154 38033 20183
tri 38033 20154 38062 20183 sw
rect 37789 20151 38062 20154
tri 37789 20150 37790 20151 ne
rect 37790 20150 38062 20151
tri 37790 20149 37791 20150 ne
rect 37791 20149 38062 20150
tri 37791 20148 37792 20149 ne
rect 37792 20148 38062 20149
tri 37792 20147 37793 20148 ne
rect 37793 20147 38062 20148
tri 37793 20146 37794 20147 ne
rect 37794 20146 38062 20147
tri 37794 20145 37795 20146 ne
rect 37795 20145 38062 20146
tri 37795 20144 37796 20145 ne
rect 37796 20144 38062 20145
tri 37796 20143 37797 20144 ne
rect 37797 20143 38062 20144
tri 37797 20142 37798 20143 ne
rect 37798 20142 38062 20143
tri 37798 20141 37799 20142 ne
rect 37799 20141 38062 20142
tri 37799 20140 37800 20141 ne
rect 37800 20140 38062 20141
tri 37800 20139 37801 20140 ne
rect 37801 20139 37938 20140
tri 37801 20138 37802 20139 ne
rect 37802 20138 37938 20139
tri 37802 20137 37803 20138 ne
rect 37803 20137 37938 20138
tri 37803 20136 37804 20137 ne
rect 37804 20136 37938 20137
tri 37804 20135 37805 20136 ne
rect 37805 20135 37938 20136
tri 37805 20134 37806 20135 ne
rect 37806 20134 37938 20135
tri 37806 20133 37807 20134 ne
rect 37807 20133 37938 20134
tri 37807 20132 37808 20133 ne
rect 37808 20132 37938 20133
tri 37808 20131 37809 20132 ne
rect 37809 20131 37938 20132
tri 37809 20130 37810 20131 ne
rect 37810 20130 37938 20131
tri 37810 20129 37811 20130 ne
rect 37811 20129 37938 20130
tri 37811 20128 37812 20129 ne
rect 37812 20128 37938 20129
tri 37812 20127 37813 20128 ne
rect 37813 20127 37938 20128
tri 37813 20126 37814 20127 ne
rect 37814 20126 37938 20127
tri 37814 20125 37815 20126 ne
rect 37815 20125 37938 20126
tri 37815 20124 37816 20125 ne
rect 37816 20124 37938 20125
tri 37816 20123 37817 20124 ne
rect 37817 20123 37938 20124
tri 37817 20122 37818 20123 ne
rect 37818 20122 37938 20123
tri 37818 20121 37819 20122 ne
rect 37819 20121 37938 20122
tri 37819 20120 37820 20121 ne
rect 37820 20120 37938 20121
tri 37820 20119 37821 20120 ne
rect 37821 20119 37938 20120
tri 37821 20118 37822 20119 ne
rect 37822 20118 37938 20119
tri 37822 20117 37823 20118 ne
rect 37823 20117 37938 20118
tri 37823 20116 37824 20117 ne
rect 37824 20116 37938 20117
tri 37824 20115 37825 20116 ne
rect 37825 20115 37938 20116
tri 37825 20114 37826 20115 ne
rect 37826 20114 37938 20115
tri 37826 20113 37827 20114 ne
rect 37827 20113 37938 20114
tri 37827 20112 37828 20113 ne
rect 37828 20112 37938 20113
tri 37828 20111 37829 20112 ne
rect 37829 20111 37938 20112
tri 37829 20110 37830 20111 ne
rect 37830 20110 37938 20111
tri 37830 20109 37831 20110 ne
rect 37831 20109 37938 20110
tri 37831 20108 37832 20109 ne
rect 37832 20108 37938 20109
tri 37832 20107 37833 20108 ne
rect 37833 20107 37938 20108
tri 37833 20106 37834 20107 ne
rect 37834 20106 37938 20107
tri 37834 20105 37835 20106 ne
rect 37835 20105 37938 20106
tri 37835 20104 37836 20105 ne
rect 37836 20104 37938 20105
tri 37836 20103 37837 20104 ne
rect 37837 20103 37938 20104
tri 37837 20102 37838 20103 ne
rect 37838 20102 37938 20103
tri 37838 20101 37839 20102 ne
rect 37839 20101 37938 20102
tri 37839 20100 37840 20101 ne
rect 37840 20100 37938 20101
tri 37840 20099 37841 20100 ne
rect 37841 20099 37938 20100
tri 37841 20098 37842 20099 ne
rect 37842 20098 37938 20099
tri 37842 20097 37843 20098 ne
rect 37843 20097 37938 20098
tri 37843 20096 37844 20097 ne
rect 37844 20096 37938 20097
tri 37844 20095 37845 20096 ne
rect 37845 20095 37938 20096
tri 37845 20094 37846 20095 ne
rect 37846 20094 37938 20095
rect 37984 20109 38062 20140
tri 38062 20109 38107 20154 sw
rect 70802 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 37984 20094 38107 20109
tri 37846 20093 37847 20094 ne
rect 37847 20093 38107 20094
tri 37847 20092 37848 20093 ne
rect 37848 20092 38107 20093
tri 37848 20091 37849 20092 ne
rect 37849 20091 38107 20092
tri 37849 20090 37850 20091 ne
rect 37850 20090 38107 20091
tri 37850 20089 37851 20090 ne
rect 37851 20089 38107 20090
tri 37851 20088 37852 20089 ne
rect 37852 20088 38107 20089
tri 37852 20087 37853 20088 ne
rect 37853 20087 38107 20088
tri 37853 20086 37854 20087 ne
rect 37854 20086 38107 20087
tri 37854 20085 37855 20086 ne
rect 37855 20085 38107 20086
tri 37855 20084 37856 20085 ne
rect 37856 20084 38107 20085
tri 37856 20083 37857 20084 ne
rect 37857 20083 38107 20084
tri 37857 20082 37858 20083 ne
rect 37858 20082 38107 20083
tri 37858 20081 37859 20082 ne
rect 37859 20081 38107 20082
tri 37859 20080 37860 20081 ne
rect 37860 20080 38107 20081
tri 37860 20079 37861 20080 ne
rect 37861 20079 38107 20080
tri 37861 20078 37862 20079 ne
rect 37862 20078 38107 20079
tri 37862 20077 37863 20078 ne
rect 37863 20077 38107 20078
tri 37863 20076 37864 20077 ne
rect 37864 20076 38107 20077
tri 37864 20075 37865 20076 ne
rect 37865 20075 38107 20076
tri 37865 20074 37866 20075 ne
rect 37866 20074 38107 20075
tri 37866 20073 37867 20074 ne
rect 37867 20073 38107 20074
tri 37867 20072 37868 20073 ne
rect 37868 20072 38107 20073
tri 37868 20071 37869 20072 ne
rect 37869 20071 38107 20072
tri 37869 20070 37870 20071 ne
rect 37870 20070 38107 20071
tri 37870 20069 37871 20070 ne
rect 37871 20069 38107 20070
tri 37871 20068 37872 20069 ne
rect 37872 20068 38107 20069
tri 37872 20067 37873 20068 ne
rect 37873 20067 38107 20068
tri 37873 20066 37874 20067 ne
rect 37874 20066 38107 20067
tri 37874 20065 37875 20066 ne
rect 37875 20065 38107 20066
tri 37875 20064 37876 20065 ne
rect 37876 20064 38107 20065
tri 38107 20064 38152 20109 sw
rect 70802 20092 71000 20150
tri 37876 20063 37877 20064 ne
rect 37877 20063 38152 20064
tri 37877 20062 37878 20063 ne
rect 37878 20062 38152 20063
tri 37878 20061 37879 20062 ne
rect 37879 20061 38152 20062
tri 37879 20060 37880 20061 ne
rect 37880 20060 38152 20061
tri 37880 20059 37881 20060 ne
rect 37881 20059 38152 20060
tri 37881 20058 37882 20059 ne
rect 37882 20058 38152 20059
tri 37882 20057 37883 20058 ne
rect 37883 20057 38152 20058
tri 37883 20056 37884 20057 ne
rect 37884 20056 38152 20057
tri 37884 20055 37885 20056 ne
rect 37885 20055 38152 20056
tri 37885 20054 37886 20055 ne
rect 37886 20054 38152 20055
tri 37886 20053 37887 20054 ne
rect 37887 20053 38152 20054
tri 37887 20052 37888 20053 ne
rect 37888 20052 38152 20053
tri 37888 20051 37889 20052 ne
rect 37889 20051 38152 20052
tri 37889 20050 37890 20051 ne
rect 37890 20050 38152 20051
tri 37890 20049 37891 20050 ne
rect 37891 20049 38152 20050
tri 37891 20048 37892 20049 ne
rect 37892 20048 38152 20049
tri 37892 20047 37893 20048 ne
rect 37893 20047 38152 20048
tri 37893 20046 37894 20047 ne
rect 37894 20046 38152 20047
tri 37894 20045 37895 20046 ne
rect 37895 20045 38152 20046
tri 37895 20044 37896 20045 ne
rect 37896 20044 38152 20045
tri 37896 20043 37897 20044 ne
rect 37897 20043 38152 20044
tri 37897 20042 37898 20043 ne
rect 37898 20042 38152 20043
tri 37898 20041 37899 20042 ne
rect 37899 20041 38152 20042
tri 37899 20040 37900 20041 ne
rect 37900 20040 38152 20041
tri 37900 20039 37901 20040 ne
rect 37901 20039 38152 20040
tri 37901 20038 37902 20039 ne
rect 37902 20038 38152 20039
tri 37902 20037 37903 20038 ne
rect 37903 20037 38152 20038
tri 37903 20036 37904 20037 ne
rect 37904 20036 38152 20037
tri 37904 20035 37905 20036 ne
rect 37905 20035 38152 20036
tri 37905 20034 37906 20035 ne
rect 37906 20034 38152 20035
tri 37906 20033 37907 20034 ne
rect 37907 20033 38152 20034
tri 37907 20032 37908 20033 ne
rect 37908 20032 38152 20033
tri 37908 20031 37909 20032 ne
rect 37909 20031 38152 20032
tri 37909 20030 37910 20031 ne
rect 37910 20030 38152 20031
tri 37910 20029 37911 20030 ne
rect 37911 20029 38152 20030
tri 37911 20028 37912 20029 ne
rect 37912 20028 38152 20029
tri 37912 20027 37913 20028 ne
rect 37913 20027 38152 20028
tri 37913 20026 37914 20027 ne
rect 37914 20026 38152 20027
tri 37914 20025 37915 20026 ne
rect 37915 20025 38152 20026
tri 37915 20024 37916 20025 ne
rect 37916 20024 38152 20025
tri 37916 20023 37917 20024 ne
rect 37917 20023 38152 20024
tri 37917 20022 37918 20023 ne
rect 37918 20022 38152 20023
tri 37918 20021 37919 20022 ne
rect 37919 20021 38152 20022
tri 37919 20020 37920 20021 ne
rect 37920 20020 38152 20021
tri 37920 20019 37921 20020 ne
rect 37921 20019 38152 20020
tri 38152 20019 38197 20064 sw
rect 70802 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37921 20018 37922 20019 ne
rect 37922 20018 38197 20019
tri 37922 20017 37923 20018 ne
rect 37923 20017 38197 20018
tri 37923 20016 37924 20017 ne
rect 37924 20016 38197 20017
tri 37924 20015 37925 20016 ne
rect 37925 20015 38197 20016
tri 37925 20014 37926 20015 ne
rect 37926 20014 38197 20015
tri 37926 20013 37927 20014 ne
rect 37927 20013 38197 20014
tri 37927 20012 37928 20013 ne
rect 37928 20012 38197 20013
tri 37928 20011 37929 20012 ne
rect 37929 20011 38197 20012
tri 37929 20010 37930 20011 ne
rect 37930 20010 38197 20011
tri 37930 20009 37931 20010 ne
rect 37931 20009 38197 20010
tri 37931 20008 37932 20009 ne
rect 37932 20008 38197 20009
tri 37932 20007 37933 20008 ne
rect 37933 20007 38070 20008
tri 37933 20006 37934 20007 ne
rect 37934 20006 38070 20007
tri 37934 20005 37935 20006 ne
rect 37935 20005 38070 20006
tri 37935 20004 37936 20005 ne
rect 37936 20004 38070 20005
tri 37936 20003 37937 20004 ne
rect 37937 20003 38070 20004
tri 37937 20002 37938 20003 ne
rect 37938 20002 38070 20003
tri 37938 20001 37939 20002 ne
rect 37939 20001 38070 20002
tri 37939 20000 37940 20001 ne
rect 37940 20000 38070 20001
tri 37940 19999 37941 20000 ne
rect 37941 19999 38070 20000
tri 37941 19998 37942 19999 ne
rect 37942 19998 38070 19999
tri 37942 19997 37943 19998 ne
rect 37943 19997 38070 19998
tri 37943 19952 37988 19997 ne
rect 37988 19962 38070 19997
rect 38116 19997 38197 20008
tri 38197 19997 38219 20019 sw
rect 38116 19974 38219 19997
tri 38219 19974 38242 19997 sw
rect 70802 19988 71000 20046
rect 38116 19962 38242 19974
rect 37988 19952 38242 19962
tri 37988 19934 38006 19952 ne
rect 38006 19934 38242 19952
tri 38006 19889 38051 19934 ne
rect 38051 19929 38242 19934
tri 38242 19929 38287 19974 sw
rect 70802 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 38051 19889 38287 19929
tri 38051 19877 38063 19889 ne
rect 38063 19884 38287 19889
tri 38287 19884 38332 19929 sw
rect 70802 19884 71000 19942
rect 38063 19877 38332 19884
tri 38063 19876 38064 19877 ne
rect 38064 19876 38332 19877
tri 38064 19875 38065 19876 ne
rect 38065 19875 38202 19876
tri 38065 19874 38066 19875 ne
rect 38066 19874 38202 19875
tri 38066 19873 38067 19874 ne
rect 38067 19873 38202 19874
tri 38067 19872 38068 19873 ne
rect 38068 19872 38202 19873
tri 38068 19871 38069 19872 ne
rect 38069 19871 38202 19872
tri 38069 19870 38070 19871 ne
rect 38070 19870 38202 19871
tri 38070 19869 38071 19870 ne
rect 38071 19869 38202 19870
tri 38071 19868 38072 19869 ne
rect 38072 19868 38202 19869
tri 38072 19867 38073 19868 ne
rect 38073 19867 38202 19868
tri 38073 19866 38074 19867 ne
rect 38074 19866 38202 19867
tri 38074 19865 38075 19866 ne
rect 38075 19865 38202 19866
tri 38075 19864 38076 19865 ne
rect 38076 19864 38202 19865
tri 38076 19863 38077 19864 ne
rect 38077 19863 38202 19864
tri 38077 19862 38078 19863 ne
rect 38078 19862 38202 19863
tri 38078 19861 38079 19862 ne
rect 38079 19861 38202 19862
tri 38079 19860 38080 19861 ne
rect 38080 19860 38202 19861
tri 38080 19859 38081 19860 ne
rect 38081 19859 38202 19860
tri 38081 19858 38082 19859 ne
rect 38082 19858 38202 19859
tri 38082 19857 38083 19858 ne
rect 38083 19857 38202 19858
tri 38083 19856 38084 19857 ne
rect 38084 19856 38202 19857
tri 38084 19855 38085 19856 ne
rect 38085 19855 38202 19856
tri 38085 19854 38086 19855 ne
rect 38086 19854 38202 19855
tri 38086 19853 38087 19854 ne
rect 38087 19853 38202 19854
tri 38087 19852 38088 19853 ne
rect 38088 19852 38202 19853
tri 38088 19851 38089 19852 ne
rect 38089 19851 38202 19852
tri 38089 19850 38090 19851 ne
rect 38090 19850 38202 19851
tri 38090 19849 38091 19850 ne
rect 38091 19849 38202 19850
tri 38091 19848 38092 19849 ne
rect 38092 19848 38202 19849
tri 38092 19847 38093 19848 ne
rect 38093 19847 38202 19848
tri 38093 19846 38094 19847 ne
rect 38094 19846 38202 19847
tri 38094 19845 38095 19846 ne
rect 38095 19845 38202 19846
tri 38095 19844 38096 19845 ne
rect 38096 19844 38202 19845
tri 38096 19843 38097 19844 ne
rect 38097 19843 38202 19844
tri 38097 19842 38098 19843 ne
rect 38098 19842 38202 19843
tri 38098 19841 38099 19842 ne
rect 38099 19841 38202 19842
tri 38099 19840 38100 19841 ne
rect 38100 19840 38202 19841
tri 38100 19839 38101 19840 ne
rect 38101 19839 38202 19840
tri 38101 19838 38102 19839 ne
rect 38102 19838 38202 19839
tri 38102 19837 38103 19838 ne
rect 38103 19837 38202 19838
tri 38103 19836 38104 19837 ne
rect 38104 19836 38202 19837
tri 38104 19835 38105 19836 ne
rect 38105 19835 38202 19836
tri 38105 19834 38106 19835 ne
rect 38106 19834 38202 19835
tri 38106 19833 38107 19834 ne
rect 38107 19833 38202 19834
tri 38107 19832 38108 19833 ne
rect 38108 19832 38202 19833
tri 38108 19831 38109 19832 ne
rect 38109 19831 38202 19832
tri 38109 19830 38110 19831 ne
rect 38110 19830 38202 19831
rect 38248 19856 38332 19876
tri 38332 19856 38360 19884 sw
rect 38248 19830 38360 19856
tri 38110 19829 38111 19830 ne
rect 38111 19829 38360 19830
tri 38111 19828 38112 19829 ne
rect 38112 19828 38360 19829
tri 38112 19827 38113 19828 ne
rect 38113 19827 38360 19828
tri 38113 19826 38114 19827 ne
rect 38114 19826 38360 19827
tri 38114 19825 38115 19826 ne
rect 38115 19825 38360 19826
tri 38115 19824 38116 19825 ne
rect 38116 19824 38360 19825
tri 38116 19823 38117 19824 ne
rect 38117 19823 38360 19824
tri 38117 19822 38118 19823 ne
rect 38118 19822 38360 19823
tri 38118 19821 38119 19822 ne
rect 38119 19821 38360 19822
tri 38119 19820 38120 19821 ne
rect 38120 19820 38360 19821
tri 38120 19819 38121 19820 ne
rect 38121 19819 38360 19820
tri 38121 19818 38122 19819 ne
rect 38122 19818 38360 19819
tri 38122 19817 38123 19818 ne
rect 38123 19817 38360 19818
tri 38123 19816 38124 19817 ne
rect 38124 19816 38360 19817
tri 38124 19815 38125 19816 ne
rect 38125 19815 38360 19816
tri 38125 19814 38126 19815 ne
rect 38126 19814 38360 19815
tri 38126 19813 38127 19814 ne
rect 38127 19813 38360 19814
tri 38127 19812 38128 19813 ne
rect 38128 19812 38360 19813
tri 38128 19811 38129 19812 ne
rect 38129 19811 38360 19812
tri 38360 19811 38405 19856 sw
rect 70802 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
tri 38129 19810 38130 19811 ne
rect 38130 19810 38405 19811
tri 38130 19809 38131 19810 ne
rect 38131 19809 38405 19810
tri 38131 19808 38132 19809 ne
rect 38132 19808 38405 19809
tri 38132 19807 38133 19808 ne
rect 38133 19807 38405 19808
tri 38133 19806 38134 19807 ne
rect 38134 19806 38405 19807
tri 38134 19805 38135 19806 ne
rect 38135 19805 38405 19806
tri 38135 19804 38136 19805 ne
rect 38136 19804 38405 19805
tri 38136 19803 38137 19804 ne
rect 38137 19803 38405 19804
tri 38137 19802 38138 19803 ne
rect 38138 19802 38405 19803
tri 38138 19801 38139 19802 ne
rect 38139 19801 38405 19802
tri 38139 19800 38140 19801 ne
rect 38140 19800 38405 19801
tri 38140 19799 38141 19800 ne
rect 38141 19799 38405 19800
tri 38141 19798 38142 19799 ne
rect 38142 19798 38405 19799
tri 38142 19797 38143 19798 ne
rect 38143 19797 38405 19798
tri 38143 19796 38144 19797 ne
rect 38144 19796 38405 19797
tri 38144 19795 38145 19796 ne
rect 38145 19795 38405 19796
tri 38145 19794 38146 19795 ne
rect 38146 19794 38405 19795
tri 38146 19793 38147 19794 ne
rect 38147 19793 38405 19794
tri 38147 19792 38148 19793 ne
rect 38148 19792 38405 19793
tri 38148 19791 38149 19792 ne
rect 38149 19791 38405 19792
tri 38149 19790 38150 19791 ne
rect 38150 19790 38405 19791
tri 38150 19789 38151 19790 ne
rect 38151 19789 38405 19790
tri 38151 19788 38152 19789 ne
rect 38152 19788 38405 19789
tri 38152 19787 38153 19788 ne
rect 38153 19787 38405 19788
tri 38153 19786 38154 19787 ne
rect 38154 19786 38405 19787
tri 38154 19785 38155 19786 ne
rect 38155 19785 38405 19786
tri 38155 19784 38156 19785 ne
rect 38156 19784 38405 19785
tri 38156 19783 38157 19784 ne
rect 38157 19783 38405 19784
tri 38157 19782 38158 19783 ne
rect 38158 19782 38405 19783
tri 38158 19781 38159 19782 ne
rect 38159 19781 38405 19782
tri 38159 19780 38160 19781 ne
rect 38160 19780 38405 19781
tri 38160 19779 38161 19780 ne
rect 38161 19779 38405 19780
tri 38161 19778 38162 19779 ne
rect 38162 19778 38405 19779
tri 38162 19777 38163 19778 ne
rect 38163 19777 38405 19778
tri 38163 19776 38164 19777 ne
rect 38164 19776 38405 19777
tri 38164 19775 38165 19776 ne
rect 38165 19775 38405 19776
tri 38165 19774 38166 19775 ne
rect 38166 19774 38405 19775
tri 38166 19773 38167 19774 ne
rect 38167 19773 38405 19774
tri 38167 19772 38168 19773 ne
rect 38168 19772 38405 19773
tri 38168 19771 38169 19772 ne
rect 38169 19771 38405 19772
tri 38169 19770 38170 19771 ne
rect 38170 19770 38405 19771
tri 38170 19769 38171 19770 ne
rect 38171 19769 38405 19770
tri 38171 19768 38172 19769 ne
rect 38172 19768 38405 19769
tri 38172 19767 38173 19768 ne
rect 38173 19767 38405 19768
tri 38173 19766 38174 19767 ne
rect 38174 19766 38405 19767
tri 38405 19766 38450 19811 sw
rect 70802 19780 71000 19838
tri 38174 19765 38175 19766 ne
rect 38175 19765 38450 19766
tri 38175 19764 38176 19765 ne
rect 38176 19764 38450 19765
tri 38176 19763 38177 19764 ne
rect 38177 19763 38450 19764
tri 38177 19762 38178 19763 ne
rect 38178 19762 38450 19763
tri 38178 19761 38179 19762 ne
rect 38179 19761 38450 19762
tri 38179 19760 38180 19761 ne
rect 38180 19760 38450 19761
tri 38180 19759 38181 19760 ne
rect 38181 19759 38450 19760
tri 38181 19758 38182 19759 ne
rect 38182 19758 38450 19759
tri 38182 19757 38183 19758 ne
rect 38183 19757 38450 19758
tri 38183 19756 38184 19757 ne
rect 38184 19756 38450 19757
tri 38184 19755 38185 19756 ne
rect 38185 19755 38450 19756
tri 38185 19754 38186 19755 ne
rect 38186 19754 38450 19755
tri 38186 19753 38187 19754 ne
rect 38187 19753 38450 19754
tri 38187 19752 38188 19753 ne
rect 38188 19752 38450 19753
tri 38188 19751 38189 19752 ne
rect 38189 19751 38450 19752
tri 38189 19750 38190 19751 ne
rect 38190 19750 38450 19751
tri 38190 19749 38191 19750 ne
rect 38191 19749 38450 19750
tri 38191 19748 38192 19749 ne
rect 38192 19748 38450 19749
tri 38192 19747 38193 19748 ne
rect 38193 19747 38450 19748
tri 38193 19746 38194 19747 ne
rect 38194 19746 38450 19747
tri 38194 19745 38195 19746 ne
rect 38195 19745 38450 19746
tri 38195 19744 38196 19745 ne
rect 38196 19744 38450 19745
tri 38196 19743 38197 19744 ne
rect 38197 19743 38334 19744
tri 38197 19742 38198 19743 ne
rect 38198 19742 38334 19743
tri 38198 19741 38199 19742 ne
rect 38199 19741 38334 19742
tri 38199 19740 38200 19741 ne
rect 38200 19740 38334 19741
tri 38200 19739 38201 19740 ne
rect 38201 19739 38334 19740
tri 38201 19738 38202 19739 ne
rect 38202 19738 38334 19739
tri 38202 19737 38203 19738 ne
rect 38203 19737 38334 19738
tri 38203 19736 38204 19737 ne
rect 38204 19736 38334 19737
tri 38204 19735 38205 19736 ne
rect 38205 19735 38334 19736
tri 38205 19734 38206 19735 ne
rect 38206 19734 38334 19735
tri 38206 19733 38207 19734 ne
rect 38207 19733 38334 19734
tri 38207 19732 38208 19733 ne
rect 38208 19732 38334 19733
tri 38208 19731 38209 19732 ne
rect 38209 19731 38334 19732
tri 38209 19730 38210 19731 ne
rect 38210 19730 38334 19731
tri 38210 19729 38211 19730 ne
rect 38211 19729 38334 19730
tri 38211 19728 38212 19729 ne
rect 38212 19728 38334 19729
tri 38212 19727 38213 19728 ne
rect 38213 19727 38334 19728
tri 38213 19726 38214 19727 ne
rect 38214 19726 38334 19727
tri 38214 19725 38215 19726 ne
rect 38215 19725 38334 19726
tri 38215 19724 38216 19725 ne
rect 38216 19724 38334 19725
tri 38216 19723 38217 19724 ne
rect 38217 19723 38334 19724
tri 38217 19722 38218 19723 ne
rect 38218 19722 38334 19723
tri 38218 19721 38219 19722 ne
rect 38219 19721 38334 19722
tri 38219 19698 38242 19721 ne
rect 38242 19698 38334 19721
rect 38380 19721 38450 19744
tri 38450 19721 38495 19766 sw
rect 70802 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 38380 19698 38495 19721
tri 38495 19698 38518 19721 sw
tri 38242 19676 38264 19698 ne
rect 38264 19676 38518 19698
tri 38264 19653 38287 19676 ne
rect 38287 19653 38518 19676
tri 38518 19653 38563 19698 sw
rect 70802 19676 71000 19734
tri 38287 19608 38332 19653 ne
rect 38332 19612 38563 19653
rect 38332 19608 38466 19612
tri 38332 19602 38338 19608 ne
rect 38338 19602 38466 19608
tri 38338 19601 38339 19602 ne
rect 38339 19601 38466 19602
tri 38339 19600 38340 19601 ne
rect 38340 19600 38466 19601
tri 38340 19599 38341 19600 ne
rect 38341 19599 38466 19600
tri 38341 19598 38342 19599 ne
rect 38342 19598 38466 19599
tri 38342 19597 38343 19598 ne
rect 38343 19597 38466 19598
tri 38343 19596 38344 19597 ne
rect 38344 19596 38466 19597
tri 38344 19595 38345 19596 ne
rect 38345 19595 38466 19596
tri 38345 19594 38346 19595 ne
rect 38346 19594 38466 19595
tri 38346 19593 38347 19594 ne
rect 38347 19593 38466 19594
tri 38347 19592 38348 19593 ne
rect 38348 19592 38466 19593
tri 38348 19591 38349 19592 ne
rect 38349 19591 38466 19592
tri 38349 19590 38350 19591 ne
rect 38350 19590 38466 19591
tri 38350 19589 38351 19590 ne
rect 38351 19589 38466 19590
tri 38351 19588 38352 19589 ne
rect 38352 19588 38466 19589
tri 38352 19587 38353 19588 ne
rect 38353 19587 38466 19588
tri 38353 19586 38354 19587 ne
rect 38354 19586 38466 19587
tri 38354 19585 38355 19586 ne
rect 38355 19585 38466 19586
tri 38355 19584 38356 19585 ne
rect 38356 19584 38466 19585
tri 38356 19583 38357 19584 ne
rect 38357 19583 38466 19584
tri 38357 19582 38358 19583 ne
rect 38358 19582 38466 19583
tri 38358 19581 38359 19582 ne
rect 38359 19581 38466 19582
tri 38359 19580 38360 19581 ne
rect 38360 19580 38466 19581
tri 38360 19579 38361 19580 ne
rect 38361 19579 38466 19580
tri 38361 19578 38362 19579 ne
rect 38362 19578 38466 19579
tri 38362 19577 38363 19578 ne
rect 38363 19577 38466 19578
tri 38363 19576 38364 19577 ne
rect 38364 19576 38466 19577
tri 38364 19575 38365 19576 ne
rect 38365 19575 38466 19576
tri 38365 19574 38366 19575 ne
rect 38366 19574 38466 19575
tri 38366 19573 38367 19574 ne
rect 38367 19573 38466 19574
tri 38367 19572 38368 19573 ne
rect 38368 19572 38466 19573
tri 38368 19571 38369 19572 ne
rect 38369 19571 38466 19572
tri 38369 19570 38370 19571 ne
rect 38370 19570 38466 19571
tri 38370 19569 38371 19570 ne
rect 38371 19569 38466 19570
tri 38371 19568 38372 19569 ne
rect 38372 19568 38466 19569
tri 38372 19567 38373 19568 ne
rect 38373 19567 38466 19568
tri 38373 19566 38374 19567 ne
rect 38374 19566 38466 19567
rect 38512 19608 38563 19612
tri 38563 19608 38608 19653 sw
rect 70802 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38512 19566 38608 19608
tri 38374 19565 38375 19566 ne
rect 38375 19565 38608 19566
tri 38375 19564 38376 19565 ne
rect 38376 19564 38608 19565
tri 38376 19563 38377 19564 ne
rect 38377 19563 38608 19564
tri 38608 19563 38653 19608 sw
rect 70802 19572 71000 19630
tri 38377 19562 38378 19563 ne
rect 38378 19562 38653 19563
tri 38378 19561 38379 19562 ne
rect 38379 19561 38653 19562
tri 38379 19560 38380 19561 ne
rect 38380 19560 38653 19561
tri 38380 19559 38381 19560 ne
rect 38381 19559 38653 19560
tri 38381 19558 38382 19559 ne
rect 38382 19558 38653 19559
tri 38382 19557 38383 19558 ne
rect 38383 19557 38653 19558
tri 38383 19556 38384 19557 ne
rect 38384 19556 38653 19557
tri 38384 19555 38385 19556 ne
rect 38385 19555 38653 19556
tri 38385 19554 38386 19555 ne
rect 38386 19554 38653 19555
tri 38386 19553 38387 19554 ne
rect 38387 19553 38653 19554
tri 38387 19552 38388 19553 ne
rect 38388 19552 38653 19553
tri 38388 19551 38389 19552 ne
rect 38389 19551 38653 19552
tri 38389 19550 38390 19551 ne
rect 38390 19550 38653 19551
tri 38390 19549 38391 19550 ne
rect 38391 19549 38653 19550
tri 38391 19548 38392 19549 ne
rect 38392 19548 38653 19549
tri 38392 19547 38393 19548 ne
rect 38393 19547 38653 19548
tri 38393 19546 38394 19547 ne
rect 38394 19546 38653 19547
tri 38394 19545 38395 19546 ne
rect 38395 19545 38653 19546
tri 38395 19544 38396 19545 ne
rect 38396 19544 38653 19545
tri 38396 19543 38397 19544 ne
rect 38397 19543 38653 19544
tri 38397 19542 38398 19543 ne
rect 38398 19542 38653 19543
tri 38398 19541 38399 19542 ne
rect 38399 19541 38653 19542
tri 38399 19540 38400 19541 ne
rect 38400 19540 38653 19541
tri 38400 19539 38401 19540 ne
rect 38401 19539 38653 19540
tri 38401 19538 38402 19539 ne
rect 38402 19538 38653 19539
tri 38402 19537 38403 19538 ne
rect 38403 19537 38653 19538
tri 38403 19536 38404 19537 ne
rect 38404 19536 38653 19537
tri 38404 19535 38405 19536 ne
rect 38405 19535 38653 19536
tri 38653 19535 38681 19563 sw
tri 38405 19534 38406 19535 ne
rect 38406 19534 38681 19535
tri 38406 19533 38407 19534 ne
rect 38407 19533 38681 19534
tri 38407 19532 38408 19533 ne
rect 38408 19532 38681 19533
tri 38408 19531 38409 19532 ne
rect 38409 19531 38681 19532
tri 38409 19530 38410 19531 ne
rect 38410 19530 38681 19531
tri 38410 19529 38411 19530 ne
rect 38411 19529 38681 19530
tri 38411 19528 38412 19529 ne
rect 38412 19528 38681 19529
tri 38412 19527 38413 19528 ne
rect 38413 19527 38681 19528
tri 38413 19526 38414 19527 ne
rect 38414 19526 38681 19527
tri 38414 19525 38415 19526 ne
rect 38415 19525 38681 19526
tri 38415 19524 38416 19525 ne
rect 38416 19524 38681 19525
tri 38416 19523 38417 19524 ne
rect 38417 19523 38681 19524
tri 38417 19522 38418 19523 ne
rect 38418 19522 38681 19523
tri 38418 19521 38419 19522 ne
rect 38419 19521 38681 19522
tri 38419 19520 38420 19521 ne
rect 38420 19520 38681 19521
tri 38420 19519 38421 19520 ne
rect 38421 19519 38681 19520
tri 38421 19518 38422 19519 ne
rect 38422 19518 38681 19519
tri 38422 19517 38423 19518 ne
rect 38423 19517 38681 19518
tri 38423 19516 38424 19517 ne
rect 38424 19516 38681 19517
tri 38424 19515 38425 19516 ne
rect 38425 19515 38681 19516
tri 38425 19514 38426 19515 ne
rect 38426 19514 38681 19515
tri 38426 19513 38427 19514 ne
rect 38427 19513 38681 19514
tri 38427 19512 38428 19513 ne
rect 38428 19512 38681 19513
tri 38428 19511 38429 19512 ne
rect 38429 19511 38681 19512
tri 38429 19510 38430 19511 ne
rect 38430 19510 38681 19511
tri 38430 19509 38431 19510 ne
rect 38431 19509 38681 19510
tri 38431 19508 38432 19509 ne
rect 38432 19508 38681 19509
tri 38432 19507 38433 19508 ne
rect 38433 19507 38681 19508
tri 38433 19506 38434 19507 ne
rect 38434 19506 38681 19507
tri 38434 19505 38435 19506 ne
rect 38435 19505 38681 19506
tri 38435 19504 38436 19505 ne
rect 38436 19504 38681 19505
tri 38436 19503 38437 19504 ne
rect 38437 19503 38681 19504
tri 38437 19502 38438 19503 ne
rect 38438 19502 38681 19503
tri 38438 19501 38439 19502 ne
rect 38439 19501 38681 19502
tri 38439 19500 38440 19501 ne
rect 38440 19500 38681 19501
tri 38440 19499 38441 19500 ne
rect 38441 19499 38681 19500
tri 38441 19498 38442 19499 ne
rect 38442 19498 38681 19499
tri 38442 19497 38443 19498 ne
rect 38443 19497 38681 19498
tri 38443 19496 38444 19497 ne
rect 38444 19496 38681 19497
tri 38444 19495 38445 19496 ne
rect 38445 19495 38681 19496
tri 38445 19494 38446 19495 ne
rect 38446 19494 38681 19495
tri 38446 19493 38447 19494 ne
rect 38447 19493 38681 19494
tri 38447 19492 38448 19493 ne
rect 38448 19492 38681 19493
tri 38448 19491 38449 19492 ne
rect 38449 19491 38681 19492
tri 38449 19490 38450 19491 ne
rect 38450 19490 38681 19491
tri 38681 19490 38726 19535 sw
rect 70802 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38450 19489 38451 19490 ne
rect 38451 19489 38726 19490
tri 38451 19488 38452 19489 ne
rect 38452 19488 38726 19489
tri 38452 19487 38453 19488 ne
rect 38453 19487 38726 19488
tri 38453 19486 38454 19487 ne
rect 38454 19486 38726 19487
tri 38454 19485 38455 19486 ne
rect 38455 19485 38726 19486
tri 38455 19484 38456 19485 ne
rect 38456 19484 38726 19485
tri 38456 19483 38457 19484 ne
rect 38457 19483 38726 19484
tri 38457 19482 38458 19483 ne
rect 38458 19482 38726 19483
tri 38458 19481 38459 19482 ne
rect 38459 19481 38726 19482
tri 38459 19480 38460 19481 ne
rect 38460 19480 38726 19481
tri 38460 19479 38461 19480 ne
rect 38461 19479 38598 19480
tri 38461 19478 38462 19479 ne
rect 38462 19478 38598 19479
tri 38462 19477 38463 19478 ne
rect 38463 19477 38598 19478
tri 38463 19476 38464 19477 ne
rect 38464 19476 38598 19477
tri 38464 19475 38465 19476 ne
rect 38465 19475 38598 19476
tri 38465 19474 38466 19475 ne
rect 38466 19474 38598 19475
tri 38466 19473 38467 19474 ne
rect 38467 19473 38598 19474
tri 38467 19472 38468 19473 ne
rect 38468 19472 38598 19473
tri 38468 19471 38469 19472 ne
rect 38469 19471 38598 19472
tri 38469 19470 38470 19471 ne
rect 38470 19470 38598 19471
tri 38470 19469 38471 19470 ne
rect 38471 19469 38598 19470
tri 38471 19468 38472 19469 ne
rect 38472 19468 38598 19469
tri 38472 19467 38473 19468 ne
rect 38473 19467 38598 19468
tri 38473 19466 38474 19467 ne
rect 38474 19466 38598 19467
tri 38474 19465 38475 19466 ne
rect 38475 19465 38598 19466
tri 38475 19464 38476 19465 ne
rect 38476 19464 38598 19465
tri 38476 19463 38477 19464 ne
rect 38477 19463 38598 19464
tri 38477 19462 38478 19463 ne
rect 38478 19462 38598 19463
tri 38478 19461 38479 19462 ne
rect 38479 19461 38598 19462
tri 38479 19460 38480 19461 ne
rect 38480 19460 38598 19461
tri 38480 19459 38481 19460 ne
rect 38481 19459 38598 19460
tri 38481 19458 38482 19459 ne
rect 38482 19458 38598 19459
tri 38482 19457 38483 19458 ne
rect 38483 19457 38598 19458
tri 38483 19456 38484 19457 ne
rect 38484 19456 38598 19457
tri 38484 19455 38485 19456 ne
rect 38485 19455 38598 19456
tri 38485 19454 38486 19455 ne
rect 38486 19454 38598 19455
tri 38486 19453 38487 19454 ne
rect 38487 19453 38598 19454
tri 38487 19452 38488 19453 ne
rect 38488 19452 38598 19453
tri 38488 19451 38489 19452 ne
rect 38489 19451 38598 19452
tri 38489 19450 38490 19451 ne
rect 38490 19450 38598 19451
tri 38490 19449 38491 19450 ne
rect 38491 19449 38598 19450
tri 38491 19448 38492 19449 ne
rect 38492 19448 38598 19449
tri 38492 19447 38493 19448 ne
rect 38493 19447 38598 19448
tri 38493 19446 38494 19447 ne
rect 38494 19446 38598 19447
tri 38494 19445 38495 19446 ne
rect 38495 19445 38598 19446
tri 38495 19400 38540 19445 ne
rect 38540 19434 38598 19445
rect 38644 19445 38726 19480
tri 38726 19445 38771 19490 sw
rect 70802 19468 71000 19526
rect 38644 19434 38771 19445
rect 38540 19400 38771 19434
tri 38771 19400 38816 19445 sw
rect 70802 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
tri 38540 19355 38585 19400 ne
rect 38585 19377 38816 19400
tri 38816 19377 38839 19400 sw
rect 38585 19355 38839 19377
tri 38585 19332 38608 19355 ne
rect 38608 19348 38839 19355
rect 38608 19332 38730 19348
tri 38608 19328 38612 19332 ne
rect 38612 19328 38730 19332
tri 38612 19327 38613 19328 ne
rect 38613 19327 38730 19328
tri 38613 19326 38614 19327 ne
rect 38614 19326 38730 19327
tri 38614 19325 38615 19326 ne
rect 38615 19325 38730 19326
tri 38615 19324 38616 19325 ne
rect 38616 19324 38730 19325
tri 38616 19323 38617 19324 ne
rect 38617 19323 38730 19324
tri 38617 19322 38618 19323 ne
rect 38618 19322 38730 19323
tri 38618 19321 38619 19322 ne
rect 38619 19321 38730 19322
tri 38619 19320 38620 19321 ne
rect 38620 19320 38730 19321
tri 38620 19319 38621 19320 ne
rect 38621 19319 38730 19320
tri 38621 19318 38622 19319 ne
rect 38622 19318 38730 19319
tri 38622 19317 38623 19318 ne
rect 38623 19317 38730 19318
tri 38623 19316 38624 19317 ne
rect 38624 19316 38730 19317
tri 38624 19315 38625 19316 ne
rect 38625 19315 38730 19316
tri 38625 19314 38626 19315 ne
rect 38626 19314 38730 19315
tri 38626 19313 38627 19314 ne
rect 38627 19313 38730 19314
tri 38627 19312 38628 19313 ne
rect 38628 19312 38730 19313
tri 38628 19311 38629 19312 ne
rect 38629 19311 38730 19312
tri 38629 19310 38630 19311 ne
rect 38630 19310 38730 19311
tri 38630 19309 38631 19310 ne
rect 38631 19309 38730 19310
tri 38631 19308 38632 19309 ne
rect 38632 19308 38730 19309
tri 38632 19307 38633 19308 ne
rect 38633 19307 38730 19308
tri 38633 19306 38634 19307 ne
rect 38634 19306 38730 19307
tri 38634 19305 38635 19306 ne
rect 38635 19305 38730 19306
tri 38635 19304 38636 19305 ne
rect 38636 19304 38730 19305
tri 38636 19303 38637 19304 ne
rect 38637 19303 38730 19304
tri 38637 19302 38638 19303 ne
rect 38638 19302 38730 19303
rect 38776 19332 38839 19348
tri 38839 19332 38884 19377 sw
rect 70802 19364 71000 19422
rect 38776 19302 38884 19332
tri 38638 19301 38639 19302 ne
rect 38639 19301 38884 19302
tri 38639 19300 38640 19301 ne
rect 38640 19300 38884 19301
tri 38640 19299 38641 19300 ne
rect 38641 19299 38884 19300
tri 38641 19298 38642 19299 ne
rect 38642 19298 38884 19299
tri 38642 19297 38643 19298 ne
rect 38643 19297 38884 19298
tri 38643 19296 38644 19297 ne
rect 38644 19296 38884 19297
tri 38644 19295 38645 19296 ne
rect 38645 19295 38884 19296
tri 38645 19294 38646 19295 ne
rect 38646 19294 38884 19295
tri 38646 19293 38647 19294 ne
rect 38647 19293 38884 19294
tri 38647 19292 38648 19293 ne
rect 38648 19292 38884 19293
tri 38648 19291 38649 19292 ne
rect 38649 19291 38884 19292
tri 38649 19290 38650 19291 ne
rect 38650 19290 38884 19291
tri 38650 19289 38651 19290 ne
rect 38651 19289 38884 19290
tri 38651 19288 38652 19289 ne
rect 38652 19288 38884 19289
tri 38652 19287 38653 19288 ne
rect 38653 19287 38884 19288
tri 38884 19287 38929 19332 sw
rect 70802 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
tri 38653 19286 38654 19287 ne
rect 38654 19286 38929 19287
tri 38654 19285 38655 19286 ne
rect 38655 19285 38929 19286
tri 38655 19284 38656 19285 ne
rect 38656 19284 38929 19285
tri 38656 19283 38657 19284 ne
rect 38657 19283 38929 19284
tri 38657 19282 38658 19283 ne
rect 38658 19282 38929 19283
tri 38658 19281 38659 19282 ne
rect 38659 19281 38929 19282
tri 38659 19280 38660 19281 ne
rect 38660 19280 38929 19281
tri 38660 19279 38661 19280 ne
rect 38661 19279 38929 19280
tri 38661 19278 38662 19279 ne
rect 38662 19278 38929 19279
tri 38662 19277 38663 19278 ne
rect 38663 19277 38929 19278
tri 38663 19276 38664 19277 ne
rect 38664 19276 38929 19277
tri 38664 19275 38665 19276 ne
rect 38665 19275 38929 19276
tri 38665 19274 38666 19275 ne
rect 38666 19274 38929 19275
tri 38666 19273 38667 19274 ne
rect 38667 19273 38929 19274
tri 38667 19272 38668 19273 ne
rect 38668 19272 38929 19273
tri 38668 19271 38669 19272 ne
rect 38669 19271 38929 19272
tri 38669 19270 38670 19271 ne
rect 38670 19270 38929 19271
tri 38670 19269 38671 19270 ne
rect 38671 19269 38929 19270
tri 38671 19268 38672 19269 ne
rect 38672 19268 38929 19269
tri 38672 19267 38673 19268 ne
rect 38673 19267 38929 19268
tri 38673 19266 38674 19267 ne
rect 38674 19266 38929 19267
tri 38674 19265 38675 19266 ne
rect 38675 19265 38929 19266
tri 38675 19264 38676 19265 ne
rect 38676 19264 38929 19265
tri 38676 19263 38677 19264 ne
rect 38677 19263 38929 19264
tri 38677 19262 38678 19263 ne
rect 38678 19262 38929 19263
tri 38678 19261 38679 19262 ne
rect 38679 19261 38929 19262
tri 38679 19260 38680 19261 ne
rect 38680 19260 38929 19261
tri 38680 19259 38681 19260 ne
rect 38681 19259 38929 19260
tri 38681 19258 38682 19259 ne
rect 38682 19258 38929 19259
tri 38682 19257 38683 19258 ne
rect 38683 19257 38929 19258
tri 38683 19256 38684 19257 ne
rect 38684 19256 38929 19257
tri 38684 19255 38685 19256 ne
rect 38685 19255 38929 19256
tri 38685 19254 38686 19255 ne
rect 38686 19254 38929 19255
tri 38686 19253 38687 19254 ne
rect 38687 19253 38929 19254
tri 38687 19252 38688 19253 ne
rect 38688 19252 38929 19253
tri 38688 19251 38689 19252 ne
rect 38689 19251 38929 19252
tri 38689 19250 38690 19251 ne
rect 38690 19250 38929 19251
tri 38690 19249 38691 19250 ne
rect 38691 19249 38929 19250
tri 38691 19248 38692 19249 ne
rect 38692 19248 38929 19249
tri 38692 19247 38693 19248 ne
rect 38693 19247 38929 19248
tri 38693 19246 38694 19247 ne
rect 38694 19246 38929 19247
tri 38694 19245 38695 19246 ne
rect 38695 19245 38929 19246
tri 38695 19244 38696 19245 ne
rect 38696 19244 38929 19245
tri 38696 19243 38697 19244 ne
rect 38697 19243 38929 19244
tri 38697 19242 38698 19243 ne
rect 38698 19242 38929 19243
tri 38929 19242 38974 19287 sw
rect 70802 19260 71000 19318
tri 38698 19241 38699 19242 ne
rect 38699 19241 38974 19242
tri 38699 19240 38700 19241 ne
rect 38700 19240 38974 19241
tri 38700 19239 38701 19240 ne
rect 38701 19239 38974 19240
tri 38701 19238 38702 19239 ne
rect 38702 19238 38974 19239
tri 38702 19237 38703 19238 ne
rect 38703 19237 38974 19238
tri 38703 19236 38704 19237 ne
rect 38704 19236 38974 19237
tri 38704 19235 38705 19236 ne
rect 38705 19235 38974 19236
tri 38705 19234 38706 19235 ne
rect 38706 19234 38974 19235
tri 38706 19233 38707 19234 ne
rect 38707 19233 38974 19234
tri 38707 19232 38708 19233 ne
rect 38708 19232 38974 19233
tri 38708 19231 38709 19232 ne
rect 38709 19231 38974 19232
tri 38709 19230 38710 19231 ne
rect 38710 19230 38974 19231
tri 38710 19229 38711 19230 ne
rect 38711 19229 38974 19230
tri 38711 19228 38712 19229 ne
rect 38712 19228 38974 19229
tri 38712 19227 38713 19228 ne
rect 38713 19227 38974 19228
tri 38713 19226 38714 19227 ne
rect 38714 19226 38974 19227
tri 38714 19225 38715 19226 ne
rect 38715 19225 38974 19226
tri 38715 19224 38716 19225 ne
rect 38716 19224 38974 19225
tri 38716 19223 38717 19224 ne
rect 38717 19223 38974 19224
tri 38717 19222 38718 19223 ne
rect 38718 19222 38974 19223
tri 38718 19221 38719 19222 ne
rect 38719 19221 38974 19222
tri 38719 19220 38720 19221 ne
rect 38720 19220 38974 19221
tri 38720 19219 38721 19220 ne
rect 38721 19219 38974 19220
tri 38721 19218 38722 19219 ne
rect 38722 19218 38974 19219
tri 38722 19217 38723 19218 ne
rect 38723 19217 38974 19218
tri 38723 19216 38724 19217 ne
rect 38724 19216 38974 19217
tri 38724 19215 38725 19216 ne
rect 38725 19215 38862 19216
tri 38725 19214 38726 19215 ne
rect 38726 19214 38862 19215
tri 38726 19213 38727 19214 ne
rect 38727 19213 38862 19214
tri 38727 19212 38728 19213 ne
rect 38728 19212 38862 19213
tri 38728 19211 38729 19212 ne
rect 38729 19211 38862 19212
tri 38729 19210 38730 19211 ne
rect 38730 19210 38862 19211
tri 38730 19209 38731 19210 ne
rect 38731 19209 38862 19210
tri 38731 19208 38732 19209 ne
rect 38732 19208 38862 19209
tri 38732 19207 38733 19208 ne
rect 38733 19207 38862 19208
tri 38733 19206 38734 19207 ne
rect 38734 19206 38862 19207
tri 38734 19205 38735 19206 ne
rect 38735 19205 38862 19206
tri 38735 19204 38736 19205 ne
rect 38736 19204 38862 19205
tri 38736 19203 38737 19204 ne
rect 38737 19203 38862 19204
tri 38737 19202 38738 19203 ne
rect 38738 19202 38862 19203
tri 38738 19201 38739 19202 ne
rect 38739 19201 38862 19202
tri 38739 19200 38740 19201 ne
rect 38740 19200 38862 19201
tri 38740 19199 38741 19200 ne
rect 38741 19199 38862 19200
tri 38741 19198 38742 19199 ne
rect 38742 19198 38862 19199
tri 38742 19197 38743 19198 ne
rect 38743 19197 38862 19198
tri 38743 19196 38744 19197 ne
rect 38744 19196 38862 19197
tri 38744 19195 38745 19196 ne
rect 38745 19195 38862 19196
tri 38745 19194 38746 19195 ne
rect 38746 19194 38862 19195
tri 38746 19193 38747 19194 ne
rect 38747 19193 38862 19194
tri 38747 19192 38748 19193 ne
rect 38748 19192 38862 19193
tri 38748 19191 38749 19192 ne
rect 38749 19191 38862 19192
tri 38749 19190 38750 19191 ne
rect 38750 19190 38862 19191
tri 38750 19189 38751 19190 ne
rect 38751 19189 38862 19190
tri 38751 19188 38752 19189 ne
rect 38752 19188 38862 19189
tri 38752 19187 38753 19188 ne
rect 38753 19187 38862 19188
tri 38753 19186 38754 19187 ne
rect 38754 19186 38862 19187
tri 38754 19185 38755 19186 ne
rect 38755 19185 38862 19186
tri 38755 19184 38756 19185 ne
rect 38756 19184 38862 19185
tri 38756 19183 38757 19184 ne
rect 38757 19183 38862 19184
tri 38757 19182 38758 19183 ne
rect 38758 19182 38862 19183
tri 38758 19181 38759 19182 ne
rect 38759 19181 38862 19182
tri 38759 19180 38760 19181 ne
rect 38760 19180 38862 19181
tri 38760 19179 38761 19180 ne
rect 38761 19179 38862 19180
tri 38761 19178 38762 19179 ne
rect 38762 19178 38862 19179
tri 38762 19177 38763 19178 ne
rect 38763 19177 38862 19178
tri 38763 19176 38764 19177 ne
rect 38764 19176 38862 19177
tri 38764 19175 38765 19176 ne
rect 38765 19175 38862 19176
tri 38765 19174 38766 19175 ne
rect 38766 19174 38862 19175
tri 38766 19173 38767 19174 ne
rect 38767 19173 38862 19174
tri 38767 19172 38768 19173 ne
rect 38768 19172 38862 19173
tri 38768 19171 38769 19172 ne
rect 38769 19171 38862 19172
tri 38769 19170 38770 19171 ne
rect 38770 19170 38862 19171
rect 38908 19214 38974 19216
tri 38974 19214 39002 19242 sw
rect 70802 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19170 39002 19214
tri 38770 19169 38771 19170 ne
rect 38771 19169 39002 19170
tri 39002 19169 39047 19214 sw
tri 38771 19124 38816 19169 ne
rect 38816 19124 39047 19169
tri 39047 19124 39092 19169 sw
rect 70802 19156 71000 19214
tri 38816 19079 38861 19124 ne
rect 38861 19084 39092 19124
rect 38861 19079 38994 19084
tri 38861 19053 38887 19079 ne
rect 38887 19053 38994 19079
tri 38887 19052 38888 19053 ne
rect 38888 19052 38994 19053
tri 38888 19051 38889 19052 ne
rect 38889 19051 38994 19052
tri 38889 19050 38890 19051 ne
rect 38890 19050 38994 19051
tri 38890 19049 38891 19050 ne
rect 38891 19049 38994 19050
tri 38891 19048 38892 19049 ne
rect 38892 19048 38994 19049
tri 38892 19047 38893 19048 ne
rect 38893 19047 38994 19048
tri 38893 19046 38894 19047 ne
rect 38894 19046 38994 19047
tri 38894 19045 38895 19046 ne
rect 38895 19045 38994 19046
tri 38895 19044 38896 19045 ne
rect 38896 19044 38994 19045
tri 38896 19043 38897 19044 ne
rect 38897 19043 38994 19044
tri 38897 19042 38898 19043 ne
rect 38898 19042 38994 19043
tri 38898 19041 38899 19042 ne
rect 38899 19041 38994 19042
tri 38899 19040 38900 19041 ne
rect 38900 19040 38994 19041
tri 38900 19039 38901 19040 ne
rect 38901 19039 38994 19040
tri 38901 19038 38902 19039 ne
rect 38902 19038 38994 19039
rect 39040 19079 39092 19084
tri 39092 19079 39137 19124 sw
rect 70802 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 39040 19056 39137 19079
tri 39137 19056 39160 19079 sw
rect 39040 19038 39160 19056
tri 38902 19037 38903 19038 ne
rect 38903 19037 39160 19038
tri 38903 19036 38904 19037 ne
rect 38904 19036 39160 19037
tri 38904 19035 38905 19036 ne
rect 38905 19035 39160 19036
tri 38905 19034 38906 19035 ne
rect 38906 19034 39160 19035
tri 38906 19033 38907 19034 ne
rect 38907 19033 39160 19034
tri 38907 19032 38908 19033 ne
rect 38908 19032 39160 19033
tri 38908 19031 38909 19032 ne
rect 38909 19031 39160 19032
tri 38909 19030 38910 19031 ne
rect 38910 19030 39160 19031
tri 38910 19029 38911 19030 ne
rect 38911 19029 39160 19030
tri 38911 19028 38912 19029 ne
rect 38912 19028 39160 19029
tri 38912 19027 38913 19028 ne
rect 38913 19027 39160 19028
tri 38913 19026 38914 19027 ne
rect 38914 19026 39160 19027
tri 38914 19025 38915 19026 ne
rect 38915 19025 39160 19026
tri 38915 19024 38916 19025 ne
rect 38916 19024 39160 19025
tri 38916 19023 38917 19024 ne
rect 38917 19023 39160 19024
tri 38917 19022 38918 19023 ne
rect 38918 19022 39160 19023
tri 38918 19021 38919 19022 ne
rect 38919 19021 39160 19022
tri 38919 19020 38920 19021 ne
rect 38920 19020 39160 19021
tri 38920 19019 38921 19020 ne
rect 38921 19019 39160 19020
tri 38921 19018 38922 19019 ne
rect 38922 19018 39160 19019
tri 38922 19017 38923 19018 ne
rect 38923 19017 39160 19018
tri 38923 19016 38924 19017 ne
rect 38924 19016 39160 19017
tri 38924 19015 38925 19016 ne
rect 38925 19015 39160 19016
tri 38925 19014 38926 19015 ne
rect 38926 19014 39160 19015
tri 38926 19013 38927 19014 ne
rect 38927 19013 39160 19014
tri 38927 19012 38928 19013 ne
rect 38928 19012 39160 19013
tri 38928 19011 38929 19012 ne
rect 38929 19011 39160 19012
tri 39160 19011 39205 19056 sw
rect 70802 19052 71000 19110
tri 38929 19010 38930 19011 ne
rect 38930 19010 39205 19011
tri 38930 19009 38931 19010 ne
rect 38931 19009 39205 19010
tri 38931 19008 38932 19009 ne
rect 38932 19008 39205 19009
tri 38932 19007 38933 19008 ne
rect 38933 19007 39205 19008
tri 38933 19006 38934 19007 ne
rect 38934 19006 39205 19007
tri 38934 19005 38935 19006 ne
rect 38935 19005 39205 19006
tri 38935 19004 38936 19005 ne
rect 38936 19004 39205 19005
tri 38936 19003 38937 19004 ne
rect 38937 19003 39205 19004
tri 38937 19002 38938 19003 ne
rect 38938 19002 39205 19003
tri 38938 19001 38939 19002 ne
rect 38939 19001 39205 19002
tri 38939 19000 38940 19001 ne
rect 38940 19000 39205 19001
tri 38940 18999 38941 19000 ne
rect 38941 18999 39205 19000
tri 38941 18998 38942 18999 ne
rect 38942 18998 39205 18999
tri 38942 18997 38943 18998 ne
rect 38943 18997 39205 18998
tri 38943 18996 38944 18997 ne
rect 38944 18996 39205 18997
tri 38944 18995 38945 18996 ne
rect 38945 18995 39205 18996
tri 38945 18994 38946 18995 ne
rect 38946 18994 39205 18995
tri 38946 18993 38947 18994 ne
rect 38947 18993 39205 18994
tri 38947 18992 38948 18993 ne
rect 38948 18992 39205 18993
tri 38948 18991 38949 18992 ne
rect 38949 18991 39205 18992
tri 38949 18990 38950 18991 ne
rect 38950 18990 39205 18991
tri 38950 18989 38951 18990 ne
rect 38951 18989 39205 18990
tri 38951 18988 38952 18989 ne
rect 38952 18988 39205 18989
tri 38952 18987 38953 18988 ne
rect 38953 18987 39205 18988
tri 38953 18986 38954 18987 ne
rect 38954 18986 39205 18987
tri 38954 18985 38955 18986 ne
rect 38955 18985 39205 18986
tri 38955 18984 38956 18985 ne
rect 38956 18984 39205 18985
tri 38956 18983 38957 18984 ne
rect 38957 18983 39205 18984
tri 38957 18982 38958 18983 ne
rect 38958 18982 39205 18983
tri 38958 18981 38959 18982 ne
rect 38959 18981 39205 18982
tri 38959 18980 38960 18981 ne
rect 38960 18980 39205 18981
tri 38960 18979 38961 18980 ne
rect 38961 18979 39205 18980
tri 38961 18978 38962 18979 ne
rect 38962 18978 39205 18979
tri 38962 18977 38963 18978 ne
rect 38963 18977 39205 18978
tri 38963 18976 38964 18977 ne
rect 38964 18976 39205 18977
tri 38964 18975 38965 18976 ne
rect 38965 18975 39205 18976
tri 38965 18974 38966 18975 ne
rect 38966 18974 39205 18975
tri 38966 18973 38967 18974 ne
rect 38967 18973 39205 18974
tri 38967 18972 38968 18973 ne
rect 38968 18972 39205 18973
tri 38968 18971 38969 18972 ne
rect 38969 18971 39205 18972
tri 38969 18970 38970 18971 ne
rect 38970 18970 39205 18971
tri 38970 18969 38971 18970 ne
rect 38971 18969 39205 18970
tri 38971 18968 38972 18969 ne
rect 38972 18968 39205 18969
tri 38972 18967 38973 18968 ne
rect 38973 18967 39205 18968
tri 38973 18966 38974 18967 ne
rect 38974 18966 39205 18967
tri 39205 18966 39250 19011 sw
rect 70802 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
tri 38974 18965 38975 18966 ne
rect 38975 18965 39250 18966
tri 38975 18964 38976 18965 ne
rect 38976 18964 39250 18965
tri 38976 18963 38977 18964 ne
rect 38977 18963 39250 18964
tri 38977 18962 38978 18963 ne
rect 38978 18962 39250 18963
tri 38978 18961 38979 18962 ne
rect 38979 18961 39250 18962
tri 38979 18960 38980 18961 ne
rect 38980 18960 39250 18961
tri 38980 18959 38981 18960 ne
rect 38981 18959 39250 18960
tri 38981 18958 38982 18959 ne
rect 38982 18958 39250 18959
tri 38982 18957 38983 18958 ne
rect 38983 18957 39250 18958
tri 38983 18956 38984 18957 ne
rect 38984 18956 39250 18957
tri 38984 18955 38985 18956 ne
rect 38985 18955 39250 18956
tri 38985 18954 38986 18955 ne
rect 38986 18954 39250 18955
tri 38986 18953 38987 18954 ne
rect 38987 18953 39250 18954
tri 38987 18952 38988 18953 ne
rect 38988 18952 39250 18953
tri 38988 18951 38989 18952 ne
rect 38989 18951 39126 18952
tri 38989 18950 38990 18951 ne
rect 38990 18950 39126 18951
tri 38990 18949 38991 18950 ne
rect 38991 18949 39126 18950
tri 38991 18948 38992 18949 ne
rect 38992 18948 39126 18949
tri 38992 18947 38993 18948 ne
rect 38993 18947 39126 18948
tri 38993 18946 38994 18947 ne
rect 38994 18946 39126 18947
tri 38994 18945 38995 18946 ne
rect 38995 18945 39126 18946
tri 38995 18944 38996 18945 ne
rect 38996 18944 39126 18945
tri 38996 18943 38997 18944 ne
rect 38997 18943 39126 18944
tri 38997 18942 38998 18943 ne
rect 38998 18942 39126 18943
tri 38998 18941 38999 18942 ne
rect 38999 18941 39126 18942
tri 38999 18940 39000 18941 ne
rect 39000 18940 39126 18941
tri 39000 18939 39001 18940 ne
rect 39001 18939 39126 18940
tri 39001 18938 39002 18939 ne
rect 39002 18938 39126 18939
tri 39002 18937 39003 18938 ne
rect 39003 18937 39126 18938
tri 39003 18936 39004 18937 ne
rect 39004 18936 39126 18937
tri 39004 18935 39005 18936 ne
rect 39005 18935 39126 18936
tri 39005 18934 39006 18935 ne
rect 39006 18934 39126 18935
tri 39006 18933 39007 18934 ne
rect 39007 18933 39126 18934
tri 39007 18932 39008 18933 ne
rect 39008 18932 39126 18933
tri 39008 18931 39009 18932 ne
rect 39009 18931 39126 18932
tri 39009 18930 39010 18931 ne
rect 39010 18930 39126 18931
tri 39010 18929 39011 18930 ne
rect 39011 18929 39126 18930
tri 39011 18928 39012 18929 ne
rect 39012 18928 39126 18929
tri 39012 18927 39013 18928 ne
rect 39013 18927 39126 18928
tri 39013 18926 39014 18927 ne
rect 39014 18926 39126 18927
tri 39014 18925 39015 18926 ne
rect 39015 18925 39126 18926
tri 39015 18924 39016 18925 ne
rect 39016 18924 39126 18925
tri 39016 18923 39017 18924 ne
rect 39017 18923 39126 18924
tri 39017 18922 39018 18923 ne
rect 39018 18922 39126 18923
tri 39018 18921 39019 18922 ne
rect 39019 18921 39126 18922
tri 39019 18920 39020 18921 ne
rect 39020 18920 39126 18921
tri 39020 18919 39021 18920 ne
rect 39021 18919 39126 18920
tri 39021 18918 39022 18919 ne
rect 39022 18918 39126 18919
tri 39022 18917 39023 18918 ne
rect 39023 18917 39126 18918
tri 39023 18916 39024 18917 ne
rect 39024 18916 39126 18917
tri 39024 18915 39025 18916 ne
rect 39025 18915 39126 18916
tri 39025 18914 39026 18915 ne
rect 39026 18914 39126 18915
tri 39026 18913 39027 18914 ne
rect 39027 18913 39126 18914
tri 39027 18912 39028 18913 ne
rect 39028 18912 39126 18913
tri 39028 18911 39029 18912 ne
rect 39029 18911 39126 18912
tri 39029 18910 39030 18911 ne
rect 39030 18910 39126 18911
tri 39030 18909 39031 18910 ne
rect 39031 18909 39126 18910
tri 39031 18908 39032 18909 ne
rect 39032 18908 39126 18909
tri 39032 18907 39033 18908 ne
rect 39033 18907 39126 18908
tri 39033 18906 39034 18907 ne
rect 39034 18906 39126 18907
rect 39172 18921 39250 18952
tri 39250 18921 39295 18966 sw
rect 70802 18948 71000 19006
rect 39172 18906 39295 18921
tri 39034 18905 39035 18906 ne
rect 39035 18905 39295 18906
tri 39035 18904 39036 18905 ne
rect 39036 18904 39295 18905
tri 39036 18903 39037 18904 ne
rect 39037 18903 39295 18904
tri 39037 18902 39038 18903 ne
rect 39038 18902 39295 18903
tri 39038 18901 39039 18902 ne
rect 39039 18901 39295 18902
tri 39039 18900 39040 18901 ne
rect 39040 18900 39295 18901
tri 39040 18899 39041 18900 ne
rect 39041 18899 39295 18900
tri 39041 18898 39042 18899 ne
rect 39042 18898 39295 18899
tri 39042 18897 39043 18898 ne
rect 39043 18897 39295 18898
tri 39043 18896 39044 18897 ne
rect 39044 18896 39295 18897
tri 39044 18895 39045 18896 ne
rect 39045 18895 39295 18896
tri 39045 18894 39046 18895 ne
rect 39046 18894 39295 18895
tri 39046 18893 39047 18894 ne
rect 39047 18893 39295 18894
tri 39295 18893 39323 18921 sw
rect 70802 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
tri 39047 18848 39092 18893 ne
rect 39092 18876 39323 18893
tri 39323 18876 39340 18893 sw
rect 39092 18848 39340 18876
tri 39092 18840 39100 18848 ne
rect 39100 18840 39340 18848
tri 39100 18795 39145 18840 ne
rect 39145 18831 39340 18840
tri 39340 18831 39385 18876 sw
rect 70802 18844 71000 18902
rect 39145 18820 39385 18831
rect 39145 18795 39258 18820
tri 39145 18779 39161 18795 ne
rect 39161 18779 39258 18795
tri 39161 18778 39162 18779 ne
rect 39162 18778 39258 18779
tri 39162 18777 39163 18778 ne
rect 39163 18777 39258 18778
tri 39163 18776 39164 18777 ne
rect 39164 18776 39258 18777
tri 39164 18775 39165 18776 ne
rect 39165 18775 39258 18776
tri 39165 18774 39166 18775 ne
rect 39166 18774 39258 18775
rect 39304 18786 39385 18820
tri 39385 18786 39430 18831 sw
rect 70802 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18774 39430 18786
tri 39166 18773 39167 18774 ne
rect 39167 18773 39430 18774
tri 39167 18772 39168 18773 ne
rect 39168 18772 39430 18773
tri 39168 18771 39169 18772 ne
rect 39169 18771 39430 18772
tri 39169 18770 39170 18771 ne
rect 39170 18770 39430 18771
tri 39170 18769 39171 18770 ne
rect 39171 18769 39430 18770
tri 39171 18768 39172 18769 ne
rect 39172 18768 39430 18769
tri 39172 18767 39173 18768 ne
rect 39173 18767 39430 18768
tri 39173 18766 39174 18767 ne
rect 39174 18766 39430 18767
tri 39174 18765 39175 18766 ne
rect 39175 18765 39430 18766
tri 39175 18764 39176 18765 ne
rect 39176 18764 39430 18765
tri 39176 18763 39177 18764 ne
rect 39177 18763 39430 18764
tri 39177 18762 39178 18763 ne
rect 39178 18762 39430 18763
tri 39178 18761 39179 18762 ne
rect 39179 18761 39430 18762
tri 39179 18760 39180 18761 ne
rect 39180 18760 39430 18761
tri 39180 18759 39181 18760 ne
rect 39181 18759 39430 18760
tri 39181 18758 39182 18759 ne
rect 39182 18758 39430 18759
tri 39182 18757 39183 18758 ne
rect 39183 18757 39430 18758
tri 39183 18756 39184 18757 ne
rect 39184 18756 39430 18757
tri 39184 18755 39185 18756 ne
rect 39185 18755 39430 18756
tri 39185 18754 39186 18755 ne
rect 39186 18754 39430 18755
tri 39186 18753 39187 18754 ne
rect 39187 18753 39430 18754
tri 39187 18752 39188 18753 ne
rect 39188 18752 39430 18753
tri 39430 18752 39464 18786 sw
tri 39188 18751 39189 18752 ne
rect 39189 18751 39464 18752
tri 39189 18750 39190 18751 ne
rect 39190 18750 39464 18751
tri 39190 18749 39191 18750 ne
rect 39191 18749 39464 18750
tri 39191 18748 39192 18749 ne
rect 39192 18748 39464 18749
tri 39192 18747 39193 18748 ne
rect 39193 18747 39464 18748
tri 39193 18746 39194 18747 ne
rect 39194 18746 39464 18747
tri 39194 18745 39195 18746 ne
rect 39195 18745 39464 18746
tri 39195 18744 39196 18745 ne
rect 39196 18744 39464 18745
tri 39196 18743 39197 18744 ne
rect 39197 18743 39464 18744
tri 39197 18742 39198 18743 ne
rect 39198 18742 39464 18743
tri 39198 18741 39199 18742 ne
rect 39199 18741 39464 18742
tri 39199 18740 39200 18741 ne
rect 39200 18740 39464 18741
tri 39200 18739 39201 18740 ne
rect 39201 18739 39464 18740
tri 39201 18738 39202 18739 ne
rect 39202 18738 39464 18739
tri 39202 18737 39203 18738 ne
rect 39203 18737 39464 18738
tri 39203 18736 39204 18737 ne
rect 39204 18736 39464 18737
tri 39204 18735 39205 18736 ne
rect 39205 18735 39464 18736
tri 39205 18734 39206 18735 ne
rect 39206 18734 39464 18735
tri 39206 18733 39207 18734 ne
rect 39207 18733 39464 18734
tri 39207 18732 39208 18733 ne
rect 39208 18732 39464 18733
tri 39208 18731 39209 18732 ne
rect 39209 18731 39464 18732
tri 39209 18730 39210 18731 ne
rect 39210 18730 39464 18731
tri 39210 18729 39211 18730 ne
rect 39211 18729 39464 18730
tri 39211 18728 39212 18729 ne
rect 39212 18728 39464 18729
tri 39212 18727 39213 18728 ne
rect 39213 18727 39464 18728
tri 39213 18726 39214 18727 ne
rect 39214 18726 39464 18727
tri 39214 18725 39215 18726 ne
rect 39215 18725 39464 18726
tri 39215 18724 39216 18725 ne
rect 39216 18724 39464 18725
tri 39216 18723 39217 18724 ne
rect 39217 18723 39464 18724
tri 39217 18722 39218 18723 ne
rect 39218 18722 39464 18723
tri 39218 18721 39219 18722 ne
rect 39219 18721 39464 18722
tri 39219 18720 39220 18721 ne
rect 39220 18720 39464 18721
tri 39220 18719 39221 18720 ne
rect 39221 18719 39464 18720
tri 39221 18718 39222 18719 ne
rect 39222 18718 39464 18719
tri 39222 18717 39223 18718 ne
rect 39223 18717 39464 18718
tri 39223 18716 39224 18717 ne
rect 39224 18716 39464 18717
tri 39224 18715 39225 18716 ne
rect 39225 18715 39464 18716
tri 39225 18714 39226 18715 ne
rect 39226 18714 39464 18715
tri 39226 18713 39227 18714 ne
rect 39227 18713 39464 18714
tri 39227 18712 39228 18713 ne
rect 39228 18712 39464 18713
tri 39228 18711 39229 18712 ne
rect 39229 18711 39464 18712
tri 39229 18710 39230 18711 ne
rect 39230 18710 39464 18711
tri 39230 18709 39231 18710 ne
rect 39231 18709 39464 18710
tri 39231 18708 39232 18709 ne
rect 39232 18708 39464 18709
tri 39232 18707 39233 18708 ne
rect 39233 18707 39464 18708
tri 39464 18707 39509 18752 sw
rect 70802 18740 71000 18798
tri 39233 18706 39234 18707 ne
rect 39234 18706 39509 18707
tri 39234 18705 39235 18706 ne
rect 39235 18705 39509 18706
tri 39235 18704 39236 18705 ne
rect 39236 18704 39509 18705
tri 39236 18703 39237 18704 ne
rect 39237 18703 39509 18704
tri 39237 18702 39238 18703 ne
rect 39238 18702 39509 18703
tri 39238 18701 39239 18702 ne
rect 39239 18701 39509 18702
tri 39239 18700 39240 18701 ne
rect 39240 18700 39509 18701
tri 39240 18699 39241 18700 ne
rect 39241 18699 39509 18700
tri 39241 18698 39242 18699 ne
rect 39242 18698 39509 18699
tri 39242 18697 39243 18698 ne
rect 39243 18697 39509 18698
tri 39243 18696 39244 18697 ne
rect 39244 18696 39509 18697
tri 39244 18695 39245 18696 ne
rect 39245 18695 39509 18696
tri 39245 18694 39246 18695 ne
rect 39246 18694 39509 18695
tri 39246 18693 39247 18694 ne
rect 39247 18693 39509 18694
tri 39247 18692 39248 18693 ne
rect 39248 18692 39509 18693
tri 39248 18691 39249 18692 ne
rect 39249 18691 39509 18692
tri 39249 18690 39250 18691 ne
rect 39250 18690 39509 18691
tri 39250 18689 39251 18690 ne
rect 39251 18689 39509 18690
tri 39251 18688 39252 18689 ne
rect 39252 18688 39509 18689
tri 39252 18687 39253 18688 ne
rect 39253 18687 39390 18688
tri 39253 18686 39254 18687 ne
rect 39254 18686 39390 18687
tri 39254 18685 39255 18686 ne
rect 39255 18685 39390 18686
tri 39255 18684 39256 18685 ne
rect 39256 18684 39390 18685
tri 39256 18683 39257 18684 ne
rect 39257 18683 39390 18684
tri 39257 18682 39258 18683 ne
rect 39258 18682 39390 18683
tri 39258 18681 39259 18682 ne
rect 39259 18681 39390 18682
tri 39259 18680 39260 18681 ne
rect 39260 18680 39390 18681
tri 39260 18679 39261 18680 ne
rect 39261 18679 39390 18680
tri 39261 18678 39262 18679 ne
rect 39262 18678 39390 18679
tri 39262 18677 39263 18678 ne
rect 39263 18677 39390 18678
tri 39263 18676 39264 18677 ne
rect 39264 18676 39390 18677
tri 39264 18675 39265 18676 ne
rect 39265 18675 39390 18676
tri 39265 18674 39266 18675 ne
rect 39266 18674 39390 18675
tri 39266 18673 39267 18674 ne
rect 39267 18673 39390 18674
tri 39267 18672 39268 18673 ne
rect 39268 18672 39390 18673
tri 39268 18671 39269 18672 ne
rect 39269 18671 39390 18672
tri 39269 18670 39270 18671 ne
rect 39270 18670 39390 18671
tri 39270 18669 39271 18670 ne
rect 39271 18669 39390 18670
tri 39271 18668 39272 18669 ne
rect 39272 18668 39390 18669
tri 39272 18667 39273 18668 ne
rect 39273 18667 39390 18668
tri 39273 18666 39274 18667 ne
rect 39274 18666 39390 18667
tri 39274 18665 39275 18666 ne
rect 39275 18665 39390 18666
tri 39275 18664 39276 18665 ne
rect 39276 18664 39390 18665
tri 39276 18663 39277 18664 ne
rect 39277 18663 39390 18664
tri 39277 18662 39278 18663 ne
rect 39278 18662 39390 18663
tri 39278 18661 39279 18662 ne
rect 39279 18661 39390 18662
tri 39279 18660 39280 18661 ne
rect 39280 18660 39390 18661
tri 39280 18659 39281 18660 ne
rect 39281 18659 39390 18660
tri 39281 18658 39282 18659 ne
rect 39282 18658 39390 18659
tri 39282 18657 39283 18658 ne
rect 39283 18657 39390 18658
tri 39283 18656 39284 18657 ne
rect 39284 18656 39390 18657
tri 39284 18655 39285 18656 ne
rect 39285 18655 39390 18656
tri 39285 18654 39286 18655 ne
rect 39286 18654 39390 18655
tri 39286 18653 39287 18654 ne
rect 39287 18653 39390 18654
tri 39287 18652 39288 18653 ne
rect 39288 18652 39390 18653
tri 39288 18651 39289 18652 ne
rect 39289 18651 39390 18652
tri 39289 18650 39290 18651 ne
rect 39290 18650 39390 18651
tri 39290 18649 39291 18650 ne
rect 39291 18649 39390 18650
tri 39291 18648 39292 18649 ne
rect 39292 18648 39390 18649
tri 39292 18647 39293 18648 ne
rect 39293 18647 39390 18648
tri 39293 18646 39294 18647 ne
rect 39294 18646 39390 18647
tri 39294 18645 39295 18646 ne
rect 39295 18645 39390 18646
tri 39295 18644 39296 18645 ne
rect 39296 18644 39390 18645
tri 39296 18643 39297 18644 ne
rect 39297 18643 39390 18644
tri 39297 18642 39298 18643 ne
rect 39298 18642 39390 18643
rect 39436 18662 39509 18688
tri 39509 18662 39554 18707 sw
rect 70802 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 39436 18642 39554 18662
tri 39298 18641 39299 18642 ne
rect 39299 18641 39554 18642
tri 39299 18640 39300 18641 ne
rect 39300 18640 39554 18641
tri 39300 18639 39301 18640 ne
rect 39301 18639 39554 18640
tri 39301 18638 39302 18639 ne
rect 39302 18638 39554 18639
tri 39302 18637 39303 18638 ne
rect 39303 18637 39554 18638
tri 39303 18636 39304 18637 ne
rect 39304 18636 39554 18637
tri 39304 18635 39305 18636 ne
rect 39305 18635 39554 18636
tri 39305 18634 39306 18635 ne
rect 39306 18634 39554 18635
tri 39306 18633 39307 18634 ne
rect 39307 18633 39554 18634
tri 39307 18632 39308 18633 ne
rect 39308 18632 39554 18633
tri 39308 18631 39309 18632 ne
rect 39309 18631 39554 18632
tri 39309 18630 39310 18631 ne
rect 39310 18630 39554 18631
tri 39310 18629 39311 18630 ne
rect 39311 18629 39554 18630
tri 39311 18628 39312 18629 ne
rect 39312 18628 39554 18629
tri 39312 18627 39313 18628 ne
rect 39313 18627 39554 18628
tri 39313 18626 39314 18627 ne
rect 39314 18626 39554 18627
tri 39314 18625 39315 18626 ne
rect 39315 18625 39554 18626
tri 39315 18624 39316 18625 ne
rect 39316 18624 39554 18625
tri 39316 18623 39317 18624 ne
rect 39317 18623 39554 18624
tri 39317 18622 39318 18623 ne
rect 39318 18622 39554 18623
tri 39318 18621 39319 18622 ne
rect 39319 18621 39554 18622
tri 39319 18620 39320 18621 ne
rect 39320 18620 39554 18621
tri 39320 18619 39321 18620 ne
rect 39321 18619 39554 18620
tri 39321 18618 39322 18619 ne
rect 39322 18618 39554 18619
tri 39322 18617 39323 18618 ne
rect 39323 18617 39554 18618
tri 39554 18617 39599 18662 sw
rect 70802 18636 71000 18694
tri 39323 18600 39340 18617 ne
rect 39340 18600 39599 18617
tri 39599 18600 39616 18617 sw
tri 39340 18572 39368 18600 ne
rect 39368 18572 39616 18600
tri 39368 18555 39385 18572 ne
rect 39385 18556 39616 18572
rect 39385 18555 39522 18556
tri 39385 18510 39430 18555 ne
rect 39430 18510 39522 18555
rect 39568 18555 39616 18556
tri 39616 18555 39661 18600 sw
rect 70802 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39568 18510 39661 18555
tri 39661 18510 39706 18555 sw
rect 70802 18532 71000 18590
tri 39430 18505 39435 18510 ne
rect 39435 18505 39706 18510
tri 39435 18504 39436 18505 ne
rect 39436 18504 39706 18505
tri 39436 18503 39437 18504 ne
rect 39437 18503 39706 18504
tri 39437 18502 39438 18503 ne
rect 39438 18502 39706 18503
tri 39438 18501 39439 18502 ne
rect 39439 18501 39706 18502
tri 39439 18500 39440 18501 ne
rect 39440 18500 39706 18501
tri 39440 18499 39441 18500 ne
rect 39441 18499 39706 18500
tri 39441 18498 39442 18499 ne
rect 39442 18498 39706 18499
tri 39442 18497 39443 18498 ne
rect 39443 18497 39706 18498
tri 39443 18496 39444 18497 ne
rect 39444 18496 39706 18497
tri 39444 18495 39445 18496 ne
rect 39445 18495 39706 18496
tri 39445 18494 39446 18495 ne
rect 39446 18494 39706 18495
tri 39446 18493 39447 18494 ne
rect 39447 18493 39706 18494
tri 39447 18492 39448 18493 ne
rect 39448 18492 39706 18493
tri 39448 18491 39449 18492 ne
rect 39449 18491 39706 18492
tri 39449 18490 39450 18491 ne
rect 39450 18490 39706 18491
tri 39450 18489 39451 18490 ne
rect 39451 18489 39706 18490
tri 39451 18488 39452 18489 ne
rect 39452 18488 39706 18489
tri 39452 18487 39453 18488 ne
rect 39453 18487 39706 18488
tri 39453 18486 39454 18487 ne
rect 39454 18486 39706 18487
tri 39454 18485 39455 18486 ne
rect 39455 18485 39706 18486
tri 39455 18484 39456 18485 ne
rect 39456 18484 39706 18485
tri 39456 18483 39457 18484 ne
rect 39457 18483 39706 18484
tri 39457 18482 39458 18483 ne
rect 39458 18482 39706 18483
tri 39458 18481 39459 18482 ne
rect 39459 18481 39706 18482
tri 39459 18480 39460 18481 ne
rect 39460 18480 39706 18481
tri 39460 18479 39461 18480 ne
rect 39461 18479 39706 18480
tri 39461 18478 39462 18479 ne
rect 39462 18478 39706 18479
tri 39462 18477 39463 18478 ne
rect 39463 18477 39706 18478
tri 39463 18476 39464 18477 ne
rect 39464 18476 39706 18477
tri 39464 18475 39465 18476 ne
rect 39465 18475 39706 18476
tri 39465 18474 39466 18475 ne
rect 39466 18474 39706 18475
tri 39466 18473 39467 18474 ne
rect 39467 18473 39706 18474
tri 39467 18472 39468 18473 ne
rect 39468 18472 39706 18473
tri 39468 18471 39469 18472 ne
rect 39469 18471 39706 18472
tri 39469 18470 39470 18471 ne
rect 39470 18470 39706 18471
tri 39470 18469 39471 18470 ne
rect 39471 18469 39706 18470
tri 39471 18468 39472 18469 ne
rect 39472 18468 39706 18469
tri 39472 18467 39473 18468 ne
rect 39473 18467 39706 18468
tri 39473 18466 39474 18467 ne
rect 39474 18466 39706 18467
tri 39474 18465 39475 18466 ne
rect 39475 18465 39706 18466
tri 39706 18465 39751 18510 sw
rect 70802 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
tri 39475 18464 39476 18465 ne
rect 39476 18464 39751 18465
tri 39476 18463 39477 18464 ne
rect 39477 18463 39751 18464
tri 39477 18462 39478 18463 ne
rect 39478 18462 39751 18463
tri 39478 18461 39479 18462 ne
rect 39479 18461 39751 18462
tri 39479 18460 39480 18461 ne
rect 39480 18460 39751 18461
tri 39480 18459 39481 18460 ne
rect 39481 18459 39751 18460
tri 39481 18458 39482 18459 ne
rect 39482 18458 39751 18459
tri 39482 18457 39483 18458 ne
rect 39483 18457 39751 18458
tri 39483 18456 39484 18457 ne
rect 39484 18456 39751 18457
tri 39484 18455 39485 18456 ne
rect 39485 18455 39751 18456
tri 39485 18454 39486 18455 ne
rect 39486 18454 39751 18455
tri 39486 18453 39487 18454 ne
rect 39487 18453 39751 18454
tri 39487 18452 39488 18453 ne
rect 39488 18452 39751 18453
tri 39488 18451 39489 18452 ne
rect 39489 18451 39751 18452
tri 39489 18450 39490 18451 ne
rect 39490 18450 39751 18451
tri 39490 18449 39491 18450 ne
rect 39491 18449 39751 18450
tri 39491 18448 39492 18449 ne
rect 39492 18448 39751 18449
tri 39492 18447 39493 18448 ne
rect 39493 18447 39751 18448
tri 39493 18446 39494 18447 ne
rect 39494 18446 39751 18447
tri 39494 18445 39495 18446 ne
rect 39495 18445 39751 18446
tri 39495 18444 39496 18445 ne
rect 39496 18444 39751 18445
tri 39496 18443 39497 18444 ne
rect 39497 18443 39751 18444
tri 39497 18442 39498 18443 ne
rect 39498 18442 39751 18443
tri 39498 18441 39499 18442 ne
rect 39499 18441 39751 18442
tri 39499 18440 39500 18441 ne
rect 39500 18440 39751 18441
tri 39500 18439 39501 18440 ne
rect 39501 18439 39751 18440
tri 39501 18438 39502 18439 ne
rect 39502 18438 39751 18439
tri 39502 18437 39503 18438 ne
rect 39503 18437 39751 18438
tri 39503 18436 39504 18437 ne
rect 39504 18436 39751 18437
tri 39504 18435 39505 18436 ne
rect 39505 18435 39751 18436
tri 39505 18434 39506 18435 ne
rect 39506 18434 39751 18435
tri 39506 18433 39507 18434 ne
rect 39507 18433 39751 18434
tri 39507 18432 39508 18433 ne
rect 39508 18432 39751 18433
tri 39508 18431 39509 18432 ne
rect 39509 18431 39751 18432
tri 39751 18431 39785 18465 sw
tri 39509 18430 39510 18431 ne
rect 39510 18430 39785 18431
tri 39510 18429 39511 18430 ne
rect 39511 18429 39785 18430
tri 39511 18428 39512 18429 ne
rect 39512 18428 39785 18429
tri 39512 18427 39513 18428 ne
rect 39513 18427 39785 18428
tri 39513 18426 39514 18427 ne
rect 39514 18426 39785 18427
tri 39514 18425 39515 18426 ne
rect 39515 18425 39785 18426
tri 39515 18424 39516 18425 ne
rect 39516 18424 39785 18425
tri 39516 18423 39517 18424 ne
rect 39517 18423 39654 18424
tri 39517 18422 39518 18423 ne
rect 39518 18422 39654 18423
tri 39518 18421 39519 18422 ne
rect 39519 18421 39654 18422
tri 39519 18420 39520 18421 ne
rect 39520 18420 39654 18421
tri 39520 18419 39521 18420 ne
rect 39521 18419 39654 18420
tri 39521 18418 39522 18419 ne
rect 39522 18418 39654 18419
tri 39522 18417 39523 18418 ne
rect 39523 18417 39654 18418
tri 39523 18416 39524 18417 ne
rect 39524 18416 39654 18417
tri 39524 18415 39525 18416 ne
rect 39525 18415 39654 18416
tri 39525 18414 39526 18415 ne
rect 39526 18414 39654 18415
tri 39526 18413 39527 18414 ne
rect 39527 18413 39654 18414
tri 39527 18412 39528 18413 ne
rect 39528 18412 39654 18413
tri 39528 18411 39529 18412 ne
rect 39529 18411 39654 18412
tri 39529 18410 39530 18411 ne
rect 39530 18410 39654 18411
tri 39530 18409 39531 18410 ne
rect 39531 18409 39654 18410
tri 39531 18408 39532 18409 ne
rect 39532 18408 39654 18409
tri 39532 18407 39533 18408 ne
rect 39533 18407 39654 18408
tri 39533 18406 39534 18407 ne
rect 39534 18406 39654 18407
tri 39534 18405 39535 18406 ne
rect 39535 18405 39654 18406
tri 39535 18404 39536 18405 ne
rect 39536 18404 39654 18405
tri 39536 18403 39537 18404 ne
rect 39537 18403 39654 18404
tri 39537 18402 39538 18403 ne
rect 39538 18402 39654 18403
tri 39538 18401 39539 18402 ne
rect 39539 18401 39654 18402
tri 39539 18400 39540 18401 ne
rect 39540 18400 39654 18401
tri 39540 18399 39541 18400 ne
rect 39541 18399 39654 18400
tri 39541 18398 39542 18399 ne
rect 39542 18398 39654 18399
tri 39542 18397 39543 18398 ne
rect 39543 18397 39654 18398
tri 39543 18396 39544 18397 ne
rect 39544 18396 39654 18397
tri 39544 18395 39545 18396 ne
rect 39545 18395 39654 18396
tri 39545 18394 39546 18395 ne
rect 39546 18394 39654 18395
tri 39546 18393 39547 18394 ne
rect 39547 18393 39654 18394
tri 39547 18392 39548 18393 ne
rect 39548 18392 39654 18393
tri 39548 18391 39549 18392 ne
rect 39549 18391 39654 18392
tri 39549 18390 39550 18391 ne
rect 39550 18390 39654 18391
tri 39550 18389 39551 18390 ne
rect 39551 18389 39654 18390
tri 39551 18388 39552 18389 ne
rect 39552 18388 39654 18389
tri 39552 18387 39553 18388 ne
rect 39553 18387 39654 18388
tri 39553 18386 39554 18387 ne
rect 39554 18386 39654 18387
tri 39554 18385 39555 18386 ne
rect 39555 18385 39654 18386
tri 39555 18384 39556 18385 ne
rect 39556 18384 39654 18385
tri 39556 18383 39557 18384 ne
rect 39557 18383 39654 18384
tri 39557 18382 39558 18383 ne
rect 39558 18382 39654 18383
tri 39558 18381 39559 18382 ne
rect 39559 18381 39654 18382
tri 39559 18380 39560 18381 ne
rect 39560 18380 39654 18381
tri 39560 18379 39561 18380 ne
rect 39561 18379 39654 18380
tri 39561 18378 39562 18379 ne
rect 39562 18378 39654 18379
rect 39700 18386 39785 18424
tri 39785 18386 39830 18431 sw
rect 70802 18428 71000 18486
rect 39700 18378 39830 18386
tri 39562 18377 39563 18378 ne
rect 39563 18377 39830 18378
tri 39563 18376 39564 18377 ne
rect 39564 18376 39830 18377
tri 39564 18375 39565 18376 ne
rect 39565 18375 39830 18376
tri 39565 18374 39566 18375 ne
rect 39566 18374 39830 18375
tri 39566 18373 39567 18374 ne
rect 39567 18373 39830 18374
tri 39567 18372 39568 18373 ne
rect 39568 18372 39830 18373
tri 39568 18371 39569 18372 ne
rect 39569 18371 39830 18372
tri 39569 18370 39570 18371 ne
rect 39570 18370 39830 18371
tri 39570 18369 39571 18370 ne
rect 39571 18369 39830 18370
tri 39571 18368 39572 18369 ne
rect 39572 18368 39830 18369
tri 39572 18367 39573 18368 ne
rect 39573 18367 39830 18368
tri 39573 18366 39574 18367 ne
rect 39574 18366 39830 18367
tri 39574 18365 39575 18366 ne
rect 39575 18365 39830 18366
tri 39575 18364 39576 18365 ne
rect 39576 18364 39830 18365
tri 39576 18363 39577 18364 ne
rect 39577 18363 39830 18364
tri 39577 18362 39578 18363 ne
rect 39578 18362 39830 18363
tri 39578 18361 39579 18362 ne
rect 39579 18361 39830 18362
tri 39579 18360 39580 18361 ne
rect 39580 18360 39830 18361
tri 39580 18359 39581 18360 ne
rect 39581 18359 39830 18360
tri 39581 18358 39582 18359 ne
rect 39582 18358 39830 18359
tri 39582 18357 39583 18358 ne
rect 39583 18357 39830 18358
tri 39583 18356 39584 18357 ne
rect 39584 18356 39830 18357
tri 39584 18355 39585 18356 ne
rect 39585 18355 39830 18356
tri 39585 18354 39586 18355 ne
rect 39586 18354 39830 18355
tri 39586 18353 39587 18354 ne
rect 39587 18353 39830 18354
tri 39587 18352 39588 18353 ne
rect 39588 18352 39830 18353
tri 39588 18351 39589 18352 ne
rect 39589 18351 39830 18352
tri 39589 18350 39590 18351 ne
rect 39590 18350 39830 18351
tri 39590 18349 39591 18350 ne
rect 39591 18349 39830 18350
tri 39591 18348 39592 18349 ne
rect 39592 18348 39830 18349
tri 39592 18347 39593 18348 ne
rect 39593 18347 39830 18348
tri 39593 18346 39594 18347 ne
rect 39594 18346 39830 18347
tri 39594 18345 39595 18346 ne
rect 39595 18345 39830 18346
tri 39595 18344 39596 18345 ne
rect 39596 18344 39830 18345
tri 39596 18343 39597 18344 ne
rect 39597 18343 39830 18344
tri 39597 18342 39598 18343 ne
rect 39598 18342 39830 18343
tri 39598 18341 39599 18342 ne
rect 39599 18341 39830 18342
tri 39830 18341 39875 18386 sw
rect 70802 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
tri 39599 18296 39644 18341 ne
rect 39644 18296 39875 18341
tri 39875 18296 39920 18341 sw
rect 70802 18324 71000 18382
tri 39644 18251 39689 18296 ne
rect 39689 18292 39920 18296
rect 39689 18251 39786 18292
tri 39689 18234 39706 18251 ne
rect 39706 18246 39786 18251
rect 39832 18279 39920 18292
tri 39920 18279 39937 18296 sw
rect 39832 18246 39937 18279
rect 39706 18234 39937 18246
tri 39937 18234 39982 18279 sw
rect 70802 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
tri 39706 18230 39710 18234 ne
rect 39710 18230 39982 18234
tri 39710 18229 39711 18230 ne
rect 39711 18229 39982 18230
tri 39711 18228 39712 18229 ne
rect 39712 18228 39982 18229
tri 39712 18227 39713 18228 ne
rect 39713 18227 39982 18228
tri 39713 18226 39714 18227 ne
rect 39714 18226 39982 18227
tri 39714 18225 39715 18226 ne
rect 39715 18225 39982 18226
tri 39715 18224 39716 18225 ne
rect 39716 18224 39982 18225
tri 39716 18223 39717 18224 ne
rect 39717 18223 39982 18224
tri 39717 18222 39718 18223 ne
rect 39718 18222 39982 18223
tri 39718 18221 39719 18222 ne
rect 39719 18221 39982 18222
tri 39719 18220 39720 18221 ne
rect 39720 18220 39982 18221
tri 39720 18219 39721 18220 ne
rect 39721 18219 39982 18220
tri 39721 18218 39722 18219 ne
rect 39722 18218 39982 18219
tri 39722 18217 39723 18218 ne
rect 39723 18217 39982 18218
tri 39723 18216 39724 18217 ne
rect 39724 18216 39982 18217
tri 39724 18215 39725 18216 ne
rect 39725 18215 39982 18216
tri 39725 18214 39726 18215 ne
rect 39726 18214 39982 18215
tri 39726 18213 39727 18214 ne
rect 39727 18213 39982 18214
tri 39727 18212 39728 18213 ne
rect 39728 18212 39982 18213
tri 39728 18211 39729 18212 ne
rect 39729 18211 39982 18212
tri 39729 18210 39730 18211 ne
rect 39730 18210 39982 18211
tri 39730 18209 39731 18210 ne
rect 39731 18209 39982 18210
tri 39731 18208 39732 18209 ne
rect 39732 18208 39982 18209
tri 39732 18207 39733 18208 ne
rect 39733 18207 39982 18208
tri 39733 18206 39734 18207 ne
rect 39734 18206 39982 18207
tri 39734 18205 39735 18206 ne
rect 39735 18205 39982 18206
tri 39735 18204 39736 18205 ne
rect 39736 18204 39982 18205
tri 39736 18203 39737 18204 ne
rect 39737 18203 39982 18204
tri 39737 18202 39738 18203 ne
rect 39738 18202 39982 18203
tri 39738 18201 39739 18202 ne
rect 39739 18201 39982 18202
tri 39739 18200 39740 18201 ne
rect 39740 18200 39982 18201
tri 39740 18199 39741 18200 ne
rect 39741 18199 39982 18200
tri 39741 18198 39742 18199 ne
rect 39742 18198 39982 18199
tri 39742 18197 39743 18198 ne
rect 39743 18197 39982 18198
tri 39743 18196 39744 18197 ne
rect 39744 18196 39982 18197
tri 39744 18195 39745 18196 ne
rect 39745 18195 39982 18196
tri 39745 18194 39746 18195 ne
rect 39746 18194 39982 18195
tri 39746 18193 39747 18194 ne
rect 39747 18193 39982 18194
tri 39747 18192 39748 18193 ne
rect 39748 18192 39982 18193
tri 39748 18191 39749 18192 ne
rect 39749 18191 39982 18192
tri 39749 18190 39750 18191 ne
rect 39750 18190 39982 18191
tri 39750 18189 39751 18190 ne
rect 39751 18189 39982 18190
tri 39982 18189 40027 18234 sw
rect 70802 18220 71000 18278
tri 39751 18188 39752 18189 ne
rect 39752 18188 40027 18189
tri 39752 18187 39753 18188 ne
rect 39753 18187 40027 18188
tri 39753 18186 39754 18187 ne
rect 39754 18186 40027 18187
tri 39754 18185 39755 18186 ne
rect 39755 18185 40027 18186
tri 39755 18184 39756 18185 ne
rect 39756 18184 40027 18185
tri 39756 18183 39757 18184 ne
rect 39757 18183 40027 18184
tri 39757 18182 39758 18183 ne
rect 39758 18182 40027 18183
tri 39758 18181 39759 18182 ne
rect 39759 18181 40027 18182
tri 39759 18180 39760 18181 ne
rect 39760 18180 40027 18181
tri 39760 18179 39761 18180 ne
rect 39761 18179 40027 18180
tri 39761 18178 39762 18179 ne
rect 39762 18178 40027 18179
tri 39762 18177 39763 18178 ne
rect 39763 18177 40027 18178
tri 39763 18176 39764 18177 ne
rect 39764 18176 40027 18177
tri 39764 18175 39765 18176 ne
rect 39765 18175 40027 18176
tri 39765 18174 39766 18175 ne
rect 39766 18174 40027 18175
tri 39766 18173 39767 18174 ne
rect 39767 18173 40027 18174
tri 39767 18172 39768 18173 ne
rect 39768 18172 40027 18173
tri 39768 18171 39769 18172 ne
rect 39769 18171 40027 18172
tri 39769 18170 39770 18171 ne
rect 39770 18170 40027 18171
tri 39770 18169 39771 18170 ne
rect 39771 18169 40027 18170
tri 39771 18168 39772 18169 ne
rect 39772 18168 40027 18169
tri 39772 18167 39773 18168 ne
rect 39773 18167 40027 18168
tri 39773 18166 39774 18167 ne
rect 39774 18166 40027 18167
tri 39774 18165 39775 18166 ne
rect 39775 18165 40027 18166
tri 39775 18164 39776 18165 ne
rect 39776 18164 40027 18165
tri 39776 18163 39777 18164 ne
rect 39777 18163 40027 18164
tri 39777 18162 39778 18163 ne
rect 39778 18162 40027 18163
tri 39778 18161 39779 18162 ne
rect 39779 18161 40027 18162
tri 39779 18160 39780 18161 ne
rect 39780 18160 40027 18161
tri 39780 18159 39781 18160 ne
rect 39781 18159 39918 18160
tri 39781 18158 39782 18159 ne
rect 39782 18158 39918 18159
tri 39782 18157 39783 18158 ne
rect 39783 18157 39918 18158
tri 39783 18156 39784 18157 ne
rect 39784 18156 39918 18157
tri 39784 18155 39785 18156 ne
rect 39785 18155 39918 18156
tri 39785 18154 39786 18155 ne
rect 39786 18154 39918 18155
tri 39786 18153 39787 18154 ne
rect 39787 18153 39918 18154
tri 39787 18152 39788 18153 ne
rect 39788 18152 39918 18153
tri 39788 18151 39789 18152 ne
rect 39789 18151 39918 18152
tri 39789 18150 39790 18151 ne
rect 39790 18150 39918 18151
tri 39790 18149 39791 18150 ne
rect 39791 18149 39918 18150
tri 39791 18148 39792 18149 ne
rect 39792 18148 39918 18149
tri 39792 18147 39793 18148 ne
rect 39793 18147 39918 18148
tri 39793 18146 39794 18147 ne
rect 39794 18146 39918 18147
tri 39794 18145 39795 18146 ne
rect 39795 18145 39918 18146
tri 39795 18144 39796 18145 ne
rect 39796 18144 39918 18145
tri 39796 18143 39797 18144 ne
rect 39797 18143 39918 18144
tri 39797 18142 39798 18143 ne
rect 39798 18142 39918 18143
tri 39798 18141 39799 18142 ne
rect 39799 18141 39918 18142
tri 39799 18140 39800 18141 ne
rect 39800 18140 39918 18141
tri 39800 18139 39801 18140 ne
rect 39801 18139 39918 18140
tri 39801 18138 39802 18139 ne
rect 39802 18138 39918 18139
tri 39802 18137 39803 18138 ne
rect 39803 18137 39918 18138
tri 39803 18136 39804 18137 ne
rect 39804 18136 39918 18137
tri 39804 18135 39805 18136 ne
rect 39805 18135 39918 18136
tri 39805 18134 39806 18135 ne
rect 39806 18134 39918 18135
tri 39806 18133 39807 18134 ne
rect 39807 18133 39918 18134
tri 39807 18132 39808 18133 ne
rect 39808 18132 39918 18133
tri 39808 18131 39809 18132 ne
rect 39809 18131 39918 18132
tri 39809 18130 39810 18131 ne
rect 39810 18130 39918 18131
tri 39810 18129 39811 18130 ne
rect 39811 18129 39918 18130
tri 39811 18128 39812 18129 ne
rect 39812 18128 39918 18129
tri 39812 18127 39813 18128 ne
rect 39813 18127 39918 18128
tri 39813 18126 39814 18127 ne
rect 39814 18126 39918 18127
tri 39814 18125 39815 18126 ne
rect 39815 18125 39918 18126
tri 39815 18124 39816 18125 ne
rect 39816 18124 39918 18125
tri 39816 18123 39817 18124 ne
rect 39817 18123 39918 18124
tri 39817 18122 39818 18123 ne
rect 39818 18122 39918 18123
tri 39818 18121 39819 18122 ne
rect 39819 18121 39918 18122
tri 39819 18120 39820 18121 ne
rect 39820 18120 39918 18121
tri 39820 18119 39821 18120 ne
rect 39821 18119 39918 18120
tri 39821 18118 39822 18119 ne
rect 39822 18118 39918 18119
tri 39822 18117 39823 18118 ne
rect 39823 18117 39918 18118
tri 39823 18116 39824 18117 ne
rect 39824 18116 39918 18117
tri 39824 18115 39825 18116 ne
rect 39825 18115 39918 18116
tri 39825 18114 39826 18115 ne
rect 39826 18114 39918 18115
rect 39964 18144 40027 18160
tri 40027 18144 40072 18189 sw
rect 70802 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 39964 18114 40072 18144
tri 39826 18113 39827 18114 ne
rect 39827 18113 40072 18114
tri 39827 18112 39828 18113 ne
rect 39828 18112 40072 18113
tri 39828 18111 39829 18112 ne
rect 39829 18111 40072 18112
tri 39829 18110 39830 18111 ne
rect 39830 18110 40072 18111
tri 40072 18110 40106 18144 sw
rect 70802 18116 71000 18174
tri 39830 18109 39831 18110 ne
rect 39831 18109 40106 18110
tri 39831 18108 39832 18109 ne
rect 39832 18108 40106 18109
tri 39832 18107 39833 18108 ne
rect 39833 18107 40106 18108
tri 39833 18106 39834 18107 ne
rect 39834 18106 40106 18107
tri 39834 18105 39835 18106 ne
rect 39835 18105 40106 18106
tri 39835 18104 39836 18105 ne
rect 39836 18104 40106 18105
tri 39836 18103 39837 18104 ne
rect 39837 18103 40106 18104
tri 39837 18102 39838 18103 ne
rect 39838 18102 40106 18103
tri 39838 18101 39839 18102 ne
rect 39839 18101 40106 18102
tri 39839 18100 39840 18101 ne
rect 39840 18100 40106 18101
tri 39840 18099 39841 18100 ne
rect 39841 18099 40106 18100
tri 39841 18098 39842 18099 ne
rect 39842 18098 40106 18099
tri 39842 18097 39843 18098 ne
rect 39843 18097 40106 18098
tri 39843 18096 39844 18097 ne
rect 39844 18096 40106 18097
tri 39844 18095 39845 18096 ne
rect 39845 18095 40106 18096
tri 39845 18094 39846 18095 ne
rect 39846 18094 40106 18095
tri 39846 18093 39847 18094 ne
rect 39847 18093 40106 18094
tri 39847 18092 39848 18093 ne
rect 39848 18092 40106 18093
tri 39848 18091 39849 18092 ne
rect 39849 18091 40106 18092
tri 39849 18090 39850 18091 ne
rect 39850 18090 40106 18091
tri 39850 18089 39851 18090 ne
rect 39851 18089 40106 18090
tri 39851 18088 39852 18089 ne
rect 39852 18088 40106 18089
tri 39852 18087 39853 18088 ne
rect 39853 18087 40106 18088
tri 39853 18086 39854 18087 ne
rect 39854 18086 40106 18087
tri 39854 18085 39855 18086 ne
rect 39855 18085 40106 18086
tri 39855 18084 39856 18085 ne
rect 39856 18084 40106 18085
tri 39856 18083 39857 18084 ne
rect 39857 18083 40106 18084
tri 39857 18082 39858 18083 ne
rect 39858 18082 40106 18083
tri 39858 18081 39859 18082 ne
rect 39859 18081 40106 18082
tri 39859 18080 39860 18081 ne
rect 39860 18080 40106 18081
tri 39860 18079 39861 18080 ne
rect 39861 18079 40106 18080
tri 39861 18078 39862 18079 ne
rect 39862 18078 40106 18079
tri 39862 18077 39863 18078 ne
rect 39863 18077 40106 18078
tri 39863 18076 39864 18077 ne
rect 39864 18076 40106 18077
tri 39864 18075 39865 18076 ne
rect 39865 18075 40106 18076
tri 39865 18074 39866 18075 ne
rect 39866 18074 40106 18075
tri 39866 18073 39867 18074 ne
rect 39867 18073 40106 18074
tri 39867 18072 39868 18073 ne
rect 39868 18072 40106 18073
tri 39868 18071 39869 18072 ne
rect 39869 18071 40106 18072
tri 39869 18070 39870 18071 ne
rect 39870 18070 40106 18071
tri 39870 18069 39871 18070 ne
rect 39871 18069 40106 18070
tri 39871 18068 39872 18069 ne
rect 39872 18068 40106 18069
tri 39872 18067 39873 18068 ne
rect 39873 18067 40106 18068
tri 39873 18066 39874 18067 ne
rect 39874 18066 40106 18067
tri 39874 18065 39875 18066 ne
rect 39875 18065 40106 18066
tri 40106 18065 40151 18110 sw
rect 70802 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39875 18020 39920 18065 ne
rect 39920 18028 40151 18065
rect 39920 18020 40050 18028
tri 39920 17975 39965 18020 ne
rect 39965 17982 40050 18020
rect 40096 18020 40151 18028
tri 40151 18020 40196 18065 sw
rect 40096 17982 40196 18020
rect 39965 17975 40196 17982
tri 40196 17975 40241 18020 sw
rect 70802 18012 71000 18070
tri 39965 17956 39984 17975 ne
rect 39984 17958 40241 17975
tri 40241 17958 40258 17975 sw
rect 70802 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 39984 17956 40258 17958
tri 39984 17955 39985 17956 ne
rect 39985 17955 40258 17956
tri 39985 17954 39986 17955 ne
rect 39986 17954 40258 17955
tri 39986 17953 39987 17954 ne
rect 39987 17953 40258 17954
tri 39987 17952 39988 17953 ne
rect 39988 17952 40258 17953
tri 39988 17951 39989 17952 ne
rect 39989 17951 40258 17952
tri 39989 17950 39990 17951 ne
rect 39990 17950 40258 17951
tri 39990 17949 39991 17950 ne
rect 39991 17949 40258 17950
tri 39991 17948 39992 17949 ne
rect 39992 17948 40258 17949
tri 39992 17947 39993 17948 ne
rect 39993 17947 40258 17948
tri 39993 17946 39994 17947 ne
rect 39994 17946 40258 17947
tri 39994 17945 39995 17946 ne
rect 39995 17945 40258 17946
tri 39995 17944 39996 17945 ne
rect 39996 17944 40258 17945
tri 39996 17943 39997 17944 ne
rect 39997 17943 40258 17944
tri 39997 17942 39998 17943 ne
rect 39998 17942 40258 17943
tri 39998 17941 39999 17942 ne
rect 39999 17941 40258 17942
tri 39999 17940 40000 17941 ne
rect 40000 17940 40258 17941
tri 40000 17939 40001 17940 ne
rect 40001 17939 40258 17940
tri 40001 17938 40002 17939 ne
rect 40002 17938 40258 17939
tri 40002 17937 40003 17938 ne
rect 40003 17937 40258 17938
tri 40003 17936 40004 17937 ne
rect 40004 17936 40258 17937
tri 40004 17935 40005 17936 ne
rect 40005 17935 40258 17936
tri 40005 17934 40006 17935 ne
rect 40006 17934 40258 17935
tri 40006 17933 40007 17934 ne
rect 40007 17933 40258 17934
tri 40007 17932 40008 17933 ne
rect 40008 17932 40258 17933
tri 40008 17931 40009 17932 ne
rect 40009 17931 40258 17932
tri 40009 17930 40010 17931 ne
rect 40010 17930 40258 17931
tri 40010 17929 40011 17930 ne
rect 40011 17929 40258 17930
tri 40011 17928 40012 17929 ne
rect 40012 17928 40258 17929
tri 40012 17927 40013 17928 ne
rect 40013 17927 40258 17928
tri 40013 17926 40014 17927 ne
rect 40014 17926 40258 17927
tri 40014 17925 40015 17926 ne
rect 40015 17925 40258 17926
tri 40015 17924 40016 17925 ne
rect 40016 17924 40258 17925
tri 40016 17923 40017 17924 ne
rect 40017 17923 40258 17924
tri 40017 17922 40018 17923 ne
rect 40018 17922 40258 17923
tri 40018 17921 40019 17922 ne
rect 40019 17921 40258 17922
tri 40019 17920 40020 17921 ne
rect 40020 17920 40258 17921
tri 40020 17919 40021 17920 ne
rect 40021 17919 40258 17920
tri 40021 17918 40022 17919 ne
rect 40022 17918 40258 17919
tri 40022 17917 40023 17918 ne
rect 40023 17917 40258 17918
tri 40023 17916 40024 17917 ne
rect 40024 17916 40258 17917
tri 40024 17915 40025 17916 ne
rect 40025 17915 40258 17916
tri 40025 17914 40026 17915 ne
rect 40026 17914 40258 17915
tri 40026 17913 40027 17914 ne
rect 40027 17913 40258 17914
tri 40258 17913 40303 17958 sw
tri 40027 17912 40028 17913 ne
rect 40028 17912 40303 17913
tri 40028 17911 40029 17912 ne
rect 40029 17911 40303 17912
tri 40029 17910 40030 17911 ne
rect 40030 17910 40303 17911
tri 40030 17909 40031 17910 ne
rect 40031 17909 40303 17910
tri 40031 17908 40032 17909 ne
rect 40032 17908 40303 17909
tri 40032 17907 40033 17908 ne
rect 40033 17907 40303 17908
tri 40033 17906 40034 17907 ne
rect 40034 17906 40303 17907
tri 40034 17905 40035 17906 ne
rect 40035 17905 40303 17906
tri 40035 17904 40036 17905 ne
rect 40036 17904 40303 17905
tri 40036 17903 40037 17904 ne
rect 40037 17903 40303 17904
tri 40037 17902 40038 17903 ne
rect 40038 17902 40303 17903
tri 40038 17901 40039 17902 ne
rect 40039 17901 40303 17902
tri 40039 17900 40040 17901 ne
rect 40040 17900 40303 17901
tri 40040 17899 40041 17900 ne
rect 40041 17899 40303 17900
tri 40041 17898 40042 17899 ne
rect 40042 17898 40303 17899
tri 40042 17897 40043 17898 ne
rect 40043 17897 40303 17898
tri 40043 17896 40044 17897 ne
rect 40044 17896 40303 17897
tri 40044 17895 40045 17896 ne
rect 40045 17895 40182 17896
tri 40045 17894 40046 17895 ne
rect 40046 17894 40182 17895
tri 40046 17893 40047 17894 ne
rect 40047 17893 40182 17894
tri 40047 17892 40048 17893 ne
rect 40048 17892 40182 17893
tri 40048 17891 40049 17892 ne
rect 40049 17891 40182 17892
tri 40049 17890 40050 17891 ne
rect 40050 17890 40182 17891
tri 40050 17889 40051 17890 ne
rect 40051 17889 40182 17890
tri 40051 17888 40052 17889 ne
rect 40052 17888 40182 17889
tri 40052 17887 40053 17888 ne
rect 40053 17887 40182 17888
tri 40053 17886 40054 17887 ne
rect 40054 17886 40182 17887
tri 40054 17885 40055 17886 ne
rect 40055 17885 40182 17886
tri 40055 17884 40056 17885 ne
rect 40056 17884 40182 17885
tri 40056 17883 40057 17884 ne
rect 40057 17883 40182 17884
tri 40057 17882 40058 17883 ne
rect 40058 17882 40182 17883
tri 40058 17881 40059 17882 ne
rect 40059 17881 40182 17882
tri 40059 17880 40060 17881 ne
rect 40060 17880 40182 17881
tri 40060 17879 40061 17880 ne
rect 40061 17879 40182 17880
tri 40061 17878 40062 17879 ne
rect 40062 17878 40182 17879
tri 40062 17877 40063 17878 ne
rect 40063 17877 40182 17878
tri 40063 17876 40064 17877 ne
rect 40064 17876 40182 17877
tri 40064 17875 40065 17876 ne
rect 40065 17875 40182 17876
tri 40065 17874 40066 17875 ne
rect 40066 17874 40182 17875
tri 40066 17873 40067 17874 ne
rect 40067 17873 40182 17874
tri 40067 17872 40068 17873 ne
rect 40068 17872 40182 17873
tri 40068 17871 40069 17872 ne
rect 40069 17871 40182 17872
tri 40069 17870 40070 17871 ne
rect 40070 17870 40182 17871
tri 40070 17869 40071 17870 ne
rect 40071 17869 40182 17870
tri 40071 17868 40072 17869 ne
rect 40072 17868 40182 17869
tri 40072 17867 40073 17868 ne
rect 40073 17867 40182 17868
tri 40073 17866 40074 17867 ne
rect 40074 17866 40182 17867
tri 40074 17865 40075 17866 ne
rect 40075 17865 40182 17866
tri 40075 17864 40076 17865 ne
rect 40076 17864 40182 17865
tri 40076 17863 40077 17864 ne
rect 40077 17863 40182 17864
tri 40077 17862 40078 17863 ne
rect 40078 17862 40182 17863
tri 40078 17861 40079 17862 ne
rect 40079 17861 40182 17862
tri 40079 17860 40080 17861 ne
rect 40080 17860 40182 17861
tri 40080 17859 40081 17860 ne
rect 40081 17859 40182 17860
tri 40081 17858 40082 17859 ne
rect 40082 17858 40182 17859
tri 40082 17857 40083 17858 ne
rect 40083 17857 40182 17858
tri 40083 17856 40084 17857 ne
rect 40084 17856 40182 17857
tri 40084 17855 40085 17856 ne
rect 40085 17855 40182 17856
tri 40085 17854 40086 17855 ne
rect 40086 17854 40182 17855
tri 40086 17853 40087 17854 ne
rect 40087 17853 40182 17854
tri 40087 17852 40088 17853 ne
rect 40088 17852 40182 17853
tri 40088 17851 40089 17852 ne
rect 40089 17851 40182 17852
tri 40089 17850 40090 17851 ne
rect 40090 17850 40182 17851
rect 40228 17868 40303 17896
tri 40303 17868 40348 17913 sw
rect 70802 17908 71000 17966
rect 40228 17850 40348 17868
tri 40090 17849 40091 17850 ne
rect 40091 17849 40348 17850
tri 40091 17848 40092 17849 ne
rect 40092 17848 40348 17849
tri 40092 17847 40093 17848 ne
rect 40093 17847 40348 17848
tri 40093 17846 40094 17847 ne
rect 40094 17846 40348 17847
tri 40094 17845 40095 17846 ne
rect 40095 17845 40348 17846
tri 40095 17844 40096 17845 ne
rect 40096 17844 40348 17845
tri 40096 17843 40097 17844 ne
rect 40097 17843 40348 17844
tri 40097 17842 40098 17843 ne
rect 40098 17842 40348 17843
tri 40098 17841 40099 17842 ne
rect 40099 17841 40348 17842
tri 40099 17840 40100 17841 ne
rect 40100 17840 40348 17841
tri 40100 17839 40101 17840 ne
rect 40101 17839 40348 17840
tri 40101 17838 40102 17839 ne
rect 40102 17838 40348 17839
tri 40102 17837 40103 17838 ne
rect 40103 17837 40348 17838
tri 40103 17836 40104 17837 ne
rect 40104 17836 40348 17837
tri 40104 17835 40105 17836 ne
rect 40105 17835 40348 17836
tri 40105 17834 40106 17835 ne
rect 40106 17834 40348 17835
tri 40106 17833 40107 17834 ne
rect 40107 17833 40348 17834
tri 40107 17832 40108 17833 ne
rect 40108 17832 40348 17833
tri 40108 17831 40109 17832 ne
rect 40109 17831 40348 17832
tri 40109 17830 40110 17831 ne
rect 40110 17830 40348 17831
tri 40110 17829 40111 17830 ne
rect 40111 17829 40348 17830
tri 40111 17828 40112 17829 ne
rect 40112 17828 40348 17829
tri 40112 17827 40113 17828 ne
rect 40113 17827 40348 17828
tri 40113 17826 40114 17827 ne
rect 40114 17826 40348 17827
tri 40114 17825 40115 17826 ne
rect 40115 17825 40348 17826
tri 40115 17824 40116 17825 ne
rect 40116 17824 40348 17825
tri 40116 17823 40117 17824 ne
rect 40117 17823 40348 17824
tri 40348 17823 40393 17868 sw
rect 70802 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
tri 40117 17822 40118 17823 ne
rect 40118 17822 40393 17823
tri 40118 17821 40119 17822 ne
rect 40119 17821 40393 17822
tri 40119 17820 40120 17821 ne
rect 40120 17820 40393 17821
tri 40120 17819 40121 17820 ne
rect 40121 17819 40393 17820
tri 40121 17818 40122 17819 ne
rect 40122 17818 40393 17819
tri 40122 17817 40123 17818 ne
rect 40123 17817 40393 17818
tri 40123 17816 40124 17817 ne
rect 40124 17816 40393 17817
tri 40124 17815 40125 17816 ne
rect 40125 17815 40393 17816
tri 40125 17814 40126 17815 ne
rect 40126 17814 40393 17815
tri 40126 17813 40127 17814 ne
rect 40127 17813 40393 17814
tri 40127 17812 40128 17813 ne
rect 40128 17812 40393 17813
tri 40128 17811 40129 17812 ne
rect 40129 17811 40393 17812
tri 40129 17810 40130 17811 ne
rect 40130 17810 40393 17811
tri 40130 17809 40131 17810 ne
rect 40131 17809 40393 17810
tri 40131 17808 40132 17809 ne
rect 40132 17808 40393 17809
tri 40132 17807 40133 17808 ne
rect 40133 17807 40393 17808
tri 40133 17806 40134 17807 ne
rect 40134 17806 40393 17807
tri 40134 17805 40135 17806 ne
rect 40135 17805 40393 17806
tri 40135 17804 40136 17805 ne
rect 40136 17804 40393 17805
tri 40136 17803 40137 17804 ne
rect 40137 17803 40393 17804
tri 40137 17802 40138 17803 ne
rect 40138 17802 40393 17803
tri 40138 17801 40139 17802 ne
rect 40139 17801 40393 17802
tri 40139 17800 40140 17801 ne
rect 40140 17800 40393 17801
tri 40140 17799 40141 17800 ne
rect 40141 17799 40393 17800
tri 40141 17798 40142 17799 ne
rect 40142 17798 40393 17799
tri 40142 17797 40143 17798 ne
rect 40143 17797 40393 17798
tri 40143 17796 40144 17797 ne
rect 40144 17796 40393 17797
tri 40144 17795 40145 17796 ne
rect 40145 17795 40393 17796
tri 40145 17794 40146 17795 ne
rect 40146 17794 40393 17795
tri 40146 17793 40147 17794 ne
rect 40147 17793 40393 17794
tri 40147 17792 40148 17793 ne
rect 40148 17792 40393 17793
tri 40148 17791 40149 17792 ne
rect 40149 17791 40393 17792
tri 40149 17790 40150 17791 ne
rect 40150 17790 40393 17791
tri 40150 17789 40151 17790 ne
rect 40151 17789 40393 17790
tri 40393 17789 40427 17823 sw
rect 70802 17804 71000 17862
tri 40151 17746 40194 17789 ne
rect 40194 17778 40427 17789
tri 40427 17778 40438 17789 sw
rect 40194 17764 40438 17778
rect 40194 17746 40314 17764
tri 40194 17701 40239 17746 ne
rect 40239 17718 40314 17746
rect 40360 17733 40438 17764
tri 40438 17733 40483 17778 sw
rect 70802 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17718 40483 17733
rect 40239 17701 40483 17718
tri 40239 17681 40259 17701 ne
rect 40259 17688 40483 17701
tri 40483 17688 40528 17733 sw
rect 70802 17700 71000 17758
rect 40259 17681 40528 17688
tri 40259 17680 40260 17681 ne
rect 40260 17680 40528 17681
tri 40260 17679 40261 17680 ne
rect 40261 17679 40528 17680
tri 40261 17678 40262 17679 ne
rect 40262 17678 40528 17679
tri 40262 17677 40263 17678 ne
rect 40263 17677 40528 17678
tri 40263 17676 40264 17677 ne
rect 40264 17676 40528 17677
tri 40264 17675 40265 17676 ne
rect 40265 17675 40528 17676
tri 40265 17674 40266 17675 ne
rect 40266 17674 40528 17675
tri 40266 17673 40267 17674 ne
rect 40267 17673 40528 17674
tri 40267 17672 40268 17673 ne
rect 40268 17672 40528 17673
tri 40268 17671 40269 17672 ne
rect 40269 17671 40528 17672
tri 40269 17670 40270 17671 ne
rect 40270 17670 40528 17671
tri 40270 17669 40271 17670 ne
rect 40271 17669 40528 17670
tri 40271 17668 40272 17669 ne
rect 40272 17668 40528 17669
tri 40272 17667 40273 17668 ne
rect 40273 17667 40528 17668
tri 40273 17666 40274 17667 ne
rect 40274 17666 40528 17667
tri 40274 17665 40275 17666 ne
rect 40275 17665 40528 17666
tri 40275 17664 40276 17665 ne
rect 40276 17664 40528 17665
tri 40276 17663 40277 17664 ne
rect 40277 17663 40528 17664
tri 40277 17662 40278 17663 ne
rect 40278 17662 40528 17663
tri 40278 17661 40279 17662 ne
rect 40279 17661 40528 17662
tri 40279 17660 40280 17661 ne
rect 40280 17660 40528 17661
tri 40280 17659 40281 17660 ne
rect 40281 17659 40528 17660
tri 40281 17658 40282 17659 ne
rect 40282 17658 40528 17659
tri 40282 17657 40283 17658 ne
rect 40283 17657 40528 17658
tri 40283 17656 40284 17657 ne
rect 40284 17656 40528 17657
tri 40284 17655 40285 17656 ne
rect 40285 17655 40528 17656
tri 40285 17654 40286 17655 ne
rect 40286 17654 40528 17655
tri 40286 17653 40287 17654 ne
rect 40287 17653 40528 17654
tri 40287 17652 40288 17653 ne
rect 40288 17652 40528 17653
tri 40288 17651 40289 17652 ne
rect 40289 17651 40528 17652
tri 40289 17650 40290 17651 ne
rect 40290 17650 40528 17651
tri 40290 17649 40291 17650 ne
rect 40291 17649 40528 17650
tri 40291 17648 40292 17649 ne
rect 40292 17648 40528 17649
tri 40528 17648 40568 17688 sw
rect 70802 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40292 17647 40293 17648 ne
rect 40293 17647 40568 17648
tri 40293 17646 40294 17647 ne
rect 40294 17646 40568 17647
tri 40294 17645 40295 17646 ne
rect 40295 17645 40568 17646
tri 40295 17644 40296 17645 ne
rect 40296 17644 40568 17645
tri 40296 17643 40297 17644 ne
rect 40297 17643 40568 17644
tri 40297 17642 40298 17643 ne
rect 40298 17642 40568 17643
tri 40298 17641 40299 17642 ne
rect 40299 17641 40568 17642
tri 40299 17640 40300 17641 ne
rect 40300 17640 40568 17641
tri 40300 17639 40301 17640 ne
rect 40301 17639 40568 17640
tri 40301 17638 40302 17639 ne
rect 40302 17638 40568 17639
tri 40302 17637 40303 17638 ne
rect 40303 17637 40568 17638
tri 40303 17636 40304 17637 ne
rect 40304 17636 40568 17637
tri 40304 17635 40305 17636 ne
rect 40305 17635 40568 17636
tri 40305 17634 40306 17635 ne
rect 40306 17634 40568 17635
tri 40306 17633 40307 17634 ne
rect 40307 17633 40568 17634
tri 40307 17632 40308 17633 ne
rect 40308 17632 40568 17633
tri 40308 17631 40309 17632 ne
rect 40309 17631 40446 17632
tri 40309 17630 40310 17631 ne
rect 40310 17630 40446 17631
tri 40310 17629 40311 17630 ne
rect 40311 17629 40446 17630
tri 40311 17628 40312 17629 ne
rect 40312 17628 40446 17629
tri 40312 17627 40313 17628 ne
rect 40313 17627 40446 17628
tri 40313 17626 40314 17627 ne
rect 40314 17626 40446 17627
tri 40314 17625 40315 17626 ne
rect 40315 17625 40446 17626
tri 40315 17624 40316 17625 ne
rect 40316 17624 40446 17625
tri 40316 17623 40317 17624 ne
rect 40317 17623 40446 17624
tri 40317 17622 40318 17623 ne
rect 40318 17622 40446 17623
tri 40318 17621 40319 17622 ne
rect 40319 17621 40446 17622
tri 40319 17620 40320 17621 ne
rect 40320 17620 40446 17621
tri 40320 17619 40321 17620 ne
rect 40321 17619 40446 17620
tri 40321 17618 40322 17619 ne
rect 40322 17618 40446 17619
tri 40322 17617 40323 17618 ne
rect 40323 17617 40446 17618
tri 40323 17616 40324 17617 ne
rect 40324 17616 40446 17617
tri 40324 17615 40325 17616 ne
rect 40325 17615 40446 17616
tri 40325 17614 40326 17615 ne
rect 40326 17614 40446 17615
tri 40326 17613 40327 17614 ne
rect 40327 17613 40446 17614
tri 40327 17612 40328 17613 ne
rect 40328 17612 40446 17613
tri 40328 17611 40329 17612 ne
rect 40329 17611 40446 17612
tri 40329 17610 40330 17611 ne
rect 40330 17610 40446 17611
tri 40330 17609 40331 17610 ne
rect 40331 17609 40446 17610
tri 40331 17608 40332 17609 ne
rect 40332 17608 40446 17609
tri 40332 17607 40333 17608 ne
rect 40333 17607 40446 17608
tri 40333 17606 40334 17607 ne
rect 40334 17606 40446 17607
tri 40334 17605 40335 17606 ne
rect 40335 17605 40446 17606
tri 40335 17604 40336 17605 ne
rect 40336 17604 40446 17605
tri 40336 17603 40337 17604 ne
rect 40337 17603 40446 17604
tri 40337 17602 40338 17603 ne
rect 40338 17602 40446 17603
tri 40338 17601 40339 17602 ne
rect 40339 17601 40446 17602
tri 40339 17600 40340 17601 ne
rect 40340 17600 40446 17601
tri 40340 17599 40341 17600 ne
rect 40341 17599 40446 17600
tri 40341 17598 40342 17599 ne
rect 40342 17598 40446 17599
tri 40342 17597 40343 17598 ne
rect 40343 17597 40446 17598
tri 40343 17596 40344 17597 ne
rect 40344 17596 40446 17597
tri 40344 17595 40345 17596 ne
rect 40345 17595 40446 17596
tri 40345 17594 40346 17595 ne
rect 40346 17594 40446 17595
tri 40346 17593 40347 17594 ne
rect 40347 17593 40446 17594
tri 40347 17592 40348 17593 ne
rect 40348 17592 40446 17593
tri 40348 17591 40349 17592 ne
rect 40349 17591 40446 17592
tri 40349 17590 40350 17591 ne
rect 40350 17590 40446 17591
tri 40350 17589 40351 17590 ne
rect 40351 17589 40446 17590
tri 40351 17588 40352 17589 ne
rect 40352 17588 40446 17589
tri 40352 17587 40353 17588 ne
rect 40353 17587 40446 17588
tri 40353 17586 40354 17587 ne
rect 40354 17586 40446 17587
rect 40492 17603 40568 17632
tri 40568 17603 40613 17648 sw
rect 40492 17586 40613 17603
tri 40354 17585 40355 17586 ne
rect 40355 17585 40613 17586
tri 40355 17584 40356 17585 ne
rect 40356 17584 40613 17585
tri 40356 17583 40357 17584 ne
rect 40357 17583 40613 17584
tri 40357 17582 40358 17583 ne
rect 40358 17582 40613 17583
tri 40358 17581 40359 17582 ne
rect 40359 17581 40613 17582
tri 40359 17580 40360 17581 ne
rect 40360 17580 40613 17581
tri 40360 17579 40361 17580 ne
rect 40361 17579 40613 17580
tri 40361 17578 40362 17579 ne
rect 40362 17578 40613 17579
tri 40362 17577 40363 17578 ne
rect 40363 17577 40613 17578
tri 40363 17576 40364 17577 ne
rect 40364 17576 40613 17577
tri 40364 17575 40365 17576 ne
rect 40365 17575 40613 17576
tri 40365 17574 40366 17575 ne
rect 40366 17574 40613 17575
tri 40366 17573 40367 17574 ne
rect 40367 17573 40613 17574
tri 40367 17572 40368 17573 ne
rect 40368 17572 40613 17573
tri 40368 17571 40369 17572 ne
rect 40369 17571 40613 17572
tri 40369 17570 40370 17571 ne
rect 40370 17570 40613 17571
tri 40370 17569 40371 17570 ne
rect 40371 17569 40613 17570
tri 40371 17568 40372 17569 ne
rect 40372 17568 40613 17569
tri 40372 17567 40373 17568 ne
rect 40373 17567 40613 17568
tri 40373 17566 40374 17567 ne
rect 40374 17566 40613 17567
tri 40374 17565 40375 17566 ne
rect 40375 17565 40613 17566
tri 40375 17564 40376 17565 ne
rect 40376 17564 40613 17565
tri 40376 17563 40377 17564 ne
rect 40377 17563 40613 17564
tri 40377 17562 40378 17563 ne
rect 40378 17562 40613 17563
tri 40378 17561 40379 17562 ne
rect 40379 17561 40613 17562
tri 40379 17560 40380 17561 ne
rect 40380 17560 40613 17561
tri 40380 17559 40381 17560 ne
rect 40381 17559 40613 17560
tri 40381 17558 40382 17559 ne
rect 40382 17558 40613 17559
tri 40613 17558 40658 17603 sw
rect 70802 17596 71000 17654
tri 40382 17557 40383 17558 ne
rect 40383 17557 40658 17558
tri 40383 17556 40384 17557 ne
rect 40384 17556 40658 17557
tri 40384 17555 40385 17556 ne
rect 40385 17555 40658 17556
tri 40385 17554 40386 17555 ne
rect 40386 17554 40658 17555
tri 40386 17553 40387 17554 ne
rect 40387 17553 40658 17554
tri 40387 17552 40388 17553 ne
rect 40388 17552 40658 17553
tri 40388 17551 40389 17552 ne
rect 40389 17551 40658 17552
tri 40389 17550 40390 17551 ne
rect 40390 17550 40658 17551
tri 40390 17549 40391 17550 ne
rect 40391 17549 40658 17550
tri 40391 17548 40392 17549 ne
rect 40392 17548 40658 17549
tri 40392 17547 40393 17548 ne
rect 40393 17547 40658 17548
tri 40393 17546 40394 17547 ne
rect 40394 17546 40658 17547
tri 40394 17545 40395 17546 ne
rect 40395 17545 40658 17546
tri 40395 17544 40396 17545 ne
rect 40396 17544 40658 17545
tri 40396 17543 40397 17544 ne
rect 40397 17543 40658 17544
tri 40397 17542 40398 17543 ne
rect 40398 17542 40658 17543
tri 40398 17541 40399 17542 ne
rect 40399 17541 40658 17542
tri 40399 17540 40400 17541 ne
rect 40400 17540 40658 17541
tri 40400 17539 40401 17540 ne
rect 40401 17539 40658 17540
tri 40401 17538 40402 17539 ne
rect 40402 17538 40658 17539
tri 40402 17537 40403 17538 ne
rect 40403 17537 40658 17538
tri 40403 17536 40404 17537 ne
rect 40404 17536 40658 17537
tri 40404 17535 40405 17536 ne
rect 40405 17535 40658 17536
tri 40405 17534 40406 17535 ne
rect 40406 17534 40658 17535
tri 40406 17533 40407 17534 ne
rect 40407 17533 40658 17534
tri 40407 17532 40408 17533 ne
rect 40408 17532 40658 17533
tri 40408 17531 40409 17532 ne
rect 40409 17531 40658 17532
tri 40409 17530 40410 17531 ne
rect 40410 17530 40658 17531
tri 40410 17529 40411 17530 ne
rect 40411 17529 40658 17530
tri 40411 17528 40412 17529 ne
rect 40412 17528 40658 17529
tri 40412 17527 40413 17528 ne
rect 40413 17527 40658 17528
tri 40413 17526 40414 17527 ne
rect 40414 17526 40658 17527
tri 40414 17525 40415 17526 ne
rect 40415 17525 40658 17526
tri 40415 17524 40416 17525 ne
rect 40416 17524 40658 17525
tri 40416 17523 40417 17524 ne
rect 40417 17523 40658 17524
tri 40417 17522 40418 17523 ne
rect 40418 17522 40658 17523
tri 40418 17521 40419 17522 ne
rect 40419 17521 40658 17522
tri 40419 17520 40420 17521 ne
rect 40420 17520 40658 17521
tri 40420 17519 40421 17520 ne
rect 40421 17519 40658 17520
tri 40421 17518 40422 17519 ne
rect 40422 17518 40658 17519
tri 40422 17517 40423 17518 ne
rect 40423 17517 40658 17518
tri 40423 17516 40424 17517 ne
rect 40424 17516 40658 17517
tri 40424 17515 40425 17516 ne
rect 40425 17515 40658 17516
tri 40425 17514 40426 17515 ne
rect 40426 17514 40658 17515
tri 40426 17513 40427 17514 ne
rect 40427 17513 40658 17514
tri 40658 17513 40703 17558 sw
rect 70802 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
tri 40427 17502 40438 17513 ne
rect 40438 17502 40703 17513
tri 40703 17502 40714 17513 sw
tri 40438 17468 40472 17502 ne
rect 40472 17500 40714 17502
rect 40472 17468 40578 17500
tri 40472 17457 40483 17468 ne
rect 40483 17457 40578 17468
tri 40483 17412 40528 17457 ne
rect 40528 17454 40578 17457
rect 40624 17457 40714 17500
tri 40714 17457 40759 17502 sw
rect 70802 17492 71000 17550
rect 40624 17454 40759 17457
rect 40528 17412 40759 17454
tri 40759 17412 40804 17457 sw
rect 70802 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
tri 40528 17407 40533 17412 ne
rect 40533 17407 40804 17412
tri 40533 17406 40534 17407 ne
rect 40534 17406 40804 17407
tri 40534 17405 40535 17406 ne
rect 40535 17405 40804 17406
tri 40535 17404 40536 17405 ne
rect 40536 17404 40804 17405
tri 40536 17403 40537 17404 ne
rect 40537 17403 40804 17404
tri 40537 17402 40538 17403 ne
rect 40538 17402 40804 17403
tri 40538 17401 40539 17402 ne
rect 40539 17401 40804 17402
tri 40539 17400 40540 17401 ne
rect 40540 17400 40804 17401
tri 40540 17399 40541 17400 ne
rect 40541 17399 40804 17400
tri 40541 17398 40542 17399 ne
rect 40542 17398 40804 17399
tri 40542 17397 40543 17398 ne
rect 40543 17397 40804 17398
tri 40543 17396 40544 17397 ne
rect 40544 17396 40804 17397
tri 40544 17395 40545 17396 ne
rect 40545 17395 40804 17396
tri 40545 17394 40546 17395 ne
rect 40546 17394 40804 17395
tri 40546 17393 40547 17394 ne
rect 40547 17393 40804 17394
tri 40547 17392 40548 17393 ne
rect 40548 17392 40804 17393
tri 40548 17391 40549 17392 ne
rect 40549 17391 40804 17392
tri 40549 17390 40550 17391 ne
rect 40550 17390 40804 17391
tri 40550 17389 40551 17390 ne
rect 40551 17389 40804 17390
tri 40551 17388 40552 17389 ne
rect 40552 17388 40804 17389
tri 40552 17387 40553 17388 ne
rect 40553 17387 40804 17388
tri 40553 17386 40554 17387 ne
rect 40554 17386 40804 17387
tri 40554 17385 40555 17386 ne
rect 40555 17385 40804 17386
tri 40555 17384 40556 17385 ne
rect 40556 17384 40804 17385
tri 40556 17383 40557 17384 ne
rect 40557 17383 40804 17384
tri 40557 17382 40558 17383 ne
rect 40558 17382 40804 17383
tri 40558 17381 40559 17382 ne
rect 40559 17381 40804 17382
tri 40559 17380 40560 17381 ne
rect 40560 17380 40804 17381
tri 40560 17379 40561 17380 ne
rect 40561 17379 40804 17380
tri 40561 17378 40562 17379 ne
rect 40562 17378 40804 17379
tri 40562 17377 40563 17378 ne
rect 40563 17377 40804 17378
tri 40563 17376 40564 17377 ne
rect 40564 17376 40804 17377
tri 40564 17375 40565 17376 ne
rect 40565 17375 40804 17376
tri 40565 17374 40566 17375 ne
rect 40566 17374 40804 17375
tri 40566 17373 40567 17374 ne
rect 40567 17373 40804 17374
tri 40567 17372 40568 17373 ne
rect 40568 17372 40804 17373
tri 40568 17371 40569 17372 ne
rect 40569 17371 40804 17372
tri 40569 17370 40570 17371 ne
rect 40570 17370 40804 17371
tri 40570 17369 40571 17370 ne
rect 40571 17369 40804 17370
tri 40571 17368 40572 17369 ne
rect 40572 17368 40804 17369
tri 40572 17367 40573 17368 ne
rect 40573 17367 40710 17368
tri 40573 17366 40574 17367 ne
rect 40574 17366 40710 17367
tri 40574 17365 40575 17366 ne
rect 40575 17365 40710 17366
tri 40575 17364 40576 17365 ne
rect 40576 17364 40710 17365
tri 40576 17363 40577 17364 ne
rect 40577 17363 40710 17364
tri 40577 17362 40578 17363 ne
rect 40578 17362 40710 17363
tri 40578 17361 40579 17362 ne
rect 40579 17361 40710 17362
tri 40579 17360 40580 17361 ne
rect 40580 17360 40710 17361
tri 40580 17359 40581 17360 ne
rect 40581 17359 40710 17360
tri 40581 17358 40582 17359 ne
rect 40582 17358 40710 17359
tri 40582 17357 40583 17358 ne
rect 40583 17357 40710 17358
tri 40583 17356 40584 17357 ne
rect 40584 17356 40710 17357
tri 40584 17355 40585 17356 ne
rect 40585 17355 40710 17356
tri 40585 17354 40586 17355 ne
rect 40586 17354 40710 17355
tri 40586 17353 40587 17354 ne
rect 40587 17353 40710 17354
tri 40587 17352 40588 17353 ne
rect 40588 17352 40710 17353
tri 40588 17351 40589 17352 ne
rect 40589 17351 40710 17352
tri 40589 17350 40590 17351 ne
rect 40590 17350 40710 17351
tri 40590 17349 40591 17350 ne
rect 40591 17349 40710 17350
tri 40591 17348 40592 17349 ne
rect 40592 17348 40710 17349
tri 40592 17347 40593 17348 ne
rect 40593 17347 40710 17348
tri 40593 17346 40594 17347 ne
rect 40594 17346 40710 17347
tri 40594 17345 40595 17346 ne
rect 40595 17345 40710 17346
tri 40595 17344 40596 17345 ne
rect 40596 17344 40710 17345
tri 40596 17343 40597 17344 ne
rect 40597 17343 40710 17344
tri 40597 17342 40598 17343 ne
rect 40598 17342 40710 17343
tri 40598 17341 40599 17342 ne
rect 40599 17341 40710 17342
tri 40599 17340 40600 17341 ne
rect 40600 17340 40710 17341
tri 40600 17339 40601 17340 ne
rect 40601 17339 40710 17340
tri 40601 17338 40602 17339 ne
rect 40602 17338 40710 17339
tri 40602 17337 40603 17338 ne
rect 40603 17337 40710 17338
tri 40603 17336 40604 17337 ne
rect 40604 17336 40710 17337
tri 40604 17335 40605 17336 ne
rect 40605 17335 40710 17336
tri 40605 17334 40606 17335 ne
rect 40606 17334 40710 17335
tri 40606 17333 40607 17334 ne
rect 40607 17333 40710 17334
tri 40607 17332 40608 17333 ne
rect 40608 17332 40710 17333
tri 40608 17331 40609 17332 ne
rect 40609 17331 40710 17332
tri 40609 17330 40610 17331 ne
rect 40610 17330 40710 17331
tri 40610 17329 40611 17330 ne
rect 40611 17329 40710 17330
tri 40611 17328 40612 17329 ne
rect 40612 17328 40710 17329
tri 40612 17327 40613 17328 ne
rect 40613 17327 40710 17328
tri 40613 17326 40614 17327 ne
rect 40614 17326 40710 17327
tri 40614 17325 40615 17326 ne
rect 40615 17325 40710 17326
tri 40615 17324 40616 17325 ne
rect 40616 17324 40710 17325
tri 40616 17323 40617 17324 ne
rect 40617 17323 40710 17324
tri 40617 17322 40618 17323 ne
rect 40618 17322 40710 17323
rect 40756 17367 40804 17368
tri 40804 17367 40849 17412 sw
rect 70802 17388 71000 17446
rect 40756 17327 40849 17367
tri 40849 17327 40889 17367 sw
rect 70802 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17322 40889 17327
tri 40618 17321 40619 17322 ne
rect 40619 17321 40889 17322
tri 40619 17320 40620 17321 ne
rect 40620 17320 40889 17321
tri 40620 17319 40621 17320 ne
rect 40621 17319 40889 17320
tri 40621 17318 40622 17319 ne
rect 40622 17318 40889 17319
tri 40622 17317 40623 17318 ne
rect 40623 17317 40889 17318
tri 40623 17316 40624 17317 ne
rect 40624 17316 40889 17317
tri 40624 17315 40625 17316 ne
rect 40625 17315 40889 17316
tri 40625 17314 40626 17315 ne
rect 40626 17314 40889 17315
tri 40626 17313 40627 17314 ne
rect 40627 17313 40889 17314
tri 40627 17312 40628 17313 ne
rect 40628 17312 40889 17313
tri 40628 17311 40629 17312 ne
rect 40629 17311 40889 17312
tri 40629 17310 40630 17311 ne
rect 40630 17310 40889 17311
tri 40630 17309 40631 17310 ne
rect 40631 17309 40889 17310
tri 40631 17308 40632 17309 ne
rect 40632 17308 40889 17309
tri 40632 17307 40633 17308 ne
rect 40633 17307 40889 17308
tri 40633 17306 40634 17307 ne
rect 40634 17306 40889 17307
tri 40634 17305 40635 17306 ne
rect 40635 17305 40889 17306
tri 40635 17304 40636 17305 ne
rect 40636 17304 40889 17305
tri 40636 17303 40637 17304 ne
rect 40637 17303 40889 17304
tri 40637 17302 40638 17303 ne
rect 40638 17302 40889 17303
tri 40638 17301 40639 17302 ne
rect 40639 17301 40889 17302
tri 40639 17300 40640 17301 ne
rect 40640 17300 40889 17301
tri 40640 17299 40641 17300 ne
rect 40641 17299 40889 17300
tri 40641 17298 40642 17299 ne
rect 40642 17298 40889 17299
tri 40642 17297 40643 17298 ne
rect 40643 17297 40889 17298
tri 40643 17296 40644 17297 ne
rect 40644 17296 40889 17297
tri 40644 17295 40645 17296 ne
rect 40645 17295 40889 17296
tri 40645 17294 40646 17295 ne
rect 40646 17294 40889 17295
tri 40646 17293 40647 17294 ne
rect 40647 17293 40889 17294
tri 40647 17292 40648 17293 ne
rect 40648 17292 40889 17293
tri 40648 17291 40649 17292 ne
rect 40649 17291 40889 17292
tri 40649 17290 40650 17291 ne
rect 40650 17290 40889 17291
tri 40650 17289 40651 17290 ne
rect 40651 17289 40889 17290
tri 40651 17288 40652 17289 ne
rect 40652 17288 40889 17289
tri 40652 17287 40653 17288 ne
rect 40653 17287 40889 17288
tri 40653 17286 40654 17287 ne
rect 40654 17286 40889 17287
tri 40654 17285 40655 17286 ne
rect 40655 17285 40889 17286
tri 40655 17284 40656 17285 ne
rect 40656 17284 40889 17285
tri 40656 17283 40657 17284 ne
rect 40657 17283 40889 17284
tri 40657 17282 40658 17283 ne
rect 40658 17282 40889 17283
tri 40889 17282 40934 17327 sw
rect 70802 17284 71000 17342
tri 40658 17281 40659 17282 ne
rect 40659 17281 40934 17282
tri 40659 17280 40660 17281 ne
rect 40660 17280 40934 17281
tri 40660 17279 40661 17280 ne
rect 40661 17279 40934 17280
tri 40661 17278 40662 17279 ne
rect 40662 17278 40934 17279
tri 40662 17277 40663 17278 ne
rect 40663 17277 40934 17278
tri 40663 17276 40664 17277 ne
rect 40664 17276 40934 17277
tri 40664 17275 40665 17276 ne
rect 40665 17275 40934 17276
tri 40665 17274 40666 17275 ne
rect 40666 17274 40934 17275
tri 40666 17273 40667 17274 ne
rect 40667 17273 40934 17274
tri 40667 17272 40668 17273 ne
rect 40668 17272 40934 17273
tri 40668 17271 40669 17272 ne
rect 40669 17271 40934 17272
tri 40669 17270 40670 17271 ne
rect 40670 17270 40934 17271
tri 40670 17269 40671 17270 ne
rect 40671 17269 40934 17270
tri 40671 17268 40672 17269 ne
rect 40672 17268 40934 17269
tri 40672 17267 40673 17268 ne
rect 40673 17267 40934 17268
tri 40673 17266 40674 17267 ne
rect 40674 17266 40934 17267
tri 40674 17265 40675 17266 ne
rect 40675 17265 40934 17266
tri 40675 17264 40676 17265 ne
rect 40676 17264 40934 17265
tri 40676 17263 40677 17264 ne
rect 40677 17263 40934 17264
tri 40677 17262 40678 17263 ne
rect 40678 17262 40934 17263
tri 40678 17261 40679 17262 ne
rect 40679 17261 40934 17262
tri 40679 17260 40680 17261 ne
rect 40680 17260 40934 17261
tri 40680 17259 40681 17260 ne
rect 40681 17259 40934 17260
tri 40681 17258 40682 17259 ne
rect 40682 17258 40934 17259
tri 40682 17257 40683 17258 ne
rect 40683 17257 40934 17258
tri 40683 17256 40684 17257 ne
rect 40684 17256 40934 17257
tri 40684 17255 40685 17256 ne
rect 40685 17255 40934 17256
tri 40685 17254 40686 17255 ne
rect 40686 17254 40934 17255
tri 40686 17253 40687 17254 ne
rect 40687 17253 40934 17254
tri 40687 17252 40688 17253 ne
rect 40688 17252 40934 17253
tri 40688 17251 40689 17252 ne
rect 40689 17251 40934 17252
tri 40689 17250 40690 17251 ne
rect 40690 17250 40934 17251
tri 40690 17249 40691 17250 ne
rect 40691 17249 40934 17250
tri 40691 17248 40692 17249 ne
rect 40692 17248 40934 17249
tri 40692 17247 40693 17248 ne
rect 40693 17247 40934 17248
tri 40693 17246 40694 17247 ne
rect 40694 17246 40934 17247
tri 40694 17245 40695 17246 ne
rect 40695 17245 40934 17246
tri 40695 17244 40696 17245 ne
rect 40696 17244 40934 17245
tri 40696 17243 40697 17244 ne
rect 40697 17243 40934 17244
tri 40697 17242 40698 17243 ne
rect 40698 17242 40934 17243
tri 40698 17241 40699 17242 ne
rect 40699 17241 40934 17242
tri 40699 17240 40700 17241 ne
rect 40700 17240 40934 17241
tri 40700 17239 40701 17240 ne
rect 40701 17239 40934 17240
tri 40701 17238 40702 17239 ne
rect 40702 17238 40934 17239
tri 40702 17237 40703 17238 ne
rect 40703 17237 40934 17238
tri 40934 17237 40979 17282 sw
rect 70802 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
tri 40703 17192 40748 17237 ne
rect 40748 17236 40979 17237
rect 40748 17192 40842 17236
tri 40748 17147 40793 17192 ne
rect 40793 17190 40842 17192
rect 40888 17192 40979 17236
tri 40979 17192 41024 17237 sw
rect 40888 17190 41024 17192
rect 40793 17181 41024 17190
tri 41024 17181 41035 17192 sw
rect 40793 17147 41035 17181
tri 40793 17136 40804 17147 ne
rect 40804 17136 41035 17147
tri 41035 17136 41080 17181 sw
rect 70802 17180 71000 17238
tri 40804 17133 40807 17136 ne
rect 40807 17133 41080 17136
tri 40807 17132 40808 17133 ne
rect 40808 17132 41080 17133
tri 40808 17131 40809 17132 ne
rect 40809 17131 41080 17132
tri 40809 17130 40810 17131 ne
rect 40810 17130 41080 17131
tri 40810 17129 40811 17130 ne
rect 40811 17129 41080 17130
tri 40811 17128 40812 17129 ne
rect 40812 17128 41080 17129
tri 40812 17127 40813 17128 ne
rect 40813 17127 41080 17128
tri 40813 17126 40814 17127 ne
rect 40814 17126 41080 17127
tri 40814 17125 40815 17126 ne
rect 40815 17125 41080 17126
tri 40815 17124 40816 17125 ne
rect 40816 17124 41080 17125
tri 40816 17123 40817 17124 ne
rect 40817 17123 41080 17124
tri 40817 17122 40818 17123 ne
rect 40818 17122 41080 17123
tri 40818 17121 40819 17122 ne
rect 40819 17121 41080 17122
tri 40819 17120 40820 17121 ne
rect 40820 17120 41080 17121
tri 40820 17119 40821 17120 ne
rect 40821 17119 41080 17120
tri 40821 17118 40822 17119 ne
rect 40822 17118 41080 17119
tri 40822 17117 40823 17118 ne
rect 40823 17117 41080 17118
tri 40823 17116 40824 17117 ne
rect 40824 17116 41080 17117
tri 40824 17115 40825 17116 ne
rect 40825 17115 41080 17116
tri 40825 17114 40826 17115 ne
rect 40826 17114 41080 17115
tri 40826 17113 40827 17114 ne
rect 40827 17113 41080 17114
tri 40827 17112 40828 17113 ne
rect 40828 17112 41080 17113
tri 40828 17111 40829 17112 ne
rect 40829 17111 41080 17112
tri 40829 17110 40830 17111 ne
rect 40830 17110 41080 17111
tri 40830 17109 40831 17110 ne
rect 40831 17109 41080 17110
tri 40831 17108 40832 17109 ne
rect 40832 17108 41080 17109
tri 40832 17107 40833 17108 ne
rect 40833 17107 41080 17108
tri 40833 17106 40834 17107 ne
rect 40834 17106 41080 17107
tri 40834 17105 40835 17106 ne
rect 40835 17105 41080 17106
tri 40835 17104 40836 17105 ne
rect 40836 17104 41080 17105
tri 40836 17103 40837 17104 ne
rect 40837 17103 40974 17104
tri 40837 17102 40838 17103 ne
rect 40838 17102 40974 17103
tri 40838 17101 40839 17102 ne
rect 40839 17101 40974 17102
tri 40839 17100 40840 17101 ne
rect 40840 17100 40974 17101
tri 40840 17099 40841 17100 ne
rect 40841 17099 40974 17100
tri 40841 17098 40842 17099 ne
rect 40842 17098 40974 17099
tri 40842 17097 40843 17098 ne
rect 40843 17097 40974 17098
tri 40843 17096 40844 17097 ne
rect 40844 17096 40974 17097
tri 40844 17095 40845 17096 ne
rect 40845 17095 40974 17096
tri 40845 17094 40846 17095 ne
rect 40846 17094 40974 17095
tri 40846 17093 40847 17094 ne
rect 40847 17093 40974 17094
tri 40847 17092 40848 17093 ne
rect 40848 17092 40974 17093
tri 40848 17091 40849 17092 ne
rect 40849 17091 40974 17092
tri 40849 17090 40850 17091 ne
rect 40850 17090 40974 17091
tri 40850 17089 40851 17090 ne
rect 40851 17089 40974 17090
tri 40851 17088 40852 17089 ne
rect 40852 17088 40974 17089
tri 40852 17087 40853 17088 ne
rect 40853 17087 40974 17088
tri 40853 17086 40854 17087 ne
rect 40854 17086 40974 17087
tri 40854 17085 40855 17086 ne
rect 40855 17085 40974 17086
tri 40855 17084 40856 17085 ne
rect 40856 17084 40974 17085
tri 40856 17083 40857 17084 ne
rect 40857 17083 40974 17084
tri 40857 17082 40858 17083 ne
rect 40858 17082 40974 17083
tri 40858 17081 40859 17082 ne
rect 40859 17081 40974 17082
tri 40859 17080 40860 17081 ne
rect 40860 17080 40974 17081
tri 40860 17079 40861 17080 ne
rect 40861 17079 40974 17080
tri 40861 17078 40862 17079 ne
rect 40862 17078 40974 17079
tri 40862 17077 40863 17078 ne
rect 40863 17077 40974 17078
tri 40863 17076 40864 17077 ne
rect 40864 17076 40974 17077
tri 40864 17075 40865 17076 ne
rect 40865 17075 40974 17076
tri 40865 17074 40866 17075 ne
rect 40866 17074 40974 17075
tri 40866 17073 40867 17074 ne
rect 40867 17073 40974 17074
tri 40867 17072 40868 17073 ne
rect 40868 17072 40974 17073
tri 40868 17071 40869 17072 ne
rect 40869 17071 40974 17072
tri 40869 17070 40870 17071 ne
rect 40870 17070 40974 17071
tri 40870 17069 40871 17070 ne
rect 40871 17069 40974 17070
tri 40871 17068 40872 17069 ne
rect 40872 17068 40974 17069
tri 40872 17067 40873 17068 ne
rect 40873 17067 40974 17068
tri 40873 17066 40874 17067 ne
rect 40874 17066 40974 17067
tri 40874 17065 40875 17066 ne
rect 40875 17065 40974 17066
tri 40875 17064 40876 17065 ne
rect 40876 17064 40974 17065
tri 40876 17063 40877 17064 ne
rect 40877 17063 40974 17064
tri 40877 17062 40878 17063 ne
rect 40878 17062 40974 17063
tri 40878 17061 40879 17062 ne
rect 40879 17061 40974 17062
tri 40879 17060 40880 17061 ne
rect 40880 17060 40974 17061
tri 40880 17059 40881 17060 ne
rect 40881 17059 40974 17060
tri 40881 17058 40882 17059 ne
rect 40882 17058 40974 17059
rect 41020 17091 41080 17104
tri 41080 17091 41125 17136 sw
rect 70802 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
rect 41020 17058 41125 17091
tri 40882 17057 40883 17058 ne
rect 40883 17057 41125 17058
tri 40883 17056 40884 17057 ne
rect 40884 17056 41125 17057
tri 40884 17055 40885 17056 ne
rect 40885 17055 41125 17056
tri 40885 17054 40886 17055 ne
rect 40886 17054 41125 17055
tri 40886 17053 40887 17054 ne
rect 40887 17053 41125 17054
tri 40887 17052 40888 17053 ne
rect 40888 17052 41125 17053
tri 40888 17051 40889 17052 ne
rect 40889 17051 41125 17052
tri 40889 17050 40890 17051 ne
rect 40890 17050 41125 17051
tri 40890 17049 40891 17050 ne
rect 40891 17049 41125 17050
tri 40891 17048 40892 17049 ne
rect 40892 17048 41125 17049
tri 40892 17047 40893 17048 ne
rect 40893 17047 41125 17048
tri 40893 17046 40894 17047 ne
rect 40894 17046 41125 17047
tri 41125 17046 41170 17091 sw
rect 70802 17076 71000 17134
tri 40894 17045 40895 17046 ne
rect 40895 17045 41170 17046
tri 40895 17044 40896 17045 ne
rect 40896 17044 41170 17045
tri 40896 17043 40897 17044 ne
rect 40897 17043 41170 17044
tri 40897 17042 40898 17043 ne
rect 40898 17042 41170 17043
tri 40898 17041 40899 17042 ne
rect 40899 17041 41170 17042
tri 40899 17040 40900 17041 ne
rect 40900 17040 41170 17041
tri 40900 17039 40901 17040 ne
rect 40901 17039 41170 17040
tri 40901 17038 40902 17039 ne
rect 40902 17038 41170 17039
tri 40902 17037 40903 17038 ne
rect 40903 17037 41170 17038
tri 40903 17036 40904 17037 ne
rect 40904 17036 41170 17037
tri 40904 17035 40905 17036 ne
rect 40905 17035 41170 17036
tri 40905 17034 40906 17035 ne
rect 40906 17034 41170 17035
tri 40906 17033 40907 17034 ne
rect 40907 17033 41170 17034
tri 40907 17032 40908 17033 ne
rect 40908 17032 41170 17033
tri 40908 17031 40909 17032 ne
rect 40909 17031 41170 17032
tri 40909 17030 40910 17031 ne
rect 40910 17030 41170 17031
tri 40910 17029 40911 17030 ne
rect 40911 17029 41170 17030
tri 40911 17028 40912 17029 ne
rect 40912 17028 41170 17029
tri 40912 17027 40913 17028 ne
rect 40913 17027 41170 17028
tri 40913 17026 40914 17027 ne
rect 40914 17026 41170 17027
tri 40914 17025 40915 17026 ne
rect 40915 17025 41170 17026
tri 40915 17024 40916 17025 ne
rect 40916 17024 41170 17025
tri 40916 17023 40917 17024 ne
rect 40917 17023 41170 17024
tri 40917 17022 40918 17023 ne
rect 40918 17022 41170 17023
tri 40918 17021 40919 17022 ne
rect 40919 17021 41170 17022
tri 40919 17020 40920 17021 ne
rect 40920 17020 41170 17021
tri 40920 17019 40921 17020 ne
rect 40921 17019 41170 17020
tri 40921 17018 40922 17019 ne
rect 40922 17018 41170 17019
tri 40922 17017 40923 17018 ne
rect 40923 17017 41170 17018
tri 40923 17016 40924 17017 ne
rect 40924 17016 41170 17017
tri 40924 17015 40925 17016 ne
rect 40925 17015 41170 17016
tri 40925 17014 40926 17015 ne
rect 40926 17014 41170 17015
tri 40926 17013 40927 17014 ne
rect 40927 17013 41170 17014
tri 40927 17012 40928 17013 ne
rect 40928 17012 41170 17013
tri 40928 17011 40929 17012 ne
rect 40929 17011 41170 17012
tri 40929 17010 40930 17011 ne
rect 40930 17010 41170 17011
tri 40930 17009 40931 17010 ne
rect 40931 17009 41170 17010
tri 40931 17008 40932 17009 ne
rect 40932 17008 41170 17009
tri 40932 17007 40933 17008 ne
rect 40933 17007 41170 17008
tri 40933 17006 40934 17007 ne
rect 40934 17006 41170 17007
tri 41170 17006 41210 17046 sw
rect 70802 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
tri 40934 17005 40935 17006 ne
rect 40935 17005 41210 17006
tri 40935 17004 40936 17005 ne
rect 40936 17004 41210 17005
tri 40936 17003 40937 17004 ne
rect 40937 17003 41210 17004
tri 40937 17002 40938 17003 ne
rect 40938 17002 41210 17003
tri 40938 17001 40939 17002 ne
rect 40939 17001 41210 17002
tri 40939 17000 40940 17001 ne
rect 40940 17000 41210 17001
tri 40940 16999 40941 17000 ne
rect 40941 16999 41210 17000
tri 40941 16998 40942 16999 ne
rect 40942 16998 41210 16999
tri 40942 16997 40943 16998 ne
rect 40943 16997 41210 16998
tri 40943 16996 40944 16997 ne
rect 40944 16996 41210 16997
tri 40944 16995 40945 16996 ne
rect 40945 16995 41210 16996
tri 40945 16994 40946 16995 ne
rect 40946 16994 41210 16995
tri 40946 16993 40947 16994 ne
rect 40947 16993 41210 16994
tri 40947 16992 40948 16993 ne
rect 40948 16992 41210 16993
tri 40948 16991 40949 16992 ne
rect 40949 16991 41210 16992
tri 40949 16990 40950 16991 ne
rect 40950 16990 41210 16991
tri 40950 16989 40951 16990 ne
rect 40951 16989 41210 16990
tri 40951 16988 40952 16989 ne
rect 40952 16988 41210 16989
tri 40952 16987 40953 16988 ne
rect 40953 16987 41210 16988
tri 40953 16986 40954 16987 ne
rect 40954 16986 41210 16987
tri 40954 16985 40955 16986 ne
rect 40955 16985 41210 16986
tri 40955 16984 40956 16985 ne
rect 40956 16984 41210 16985
tri 40956 16983 40957 16984 ne
rect 40957 16983 41210 16984
tri 40957 16982 40958 16983 ne
rect 40958 16982 41210 16983
tri 40958 16981 40959 16982 ne
rect 40959 16981 41210 16982
tri 40959 16980 40960 16981 ne
rect 40960 16980 41210 16981
tri 40960 16979 40961 16980 ne
rect 40961 16979 41210 16980
tri 40961 16978 40962 16979 ne
rect 40962 16978 41210 16979
tri 40962 16977 40963 16978 ne
rect 40963 16977 41210 16978
tri 40963 16976 40964 16977 ne
rect 40964 16976 41210 16977
tri 40964 16975 40965 16976 ne
rect 40965 16975 41210 16976
tri 40965 16974 40966 16975 ne
rect 40966 16974 41210 16975
tri 40966 16973 40967 16974 ne
rect 40967 16973 41210 16974
tri 40967 16972 40968 16973 ne
rect 40968 16972 41210 16973
tri 40968 16971 40969 16972 ne
rect 40969 16971 41106 16972
tri 40969 16970 40970 16971 ne
rect 40970 16970 41106 16971
tri 40970 16969 40971 16970 ne
rect 40971 16969 41106 16970
tri 40971 16968 40972 16969 ne
rect 40972 16968 41106 16969
tri 40972 16967 40973 16968 ne
rect 40973 16967 41106 16968
tri 40973 16966 40974 16967 ne
rect 40974 16966 41106 16967
tri 40974 16965 40975 16966 ne
rect 40975 16965 41106 16966
tri 40975 16964 40976 16965 ne
rect 40976 16964 41106 16965
tri 40976 16963 40977 16964 ne
rect 40977 16963 41106 16964
tri 40977 16962 40978 16963 ne
rect 40978 16962 41106 16963
tri 40978 16961 40979 16962 ne
rect 40979 16961 41106 16962
tri 40979 16916 41024 16961 ne
rect 41024 16926 41106 16961
rect 41152 16961 41210 16972
tri 41210 16961 41255 17006 sw
rect 70802 16972 71000 17030
rect 41152 16926 41255 16961
rect 41024 16916 41255 16926
tri 41255 16916 41300 16961 sw
rect 70802 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41024 16871 41069 16916 ne
rect 41069 16871 41300 16916
tri 41300 16871 41345 16916 sw
tri 41069 16858 41082 16871 ne
rect 41082 16860 41345 16871
tri 41345 16860 41356 16871 sw
rect 70802 16868 71000 16926
rect 41082 16858 41356 16860
tri 41082 16857 41083 16858 ne
rect 41083 16857 41356 16858
tri 41083 16856 41084 16857 ne
rect 41084 16856 41356 16857
tri 41084 16855 41085 16856 ne
rect 41085 16855 41356 16856
tri 41085 16854 41086 16855 ne
rect 41086 16854 41356 16855
tri 41086 16853 41087 16854 ne
rect 41087 16853 41356 16854
tri 41087 16852 41088 16853 ne
rect 41088 16852 41356 16853
tri 41088 16851 41089 16852 ne
rect 41089 16851 41356 16852
tri 41089 16850 41090 16851 ne
rect 41090 16850 41356 16851
tri 41090 16849 41091 16850 ne
rect 41091 16849 41356 16850
tri 41091 16848 41092 16849 ne
rect 41092 16848 41356 16849
tri 41092 16847 41093 16848 ne
rect 41093 16847 41356 16848
tri 41093 16846 41094 16847 ne
rect 41094 16846 41356 16847
tri 41094 16845 41095 16846 ne
rect 41095 16845 41356 16846
tri 41095 16844 41096 16845 ne
rect 41096 16844 41356 16845
tri 41096 16843 41097 16844 ne
rect 41097 16843 41356 16844
tri 41097 16842 41098 16843 ne
rect 41098 16842 41356 16843
tri 41098 16841 41099 16842 ne
rect 41099 16841 41356 16842
tri 41099 16840 41100 16841 ne
rect 41100 16840 41356 16841
tri 41100 16839 41101 16840 ne
rect 41101 16839 41238 16840
tri 41101 16838 41102 16839 ne
rect 41102 16838 41238 16839
tri 41102 16837 41103 16838 ne
rect 41103 16837 41238 16838
tri 41103 16836 41104 16837 ne
rect 41104 16836 41238 16837
tri 41104 16835 41105 16836 ne
rect 41105 16835 41238 16836
tri 41105 16834 41106 16835 ne
rect 41106 16834 41238 16835
tri 41106 16833 41107 16834 ne
rect 41107 16833 41238 16834
tri 41107 16832 41108 16833 ne
rect 41108 16832 41238 16833
tri 41108 16831 41109 16832 ne
rect 41109 16831 41238 16832
tri 41109 16830 41110 16831 ne
rect 41110 16830 41238 16831
tri 41110 16829 41111 16830 ne
rect 41111 16829 41238 16830
tri 41111 16828 41112 16829 ne
rect 41112 16828 41238 16829
tri 41112 16827 41113 16828 ne
rect 41113 16827 41238 16828
tri 41113 16826 41114 16827 ne
rect 41114 16826 41238 16827
tri 41114 16825 41115 16826 ne
rect 41115 16825 41238 16826
tri 41115 16824 41116 16825 ne
rect 41116 16824 41238 16825
tri 41116 16823 41117 16824 ne
rect 41117 16823 41238 16824
tri 41117 16822 41118 16823 ne
rect 41118 16822 41238 16823
tri 41118 16821 41119 16822 ne
rect 41119 16821 41238 16822
tri 41119 16820 41120 16821 ne
rect 41120 16820 41238 16821
tri 41120 16819 41121 16820 ne
rect 41121 16819 41238 16820
tri 41121 16818 41122 16819 ne
rect 41122 16818 41238 16819
tri 41122 16817 41123 16818 ne
rect 41123 16817 41238 16818
tri 41123 16816 41124 16817 ne
rect 41124 16816 41238 16817
tri 41124 16815 41125 16816 ne
rect 41125 16815 41238 16816
tri 41125 16814 41126 16815 ne
rect 41126 16814 41238 16815
tri 41126 16813 41127 16814 ne
rect 41127 16813 41238 16814
tri 41127 16812 41128 16813 ne
rect 41128 16812 41238 16813
tri 41128 16811 41129 16812 ne
rect 41129 16811 41238 16812
tri 41129 16810 41130 16811 ne
rect 41130 16810 41238 16811
tri 41130 16809 41131 16810 ne
rect 41131 16809 41238 16810
tri 41131 16808 41132 16809 ne
rect 41132 16808 41238 16809
tri 41132 16807 41133 16808 ne
rect 41133 16807 41238 16808
tri 41133 16806 41134 16807 ne
rect 41134 16806 41238 16807
tri 41134 16805 41135 16806 ne
rect 41135 16805 41238 16806
tri 41135 16804 41136 16805 ne
rect 41136 16804 41238 16805
tri 41136 16803 41137 16804 ne
rect 41137 16803 41238 16804
tri 41137 16802 41138 16803 ne
rect 41138 16802 41238 16803
tri 41138 16801 41139 16802 ne
rect 41139 16801 41238 16802
tri 41139 16800 41140 16801 ne
rect 41140 16800 41238 16801
tri 41140 16799 41141 16800 ne
rect 41141 16799 41238 16800
tri 41141 16798 41142 16799 ne
rect 41142 16798 41238 16799
tri 41142 16797 41143 16798 ne
rect 41143 16797 41238 16798
tri 41143 16796 41144 16797 ne
rect 41144 16796 41238 16797
tri 41144 16795 41145 16796 ne
rect 41145 16795 41238 16796
tri 41145 16794 41146 16795 ne
rect 41146 16794 41238 16795
rect 41284 16815 41356 16840
tri 41356 16815 41401 16860 sw
rect 70802 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16794 41401 16815
tri 41146 16793 41147 16794 ne
rect 41147 16793 41401 16794
tri 41147 16792 41148 16793 ne
rect 41148 16792 41401 16793
tri 41148 16791 41149 16792 ne
rect 41149 16791 41401 16792
tri 41149 16790 41150 16791 ne
rect 41150 16790 41401 16791
tri 41150 16789 41151 16790 ne
rect 41151 16789 41401 16790
tri 41151 16788 41152 16789 ne
rect 41152 16788 41401 16789
tri 41152 16787 41153 16788 ne
rect 41153 16787 41401 16788
tri 41153 16786 41154 16787 ne
rect 41154 16786 41401 16787
tri 41154 16785 41155 16786 ne
rect 41155 16785 41401 16786
tri 41155 16784 41156 16785 ne
rect 41156 16784 41401 16785
tri 41156 16783 41157 16784 ne
rect 41157 16783 41401 16784
tri 41157 16782 41158 16783 ne
rect 41158 16782 41401 16783
tri 41158 16781 41159 16782 ne
rect 41159 16781 41401 16782
tri 41159 16780 41160 16781 ne
rect 41160 16780 41401 16781
tri 41160 16779 41161 16780 ne
rect 41161 16779 41401 16780
tri 41161 16778 41162 16779 ne
rect 41162 16778 41401 16779
tri 41162 16777 41163 16778 ne
rect 41163 16777 41401 16778
tri 41163 16776 41164 16777 ne
rect 41164 16776 41401 16777
tri 41164 16775 41165 16776 ne
rect 41165 16775 41401 16776
tri 41165 16774 41166 16775 ne
rect 41166 16774 41401 16775
tri 41166 16773 41167 16774 ne
rect 41167 16773 41401 16774
tri 41167 16772 41168 16773 ne
rect 41168 16772 41401 16773
tri 41168 16771 41169 16772 ne
rect 41169 16771 41401 16772
tri 41169 16770 41170 16771 ne
rect 41170 16770 41401 16771
tri 41401 16770 41446 16815 sw
tri 41170 16769 41171 16770 ne
rect 41171 16769 41446 16770
tri 41171 16768 41172 16769 ne
rect 41172 16768 41446 16769
tri 41172 16767 41173 16768 ne
rect 41173 16767 41446 16768
tri 41173 16766 41174 16767 ne
rect 41174 16766 41446 16767
tri 41174 16765 41175 16766 ne
rect 41175 16765 41446 16766
tri 41175 16764 41176 16765 ne
rect 41176 16764 41446 16765
tri 41176 16763 41177 16764 ne
rect 41177 16763 41446 16764
tri 41177 16762 41178 16763 ne
rect 41178 16762 41446 16763
tri 41178 16761 41179 16762 ne
rect 41179 16761 41446 16762
tri 41179 16760 41180 16761 ne
rect 41180 16760 41446 16761
tri 41180 16759 41181 16760 ne
rect 41181 16759 41446 16760
tri 41181 16758 41182 16759 ne
rect 41182 16758 41446 16759
tri 41182 16757 41183 16758 ne
rect 41183 16757 41446 16758
tri 41183 16756 41184 16757 ne
rect 41184 16756 41446 16757
tri 41184 16755 41185 16756 ne
rect 41185 16755 41446 16756
tri 41185 16754 41186 16755 ne
rect 41186 16754 41446 16755
tri 41186 16753 41187 16754 ne
rect 41187 16753 41446 16754
tri 41187 16752 41188 16753 ne
rect 41188 16752 41446 16753
tri 41188 16751 41189 16752 ne
rect 41189 16751 41446 16752
tri 41189 16750 41190 16751 ne
rect 41190 16750 41446 16751
tri 41190 16749 41191 16750 ne
rect 41191 16749 41446 16750
tri 41191 16748 41192 16749 ne
rect 41192 16748 41446 16749
tri 41192 16747 41193 16748 ne
rect 41193 16747 41446 16748
tri 41193 16746 41194 16747 ne
rect 41194 16746 41446 16747
tri 41194 16745 41195 16746 ne
rect 41195 16745 41446 16746
tri 41195 16744 41196 16745 ne
rect 41196 16744 41446 16745
tri 41196 16743 41197 16744 ne
rect 41197 16743 41446 16744
tri 41197 16742 41198 16743 ne
rect 41198 16742 41446 16743
tri 41198 16741 41199 16742 ne
rect 41199 16741 41446 16742
tri 41199 16740 41200 16741 ne
rect 41200 16740 41446 16741
tri 41200 16739 41201 16740 ne
rect 41201 16739 41446 16740
tri 41201 16738 41202 16739 ne
rect 41202 16738 41446 16739
tri 41202 16737 41203 16738 ne
rect 41203 16737 41446 16738
tri 41203 16736 41204 16737 ne
rect 41204 16736 41446 16737
tri 41204 16735 41205 16736 ne
rect 41205 16735 41446 16736
tri 41205 16734 41206 16735 ne
rect 41206 16734 41446 16735
tri 41206 16733 41207 16734 ne
rect 41207 16733 41446 16734
tri 41207 16732 41208 16733 ne
rect 41208 16732 41446 16733
tri 41208 16731 41209 16732 ne
rect 41209 16731 41446 16732
tri 41209 16730 41210 16731 ne
rect 41210 16730 41446 16731
tri 41210 16729 41211 16730 ne
rect 41211 16729 41446 16730
tri 41211 16728 41212 16729 ne
rect 41212 16728 41446 16729
tri 41212 16727 41213 16728 ne
rect 41213 16727 41446 16728
tri 41213 16726 41214 16727 ne
rect 41214 16726 41446 16727
tri 41214 16725 41215 16726 ne
rect 41215 16725 41446 16726
tri 41446 16725 41491 16770 sw
rect 70802 16764 71000 16822
tri 41215 16724 41216 16725 ne
rect 41216 16724 41491 16725
tri 41216 16723 41217 16724 ne
rect 41217 16723 41491 16724
tri 41217 16722 41218 16723 ne
rect 41218 16722 41491 16723
tri 41218 16721 41219 16722 ne
rect 41219 16721 41491 16722
tri 41219 16720 41220 16721 ne
rect 41220 16720 41491 16721
tri 41220 16719 41221 16720 ne
rect 41221 16719 41491 16720
tri 41221 16718 41222 16719 ne
rect 41222 16718 41491 16719
tri 41222 16717 41223 16718 ne
rect 41223 16717 41491 16718
tri 41223 16716 41224 16717 ne
rect 41224 16716 41491 16717
tri 41224 16715 41225 16716 ne
rect 41225 16715 41491 16716
tri 41225 16714 41226 16715 ne
rect 41226 16714 41491 16715
tri 41226 16713 41227 16714 ne
rect 41227 16713 41491 16714
tri 41227 16712 41228 16713 ne
rect 41228 16712 41491 16713
tri 41228 16711 41229 16712 ne
rect 41229 16711 41491 16712
tri 41229 16710 41230 16711 ne
rect 41230 16710 41491 16711
tri 41230 16709 41231 16710 ne
rect 41231 16709 41491 16710
tri 41231 16708 41232 16709 ne
rect 41232 16708 41491 16709
tri 41232 16707 41233 16708 ne
rect 41233 16707 41370 16708
tri 41233 16706 41234 16707 ne
rect 41234 16706 41370 16707
tri 41234 16705 41235 16706 ne
rect 41235 16705 41370 16706
tri 41235 16704 41236 16705 ne
rect 41236 16704 41370 16705
tri 41236 16703 41237 16704 ne
rect 41237 16703 41370 16704
tri 41237 16702 41238 16703 ne
rect 41238 16702 41370 16703
tri 41238 16701 41239 16702 ne
rect 41239 16701 41370 16702
tri 41239 16700 41240 16701 ne
rect 41240 16700 41370 16701
tri 41240 16699 41241 16700 ne
rect 41241 16699 41370 16700
tri 41241 16698 41242 16699 ne
rect 41242 16698 41370 16699
tri 41242 16697 41243 16698 ne
rect 41243 16697 41370 16698
tri 41243 16696 41244 16697 ne
rect 41244 16696 41370 16697
tri 41244 16695 41245 16696 ne
rect 41245 16695 41370 16696
tri 41245 16694 41246 16695 ne
rect 41246 16694 41370 16695
tri 41246 16693 41247 16694 ne
rect 41247 16693 41370 16694
tri 41247 16692 41248 16693 ne
rect 41248 16692 41370 16693
tri 41248 16691 41249 16692 ne
rect 41249 16691 41370 16692
tri 41249 16690 41250 16691 ne
rect 41250 16690 41370 16691
tri 41250 16689 41251 16690 ne
rect 41251 16689 41370 16690
tri 41251 16688 41252 16689 ne
rect 41252 16688 41370 16689
tri 41252 16687 41253 16688 ne
rect 41253 16687 41370 16688
tri 41253 16686 41254 16687 ne
rect 41254 16686 41370 16687
tri 41254 16685 41255 16686 ne
rect 41255 16685 41370 16686
tri 41255 16651 41289 16685 ne
rect 41289 16662 41370 16685
rect 41416 16685 41491 16708
tri 41491 16685 41531 16725 sw
rect 70802 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 41416 16680 41531 16685
tri 41531 16680 41536 16685 sw
rect 41416 16662 41536 16680
rect 41289 16651 41536 16662
tri 41289 16606 41334 16651 ne
rect 41334 16635 41536 16651
tri 41536 16635 41581 16680 sw
rect 70802 16660 71000 16718
rect 41334 16606 41581 16635
tri 41334 16584 41356 16606 ne
rect 41356 16590 41581 16606
tri 41581 16590 41626 16635 sw
rect 70802 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41356 16584 41626 16590
tri 41356 16583 41357 16584 ne
rect 41357 16583 41626 16584
tri 41357 16582 41358 16583 ne
rect 41358 16582 41626 16583
tri 41358 16581 41359 16582 ne
rect 41359 16581 41626 16582
tri 41359 16580 41360 16581 ne
rect 41360 16580 41626 16581
tri 41360 16579 41361 16580 ne
rect 41361 16579 41626 16580
tri 41361 16578 41362 16579 ne
rect 41362 16578 41626 16579
tri 41362 16577 41363 16578 ne
rect 41363 16577 41626 16578
tri 41363 16576 41364 16577 ne
rect 41364 16576 41626 16577
tri 41364 16575 41365 16576 ne
rect 41365 16575 41502 16576
tri 41365 16574 41366 16575 ne
rect 41366 16574 41502 16575
tri 41366 16573 41367 16574 ne
rect 41367 16573 41502 16574
tri 41367 16572 41368 16573 ne
rect 41368 16572 41502 16573
tri 41368 16571 41369 16572 ne
rect 41369 16571 41502 16572
tri 41369 16570 41370 16571 ne
rect 41370 16570 41502 16571
tri 41370 16569 41371 16570 ne
rect 41371 16569 41502 16570
tri 41371 16568 41372 16569 ne
rect 41372 16568 41502 16569
tri 41372 16567 41373 16568 ne
rect 41373 16567 41502 16568
tri 41373 16566 41374 16567 ne
rect 41374 16566 41502 16567
tri 41374 16565 41375 16566 ne
rect 41375 16565 41502 16566
tri 41375 16564 41376 16565 ne
rect 41376 16564 41502 16565
tri 41376 16563 41377 16564 ne
rect 41377 16563 41502 16564
tri 41377 16562 41378 16563 ne
rect 41378 16562 41502 16563
tri 41378 16561 41379 16562 ne
rect 41379 16561 41502 16562
tri 41379 16560 41380 16561 ne
rect 41380 16560 41502 16561
tri 41380 16559 41381 16560 ne
rect 41381 16559 41502 16560
tri 41381 16558 41382 16559 ne
rect 41382 16558 41502 16559
tri 41382 16557 41383 16558 ne
rect 41383 16557 41502 16558
tri 41383 16556 41384 16557 ne
rect 41384 16556 41502 16557
tri 41384 16555 41385 16556 ne
rect 41385 16555 41502 16556
tri 41385 16554 41386 16555 ne
rect 41386 16554 41502 16555
tri 41386 16553 41387 16554 ne
rect 41387 16553 41502 16554
tri 41387 16552 41388 16553 ne
rect 41388 16552 41502 16553
tri 41388 16551 41389 16552 ne
rect 41389 16551 41502 16552
tri 41389 16550 41390 16551 ne
rect 41390 16550 41502 16551
tri 41390 16549 41391 16550 ne
rect 41391 16549 41502 16550
tri 41391 16548 41392 16549 ne
rect 41392 16548 41502 16549
tri 41392 16547 41393 16548 ne
rect 41393 16547 41502 16548
tri 41393 16546 41394 16547 ne
rect 41394 16546 41502 16547
tri 41394 16545 41395 16546 ne
rect 41395 16545 41502 16546
tri 41395 16544 41396 16545 ne
rect 41396 16544 41502 16545
tri 41396 16543 41397 16544 ne
rect 41397 16543 41502 16544
tri 41397 16542 41398 16543 ne
rect 41398 16542 41502 16543
tri 41398 16541 41399 16542 ne
rect 41399 16541 41502 16542
tri 41399 16540 41400 16541 ne
rect 41400 16540 41502 16541
tri 41400 16539 41401 16540 ne
rect 41401 16539 41502 16540
tri 41401 16538 41402 16539 ne
rect 41402 16538 41502 16539
tri 41402 16537 41403 16538 ne
rect 41403 16537 41502 16538
tri 41403 16536 41404 16537 ne
rect 41404 16536 41502 16537
tri 41404 16535 41405 16536 ne
rect 41405 16535 41502 16536
tri 41405 16534 41406 16535 ne
rect 41406 16534 41502 16535
tri 41406 16533 41407 16534 ne
rect 41407 16533 41502 16534
tri 41407 16532 41408 16533 ne
rect 41408 16532 41502 16533
tri 41408 16531 41409 16532 ne
rect 41409 16531 41502 16532
tri 41409 16530 41410 16531 ne
rect 41410 16530 41502 16531
rect 41548 16545 41626 16576
tri 41626 16545 41671 16590 sw
rect 70802 16556 71000 16614
rect 41548 16544 41671 16545
tri 41671 16544 41672 16545 sw
rect 41548 16530 41672 16544
tri 41410 16529 41411 16530 ne
rect 41411 16529 41672 16530
tri 41411 16528 41412 16529 ne
rect 41412 16528 41672 16529
tri 41412 16527 41413 16528 ne
rect 41413 16527 41672 16528
tri 41413 16526 41414 16527 ne
rect 41414 16526 41672 16527
tri 41414 16525 41415 16526 ne
rect 41415 16525 41672 16526
tri 41415 16524 41416 16525 ne
rect 41416 16524 41672 16525
tri 41416 16523 41417 16524 ne
rect 41417 16523 41672 16524
tri 41417 16522 41418 16523 ne
rect 41418 16522 41672 16523
tri 41418 16521 41419 16522 ne
rect 41419 16521 41672 16522
tri 41419 16520 41420 16521 ne
rect 41420 16520 41672 16521
tri 41420 16519 41421 16520 ne
rect 41421 16519 41672 16520
tri 41421 16518 41422 16519 ne
rect 41422 16518 41672 16519
tri 41422 16517 41423 16518 ne
rect 41423 16517 41672 16518
tri 41423 16516 41424 16517 ne
rect 41424 16516 41672 16517
tri 41424 16515 41425 16516 ne
rect 41425 16515 41672 16516
tri 41425 16514 41426 16515 ne
rect 41426 16514 41672 16515
tri 41426 16513 41427 16514 ne
rect 41427 16513 41672 16514
tri 41427 16512 41428 16513 ne
rect 41428 16512 41672 16513
tri 41428 16511 41429 16512 ne
rect 41429 16511 41672 16512
tri 41429 16510 41430 16511 ne
rect 41430 16510 41672 16511
tri 41430 16509 41431 16510 ne
rect 41431 16509 41672 16510
tri 41431 16508 41432 16509 ne
rect 41432 16508 41672 16509
tri 41432 16507 41433 16508 ne
rect 41433 16507 41672 16508
tri 41433 16506 41434 16507 ne
rect 41434 16506 41672 16507
tri 41434 16505 41435 16506 ne
rect 41435 16505 41672 16506
tri 41435 16504 41436 16505 ne
rect 41436 16504 41672 16505
tri 41436 16503 41437 16504 ne
rect 41437 16503 41672 16504
tri 41437 16502 41438 16503 ne
rect 41438 16502 41672 16503
tri 41438 16501 41439 16502 ne
rect 41439 16501 41672 16502
tri 41439 16500 41440 16501 ne
rect 41440 16500 41672 16501
tri 41440 16499 41441 16500 ne
rect 41441 16499 41672 16500
tri 41672 16499 41717 16544 sw
rect 70802 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41441 16498 41442 16499 ne
rect 41442 16498 41717 16499
tri 41442 16497 41443 16498 ne
rect 41443 16497 41717 16498
tri 41443 16496 41444 16497 ne
rect 41444 16496 41717 16497
tri 41444 16495 41445 16496 ne
rect 41445 16495 41717 16496
tri 41445 16494 41446 16495 ne
rect 41446 16494 41717 16495
tri 41446 16493 41447 16494 ne
rect 41447 16493 41717 16494
tri 41447 16492 41448 16493 ne
rect 41448 16492 41717 16493
tri 41448 16491 41449 16492 ne
rect 41449 16491 41717 16492
tri 41449 16490 41450 16491 ne
rect 41450 16490 41717 16491
tri 41450 16489 41451 16490 ne
rect 41451 16489 41717 16490
tri 41451 16488 41452 16489 ne
rect 41452 16488 41717 16489
tri 41452 16487 41453 16488 ne
rect 41453 16487 41717 16488
tri 41453 16486 41454 16487 ne
rect 41454 16486 41717 16487
tri 41454 16485 41455 16486 ne
rect 41455 16485 41717 16486
tri 41455 16484 41456 16485 ne
rect 41456 16484 41717 16485
tri 41456 16483 41457 16484 ne
rect 41457 16483 41717 16484
tri 41457 16482 41458 16483 ne
rect 41458 16482 41717 16483
tri 41458 16481 41459 16482 ne
rect 41459 16481 41717 16482
tri 41459 16480 41460 16481 ne
rect 41460 16480 41717 16481
tri 41460 16479 41461 16480 ne
rect 41461 16479 41717 16480
tri 41461 16478 41462 16479 ne
rect 41462 16478 41717 16479
tri 41462 16477 41463 16478 ne
rect 41463 16477 41717 16478
tri 41463 16476 41464 16477 ne
rect 41464 16476 41717 16477
tri 41464 16475 41465 16476 ne
rect 41465 16475 41717 16476
tri 41465 16474 41466 16475 ne
rect 41466 16474 41717 16475
tri 41466 16473 41467 16474 ne
rect 41467 16473 41717 16474
tri 41467 16472 41468 16473 ne
rect 41468 16472 41717 16473
tri 41468 16471 41469 16472 ne
rect 41469 16471 41717 16472
tri 41469 16470 41470 16471 ne
rect 41470 16470 41717 16471
tri 41470 16469 41471 16470 ne
rect 41471 16469 41717 16470
tri 41471 16468 41472 16469 ne
rect 41472 16468 41717 16469
tri 41472 16467 41473 16468 ne
rect 41473 16467 41717 16468
tri 41473 16466 41474 16467 ne
rect 41474 16466 41717 16467
tri 41474 16465 41475 16466 ne
rect 41475 16465 41717 16466
tri 41475 16464 41476 16465 ne
rect 41476 16464 41717 16465
tri 41476 16463 41477 16464 ne
rect 41477 16463 41717 16464
tri 41477 16462 41478 16463 ne
rect 41478 16462 41717 16463
tri 41478 16461 41479 16462 ne
rect 41479 16461 41717 16462
tri 41479 16460 41480 16461 ne
rect 41480 16460 41717 16461
tri 41480 16459 41481 16460 ne
rect 41481 16459 41717 16460
tri 41481 16458 41482 16459 ne
rect 41482 16458 41717 16459
tri 41482 16457 41483 16458 ne
rect 41483 16457 41717 16458
tri 41483 16456 41484 16457 ne
rect 41484 16456 41717 16457
tri 41484 16455 41485 16456 ne
rect 41485 16455 41717 16456
tri 41485 16454 41486 16455 ne
rect 41486 16454 41717 16455
tri 41717 16454 41762 16499 sw
tri 41486 16453 41487 16454 ne
rect 41487 16453 41762 16454
tri 41487 16452 41488 16453 ne
rect 41488 16452 41762 16453
tri 41488 16451 41489 16452 ne
rect 41489 16451 41762 16452
tri 41489 16450 41490 16451 ne
rect 41490 16450 41762 16451
tri 41490 16449 41491 16450 ne
rect 41491 16449 41762 16450
tri 41491 16448 41492 16449 ne
rect 41492 16448 41762 16449
tri 41492 16447 41493 16448 ne
rect 41493 16447 41762 16448
tri 41493 16446 41494 16447 ne
rect 41494 16446 41762 16447
tri 41494 16445 41495 16446 ne
rect 41495 16445 41762 16446
tri 41495 16444 41496 16445 ne
rect 41496 16444 41762 16445
tri 41496 16443 41497 16444 ne
rect 41497 16443 41634 16444
tri 41497 16442 41498 16443 ne
rect 41498 16442 41634 16443
tri 41498 16441 41499 16442 ne
rect 41499 16441 41634 16442
tri 41499 16440 41500 16441 ne
rect 41500 16440 41634 16441
tri 41500 16439 41501 16440 ne
rect 41501 16439 41634 16440
tri 41501 16438 41502 16439 ne
rect 41502 16438 41634 16439
tri 41502 16437 41503 16438 ne
rect 41503 16437 41634 16438
tri 41503 16436 41504 16437 ne
rect 41504 16436 41634 16437
tri 41504 16435 41505 16436 ne
rect 41505 16435 41634 16436
tri 41505 16434 41506 16435 ne
rect 41506 16434 41634 16435
tri 41506 16433 41507 16434 ne
rect 41507 16433 41634 16434
tri 41507 16432 41508 16433 ne
rect 41508 16432 41634 16433
tri 41508 16431 41509 16432 ne
rect 41509 16431 41634 16432
tri 41509 16430 41510 16431 ne
rect 41510 16430 41634 16431
tri 41510 16429 41511 16430 ne
rect 41511 16429 41634 16430
tri 41511 16428 41512 16429 ne
rect 41512 16428 41634 16429
tri 41512 16427 41513 16428 ne
rect 41513 16427 41634 16428
tri 41513 16426 41514 16427 ne
rect 41514 16426 41634 16427
tri 41514 16425 41515 16426 ne
rect 41515 16425 41634 16426
tri 41515 16424 41516 16425 ne
rect 41516 16424 41634 16425
tri 41516 16423 41517 16424 ne
rect 41517 16423 41634 16424
tri 41517 16422 41518 16423 ne
rect 41518 16422 41634 16423
tri 41518 16421 41519 16422 ne
rect 41519 16421 41634 16422
tri 41519 16420 41520 16421 ne
rect 41520 16420 41634 16421
tri 41520 16419 41521 16420 ne
rect 41521 16419 41634 16420
tri 41521 16418 41522 16419 ne
rect 41522 16418 41634 16419
tri 41522 16417 41523 16418 ne
rect 41523 16417 41634 16418
tri 41523 16416 41524 16417 ne
rect 41524 16416 41634 16417
tri 41524 16415 41525 16416 ne
rect 41525 16415 41634 16416
tri 41525 16414 41526 16415 ne
rect 41526 16414 41634 16415
tri 41526 16413 41527 16414 ne
rect 41527 16413 41634 16414
tri 41527 16412 41528 16413 ne
rect 41528 16412 41634 16413
tri 41528 16411 41529 16412 ne
rect 41529 16411 41634 16412
tri 41529 16410 41530 16411 ne
rect 41530 16410 41634 16411
tri 41530 16409 41531 16410 ne
rect 41531 16409 41634 16410
tri 41531 16404 41536 16409 ne
rect 41536 16404 41634 16409
tri 41536 16364 41576 16404 ne
rect 41576 16398 41634 16404
rect 41680 16409 41762 16444
tri 41762 16409 41807 16454 sw
rect 70802 16452 71000 16510
rect 41680 16404 41807 16409
tri 41807 16404 41812 16409 sw
rect 70802 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 41680 16398 41812 16404
rect 41576 16364 41812 16398
tri 41576 16359 41581 16364 ne
rect 41581 16359 41812 16364
tri 41812 16359 41857 16404 sw
tri 41581 16314 41626 16359 ne
rect 41626 16314 41857 16359
tri 41857 16314 41902 16359 sw
rect 70802 16348 71000 16406
tri 41626 16309 41631 16314 ne
rect 41631 16312 41902 16314
rect 41631 16309 41766 16312
tri 41631 16308 41632 16309 ne
rect 41632 16308 41766 16309
tri 41632 16307 41633 16308 ne
rect 41633 16307 41766 16308
tri 41633 16306 41634 16307 ne
rect 41634 16306 41766 16307
tri 41634 16305 41635 16306 ne
rect 41635 16305 41766 16306
tri 41635 16304 41636 16305 ne
rect 41636 16304 41766 16305
tri 41636 16303 41637 16304 ne
rect 41637 16303 41766 16304
tri 41637 16302 41638 16303 ne
rect 41638 16302 41766 16303
tri 41638 16301 41639 16302 ne
rect 41639 16301 41766 16302
tri 41639 16300 41640 16301 ne
rect 41640 16300 41766 16301
tri 41640 16299 41641 16300 ne
rect 41641 16299 41766 16300
tri 41641 16298 41642 16299 ne
rect 41642 16298 41766 16299
tri 41642 16297 41643 16298 ne
rect 41643 16297 41766 16298
tri 41643 16296 41644 16297 ne
rect 41644 16296 41766 16297
tri 41644 16295 41645 16296 ne
rect 41645 16295 41766 16296
tri 41645 16294 41646 16295 ne
rect 41646 16294 41766 16295
tri 41646 16293 41647 16294 ne
rect 41647 16293 41766 16294
tri 41647 16292 41648 16293 ne
rect 41648 16292 41766 16293
tri 41648 16291 41649 16292 ne
rect 41649 16291 41766 16292
tri 41649 16290 41650 16291 ne
rect 41650 16290 41766 16291
tri 41650 16289 41651 16290 ne
rect 41651 16289 41766 16290
tri 41651 16288 41652 16289 ne
rect 41652 16288 41766 16289
tri 41652 16287 41653 16288 ne
rect 41653 16287 41766 16288
tri 41653 16286 41654 16287 ne
rect 41654 16286 41766 16287
tri 41654 16285 41655 16286 ne
rect 41655 16285 41766 16286
tri 41655 16284 41656 16285 ne
rect 41656 16284 41766 16285
tri 41656 16283 41657 16284 ne
rect 41657 16283 41766 16284
tri 41657 16282 41658 16283 ne
rect 41658 16282 41766 16283
tri 41658 16281 41659 16282 ne
rect 41659 16281 41766 16282
tri 41659 16280 41660 16281 ne
rect 41660 16280 41766 16281
tri 41660 16279 41661 16280 ne
rect 41661 16279 41766 16280
tri 41661 16278 41662 16279 ne
rect 41662 16278 41766 16279
tri 41662 16277 41663 16278 ne
rect 41663 16277 41766 16278
tri 41663 16276 41664 16277 ne
rect 41664 16276 41766 16277
tri 41664 16275 41665 16276 ne
rect 41665 16275 41766 16276
tri 41665 16274 41666 16275 ne
rect 41666 16274 41766 16275
tri 41666 16273 41667 16274 ne
rect 41667 16273 41766 16274
tri 41667 16272 41668 16273 ne
rect 41668 16272 41766 16273
tri 41668 16271 41669 16272 ne
rect 41669 16271 41766 16272
tri 41669 16270 41670 16271 ne
rect 41670 16270 41766 16271
tri 41670 16269 41671 16270 ne
rect 41671 16269 41766 16270
tri 41671 16268 41672 16269 ne
rect 41672 16268 41766 16269
tri 41672 16267 41673 16268 ne
rect 41673 16267 41766 16268
tri 41673 16266 41674 16267 ne
rect 41674 16266 41766 16267
rect 41812 16269 41902 16312
tri 41902 16269 41947 16314 sw
rect 70802 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16266 41947 16269
tri 41674 16265 41675 16266 ne
rect 41675 16265 41947 16266
tri 41675 16264 41676 16265 ne
rect 41676 16264 41947 16265
tri 41676 16263 41677 16264 ne
rect 41677 16263 41947 16264
tri 41677 16262 41678 16263 ne
rect 41678 16262 41947 16263
tri 41678 16261 41679 16262 ne
rect 41679 16261 41947 16262
tri 41679 16260 41680 16261 ne
rect 41680 16260 41947 16261
tri 41680 16259 41681 16260 ne
rect 41681 16259 41947 16260
tri 41681 16258 41682 16259 ne
rect 41682 16258 41947 16259
tri 41682 16257 41683 16258 ne
rect 41683 16257 41947 16258
tri 41683 16256 41684 16257 ne
rect 41684 16256 41947 16257
tri 41684 16255 41685 16256 ne
rect 41685 16255 41947 16256
tri 41685 16254 41686 16255 ne
rect 41686 16254 41947 16255
tri 41686 16253 41687 16254 ne
rect 41687 16253 41947 16254
tri 41687 16252 41688 16253 ne
rect 41688 16252 41947 16253
tri 41688 16251 41689 16252 ne
rect 41689 16251 41947 16252
tri 41689 16250 41690 16251 ne
rect 41690 16250 41947 16251
tri 41690 16249 41691 16250 ne
rect 41691 16249 41947 16250
tri 41691 16248 41692 16249 ne
rect 41692 16248 41947 16249
tri 41692 16247 41693 16248 ne
rect 41693 16247 41947 16248
tri 41693 16246 41694 16247 ne
rect 41694 16246 41947 16247
tri 41694 16245 41695 16246 ne
rect 41695 16245 41947 16246
tri 41695 16244 41696 16245 ne
rect 41696 16244 41947 16245
tri 41696 16243 41697 16244 ne
rect 41697 16243 41947 16244
tri 41697 16242 41698 16243 ne
rect 41698 16242 41947 16243
tri 41698 16241 41699 16242 ne
rect 41699 16241 41947 16242
tri 41699 16240 41700 16241 ne
rect 41700 16240 41947 16241
tri 41700 16239 41701 16240 ne
rect 41701 16239 41947 16240
tri 41701 16238 41702 16239 ne
rect 41702 16238 41947 16239
tri 41702 16237 41703 16238 ne
rect 41703 16237 41947 16238
tri 41703 16236 41704 16237 ne
rect 41704 16236 41947 16237
tri 41704 16235 41705 16236 ne
rect 41705 16235 41947 16236
tri 41705 16234 41706 16235 ne
rect 41706 16234 41947 16235
tri 41706 16233 41707 16234 ne
rect 41707 16233 41947 16234
tri 41707 16232 41708 16233 ne
rect 41708 16232 41947 16233
tri 41708 16231 41709 16232 ne
rect 41709 16231 41947 16232
tri 41709 16230 41710 16231 ne
rect 41710 16230 41947 16231
tri 41710 16229 41711 16230 ne
rect 41711 16229 41947 16230
tri 41711 16228 41712 16229 ne
rect 41712 16228 41947 16229
tri 41712 16227 41713 16228 ne
rect 41713 16227 41947 16228
tri 41713 16226 41714 16227 ne
rect 41714 16226 41947 16227
tri 41714 16225 41715 16226 ne
rect 41715 16225 41947 16226
tri 41715 16224 41716 16225 ne
rect 41716 16224 41947 16225
tri 41947 16224 41992 16269 sw
rect 70802 16244 71000 16302
tri 41716 16223 41717 16224 ne
rect 41717 16223 41992 16224
tri 41992 16223 41993 16224 sw
tri 41717 16222 41718 16223 ne
rect 41718 16222 41993 16223
tri 41718 16221 41719 16222 ne
rect 41719 16221 41993 16222
tri 41719 16220 41720 16221 ne
rect 41720 16220 41993 16221
tri 41720 16219 41721 16220 ne
rect 41721 16219 41993 16220
tri 41721 16218 41722 16219 ne
rect 41722 16218 41993 16219
tri 41722 16217 41723 16218 ne
rect 41723 16217 41993 16218
tri 41723 16216 41724 16217 ne
rect 41724 16216 41993 16217
tri 41724 16215 41725 16216 ne
rect 41725 16215 41993 16216
tri 41725 16214 41726 16215 ne
rect 41726 16214 41993 16215
tri 41726 16213 41727 16214 ne
rect 41727 16213 41993 16214
tri 41727 16212 41728 16213 ne
rect 41728 16212 41993 16213
tri 41728 16211 41729 16212 ne
rect 41729 16211 41993 16212
tri 41729 16210 41730 16211 ne
rect 41730 16210 41993 16211
tri 41730 16209 41731 16210 ne
rect 41731 16209 41993 16210
tri 41731 16208 41732 16209 ne
rect 41732 16208 41993 16209
tri 41732 16207 41733 16208 ne
rect 41733 16207 41993 16208
tri 41733 16206 41734 16207 ne
rect 41734 16206 41993 16207
tri 41734 16205 41735 16206 ne
rect 41735 16205 41993 16206
tri 41735 16204 41736 16205 ne
rect 41736 16204 41993 16205
tri 41736 16203 41737 16204 ne
rect 41737 16203 41993 16204
tri 41737 16202 41738 16203 ne
rect 41738 16202 41993 16203
tri 41738 16201 41739 16202 ne
rect 41739 16201 41993 16202
tri 41739 16200 41740 16201 ne
rect 41740 16200 41993 16201
tri 41740 16199 41741 16200 ne
rect 41741 16199 41993 16200
tri 41741 16198 41742 16199 ne
rect 41742 16198 41993 16199
tri 41742 16197 41743 16198 ne
rect 41743 16197 41993 16198
tri 41743 16196 41744 16197 ne
rect 41744 16196 41993 16197
tri 41744 16195 41745 16196 ne
rect 41745 16195 41993 16196
tri 41745 16194 41746 16195 ne
rect 41746 16194 41993 16195
tri 41746 16193 41747 16194 ne
rect 41747 16193 41993 16194
tri 41747 16192 41748 16193 ne
rect 41748 16192 41993 16193
tri 41748 16191 41749 16192 ne
rect 41749 16191 41993 16192
tri 41749 16190 41750 16191 ne
rect 41750 16190 41993 16191
tri 41750 16189 41751 16190 ne
rect 41751 16189 41993 16190
tri 41751 16188 41752 16189 ne
rect 41752 16188 41993 16189
tri 41752 16187 41753 16188 ne
rect 41753 16187 41993 16188
tri 41753 16186 41754 16187 ne
rect 41754 16186 41993 16187
tri 41754 16185 41755 16186 ne
rect 41755 16185 41993 16186
tri 41755 16184 41756 16185 ne
rect 41756 16184 41993 16185
tri 41756 16183 41757 16184 ne
rect 41757 16183 41993 16184
tri 41757 16182 41758 16183 ne
rect 41758 16182 41993 16183
tri 41758 16181 41759 16182 ne
rect 41759 16181 41993 16182
tri 41759 16180 41760 16181 ne
rect 41760 16180 41993 16181
tri 41760 16179 41761 16180 ne
rect 41761 16179 41898 16180
tri 41761 16178 41762 16179 ne
rect 41762 16178 41898 16179
tri 41762 16177 41763 16178 ne
rect 41763 16177 41898 16178
tri 41763 16176 41764 16177 ne
rect 41764 16176 41898 16177
tri 41764 16175 41765 16176 ne
rect 41765 16175 41898 16176
tri 41765 16174 41766 16175 ne
rect 41766 16174 41898 16175
tri 41766 16173 41767 16174 ne
rect 41767 16173 41898 16174
tri 41767 16172 41768 16173 ne
rect 41768 16172 41898 16173
tri 41768 16171 41769 16172 ne
rect 41769 16171 41898 16172
tri 41769 16170 41770 16171 ne
rect 41770 16170 41898 16171
tri 41770 16169 41771 16170 ne
rect 41771 16169 41898 16170
tri 41771 16168 41772 16169 ne
rect 41772 16168 41898 16169
tri 41772 16167 41773 16168 ne
rect 41773 16167 41898 16168
tri 41773 16166 41774 16167 ne
rect 41774 16166 41898 16167
tri 41774 16165 41775 16166 ne
rect 41775 16165 41898 16166
tri 41775 16164 41776 16165 ne
rect 41776 16164 41898 16165
tri 41776 16163 41777 16164 ne
rect 41777 16163 41898 16164
tri 41777 16162 41778 16163 ne
rect 41778 16162 41898 16163
tri 41778 16161 41779 16162 ne
rect 41779 16161 41898 16162
tri 41779 16160 41780 16161 ne
rect 41780 16160 41898 16161
tri 41780 16159 41781 16160 ne
rect 41781 16159 41898 16160
tri 41781 16158 41782 16159 ne
rect 41782 16158 41898 16159
tri 41782 16157 41783 16158 ne
rect 41783 16157 41898 16158
tri 41783 16156 41784 16157 ne
rect 41784 16156 41898 16157
tri 41784 16155 41785 16156 ne
rect 41785 16155 41898 16156
tri 41785 16154 41786 16155 ne
rect 41786 16154 41898 16155
tri 41786 16153 41787 16154 ne
rect 41787 16153 41898 16154
tri 41787 16152 41788 16153 ne
rect 41788 16152 41898 16153
tri 41788 16151 41789 16152 ne
rect 41789 16151 41898 16152
tri 41789 16150 41790 16151 ne
rect 41790 16150 41898 16151
tri 41790 16149 41791 16150 ne
rect 41791 16149 41898 16150
tri 41791 16148 41792 16149 ne
rect 41792 16148 41898 16149
tri 41792 16147 41793 16148 ne
rect 41793 16147 41898 16148
tri 41793 16146 41794 16147 ne
rect 41794 16146 41898 16147
tri 41794 16145 41795 16146 ne
rect 41795 16145 41898 16146
tri 41795 16144 41796 16145 ne
rect 41796 16144 41898 16145
tri 41796 16143 41797 16144 ne
rect 41797 16143 41898 16144
tri 41797 16142 41798 16143 ne
rect 41798 16142 41898 16143
tri 41798 16141 41799 16142 ne
rect 41799 16141 41898 16142
tri 41799 16140 41800 16141 ne
rect 41800 16140 41898 16141
tri 41800 16139 41801 16140 ne
rect 41801 16139 41898 16140
tri 41801 16138 41802 16139 ne
rect 41802 16138 41898 16139
tri 41802 16137 41803 16138 ne
rect 41803 16137 41898 16138
tri 41803 16136 41804 16137 ne
rect 41804 16136 41898 16137
tri 41804 16135 41805 16136 ne
rect 41805 16135 41898 16136
tri 41805 16134 41806 16135 ne
rect 41806 16134 41898 16135
rect 41944 16178 41993 16180
tri 41993 16178 42038 16223 sw
rect 70802 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 41944 16134 42038 16178
tri 41806 16133 41807 16134 ne
rect 41807 16133 42038 16134
tri 42038 16133 42083 16178 sw
rect 70802 16140 71000 16198
tri 41807 16088 41852 16133 ne
rect 41852 16088 42083 16133
tri 42083 16088 42128 16133 sw
rect 70802 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41852 16043 41897 16088 ne
rect 41897 16083 42128 16088
tri 42128 16083 42133 16088 sw
rect 41897 16048 42133 16083
rect 41897 16043 42030 16048
tri 41897 16038 41902 16043 ne
rect 41902 16038 42030 16043
tri 41902 16035 41905 16038 ne
rect 41905 16035 42030 16038
tri 41905 16034 41906 16035 ne
rect 41906 16034 42030 16035
tri 41906 16033 41907 16034 ne
rect 41907 16033 42030 16034
tri 41907 16032 41908 16033 ne
rect 41908 16032 42030 16033
tri 41908 16031 41909 16032 ne
rect 41909 16031 42030 16032
tri 41909 16030 41910 16031 ne
rect 41910 16030 42030 16031
tri 41910 16029 41911 16030 ne
rect 41911 16029 42030 16030
tri 41911 16028 41912 16029 ne
rect 41912 16028 42030 16029
tri 41912 16027 41913 16028 ne
rect 41913 16027 42030 16028
tri 41913 16026 41914 16027 ne
rect 41914 16026 42030 16027
tri 41914 16025 41915 16026 ne
rect 41915 16025 42030 16026
tri 41915 16024 41916 16025 ne
rect 41916 16024 42030 16025
tri 41916 16023 41917 16024 ne
rect 41917 16023 42030 16024
tri 41917 16022 41918 16023 ne
rect 41918 16022 42030 16023
tri 41918 16021 41919 16022 ne
rect 41919 16021 42030 16022
tri 41919 16020 41920 16021 ne
rect 41920 16020 42030 16021
tri 41920 16019 41921 16020 ne
rect 41921 16019 42030 16020
tri 41921 16018 41922 16019 ne
rect 41922 16018 42030 16019
tri 41922 16017 41923 16018 ne
rect 41923 16017 42030 16018
tri 41923 16016 41924 16017 ne
rect 41924 16016 42030 16017
tri 41924 16015 41925 16016 ne
rect 41925 16015 42030 16016
tri 41925 16014 41926 16015 ne
rect 41926 16014 42030 16015
tri 41926 16013 41927 16014 ne
rect 41927 16013 42030 16014
tri 41927 16012 41928 16013 ne
rect 41928 16012 42030 16013
tri 41928 16011 41929 16012 ne
rect 41929 16011 42030 16012
tri 41929 16010 41930 16011 ne
rect 41930 16010 42030 16011
tri 41930 16009 41931 16010 ne
rect 41931 16009 42030 16010
tri 41931 16008 41932 16009 ne
rect 41932 16008 42030 16009
tri 41932 16007 41933 16008 ne
rect 41933 16007 42030 16008
tri 41933 16006 41934 16007 ne
rect 41934 16006 42030 16007
tri 41934 16005 41935 16006 ne
rect 41935 16005 42030 16006
tri 41935 16004 41936 16005 ne
rect 41936 16004 42030 16005
tri 41936 16003 41937 16004 ne
rect 41937 16003 42030 16004
tri 41937 16002 41938 16003 ne
rect 41938 16002 42030 16003
rect 42076 16038 42133 16048
tri 42133 16038 42178 16083 sw
rect 42076 16002 42178 16038
tri 41938 16001 41939 16002 ne
rect 41939 16001 42178 16002
tri 41939 16000 41940 16001 ne
rect 41940 16000 42178 16001
tri 41940 15999 41941 16000 ne
rect 41941 15999 42178 16000
tri 41941 15998 41942 15999 ne
rect 41942 15998 42178 15999
tri 41942 15997 41943 15998 ne
rect 41943 15997 42178 15998
tri 41943 15996 41944 15997 ne
rect 41944 15996 42178 15997
tri 41944 15995 41945 15996 ne
rect 41945 15995 42178 15996
tri 41945 15994 41946 15995 ne
rect 41946 15994 42178 15995
tri 41946 15993 41947 15994 ne
rect 41947 15993 42178 15994
tri 42178 15993 42223 16038 sw
rect 70802 16036 71000 16094
tri 41947 15992 41948 15993 ne
rect 41948 15992 42223 15993
tri 41948 15991 41949 15992 ne
rect 41949 15991 42223 15992
tri 41949 15990 41950 15991 ne
rect 41950 15990 42223 15991
tri 41950 15989 41951 15990 ne
rect 41951 15989 42223 15990
tri 41951 15988 41952 15989 ne
rect 41952 15988 42223 15989
tri 41952 15987 41953 15988 ne
rect 41953 15987 42223 15988
tri 41953 15986 41954 15987 ne
rect 41954 15986 42223 15987
tri 41954 15985 41955 15986 ne
rect 41955 15985 42223 15986
tri 41955 15984 41956 15985 ne
rect 41956 15984 42223 15985
tri 41956 15983 41957 15984 ne
rect 41957 15983 42223 15984
tri 41957 15982 41958 15983 ne
rect 41958 15982 42223 15983
tri 41958 15981 41959 15982 ne
rect 41959 15981 42223 15982
tri 41959 15980 41960 15981 ne
rect 41960 15980 42223 15981
tri 41960 15979 41961 15980 ne
rect 41961 15979 42223 15980
tri 41961 15978 41962 15979 ne
rect 41962 15978 42223 15979
tri 41962 15977 41963 15978 ne
rect 41963 15977 42223 15978
tri 41963 15976 41964 15977 ne
rect 41964 15976 42223 15977
tri 41964 15975 41965 15976 ne
rect 41965 15975 42223 15976
tri 41965 15974 41966 15975 ne
rect 41966 15974 42223 15975
tri 41966 15973 41967 15974 ne
rect 41967 15973 42223 15974
tri 41967 15972 41968 15973 ne
rect 41968 15972 42223 15973
tri 41968 15971 41969 15972 ne
rect 41969 15971 42223 15972
tri 41969 15970 41970 15971 ne
rect 41970 15970 42223 15971
tri 41970 15969 41971 15970 ne
rect 41971 15969 42223 15970
tri 41971 15968 41972 15969 ne
rect 41972 15968 42223 15969
tri 41972 15967 41973 15968 ne
rect 41973 15967 42223 15968
tri 41973 15966 41974 15967 ne
rect 41974 15966 42223 15967
tri 41974 15965 41975 15966 ne
rect 41975 15965 42223 15966
tri 41975 15964 41976 15965 ne
rect 41976 15964 42223 15965
tri 41976 15963 41977 15964 ne
rect 41977 15963 42223 15964
tri 41977 15962 41978 15963 ne
rect 41978 15962 42223 15963
tri 41978 15961 41979 15962 ne
rect 41979 15961 42223 15962
tri 41979 15960 41980 15961 ne
rect 41980 15960 42223 15961
tri 41980 15959 41981 15960 ne
rect 41981 15959 42223 15960
tri 41981 15958 41982 15959 ne
rect 41982 15958 42223 15959
tri 41982 15957 41983 15958 ne
rect 41983 15957 42223 15958
tri 41983 15956 41984 15957 ne
rect 41984 15956 42223 15957
tri 41984 15955 41985 15956 ne
rect 41985 15955 42223 15956
tri 41985 15954 41986 15955 ne
rect 41986 15954 42223 15955
tri 41986 15953 41987 15954 ne
rect 41987 15953 42223 15954
tri 41987 15952 41988 15953 ne
rect 41988 15952 42223 15953
tri 41988 15951 41989 15952 ne
rect 41989 15951 42223 15952
tri 41989 15950 41990 15951 ne
rect 41990 15950 42223 15951
tri 41990 15949 41991 15950 ne
rect 41991 15949 42223 15950
tri 41991 15948 41992 15949 ne
rect 41992 15948 42223 15949
tri 42223 15948 42268 15993 sw
rect 70802 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
tri 41992 15947 41993 15948 ne
rect 41993 15947 42268 15948
tri 41993 15946 41994 15947 ne
rect 41994 15946 42268 15947
tri 41994 15945 41995 15946 ne
rect 41995 15945 42268 15946
tri 41995 15944 41996 15945 ne
rect 41996 15944 42268 15945
tri 41996 15943 41997 15944 ne
rect 41997 15943 42268 15944
tri 41997 15942 41998 15943 ne
rect 41998 15942 42268 15943
tri 41998 15941 41999 15942 ne
rect 41999 15941 42268 15942
tri 41999 15940 42000 15941 ne
rect 42000 15940 42268 15941
tri 42000 15939 42001 15940 ne
rect 42001 15939 42268 15940
tri 42001 15938 42002 15939 ne
rect 42002 15938 42268 15939
tri 42002 15937 42003 15938 ne
rect 42003 15937 42268 15938
tri 42003 15936 42004 15937 ne
rect 42004 15936 42268 15937
tri 42004 15935 42005 15936 ne
rect 42005 15935 42268 15936
tri 42005 15934 42006 15935 ne
rect 42006 15934 42268 15935
tri 42006 15933 42007 15934 ne
rect 42007 15933 42268 15934
tri 42007 15932 42008 15933 ne
rect 42008 15932 42268 15933
tri 42008 15931 42009 15932 ne
rect 42009 15931 42268 15932
tri 42009 15930 42010 15931 ne
rect 42010 15930 42268 15931
tri 42010 15929 42011 15930 ne
rect 42011 15929 42268 15930
tri 42011 15928 42012 15929 ne
rect 42012 15928 42268 15929
tri 42012 15927 42013 15928 ne
rect 42013 15927 42268 15928
tri 42013 15926 42014 15927 ne
rect 42014 15926 42268 15927
tri 42014 15925 42015 15926 ne
rect 42015 15925 42268 15926
tri 42015 15924 42016 15925 ne
rect 42016 15924 42268 15925
tri 42016 15923 42017 15924 ne
rect 42017 15923 42268 15924
tri 42017 15922 42018 15923 ne
rect 42018 15922 42268 15923
tri 42018 15921 42019 15922 ne
rect 42019 15921 42268 15922
tri 42019 15920 42020 15921 ne
rect 42020 15920 42268 15921
tri 42020 15919 42021 15920 ne
rect 42021 15919 42268 15920
tri 42021 15918 42022 15919 ne
rect 42022 15918 42268 15919
tri 42022 15917 42023 15918 ne
rect 42023 15917 42268 15918
tri 42023 15916 42024 15917 ne
rect 42024 15916 42268 15917
tri 42024 15915 42025 15916 ne
rect 42025 15915 42162 15916
tri 42025 15914 42026 15915 ne
rect 42026 15914 42162 15915
tri 42026 15913 42027 15914 ne
rect 42027 15913 42162 15914
tri 42027 15912 42028 15913 ne
rect 42028 15912 42162 15913
tri 42028 15911 42029 15912 ne
rect 42029 15911 42162 15912
tri 42029 15910 42030 15911 ne
rect 42030 15910 42162 15911
tri 42030 15909 42031 15910 ne
rect 42031 15909 42162 15910
tri 42031 15908 42032 15909 ne
rect 42032 15908 42162 15909
tri 42032 15907 42033 15908 ne
rect 42033 15907 42162 15908
tri 42033 15906 42034 15907 ne
rect 42034 15906 42162 15907
tri 42034 15905 42035 15906 ne
rect 42035 15905 42162 15906
tri 42035 15904 42036 15905 ne
rect 42036 15904 42162 15905
tri 42036 15903 42037 15904 ne
rect 42037 15903 42162 15904
tri 42037 15902 42038 15903 ne
rect 42038 15902 42162 15903
tri 42038 15901 42039 15902 ne
rect 42039 15901 42162 15902
tri 42039 15900 42040 15901 ne
rect 42040 15900 42162 15901
tri 42040 15899 42041 15900 ne
rect 42041 15899 42162 15900
tri 42041 15898 42042 15899 ne
rect 42042 15898 42162 15899
tri 42042 15897 42043 15898 ne
rect 42043 15897 42162 15898
tri 42043 15896 42044 15897 ne
rect 42044 15896 42162 15897
tri 42044 15895 42045 15896 ne
rect 42045 15895 42162 15896
tri 42045 15894 42046 15895 ne
rect 42046 15894 42162 15895
tri 42046 15893 42047 15894 ne
rect 42047 15893 42162 15894
tri 42047 15892 42048 15893 ne
rect 42048 15892 42162 15893
tri 42048 15891 42049 15892 ne
rect 42049 15891 42162 15892
tri 42049 15890 42050 15891 ne
rect 42050 15890 42162 15891
tri 42050 15889 42051 15890 ne
rect 42051 15889 42162 15890
tri 42051 15888 42052 15889 ne
rect 42052 15888 42162 15889
tri 42052 15887 42053 15888 ne
rect 42053 15887 42162 15888
tri 42053 15886 42054 15887 ne
rect 42054 15886 42162 15887
tri 42054 15885 42055 15886 ne
rect 42055 15885 42162 15886
tri 42055 15884 42056 15885 ne
rect 42056 15884 42162 15885
tri 42056 15883 42057 15884 ne
rect 42057 15883 42162 15884
tri 42057 15882 42058 15883 ne
rect 42058 15882 42162 15883
tri 42058 15881 42059 15882 ne
rect 42059 15881 42162 15882
tri 42059 15880 42060 15881 ne
rect 42060 15880 42162 15881
tri 42060 15879 42061 15880 ne
rect 42061 15879 42162 15880
tri 42061 15878 42062 15879 ne
rect 42062 15878 42162 15879
tri 42062 15877 42063 15878 ne
rect 42063 15877 42162 15878
tri 42063 15876 42064 15877 ne
rect 42064 15876 42162 15877
tri 42064 15875 42065 15876 ne
rect 42065 15875 42162 15876
tri 42065 15874 42066 15875 ne
rect 42066 15874 42162 15875
tri 42066 15873 42067 15874 ne
rect 42067 15873 42162 15874
tri 42067 15872 42068 15873 ne
rect 42068 15872 42162 15873
tri 42068 15871 42069 15872 ne
rect 42069 15871 42162 15872
tri 42069 15870 42070 15871 ne
rect 42070 15870 42162 15871
rect 42208 15903 42268 15916
tri 42268 15903 42313 15948 sw
rect 70802 15932 71000 15990
rect 42208 15902 42313 15903
tri 42313 15902 42314 15903 sw
rect 42208 15870 42314 15902
tri 42070 15869 42071 15870 ne
rect 42071 15869 42314 15870
tri 42071 15868 42072 15869 ne
rect 42072 15868 42314 15869
tri 42072 15867 42073 15868 ne
rect 42073 15867 42314 15868
tri 42073 15866 42074 15867 ne
rect 42074 15866 42314 15867
tri 42074 15865 42075 15866 ne
rect 42075 15865 42314 15866
tri 42075 15864 42076 15865 ne
rect 42076 15864 42314 15865
tri 42076 15863 42077 15864 ne
rect 42077 15863 42314 15864
tri 42077 15862 42078 15863 ne
rect 42078 15862 42314 15863
tri 42078 15861 42079 15862 ne
rect 42079 15861 42314 15862
tri 42079 15860 42080 15861 ne
rect 42080 15860 42314 15861
tri 42080 15859 42081 15860 ne
rect 42081 15859 42314 15860
tri 42081 15858 42082 15859 ne
rect 42082 15858 42314 15859
tri 42082 15857 42083 15858 ne
rect 42083 15857 42314 15858
tri 42314 15857 42359 15902 sw
rect 70802 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
tri 42083 15812 42128 15857 ne
rect 42128 15812 42359 15857
tri 42359 15812 42404 15857 sw
rect 70802 15828 71000 15886
tri 42128 15767 42173 15812 ne
rect 42173 15784 42404 15812
rect 42173 15767 42294 15784
tri 42173 15761 42179 15767 ne
rect 42179 15761 42294 15767
tri 42179 15760 42180 15761 ne
rect 42180 15760 42294 15761
tri 42180 15759 42181 15760 ne
rect 42181 15759 42294 15760
tri 42181 15758 42182 15759 ne
rect 42182 15758 42294 15759
tri 42182 15757 42183 15758 ne
rect 42183 15757 42294 15758
tri 42183 15756 42184 15757 ne
rect 42184 15756 42294 15757
tri 42184 15755 42185 15756 ne
rect 42185 15755 42294 15756
tri 42185 15754 42186 15755 ne
rect 42186 15754 42294 15755
tri 42186 15753 42187 15754 ne
rect 42187 15753 42294 15754
tri 42187 15752 42188 15753 ne
rect 42188 15752 42294 15753
tri 42188 15751 42189 15752 ne
rect 42189 15751 42294 15752
tri 42189 15750 42190 15751 ne
rect 42190 15750 42294 15751
tri 42190 15749 42191 15750 ne
rect 42191 15749 42294 15750
tri 42191 15748 42192 15749 ne
rect 42192 15748 42294 15749
tri 42192 15747 42193 15748 ne
rect 42193 15747 42294 15748
tri 42193 15746 42194 15747 ne
rect 42194 15746 42294 15747
tri 42194 15745 42195 15746 ne
rect 42195 15745 42294 15746
tri 42195 15744 42196 15745 ne
rect 42196 15744 42294 15745
tri 42196 15743 42197 15744 ne
rect 42197 15743 42294 15744
tri 42197 15742 42198 15743 ne
rect 42198 15742 42294 15743
tri 42198 15741 42199 15742 ne
rect 42199 15741 42294 15742
tri 42199 15740 42200 15741 ne
rect 42200 15740 42294 15741
tri 42200 15739 42201 15740 ne
rect 42201 15739 42294 15740
tri 42201 15738 42202 15739 ne
rect 42202 15738 42294 15739
rect 42340 15767 42404 15784
tri 42404 15767 42449 15812 sw
rect 70802 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15762 42449 15767
tri 42449 15762 42454 15767 sw
rect 42340 15738 42454 15762
tri 42202 15737 42203 15738 ne
rect 42203 15737 42454 15738
tri 42203 15736 42204 15737 ne
rect 42204 15736 42454 15737
tri 42204 15735 42205 15736 ne
rect 42205 15735 42454 15736
tri 42205 15734 42206 15735 ne
rect 42206 15734 42454 15735
tri 42206 15733 42207 15734 ne
rect 42207 15733 42454 15734
tri 42207 15732 42208 15733 ne
rect 42208 15732 42454 15733
tri 42208 15731 42209 15732 ne
rect 42209 15731 42454 15732
tri 42209 15730 42210 15731 ne
rect 42210 15730 42454 15731
tri 42210 15729 42211 15730 ne
rect 42211 15729 42454 15730
tri 42211 15728 42212 15729 ne
rect 42212 15728 42454 15729
tri 42212 15727 42213 15728 ne
rect 42213 15727 42454 15728
tri 42213 15726 42214 15727 ne
rect 42214 15726 42454 15727
tri 42214 15725 42215 15726 ne
rect 42215 15725 42454 15726
tri 42215 15724 42216 15725 ne
rect 42216 15724 42454 15725
tri 42216 15723 42217 15724 ne
rect 42217 15723 42454 15724
tri 42217 15722 42218 15723 ne
rect 42218 15722 42454 15723
tri 42218 15721 42219 15722 ne
rect 42219 15721 42454 15722
tri 42219 15720 42220 15721 ne
rect 42220 15720 42454 15721
tri 42220 15719 42221 15720 ne
rect 42221 15719 42454 15720
tri 42221 15718 42222 15719 ne
rect 42222 15718 42454 15719
tri 42222 15717 42223 15718 ne
rect 42223 15717 42454 15718
tri 42454 15717 42499 15762 sw
rect 70802 15724 71000 15782
tri 42223 15716 42224 15717 ne
rect 42224 15716 42499 15717
tri 42224 15715 42225 15716 ne
rect 42225 15715 42499 15716
tri 42225 15714 42226 15715 ne
rect 42226 15714 42499 15715
tri 42226 15713 42227 15714 ne
rect 42227 15713 42499 15714
tri 42227 15712 42228 15713 ne
rect 42228 15712 42499 15713
tri 42228 15711 42229 15712 ne
rect 42229 15711 42499 15712
tri 42229 15710 42230 15711 ne
rect 42230 15710 42499 15711
tri 42230 15709 42231 15710 ne
rect 42231 15709 42499 15710
tri 42231 15708 42232 15709 ne
rect 42232 15708 42499 15709
tri 42232 15707 42233 15708 ne
rect 42233 15707 42499 15708
tri 42233 15706 42234 15707 ne
rect 42234 15706 42499 15707
tri 42234 15705 42235 15706 ne
rect 42235 15705 42499 15706
tri 42235 15704 42236 15705 ne
rect 42236 15704 42499 15705
tri 42236 15703 42237 15704 ne
rect 42237 15703 42499 15704
tri 42237 15702 42238 15703 ne
rect 42238 15702 42499 15703
tri 42238 15701 42239 15702 ne
rect 42239 15701 42499 15702
tri 42239 15700 42240 15701 ne
rect 42240 15700 42499 15701
tri 42240 15699 42241 15700 ne
rect 42241 15699 42499 15700
tri 42241 15698 42242 15699 ne
rect 42242 15698 42499 15699
tri 42242 15697 42243 15698 ne
rect 42243 15697 42499 15698
tri 42243 15696 42244 15697 ne
rect 42244 15696 42499 15697
tri 42244 15695 42245 15696 ne
rect 42245 15695 42499 15696
tri 42245 15694 42246 15695 ne
rect 42246 15694 42499 15695
tri 42246 15693 42247 15694 ne
rect 42247 15693 42499 15694
tri 42247 15692 42248 15693 ne
rect 42248 15692 42499 15693
tri 42248 15691 42249 15692 ne
rect 42249 15691 42499 15692
tri 42249 15690 42250 15691 ne
rect 42250 15690 42499 15691
tri 42250 15689 42251 15690 ne
rect 42251 15689 42499 15690
tri 42251 15688 42252 15689 ne
rect 42252 15688 42499 15689
tri 42252 15687 42253 15688 ne
rect 42253 15687 42499 15688
tri 42253 15686 42254 15687 ne
rect 42254 15686 42499 15687
tri 42254 15685 42255 15686 ne
rect 42255 15685 42499 15686
tri 42255 15684 42256 15685 ne
rect 42256 15684 42499 15685
tri 42256 15683 42257 15684 ne
rect 42257 15683 42499 15684
tri 42257 15682 42258 15683 ne
rect 42258 15682 42499 15683
tri 42258 15681 42259 15682 ne
rect 42259 15681 42499 15682
tri 42259 15680 42260 15681 ne
rect 42260 15680 42499 15681
tri 42260 15679 42261 15680 ne
rect 42261 15679 42499 15680
tri 42261 15678 42262 15679 ne
rect 42262 15678 42499 15679
tri 42262 15677 42263 15678 ne
rect 42263 15677 42499 15678
tri 42263 15676 42264 15677 ne
rect 42264 15676 42499 15677
tri 42264 15675 42265 15676 ne
rect 42265 15675 42499 15676
tri 42265 15674 42266 15675 ne
rect 42266 15674 42499 15675
tri 42266 15673 42267 15674 ne
rect 42267 15673 42499 15674
tri 42267 15672 42268 15673 ne
rect 42268 15672 42499 15673
tri 42499 15672 42544 15717 sw
rect 70802 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
tri 42268 15671 42269 15672 ne
rect 42269 15671 42544 15672
tri 42269 15670 42270 15671 ne
rect 42270 15670 42544 15671
tri 42270 15669 42271 15670 ne
rect 42271 15669 42544 15670
tri 42271 15668 42272 15669 ne
rect 42272 15668 42544 15669
tri 42272 15667 42273 15668 ne
rect 42273 15667 42544 15668
tri 42273 15666 42274 15667 ne
rect 42274 15666 42544 15667
tri 42274 15665 42275 15666 ne
rect 42275 15665 42544 15666
tri 42275 15664 42276 15665 ne
rect 42276 15664 42544 15665
tri 42276 15663 42277 15664 ne
rect 42277 15663 42544 15664
tri 42277 15662 42278 15663 ne
rect 42278 15662 42544 15663
tri 42278 15661 42279 15662 ne
rect 42279 15661 42544 15662
tri 42279 15660 42280 15661 ne
rect 42280 15660 42544 15661
tri 42280 15659 42281 15660 ne
rect 42281 15659 42544 15660
tri 42281 15658 42282 15659 ne
rect 42282 15658 42544 15659
tri 42282 15657 42283 15658 ne
rect 42283 15657 42544 15658
tri 42283 15656 42284 15657 ne
rect 42284 15656 42544 15657
tri 42284 15655 42285 15656 ne
rect 42285 15655 42544 15656
tri 42285 15654 42286 15655 ne
rect 42286 15654 42544 15655
tri 42286 15653 42287 15654 ne
rect 42287 15653 42544 15654
tri 42287 15652 42288 15653 ne
rect 42288 15652 42544 15653
tri 42288 15651 42289 15652 ne
rect 42289 15651 42426 15652
tri 42289 15650 42290 15651 ne
rect 42290 15650 42426 15651
tri 42290 15649 42291 15650 ne
rect 42291 15649 42426 15650
tri 42291 15648 42292 15649 ne
rect 42292 15648 42426 15649
tri 42292 15647 42293 15648 ne
rect 42293 15647 42426 15648
tri 42293 15646 42294 15647 ne
rect 42294 15646 42426 15647
tri 42294 15645 42295 15646 ne
rect 42295 15645 42426 15646
tri 42295 15644 42296 15645 ne
rect 42296 15644 42426 15645
tri 42296 15643 42297 15644 ne
rect 42297 15643 42426 15644
tri 42297 15642 42298 15643 ne
rect 42298 15642 42426 15643
tri 42298 15641 42299 15642 ne
rect 42299 15641 42426 15642
tri 42299 15640 42300 15641 ne
rect 42300 15640 42426 15641
tri 42300 15639 42301 15640 ne
rect 42301 15639 42426 15640
tri 42301 15638 42302 15639 ne
rect 42302 15638 42426 15639
tri 42302 15637 42303 15638 ne
rect 42303 15637 42426 15638
tri 42303 15636 42304 15637 ne
rect 42304 15636 42426 15637
tri 42304 15635 42305 15636 ne
rect 42305 15635 42426 15636
tri 42305 15634 42306 15635 ne
rect 42306 15634 42426 15635
tri 42306 15633 42307 15634 ne
rect 42307 15633 42426 15634
tri 42307 15632 42308 15633 ne
rect 42308 15632 42426 15633
tri 42308 15631 42309 15632 ne
rect 42309 15631 42426 15632
tri 42309 15630 42310 15631 ne
rect 42310 15630 42426 15631
tri 42310 15629 42311 15630 ne
rect 42311 15629 42426 15630
tri 42311 15628 42312 15629 ne
rect 42312 15628 42426 15629
tri 42312 15627 42313 15628 ne
rect 42313 15627 42426 15628
tri 42313 15626 42314 15627 ne
rect 42314 15626 42426 15627
tri 42314 15625 42315 15626 ne
rect 42315 15625 42426 15626
tri 42315 15624 42316 15625 ne
rect 42316 15624 42426 15625
tri 42316 15623 42317 15624 ne
rect 42317 15623 42426 15624
tri 42317 15622 42318 15623 ne
rect 42318 15622 42426 15623
tri 42318 15621 42319 15622 ne
rect 42319 15621 42426 15622
tri 42319 15620 42320 15621 ne
rect 42320 15620 42426 15621
tri 42320 15619 42321 15620 ne
rect 42321 15619 42426 15620
tri 42321 15618 42322 15619 ne
rect 42322 15618 42426 15619
tri 42322 15617 42323 15618 ne
rect 42323 15617 42426 15618
tri 42323 15616 42324 15617 ne
rect 42324 15616 42426 15617
tri 42324 15615 42325 15616 ne
rect 42325 15615 42426 15616
tri 42325 15614 42326 15615 ne
rect 42326 15614 42426 15615
tri 42326 15613 42327 15614 ne
rect 42327 15613 42426 15614
tri 42327 15612 42328 15613 ne
rect 42328 15612 42426 15613
tri 42328 15611 42329 15612 ne
rect 42329 15611 42426 15612
tri 42329 15610 42330 15611 ne
rect 42330 15610 42426 15611
tri 42330 15609 42331 15610 ne
rect 42331 15609 42426 15610
tri 42331 15608 42332 15609 ne
rect 42332 15608 42426 15609
tri 42332 15607 42333 15608 ne
rect 42333 15607 42426 15608
tri 42333 15606 42334 15607 ne
rect 42334 15606 42426 15607
rect 42472 15627 42544 15652
tri 42544 15627 42589 15672 sw
rect 42472 15606 42589 15627
tri 42334 15605 42335 15606 ne
rect 42335 15605 42589 15606
tri 42335 15604 42336 15605 ne
rect 42336 15604 42589 15605
tri 42336 15603 42337 15604 ne
rect 42337 15603 42589 15604
tri 42337 15602 42338 15603 ne
rect 42338 15602 42589 15603
tri 42338 15601 42339 15602 ne
rect 42339 15601 42589 15602
tri 42339 15600 42340 15601 ne
rect 42340 15600 42589 15601
tri 42340 15599 42341 15600 ne
rect 42341 15599 42589 15600
tri 42341 15598 42342 15599 ne
rect 42342 15598 42589 15599
tri 42342 15597 42343 15598 ne
rect 42343 15597 42589 15598
tri 42343 15596 42344 15597 ne
rect 42344 15596 42589 15597
tri 42344 15595 42345 15596 ne
rect 42345 15595 42589 15596
tri 42345 15594 42346 15595 ne
rect 42346 15594 42589 15595
tri 42346 15593 42347 15594 ne
rect 42347 15593 42589 15594
tri 42347 15592 42348 15593 ne
rect 42348 15592 42589 15593
tri 42348 15591 42349 15592 ne
rect 42349 15591 42589 15592
tri 42349 15590 42350 15591 ne
rect 42350 15590 42589 15591
tri 42350 15589 42351 15590 ne
rect 42351 15589 42589 15590
tri 42351 15588 42352 15589 ne
rect 42352 15588 42589 15589
tri 42352 15587 42353 15588 ne
rect 42353 15587 42589 15588
tri 42353 15586 42354 15587 ne
rect 42354 15586 42589 15587
tri 42354 15585 42355 15586 ne
rect 42355 15585 42589 15586
tri 42355 15584 42356 15585 ne
rect 42356 15584 42589 15585
tri 42356 15583 42357 15584 ne
rect 42357 15583 42589 15584
tri 42357 15582 42358 15583 ne
rect 42358 15582 42589 15583
tri 42589 15582 42634 15627 sw
rect 70802 15620 71000 15678
tri 42358 15581 42359 15582 ne
rect 42359 15581 42634 15582
tri 42634 15581 42635 15582 sw
tri 42359 15557 42383 15581 ne
rect 42383 15557 42635 15581
tri 42383 15512 42428 15557 ne
rect 42428 15536 42635 15557
tri 42635 15536 42680 15581 sw
rect 70802 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
rect 42428 15520 42680 15536
rect 42428 15512 42558 15520
tri 42428 15486 42454 15512 ne
rect 42454 15486 42558 15512
tri 42454 15485 42455 15486 ne
rect 42455 15485 42558 15486
tri 42455 15484 42456 15485 ne
rect 42456 15484 42558 15485
tri 42456 15483 42457 15484 ne
rect 42457 15483 42558 15484
tri 42457 15482 42458 15483 ne
rect 42458 15482 42558 15483
tri 42458 15481 42459 15482 ne
rect 42459 15481 42558 15482
tri 42459 15480 42460 15481 ne
rect 42460 15480 42558 15481
tri 42460 15479 42461 15480 ne
rect 42461 15479 42558 15480
tri 42461 15478 42462 15479 ne
rect 42462 15478 42558 15479
tri 42462 15477 42463 15478 ne
rect 42463 15477 42558 15478
tri 42463 15476 42464 15477 ne
rect 42464 15476 42558 15477
tri 42464 15475 42465 15476 ne
rect 42465 15475 42558 15476
tri 42465 15474 42466 15475 ne
rect 42466 15474 42558 15475
rect 42604 15491 42680 15520
tri 42680 15491 42725 15536 sw
rect 70802 15516 71000 15574
rect 42604 15474 42725 15491
tri 42466 15473 42467 15474 ne
rect 42467 15473 42725 15474
tri 42467 15472 42468 15473 ne
rect 42468 15472 42725 15473
tri 42468 15471 42469 15472 ne
rect 42469 15471 42725 15472
tri 42469 15470 42470 15471 ne
rect 42470 15470 42725 15471
tri 42470 15469 42471 15470 ne
rect 42471 15469 42725 15470
tri 42471 15468 42472 15469 ne
rect 42472 15468 42725 15469
tri 42472 15467 42473 15468 ne
rect 42473 15467 42725 15468
tri 42473 15466 42474 15467 ne
rect 42474 15466 42725 15467
tri 42474 15465 42475 15466 ne
rect 42475 15465 42725 15466
tri 42475 15464 42476 15465 ne
rect 42476 15464 42725 15465
tri 42476 15463 42477 15464 ne
rect 42477 15463 42725 15464
tri 42477 15462 42478 15463 ne
rect 42478 15462 42725 15463
tri 42478 15461 42479 15462 ne
rect 42479 15461 42725 15462
tri 42479 15460 42480 15461 ne
rect 42480 15460 42725 15461
tri 42480 15459 42481 15460 ne
rect 42481 15459 42725 15460
tri 42481 15458 42482 15459 ne
rect 42482 15458 42725 15459
tri 42482 15457 42483 15458 ne
rect 42483 15457 42725 15458
tri 42483 15456 42484 15457 ne
rect 42484 15456 42725 15457
tri 42484 15455 42485 15456 ne
rect 42485 15455 42725 15456
tri 42485 15454 42486 15455 ne
rect 42486 15454 42725 15455
tri 42486 15453 42487 15454 ne
rect 42487 15453 42725 15454
tri 42487 15452 42488 15453 ne
rect 42488 15452 42725 15453
tri 42488 15451 42489 15452 ne
rect 42489 15451 42725 15452
tri 42489 15450 42490 15451 ne
rect 42490 15450 42725 15451
tri 42490 15449 42491 15450 ne
rect 42491 15449 42725 15450
tri 42491 15448 42492 15449 ne
rect 42492 15448 42725 15449
tri 42492 15447 42493 15448 ne
rect 42493 15447 42725 15448
tri 42493 15446 42494 15447 ne
rect 42494 15446 42725 15447
tri 42725 15446 42770 15491 sw
rect 70802 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
tri 42494 15445 42495 15446 ne
rect 42495 15445 42770 15446
tri 42495 15444 42496 15445 ne
rect 42496 15444 42770 15445
tri 42496 15443 42497 15444 ne
rect 42497 15443 42770 15444
tri 42497 15442 42498 15443 ne
rect 42498 15442 42770 15443
tri 42498 15441 42499 15442 ne
rect 42499 15441 42770 15442
tri 42499 15440 42500 15441 ne
rect 42500 15440 42770 15441
tri 42770 15440 42776 15446 sw
tri 42500 15439 42501 15440 ne
rect 42501 15439 42776 15440
tri 42501 15438 42502 15439 ne
rect 42502 15438 42776 15439
tri 42502 15437 42503 15438 ne
rect 42503 15437 42776 15438
tri 42503 15436 42504 15437 ne
rect 42504 15436 42776 15437
tri 42504 15435 42505 15436 ne
rect 42505 15435 42776 15436
tri 42505 15434 42506 15435 ne
rect 42506 15434 42776 15435
tri 42506 15433 42507 15434 ne
rect 42507 15433 42776 15434
tri 42507 15432 42508 15433 ne
rect 42508 15432 42776 15433
tri 42508 15431 42509 15432 ne
rect 42509 15431 42776 15432
tri 42509 15430 42510 15431 ne
rect 42510 15430 42776 15431
tri 42510 15429 42511 15430 ne
rect 42511 15429 42776 15430
tri 42511 15428 42512 15429 ne
rect 42512 15428 42776 15429
tri 42512 15427 42513 15428 ne
rect 42513 15427 42776 15428
tri 42513 15426 42514 15427 ne
rect 42514 15426 42776 15427
tri 42514 15425 42515 15426 ne
rect 42515 15425 42776 15426
tri 42515 15424 42516 15425 ne
rect 42516 15424 42776 15425
tri 42516 15423 42517 15424 ne
rect 42517 15423 42776 15424
tri 42517 15422 42518 15423 ne
rect 42518 15422 42776 15423
tri 42518 15421 42519 15422 ne
rect 42519 15421 42776 15422
tri 42519 15420 42520 15421 ne
rect 42520 15420 42776 15421
tri 42520 15419 42521 15420 ne
rect 42521 15419 42776 15420
tri 42521 15418 42522 15419 ne
rect 42522 15418 42776 15419
tri 42522 15417 42523 15418 ne
rect 42523 15417 42776 15418
tri 42523 15416 42524 15417 ne
rect 42524 15416 42776 15417
tri 42524 15415 42525 15416 ne
rect 42525 15415 42776 15416
tri 42525 15414 42526 15415 ne
rect 42526 15414 42776 15415
tri 42526 15413 42527 15414 ne
rect 42527 15413 42776 15414
tri 42527 15412 42528 15413 ne
rect 42528 15412 42776 15413
tri 42528 15411 42529 15412 ne
rect 42529 15411 42776 15412
tri 42529 15410 42530 15411 ne
rect 42530 15410 42776 15411
tri 42530 15409 42531 15410 ne
rect 42531 15409 42776 15410
tri 42531 15408 42532 15409 ne
rect 42532 15408 42776 15409
tri 42532 15407 42533 15408 ne
rect 42533 15407 42776 15408
tri 42533 15406 42534 15407 ne
rect 42534 15406 42776 15407
tri 42534 15405 42535 15406 ne
rect 42535 15405 42776 15406
tri 42535 15404 42536 15405 ne
rect 42536 15404 42776 15405
tri 42536 15403 42537 15404 ne
rect 42537 15403 42776 15404
tri 42537 15402 42538 15403 ne
rect 42538 15402 42776 15403
tri 42538 15401 42539 15402 ne
rect 42539 15401 42776 15402
tri 42539 15400 42540 15401 ne
rect 42540 15400 42776 15401
tri 42540 15399 42541 15400 ne
rect 42541 15399 42776 15400
tri 42541 15398 42542 15399 ne
rect 42542 15398 42776 15399
tri 42542 15397 42543 15398 ne
rect 42543 15397 42776 15398
tri 42543 15396 42544 15397 ne
rect 42544 15396 42776 15397
tri 42544 15395 42545 15396 ne
rect 42545 15395 42776 15396
tri 42776 15395 42821 15440 sw
rect 70802 15412 71000 15470
tri 42545 15394 42546 15395 ne
rect 42546 15394 42821 15395
tri 42546 15393 42547 15394 ne
rect 42547 15393 42821 15394
tri 42547 15392 42548 15393 ne
rect 42548 15392 42821 15393
tri 42548 15391 42549 15392 ne
rect 42549 15391 42821 15392
tri 42549 15390 42550 15391 ne
rect 42550 15390 42821 15391
tri 42550 15389 42551 15390 ne
rect 42551 15389 42821 15390
tri 42551 15388 42552 15389 ne
rect 42552 15388 42821 15389
tri 42552 15387 42553 15388 ne
rect 42553 15387 42690 15388
tri 42553 15386 42554 15387 ne
rect 42554 15386 42690 15387
tri 42554 15385 42555 15386 ne
rect 42555 15385 42690 15386
tri 42555 15384 42556 15385 ne
rect 42556 15384 42690 15385
tri 42556 15383 42557 15384 ne
rect 42557 15383 42690 15384
tri 42557 15382 42558 15383 ne
rect 42558 15382 42690 15383
tri 42558 15381 42559 15382 ne
rect 42559 15381 42690 15382
tri 42559 15380 42560 15381 ne
rect 42560 15380 42690 15381
tri 42560 15379 42561 15380 ne
rect 42561 15379 42690 15380
tri 42561 15378 42562 15379 ne
rect 42562 15378 42690 15379
tri 42562 15377 42563 15378 ne
rect 42563 15377 42690 15378
tri 42563 15376 42564 15377 ne
rect 42564 15376 42690 15377
tri 42564 15375 42565 15376 ne
rect 42565 15375 42690 15376
tri 42565 15374 42566 15375 ne
rect 42566 15374 42690 15375
tri 42566 15373 42567 15374 ne
rect 42567 15373 42690 15374
tri 42567 15372 42568 15373 ne
rect 42568 15372 42690 15373
tri 42568 15371 42569 15372 ne
rect 42569 15371 42690 15372
tri 42569 15370 42570 15371 ne
rect 42570 15370 42690 15371
tri 42570 15369 42571 15370 ne
rect 42571 15369 42690 15370
tri 42571 15368 42572 15369 ne
rect 42572 15368 42690 15369
tri 42572 15367 42573 15368 ne
rect 42573 15367 42690 15368
tri 42573 15366 42574 15367 ne
rect 42574 15366 42690 15367
tri 42574 15365 42575 15366 ne
rect 42575 15365 42690 15366
tri 42575 15364 42576 15365 ne
rect 42576 15364 42690 15365
tri 42576 15363 42577 15364 ne
rect 42577 15363 42690 15364
tri 42577 15362 42578 15363 ne
rect 42578 15362 42690 15363
tri 42578 15361 42579 15362 ne
rect 42579 15361 42690 15362
tri 42579 15360 42580 15361 ne
rect 42580 15360 42690 15361
tri 42580 15359 42581 15360 ne
rect 42581 15359 42690 15360
tri 42581 15358 42582 15359 ne
rect 42582 15358 42690 15359
tri 42582 15357 42583 15358 ne
rect 42583 15357 42690 15358
tri 42583 15356 42584 15357 ne
rect 42584 15356 42690 15357
tri 42584 15355 42585 15356 ne
rect 42585 15355 42690 15356
tri 42585 15354 42586 15355 ne
rect 42586 15354 42690 15355
tri 42586 15353 42587 15354 ne
rect 42587 15353 42690 15354
tri 42587 15352 42588 15353 ne
rect 42588 15352 42690 15353
tri 42588 15351 42589 15352 ne
rect 42589 15351 42690 15352
tri 42589 15350 42590 15351 ne
rect 42590 15350 42690 15351
tri 42590 15349 42591 15350 ne
rect 42591 15349 42690 15350
tri 42591 15348 42592 15349 ne
rect 42592 15348 42690 15349
tri 42592 15347 42593 15348 ne
rect 42593 15347 42690 15348
tri 42593 15346 42594 15347 ne
rect 42594 15346 42690 15347
tri 42594 15345 42595 15346 ne
rect 42595 15345 42690 15346
tri 42595 15344 42596 15345 ne
rect 42596 15344 42690 15345
tri 42596 15343 42597 15344 ne
rect 42597 15343 42690 15344
tri 42597 15342 42598 15343 ne
rect 42598 15342 42690 15343
rect 42736 15350 42821 15388
tri 42821 15350 42866 15395 sw
rect 70802 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15342 42866 15350
tri 42598 15341 42599 15342 ne
rect 42599 15341 42866 15342
tri 42599 15340 42600 15341 ne
rect 42600 15340 42866 15341
tri 42600 15339 42601 15340 ne
rect 42601 15339 42866 15340
tri 42601 15338 42602 15339 ne
rect 42602 15338 42866 15339
tri 42602 15337 42603 15338 ne
rect 42603 15337 42866 15338
tri 42603 15336 42604 15337 ne
rect 42604 15336 42866 15337
tri 42604 15335 42605 15336 ne
rect 42605 15335 42866 15336
tri 42605 15334 42606 15335 ne
rect 42606 15334 42866 15335
tri 42606 15333 42607 15334 ne
rect 42607 15333 42866 15334
tri 42607 15332 42608 15333 ne
rect 42608 15332 42866 15333
tri 42608 15331 42609 15332 ne
rect 42609 15331 42866 15332
tri 42609 15330 42610 15331 ne
rect 42610 15330 42866 15331
tri 42610 15329 42611 15330 ne
rect 42611 15329 42866 15330
tri 42611 15328 42612 15329 ne
rect 42612 15328 42866 15329
tri 42612 15327 42613 15328 ne
rect 42613 15327 42866 15328
tri 42613 15326 42614 15327 ne
rect 42614 15326 42866 15327
tri 42614 15325 42615 15326 ne
rect 42615 15325 42866 15326
tri 42615 15324 42616 15325 ne
rect 42616 15324 42866 15325
tri 42616 15323 42617 15324 ne
rect 42617 15323 42866 15324
tri 42617 15322 42618 15323 ne
rect 42618 15322 42866 15323
tri 42618 15321 42619 15322 ne
rect 42619 15321 42866 15322
tri 42619 15320 42620 15321 ne
rect 42620 15320 42866 15321
tri 42620 15319 42621 15320 ne
rect 42621 15319 42866 15320
tri 42621 15318 42622 15319 ne
rect 42622 15318 42866 15319
tri 42622 15317 42623 15318 ne
rect 42623 15317 42866 15318
tri 42623 15316 42624 15317 ne
rect 42624 15316 42866 15317
tri 42624 15315 42625 15316 ne
rect 42625 15315 42866 15316
tri 42625 15314 42626 15315 ne
rect 42626 15314 42866 15315
tri 42626 15313 42627 15314 ne
rect 42627 15313 42866 15314
tri 42627 15312 42628 15313 ne
rect 42628 15312 42866 15313
tri 42628 15311 42629 15312 ne
rect 42629 15311 42866 15312
tri 42629 15310 42630 15311 ne
rect 42630 15310 42866 15311
tri 42630 15309 42631 15310 ne
rect 42631 15309 42866 15310
tri 42631 15308 42632 15309 ne
rect 42632 15308 42866 15309
tri 42632 15307 42633 15308 ne
rect 42633 15307 42866 15308
tri 42633 15306 42634 15307 ne
rect 42634 15306 42866 15307
tri 42634 15305 42635 15306 ne
rect 42635 15305 42866 15306
tri 42866 15305 42911 15350 sw
rect 70802 15308 71000 15366
tri 42635 15261 42679 15305 ne
rect 42679 15261 42911 15305
tri 42911 15261 42955 15305 sw
rect 70802 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
tri 42679 15216 42724 15261 ne
rect 42724 15256 42955 15261
rect 42724 15216 42822 15256
tri 42724 15212 42728 15216 ne
rect 42728 15212 42822 15216
tri 42728 15211 42729 15212 ne
rect 42729 15211 42822 15212
tri 42729 15210 42730 15211 ne
rect 42730 15210 42822 15211
rect 42868 15216 42955 15256
tri 42955 15216 43000 15261 sw
rect 42868 15210 43000 15216
tri 42730 15209 42731 15210 ne
rect 42731 15209 43000 15210
tri 42731 15208 42732 15209 ne
rect 42732 15208 43000 15209
tri 42732 15207 42733 15208 ne
rect 42733 15207 43000 15208
tri 42733 15206 42734 15207 ne
rect 42734 15206 43000 15207
tri 42734 15205 42735 15206 ne
rect 42735 15205 43000 15206
tri 42735 15204 42736 15205 ne
rect 42736 15204 43000 15205
tri 42736 15203 42737 15204 ne
rect 42737 15203 43000 15204
tri 42737 15202 42738 15203 ne
rect 42738 15202 43000 15203
tri 42738 15201 42739 15202 ne
rect 42739 15201 43000 15202
tri 42739 15200 42740 15201 ne
rect 42740 15200 43000 15201
tri 42740 15199 42741 15200 ne
rect 42741 15199 43000 15200
tri 42741 15198 42742 15199 ne
rect 42742 15198 43000 15199
tri 42742 15197 42743 15198 ne
rect 42743 15197 43000 15198
tri 42743 15196 42744 15197 ne
rect 42744 15196 43000 15197
tri 42744 15195 42745 15196 ne
rect 42745 15195 43000 15196
tri 42745 15194 42746 15195 ne
rect 42746 15194 43000 15195
tri 42746 15193 42747 15194 ne
rect 42747 15193 43000 15194
tri 42747 15192 42748 15193 ne
rect 42748 15192 43000 15193
tri 42748 15191 42749 15192 ne
rect 42749 15191 43000 15192
tri 42749 15190 42750 15191 ne
rect 42750 15190 43000 15191
tri 42750 15189 42751 15190 ne
rect 42751 15189 43000 15190
tri 42751 15188 42752 15189 ne
rect 42752 15188 43000 15189
tri 42752 15187 42753 15188 ne
rect 42753 15187 43000 15188
tri 42753 15186 42754 15187 ne
rect 42754 15186 43000 15187
tri 42754 15185 42755 15186 ne
rect 42755 15185 43000 15186
tri 42755 15184 42756 15185 ne
rect 42756 15184 43000 15185
tri 42756 15183 42757 15184 ne
rect 42757 15183 43000 15184
tri 42757 15182 42758 15183 ne
rect 42758 15182 43000 15183
tri 42758 15181 42759 15182 ne
rect 42759 15181 43000 15182
tri 42759 15180 42760 15181 ne
rect 42760 15180 43000 15181
tri 42760 15179 42761 15180 ne
rect 42761 15179 43000 15180
tri 42761 15178 42762 15179 ne
rect 42762 15178 43000 15179
tri 42762 15177 42763 15178 ne
rect 42763 15177 43000 15178
tri 42763 15176 42764 15177 ne
rect 42764 15176 43000 15177
tri 42764 15175 42765 15176 ne
rect 42765 15175 43000 15176
tri 42765 15174 42766 15175 ne
rect 42766 15174 43000 15175
tri 42766 15173 42767 15174 ne
rect 42767 15173 43000 15174
tri 42767 15172 42768 15173 ne
rect 42768 15172 43000 15173
tri 42768 15171 42769 15172 ne
rect 42769 15171 43000 15172
tri 43000 15171 43045 15216 sw
rect 70802 15204 71000 15262
tri 42769 15170 42770 15171 ne
rect 42770 15170 43045 15171
tri 42770 15169 42771 15170 ne
rect 42771 15169 43045 15170
tri 42771 15168 42772 15169 ne
rect 42772 15168 43045 15169
tri 42772 15167 42773 15168 ne
rect 42773 15167 43045 15168
tri 42773 15166 42774 15167 ne
rect 42774 15166 43045 15167
tri 42774 15165 42775 15166 ne
rect 42775 15165 43045 15166
tri 42775 15164 42776 15165 ne
rect 42776 15164 43045 15165
tri 42776 15163 42777 15164 ne
rect 42777 15163 43045 15164
tri 42777 15162 42778 15163 ne
rect 42778 15162 43045 15163
tri 42778 15161 42779 15162 ne
rect 42779 15161 43045 15162
tri 42779 15160 42780 15161 ne
rect 42780 15160 43045 15161
tri 42780 15159 42781 15160 ne
rect 42781 15159 43045 15160
tri 42781 15158 42782 15159 ne
rect 42782 15158 43045 15159
tri 42782 15157 42783 15158 ne
rect 42783 15157 43045 15158
tri 42783 15156 42784 15157 ne
rect 42784 15156 43045 15157
tri 42784 15155 42785 15156 ne
rect 42785 15155 43045 15156
tri 42785 15154 42786 15155 ne
rect 42786 15154 43045 15155
tri 42786 15153 42787 15154 ne
rect 42787 15153 43045 15154
tri 42787 15152 42788 15153 ne
rect 42788 15152 43045 15153
tri 42788 15151 42789 15152 ne
rect 42789 15151 43045 15152
tri 42789 15150 42790 15151 ne
rect 42790 15150 43045 15151
tri 42790 15149 42791 15150 ne
rect 42791 15149 43045 15150
tri 42791 15148 42792 15149 ne
rect 42792 15148 43045 15149
tri 42792 15147 42793 15148 ne
rect 42793 15147 43045 15148
tri 42793 15146 42794 15147 ne
rect 42794 15146 43045 15147
tri 42794 15145 42795 15146 ne
rect 42795 15145 43045 15146
tri 42795 15144 42796 15145 ne
rect 42796 15144 43045 15145
tri 42796 15143 42797 15144 ne
rect 42797 15143 43045 15144
tri 42797 15142 42798 15143 ne
rect 42798 15142 43045 15143
tri 42798 15141 42799 15142 ne
rect 42799 15141 43045 15142
tri 42799 15140 42800 15141 ne
rect 42800 15140 43045 15141
tri 42800 15139 42801 15140 ne
rect 42801 15139 43045 15140
tri 42801 15138 42802 15139 ne
rect 42802 15138 43045 15139
tri 42802 15137 42803 15138 ne
rect 42803 15137 43045 15138
tri 42803 15136 42804 15137 ne
rect 42804 15136 43045 15137
tri 42804 15135 42805 15136 ne
rect 42805 15135 43045 15136
tri 42805 15134 42806 15135 ne
rect 42806 15134 43045 15135
tri 42806 15133 42807 15134 ne
rect 42807 15133 43045 15134
tri 42807 15132 42808 15133 ne
rect 42808 15132 43045 15133
tri 42808 15131 42809 15132 ne
rect 42809 15131 43045 15132
tri 42809 15130 42810 15131 ne
rect 42810 15130 43045 15131
tri 42810 15129 42811 15130 ne
rect 42811 15129 43045 15130
tri 42811 15128 42812 15129 ne
rect 42812 15128 43045 15129
tri 42812 15127 42813 15128 ne
rect 42813 15127 43045 15128
tri 42813 15126 42814 15127 ne
rect 42814 15126 43045 15127
tri 43045 15126 43090 15171 sw
rect 70802 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42814 15125 42815 15126 ne
rect 42815 15125 43090 15126
tri 42815 15124 42816 15125 ne
rect 42816 15124 43090 15125
tri 42816 15123 42817 15124 ne
rect 42817 15123 42954 15124
tri 42817 15122 42818 15123 ne
rect 42818 15122 42954 15123
tri 42818 15121 42819 15122 ne
rect 42819 15121 42954 15122
tri 42819 15120 42820 15121 ne
rect 42820 15120 42954 15121
tri 42820 15119 42821 15120 ne
rect 42821 15119 42954 15120
tri 42821 15118 42822 15119 ne
rect 42822 15118 42954 15119
tri 42822 15117 42823 15118 ne
rect 42823 15117 42954 15118
tri 42823 15116 42824 15117 ne
rect 42824 15116 42954 15117
tri 42824 15115 42825 15116 ne
rect 42825 15115 42954 15116
tri 42825 15114 42826 15115 ne
rect 42826 15114 42954 15115
tri 42826 15113 42827 15114 ne
rect 42827 15113 42954 15114
tri 42827 15112 42828 15113 ne
rect 42828 15112 42954 15113
tri 42828 15111 42829 15112 ne
rect 42829 15111 42954 15112
tri 42829 15110 42830 15111 ne
rect 42830 15110 42954 15111
tri 42830 15109 42831 15110 ne
rect 42831 15109 42954 15110
tri 42831 15108 42832 15109 ne
rect 42832 15108 42954 15109
tri 42832 15107 42833 15108 ne
rect 42833 15107 42954 15108
tri 42833 15106 42834 15107 ne
rect 42834 15106 42954 15107
tri 42834 15105 42835 15106 ne
rect 42835 15105 42954 15106
tri 42835 15104 42836 15105 ne
rect 42836 15104 42954 15105
tri 42836 15103 42837 15104 ne
rect 42837 15103 42954 15104
tri 42837 15102 42838 15103 ne
rect 42838 15102 42954 15103
tri 42838 15101 42839 15102 ne
rect 42839 15101 42954 15102
tri 42839 15100 42840 15101 ne
rect 42840 15100 42954 15101
tri 42840 15099 42841 15100 ne
rect 42841 15099 42954 15100
tri 42841 15098 42842 15099 ne
rect 42842 15098 42954 15099
tri 42842 15097 42843 15098 ne
rect 42843 15097 42954 15098
tri 42843 15096 42844 15097 ne
rect 42844 15096 42954 15097
tri 42844 15095 42845 15096 ne
rect 42845 15095 42954 15096
tri 42845 15094 42846 15095 ne
rect 42846 15094 42954 15095
tri 42846 15093 42847 15094 ne
rect 42847 15093 42954 15094
tri 42847 15092 42848 15093 ne
rect 42848 15092 42954 15093
tri 42848 15091 42849 15092 ne
rect 42849 15091 42954 15092
tri 42849 15090 42850 15091 ne
rect 42850 15090 42954 15091
tri 42850 15089 42851 15090 ne
rect 42851 15089 42954 15090
tri 42851 15088 42852 15089 ne
rect 42852 15088 42954 15089
tri 42852 15087 42853 15088 ne
rect 42853 15087 42954 15088
tri 42853 15086 42854 15087 ne
rect 42854 15086 42954 15087
tri 42854 15085 42855 15086 ne
rect 42855 15085 42954 15086
tri 42855 15084 42856 15085 ne
rect 42856 15084 42954 15085
tri 42856 15083 42857 15084 ne
rect 42857 15083 42954 15084
tri 42857 15082 42858 15083 ne
rect 42858 15082 42954 15083
tri 42858 15081 42859 15082 ne
rect 42859 15081 42954 15082
tri 42859 15080 42860 15081 ne
rect 42860 15080 42954 15081
tri 42860 15079 42861 15080 ne
rect 42861 15079 42954 15080
tri 42861 15078 42862 15079 ne
rect 42862 15078 42954 15079
rect 43000 15119 43090 15124
tri 43090 15119 43097 15126 sw
rect 43000 15078 43097 15119
tri 42862 15077 42863 15078 ne
rect 42863 15077 43097 15078
tri 42863 15076 42864 15077 ne
rect 42864 15076 43097 15077
tri 42864 15075 42865 15076 ne
rect 42865 15075 43097 15076
tri 42865 15074 42866 15075 ne
rect 42866 15074 43097 15075
tri 43097 15074 43142 15119 sw
rect 70802 15100 71000 15158
tri 42866 15073 42867 15074 ne
rect 42867 15073 43142 15074
tri 42867 15072 42868 15073 ne
rect 42868 15072 43142 15073
tri 42868 15071 42869 15072 ne
rect 42869 15071 43142 15072
tri 42869 15070 42870 15071 ne
rect 42870 15070 43142 15071
tri 42870 15069 42871 15070 ne
rect 42871 15069 43142 15070
tri 42871 15068 42872 15069 ne
rect 42872 15068 43142 15069
tri 42872 15067 42873 15068 ne
rect 42873 15067 43142 15068
tri 42873 15066 42874 15067 ne
rect 42874 15066 43142 15067
tri 42874 15065 42875 15066 ne
rect 42875 15065 43142 15066
tri 42875 15064 42876 15065 ne
rect 42876 15064 43142 15065
tri 42876 15063 42877 15064 ne
rect 42877 15063 43142 15064
tri 42877 15062 42878 15063 ne
rect 42878 15062 43142 15063
tri 42878 15061 42879 15062 ne
rect 42879 15061 43142 15062
tri 42879 15060 42880 15061 ne
rect 42880 15060 43142 15061
tri 42880 15059 42881 15060 ne
rect 42881 15059 43142 15060
tri 42881 15058 42882 15059 ne
rect 42882 15058 43142 15059
tri 42882 15057 42883 15058 ne
rect 42883 15057 43142 15058
tri 42883 15056 42884 15057 ne
rect 42884 15056 43142 15057
tri 42884 15055 42885 15056 ne
rect 42885 15055 43142 15056
tri 42885 15054 42886 15055 ne
rect 42886 15054 43142 15055
tri 42886 15053 42887 15054 ne
rect 42887 15053 43142 15054
tri 42887 15052 42888 15053 ne
rect 42888 15052 43142 15053
tri 42888 15051 42889 15052 ne
rect 42889 15051 43142 15052
tri 42889 15050 42890 15051 ne
rect 42890 15050 43142 15051
tri 42890 15049 42891 15050 ne
rect 42891 15049 43142 15050
tri 42891 15048 42892 15049 ne
rect 42892 15048 43142 15049
tri 42892 15047 42893 15048 ne
rect 42893 15047 43142 15048
tri 42893 15046 42894 15047 ne
rect 42894 15046 43142 15047
tri 42894 15045 42895 15046 ne
rect 42895 15045 43142 15046
tri 42895 15044 42896 15045 ne
rect 42896 15044 43142 15045
tri 42896 15043 42897 15044 ne
rect 42897 15043 43142 15044
tri 42897 15042 42898 15043 ne
rect 42898 15042 43142 15043
tri 42898 15041 42899 15042 ne
rect 42899 15041 43142 15042
tri 42899 15040 42900 15041 ne
rect 42900 15040 43142 15041
tri 42900 15039 42901 15040 ne
rect 42901 15039 43142 15040
tri 42901 15038 42902 15039 ne
rect 42902 15038 43142 15039
tri 42902 15037 42903 15038 ne
rect 42903 15037 43142 15038
tri 42903 15036 42904 15037 ne
rect 42904 15036 43142 15037
tri 42904 15035 42905 15036 ne
rect 42905 15035 43142 15036
tri 42905 15034 42906 15035 ne
rect 42906 15034 43142 15035
tri 42906 15033 42907 15034 ne
rect 42907 15033 43142 15034
tri 42907 15032 42908 15033 ne
rect 42908 15032 43142 15033
tri 42908 15031 42909 15032 ne
rect 42909 15031 43142 15032
tri 42909 15030 42910 15031 ne
rect 42910 15030 43142 15031
tri 42910 15029 42911 15030 ne
rect 42911 15029 43142 15030
tri 43142 15029 43187 15074 sw
rect 70802 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42911 14984 42956 15029 ne
rect 42956 14992 43187 15029
rect 42956 14984 43086 14992
tri 42956 14940 43000 14984 ne
rect 43000 14946 43086 14984
rect 43132 14984 43187 14992
tri 43187 14984 43232 15029 sw
rect 70802 14996 71000 15054
rect 43132 14946 43232 14984
rect 43000 14940 43232 14946
tri 43232 14940 43276 14984 sw
rect 70802 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
tri 43000 14939 43001 14940 ne
rect 43001 14939 43276 14940
tri 43001 14937 43003 14939 ne
rect 43003 14937 43276 14939
tri 43003 14936 43004 14937 ne
rect 43004 14936 43276 14937
tri 43004 14935 43005 14936 ne
rect 43005 14935 43276 14936
tri 43005 14934 43006 14935 ne
rect 43006 14934 43276 14935
tri 43006 14933 43007 14934 ne
rect 43007 14933 43276 14934
tri 43007 14932 43008 14933 ne
rect 43008 14932 43276 14933
tri 43008 14931 43009 14932 ne
rect 43009 14931 43276 14932
tri 43009 14930 43010 14931 ne
rect 43010 14930 43276 14931
tri 43010 14929 43011 14930 ne
rect 43011 14929 43276 14930
tri 43011 14928 43012 14929 ne
rect 43012 14928 43276 14929
tri 43012 14927 43013 14928 ne
rect 43013 14927 43276 14928
tri 43013 14926 43014 14927 ne
rect 43014 14926 43276 14927
tri 43014 14925 43015 14926 ne
rect 43015 14925 43276 14926
tri 43015 14924 43016 14925 ne
rect 43016 14924 43276 14925
tri 43016 14923 43017 14924 ne
rect 43017 14923 43276 14924
tri 43017 14922 43018 14923 ne
rect 43018 14922 43276 14923
tri 43018 14921 43019 14922 ne
rect 43019 14921 43276 14922
tri 43019 14920 43020 14921 ne
rect 43020 14920 43276 14921
tri 43020 14919 43021 14920 ne
rect 43021 14919 43276 14920
tri 43021 14918 43022 14919 ne
rect 43022 14918 43276 14919
tri 43022 14917 43023 14918 ne
rect 43023 14917 43276 14918
tri 43023 14916 43024 14917 ne
rect 43024 14916 43276 14917
tri 43024 14915 43025 14916 ne
rect 43025 14915 43276 14916
tri 43025 14914 43026 14915 ne
rect 43026 14914 43276 14915
tri 43026 14913 43027 14914 ne
rect 43027 14913 43276 14914
tri 43027 14912 43028 14913 ne
rect 43028 14912 43276 14913
tri 43028 14911 43029 14912 ne
rect 43029 14911 43276 14912
tri 43029 14910 43030 14911 ne
rect 43030 14910 43276 14911
tri 43030 14909 43031 14910 ne
rect 43031 14909 43276 14910
tri 43031 14908 43032 14909 ne
rect 43032 14908 43276 14909
tri 43032 14907 43033 14908 ne
rect 43033 14907 43276 14908
tri 43033 14906 43034 14907 ne
rect 43034 14906 43276 14907
tri 43034 14905 43035 14906 ne
rect 43035 14905 43276 14906
tri 43035 14904 43036 14905 ne
rect 43036 14904 43276 14905
tri 43036 14903 43037 14904 ne
rect 43037 14903 43276 14904
tri 43037 14902 43038 14903 ne
rect 43038 14902 43276 14903
tri 43038 14901 43039 14902 ne
rect 43039 14901 43276 14902
tri 43039 14900 43040 14901 ne
rect 43040 14900 43276 14901
tri 43040 14899 43041 14900 ne
rect 43041 14899 43276 14900
tri 43041 14898 43042 14899 ne
rect 43042 14898 43276 14899
tri 43042 14897 43043 14898 ne
rect 43043 14897 43276 14898
tri 43043 14896 43044 14897 ne
rect 43044 14896 43276 14897
tri 43044 14895 43045 14896 ne
rect 43045 14895 43276 14896
tri 43276 14895 43321 14940 sw
tri 43045 14894 43046 14895 ne
rect 43046 14894 43321 14895
tri 43046 14893 43047 14894 ne
rect 43047 14893 43321 14894
tri 43047 14892 43048 14893 ne
rect 43048 14892 43321 14893
tri 43048 14891 43049 14892 ne
rect 43049 14891 43321 14892
tri 43049 14890 43050 14891 ne
rect 43050 14890 43321 14891
tri 43050 14889 43051 14890 ne
rect 43051 14889 43321 14890
tri 43051 14888 43052 14889 ne
rect 43052 14888 43321 14889
tri 43052 14887 43053 14888 ne
rect 43053 14887 43321 14888
tri 43053 14886 43054 14887 ne
rect 43054 14886 43321 14887
tri 43054 14885 43055 14886 ne
rect 43055 14885 43321 14886
tri 43055 14884 43056 14885 ne
rect 43056 14884 43321 14885
tri 43056 14883 43057 14884 ne
rect 43057 14883 43321 14884
tri 43057 14882 43058 14883 ne
rect 43058 14882 43321 14883
tri 43058 14881 43059 14882 ne
rect 43059 14881 43321 14882
tri 43059 14880 43060 14881 ne
rect 43060 14880 43321 14881
tri 43060 14879 43061 14880 ne
rect 43061 14879 43321 14880
tri 43061 14878 43062 14879 ne
rect 43062 14878 43321 14879
tri 43062 14877 43063 14878 ne
rect 43063 14877 43321 14878
tri 43063 14876 43064 14877 ne
rect 43064 14876 43321 14877
tri 43064 14875 43065 14876 ne
rect 43065 14875 43321 14876
tri 43065 14874 43066 14875 ne
rect 43066 14874 43321 14875
tri 43066 14873 43067 14874 ne
rect 43067 14873 43321 14874
tri 43067 14872 43068 14873 ne
rect 43068 14872 43321 14873
tri 43068 14871 43069 14872 ne
rect 43069 14871 43321 14872
tri 43069 14870 43070 14871 ne
rect 43070 14870 43321 14871
tri 43070 14869 43071 14870 ne
rect 43071 14869 43321 14870
tri 43071 14868 43072 14869 ne
rect 43072 14868 43321 14869
tri 43072 14867 43073 14868 ne
rect 43073 14867 43321 14868
tri 43073 14866 43074 14867 ne
rect 43074 14866 43321 14867
tri 43074 14865 43075 14866 ne
rect 43075 14865 43321 14866
tri 43075 14864 43076 14865 ne
rect 43076 14864 43321 14865
tri 43076 14863 43077 14864 ne
rect 43077 14863 43321 14864
tri 43077 14862 43078 14863 ne
rect 43078 14862 43321 14863
tri 43078 14861 43079 14862 ne
rect 43079 14861 43321 14862
tri 43079 14860 43080 14861 ne
rect 43080 14860 43321 14861
tri 43080 14859 43081 14860 ne
rect 43081 14859 43218 14860
tri 43081 14858 43082 14859 ne
rect 43082 14858 43218 14859
tri 43082 14857 43083 14858 ne
rect 43083 14857 43218 14858
tri 43083 14856 43084 14857 ne
rect 43084 14856 43218 14857
tri 43084 14855 43085 14856 ne
rect 43085 14855 43218 14856
tri 43085 14854 43086 14855 ne
rect 43086 14854 43218 14855
tri 43086 14853 43087 14854 ne
rect 43087 14853 43218 14854
tri 43087 14852 43088 14853 ne
rect 43088 14852 43218 14853
tri 43088 14851 43089 14852 ne
rect 43089 14851 43218 14852
tri 43089 14850 43090 14851 ne
rect 43090 14850 43218 14851
tri 43090 14849 43091 14850 ne
rect 43091 14849 43218 14850
tri 43091 14848 43092 14849 ne
rect 43092 14848 43218 14849
tri 43092 14847 43093 14848 ne
rect 43093 14847 43218 14848
tri 43093 14846 43094 14847 ne
rect 43094 14846 43218 14847
tri 43094 14845 43095 14846 ne
rect 43095 14845 43218 14846
tri 43095 14844 43096 14845 ne
rect 43096 14844 43218 14845
tri 43096 14843 43097 14844 ne
rect 43097 14843 43218 14844
tri 43097 14842 43098 14843 ne
rect 43098 14842 43218 14843
tri 43098 14841 43099 14842 ne
rect 43099 14841 43218 14842
tri 43099 14840 43100 14841 ne
rect 43100 14840 43218 14841
tri 43100 14839 43101 14840 ne
rect 43101 14839 43218 14840
tri 43101 14838 43102 14839 ne
rect 43102 14838 43218 14839
tri 43102 14837 43103 14838 ne
rect 43103 14837 43218 14838
tri 43103 14836 43104 14837 ne
rect 43104 14836 43218 14837
tri 43104 14835 43105 14836 ne
rect 43105 14835 43218 14836
tri 43105 14834 43106 14835 ne
rect 43106 14834 43218 14835
tri 43106 14833 43107 14834 ne
rect 43107 14833 43218 14834
tri 43107 14832 43108 14833 ne
rect 43108 14832 43218 14833
tri 43108 14831 43109 14832 ne
rect 43109 14831 43218 14832
tri 43109 14830 43110 14831 ne
rect 43110 14830 43218 14831
tri 43110 14829 43111 14830 ne
rect 43111 14829 43218 14830
tri 43111 14828 43112 14829 ne
rect 43112 14828 43218 14829
tri 43112 14827 43113 14828 ne
rect 43113 14827 43218 14828
tri 43113 14826 43114 14827 ne
rect 43114 14826 43218 14827
tri 43114 14825 43115 14826 ne
rect 43115 14825 43218 14826
tri 43115 14824 43116 14825 ne
rect 43116 14824 43218 14825
tri 43116 14823 43117 14824 ne
rect 43117 14823 43218 14824
tri 43117 14822 43118 14823 ne
rect 43118 14822 43218 14823
tri 43118 14821 43119 14822 ne
rect 43119 14821 43218 14822
tri 43119 14820 43120 14821 ne
rect 43120 14820 43218 14821
tri 43120 14819 43121 14820 ne
rect 43121 14819 43218 14820
tri 43121 14818 43122 14819 ne
rect 43122 14818 43218 14819
tri 43122 14817 43123 14818 ne
rect 43123 14817 43218 14818
tri 43123 14816 43124 14817 ne
rect 43124 14816 43218 14817
tri 43124 14815 43125 14816 ne
rect 43125 14815 43218 14816
tri 43125 14814 43126 14815 ne
rect 43126 14814 43218 14815
rect 43264 14850 43321 14860
tri 43321 14850 43366 14895 sw
rect 70802 14892 71000 14950
rect 43264 14814 43366 14850
tri 43126 14813 43127 14814 ne
rect 43127 14813 43366 14814
tri 43127 14812 43128 14813 ne
rect 43128 14812 43366 14813
tri 43128 14811 43129 14812 ne
rect 43129 14811 43366 14812
tri 43129 14810 43130 14811 ne
rect 43130 14810 43366 14811
tri 43130 14809 43131 14810 ne
rect 43131 14809 43366 14810
tri 43131 14808 43132 14809 ne
rect 43132 14808 43366 14809
tri 43132 14807 43133 14808 ne
rect 43133 14807 43366 14808
tri 43133 14806 43134 14807 ne
rect 43134 14806 43366 14807
tri 43134 14805 43135 14806 ne
rect 43135 14805 43366 14806
tri 43366 14805 43411 14850 sw
rect 70802 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
tri 43135 14804 43136 14805 ne
rect 43136 14804 43411 14805
tri 43136 14803 43137 14804 ne
rect 43137 14803 43411 14804
tri 43137 14802 43138 14803 ne
rect 43138 14802 43411 14803
tri 43138 14801 43139 14802 ne
rect 43139 14801 43411 14802
tri 43139 14800 43140 14801 ne
rect 43140 14800 43411 14801
tri 43140 14799 43141 14800 ne
rect 43141 14799 43411 14800
tri 43141 14798 43142 14799 ne
rect 43142 14798 43411 14799
tri 43411 14798 43418 14805 sw
tri 43142 14797 43143 14798 ne
rect 43143 14797 43418 14798
tri 43143 14796 43144 14797 ne
rect 43144 14796 43418 14797
tri 43144 14795 43145 14796 ne
rect 43145 14795 43418 14796
tri 43145 14794 43146 14795 ne
rect 43146 14794 43418 14795
tri 43146 14793 43147 14794 ne
rect 43147 14793 43418 14794
tri 43147 14792 43148 14793 ne
rect 43148 14792 43418 14793
tri 43148 14791 43149 14792 ne
rect 43149 14791 43418 14792
tri 43149 14790 43150 14791 ne
rect 43150 14790 43418 14791
tri 43150 14789 43151 14790 ne
rect 43151 14789 43418 14790
tri 43151 14788 43152 14789 ne
rect 43152 14788 43418 14789
tri 43152 14787 43153 14788 ne
rect 43153 14787 43418 14788
tri 43153 14786 43154 14787 ne
rect 43154 14786 43418 14787
tri 43154 14785 43155 14786 ne
rect 43155 14785 43418 14786
tri 43155 14784 43156 14785 ne
rect 43156 14784 43418 14785
tri 43156 14783 43157 14784 ne
rect 43157 14783 43418 14784
tri 43157 14782 43158 14783 ne
rect 43158 14782 43418 14783
tri 43158 14781 43159 14782 ne
rect 43159 14781 43418 14782
tri 43159 14780 43160 14781 ne
rect 43160 14780 43418 14781
tri 43160 14779 43161 14780 ne
rect 43161 14779 43418 14780
tri 43161 14778 43162 14779 ne
rect 43162 14778 43418 14779
tri 43162 14777 43163 14778 ne
rect 43163 14777 43418 14778
tri 43163 14776 43164 14777 ne
rect 43164 14776 43418 14777
tri 43164 14775 43165 14776 ne
rect 43165 14775 43418 14776
tri 43165 14774 43166 14775 ne
rect 43166 14774 43418 14775
tri 43166 14773 43167 14774 ne
rect 43167 14773 43418 14774
tri 43167 14772 43168 14773 ne
rect 43168 14772 43418 14773
tri 43168 14771 43169 14772 ne
rect 43169 14771 43418 14772
tri 43169 14770 43170 14771 ne
rect 43170 14770 43418 14771
tri 43170 14769 43171 14770 ne
rect 43171 14769 43418 14770
tri 43171 14768 43172 14769 ne
rect 43172 14768 43418 14769
tri 43172 14767 43173 14768 ne
rect 43173 14767 43418 14768
tri 43173 14766 43174 14767 ne
rect 43174 14766 43418 14767
tri 43174 14765 43175 14766 ne
rect 43175 14765 43418 14766
tri 43175 14764 43176 14765 ne
rect 43176 14764 43418 14765
tri 43176 14763 43177 14764 ne
rect 43177 14763 43418 14764
tri 43177 14762 43178 14763 ne
rect 43178 14762 43418 14763
tri 43178 14761 43179 14762 ne
rect 43179 14761 43418 14762
tri 43179 14760 43180 14761 ne
rect 43180 14760 43418 14761
tri 43180 14759 43181 14760 ne
rect 43181 14759 43418 14760
tri 43181 14758 43182 14759 ne
rect 43182 14758 43418 14759
tri 43182 14757 43183 14758 ne
rect 43183 14757 43418 14758
tri 43183 14756 43184 14757 ne
rect 43184 14756 43418 14757
tri 43184 14755 43185 14756 ne
rect 43185 14755 43418 14756
tri 43185 14754 43186 14755 ne
rect 43186 14754 43418 14755
tri 43186 14753 43187 14754 ne
rect 43187 14753 43418 14754
tri 43418 14753 43463 14798 sw
rect 70802 14788 71000 14846
tri 43187 14708 43232 14753 ne
rect 43232 14728 43463 14753
rect 43232 14708 43350 14728
tri 43232 14663 43277 14708 ne
rect 43277 14682 43350 14708
rect 43396 14708 43463 14728
tri 43463 14708 43508 14753 sw
rect 70802 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
rect 43396 14682 43508 14708
rect 43277 14663 43508 14682
tri 43508 14663 43553 14708 sw
rect 70802 14684 71000 14742
tri 43277 14662 43278 14663 ne
rect 43278 14662 43553 14663
tri 43278 14661 43279 14662 ne
rect 43279 14661 43553 14662
tri 43279 14660 43280 14661 ne
rect 43280 14660 43553 14661
tri 43280 14659 43281 14660 ne
rect 43281 14659 43553 14660
tri 43281 14658 43282 14659 ne
rect 43282 14658 43553 14659
tri 43282 14657 43283 14658 ne
rect 43283 14657 43553 14658
tri 43283 14656 43284 14657 ne
rect 43284 14656 43553 14657
tri 43284 14655 43285 14656 ne
rect 43285 14655 43553 14656
tri 43285 14654 43286 14655 ne
rect 43286 14654 43553 14655
tri 43286 14653 43287 14654 ne
rect 43287 14653 43553 14654
tri 43287 14652 43288 14653 ne
rect 43288 14652 43553 14653
tri 43288 14651 43289 14652 ne
rect 43289 14651 43553 14652
tri 43289 14650 43290 14651 ne
rect 43290 14650 43553 14651
tri 43290 14649 43291 14650 ne
rect 43291 14649 43553 14650
tri 43291 14648 43292 14649 ne
rect 43292 14648 43553 14649
tri 43292 14647 43293 14648 ne
rect 43293 14647 43553 14648
tri 43293 14646 43294 14647 ne
rect 43294 14646 43553 14647
tri 43294 14645 43295 14646 ne
rect 43295 14645 43553 14646
tri 43295 14644 43296 14645 ne
rect 43296 14644 43553 14645
tri 43296 14643 43297 14644 ne
rect 43297 14643 43553 14644
tri 43297 14642 43298 14643 ne
rect 43298 14642 43553 14643
tri 43298 14641 43299 14642 ne
rect 43299 14641 43553 14642
tri 43299 14640 43300 14641 ne
rect 43300 14640 43553 14641
tri 43300 14639 43301 14640 ne
rect 43301 14639 43553 14640
tri 43301 14638 43302 14639 ne
rect 43302 14638 43553 14639
tri 43302 14637 43303 14638 ne
rect 43303 14637 43553 14638
tri 43303 14636 43304 14637 ne
rect 43304 14636 43553 14637
tri 43304 14635 43305 14636 ne
rect 43305 14635 43553 14636
tri 43305 14634 43306 14635 ne
rect 43306 14634 43553 14635
tri 43306 14633 43307 14634 ne
rect 43307 14633 43553 14634
tri 43307 14632 43308 14633 ne
rect 43308 14632 43553 14633
tri 43308 14631 43309 14632 ne
rect 43309 14631 43553 14632
tri 43309 14630 43310 14631 ne
rect 43310 14630 43553 14631
tri 43310 14629 43311 14630 ne
rect 43311 14629 43553 14630
tri 43311 14628 43312 14629 ne
rect 43312 14628 43553 14629
tri 43312 14627 43313 14628 ne
rect 43313 14627 43553 14628
tri 43313 14626 43314 14627 ne
rect 43314 14626 43553 14627
tri 43314 14625 43315 14626 ne
rect 43315 14625 43553 14626
tri 43315 14624 43316 14625 ne
rect 43316 14624 43553 14625
tri 43316 14623 43317 14624 ne
rect 43317 14623 43553 14624
tri 43317 14622 43318 14623 ne
rect 43318 14622 43553 14623
tri 43318 14621 43319 14622 ne
rect 43319 14621 43553 14622
tri 43319 14620 43320 14621 ne
rect 43320 14620 43553 14621
tri 43320 14619 43321 14620 ne
rect 43321 14619 43553 14620
tri 43553 14619 43597 14663 sw
rect 70802 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43321 14618 43322 14619 ne
rect 43322 14618 43597 14619
tri 43322 14617 43323 14618 ne
rect 43323 14617 43597 14618
tri 43323 14616 43324 14617 ne
rect 43324 14616 43597 14617
tri 43324 14615 43325 14616 ne
rect 43325 14615 43597 14616
tri 43325 14614 43326 14615 ne
rect 43326 14614 43597 14615
tri 43326 14613 43327 14614 ne
rect 43327 14613 43597 14614
tri 43327 14612 43328 14613 ne
rect 43328 14612 43597 14613
tri 43328 14611 43329 14612 ne
rect 43329 14611 43597 14612
tri 43329 14610 43330 14611 ne
rect 43330 14610 43597 14611
tri 43330 14609 43331 14610 ne
rect 43331 14609 43597 14610
tri 43331 14608 43332 14609 ne
rect 43332 14608 43597 14609
tri 43332 14607 43333 14608 ne
rect 43333 14607 43597 14608
tri 43333 14606 43334 14607 ne
rect 43334 14606 43597 14607
tri 43334 14605 43335 14606 ne
rect 43335 14605 43597 14606
tri 43335 14604 43336 14605 ne
rect 43336 14604 43597 14605
tri 43336 14603 43337 14604 ne
rect 43337 14603 43597 14604
tri 43337 14602 43338 14603 ne
rect 43338 14602 43597 14603
tri 43338 14601 43339 14602 ne
rect 43339 14601 43597 14602
tri 43339 14600 43340 14601 ne
rect 43340 14600 43597 14601
tri 43340 14599 43341 14600 ne
rect 43341 14599 43597 14600
tri 43341 14598 43342 14599 ne
rect 43342 14598 43597 14599
tri 43342 14597 43343 14598 ne
rect 43343 14597 43597 14598
tri 43343 14596 43344 14597 ne
rect 43344 14596 43597 14597
tri 43344 14595 43345 14596 ne
rect 43345 14595 43482 14596
tri 43345 14594 43346 14595 ne
rect 43346 14594 43482 14595
tri 43346 14593 43347 14594 ne
rect 43347 14593 43482 14594
tri 43347 14592 43348 14593 ne
rect 43348 14592 43482 14593
tri 43348 14591 43349 14592 ne
rect 43349 14591 43482 14592
tri 43349 14590 43350 14591 ne
rect 43350 14590 43482 14591
tri 43350 14589 43351 14590 ne
rect 43351 14589 43482 14590
tri 43351 14588 43352 14589 ne
rect 43352 14588 43482 14589
tri 43352 14587 43353 14588 ne
rect 43353 14587 43482 14588
tri 43353 14586 43354 14587 ne
rect 43354 14586 43482 14587
tri 43354 14585 43355 14586 ne
rect 43355 14585 43482 14586
tri 43355 14584 43356 14585 ne
rect 43356 14584 43482 14585
tri 43356 14583 43357 14584 ne
rect 43357 14583 43482 14584
tri 43357 14582 43358 14583 ne
rect 43358 14582 43482 14583
tri 43358 14581 43359 14582 ne
rect 43359 14581 43482 14582
tri 43359 14580 43360 14581 ne
rect 43360 14580 43482 14581
tri 43360 14579 43361 14580 ne
rect 43361 14579 43482 14580
tri 43361 14578 43362 14579 ne
rect 43362 14578 43482 14579
tri 43362 14577 43363 14578 ne
rect 43363 14577 43482 14578
tri 43363 14576 43364 14577 ne
rect 43364 14576 43482 14577
tri 43364 14575 43365 14576 ne
rect 43365 14575 43482 14576
tri 43365 14574 43366 14575 ne
rect 43366 14574 43482 14575
tri 43366 14573 43367 14574 ne
rect 43367 14573 43482 14574
tri 43367 14572 43368 14573 ne
rect 43368 14572 43482 14573
tri 43368 14571 43369 14572 ne
rect 43369 14571 43482 14572
tri 43369 14570 43370 14571 ne
rect 43370 14570 43482 14571
tri 43370 14569 43371 14570 ne
rect 43371 14569 43482 14570
tri 43371 14568 43372 14569 ne
rect 43372 14568 43482 14569
tri 43372 14567 43373 14568 ne
rect 43373 14567 43482 14568
tri 43373 14566 43374 14567 ne
rect 43374 14566 43482 14567
tri 43374 14565 43375 14566 ne
rect 43375 14565 43482 14566
tri 43375 14564 43376 14565 ne
rect 43376 14564 43482 14565
tri 43376 14563 43377 14564 ne
rect 43377 14563 43482 14564
tri 43377 14562 43378 14563 ne
rect 43378 14562 43482 14563
tri 43378 14561 43379 14562 ne
rect 43379 14561 43482 14562
tri 43379 14560 43380 14561 ne
rect 43380 14560 43482 14561
tri 43380 14559 43381 14560 ne
rect 43381 14559 43482 14560
tri 43381 14558 43382 14559 ne
rect 43382 14558 43482 14559
tri 43382 14557 43383 14558 ne
rect 43383 14557 43482 14558
tri 43383 14556 43384 14557 ne
rect 43384 14556 43482 14557
tri 43384 14555 43385 14556 ne
rect 43385 14555 43482 14556
tri 43385 14554 43386 14555 ne
rect 43386 14554 43482 14555
tri 43386 14553 43387 14554 ne
rect 43387 14553 43482 14554
tri 43387 14552 43388 14553 ne
rect 43388 14552 43482 14553
tri 43388 14551 43389 14552 ne
rect 43389 14551 43482 14552
tri 43389 14550 43390 14551 ne
rect 43390 14550 43482 14551
rect 43528 14574 43597 14596
tri 43597 14574 43642 14619 sw
rect 70802 14580 71000 14638
rect 43528 14550 43642 14574
tri 43390 14549 43391 14550 ne
rect 43391 14549 43642 14550
tri 43391 14548 43392 14549 ne
rect 43392 14548 43642 14549
tri 43392 14547 43393 14548 ne
rect 43393 14547 43642 14548
tri 43393 14546 43394 14547 ne
rect 43394 14546 43642 14547
tri 43394 14545 43395 14546 ne
rect 43395 14545 43642 14546
tri 43395 14544 43396 14545 ne
rect 43396 14544 43642 14545
tri 43396 14543 43397 14544 ne
rect 43397 14543 43642 14544
tri 43397 14542 43398 14543 ne
rect 43398 14542 43642 14543
tri 43398 14541 43399 14542 ne
rect 43399 14541 43642 14542
tri 43399 14540 43400 14541 ne
rect 43400 14540 43642 14541
tri 43400 14539 43401 14540 ne
rect 43401 14539 43642 14540
tri 43401 14538 43402 14539 ne
rect 43402 14538 43642 14539
tri 43402 14537 43403 14538 ne
rect 43403 14537 43642 14538
tri 43403 14536 43404 14537 ne
rect 43404 14536 43642 14537
tri 43404 14535 43405 14536 ne
rect 43405 14535 43642 14536
tri 43405 14534 43406 14535 ne
rect 43406 14534 43642 14535
tri 43406 14533 43407 14534 ne
rect 43407 14533 43642 14534
tri 43407 14532 43408 14533 ne
rect 43408 14532 43642 14533
tri 43408 14531 43409 14532 ne
rect 43409 14531 43642 14532
tri 43409 14530 43410 14531 ne
rect 43410 14530 43642 14531
tri 43410 14529 43411 14530 ne
rect 43411 14529 43642 14530
tri 43642 14529 43687 14574 sw
rect 70802 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
tri 43411 14528 43412 14529 ne
rect 43412 14528 43687 14529
tri 43412 14527 43413 14528 ne
rect 43413 14527 43687 14528
tri 43413 14526 43414 14527 ne
rect 43414 14526 43687 14527
tri 43414 14525 43415 14526 ne
rect 43415 14525 43687 14526
tri 43415 14524 43416 14525 ne
rect 43416 14524 43687 14525
tri 43416 14523 43417 14524 ne
rect 43417 14523 43687 14524
tri 43417 14522 43418 14523 ne
rect 43418 14522 43687 14523
tri 43418 14521 43419 14522 ne
rect 43419 14521 43687 14522
tri 43419 14520 43420 14521 ne
rect 43420 14520 43687 14521
tri 43420 14519 43421 14520 ne
rect 43421 14519 43687 14520
tri 43421 14518 43422 14519 ne
rect 43422 14518 43687 14519
tri 43422 14517 43423 14518 ne
rect 43423 14517 43687 14518
tri 43423 14516 43424 14517 ne
rect 43424 14516 43687 14517
tri 43424 14515 43425 14516 ne
rect 43425 14515 43687 14516
tri 43425 14514 43426 14515 ne
rect 43426 14514 43687 14515
tri 43426 14513 43427 14514 ne
rect 43427 14513 43687 14514
tri 43427 14512 43428 14513 ne
rect 43428 14512 43687 14513
tri 43428 14511 43429 14512 ne
rect 43429 14511 43687 14512
tri 43429 14510 43430 14511 ne
rect 43430 14510 43687 14511
tri 43430 14509 43431 14510 ne
rect 43431 14509 43687 14510
tri 43431 14508 43432 14509 ne
rect 43432 14508 43687 14509
tri 43432 14507 43433 14508 ne
rect 43433 14507 43687 14508
tri 43433 14506 43434 14507 ne
rect 43434 14506 43687 14507
tri 43434 14505 43435 14506 ne
rect 43435 14505 43687 14506
tri 43435 14504 43436 14505 ne
rect 43436 14504 43687 14505
tri 43436 14503 43437 14504 ne
rect 43437 14503 43687 14504
tri 43437 14502 43438 14503 ne
rect 43438 14502 43687 14503
tri 43438 14501 43439 14502 ne
rect 43439 14501 43687 14502
tri 43439 14500 43440 14501 ne
rect 43440 14500 43687 14501
tri 43440 14499 43441 14500 ne
rect 43441 14499 43687 14500
tri 43441 14498 43442 14499 ne
rect 43442 14498 43687 14499
tri 43442 14497 43443 14498 ne
rect 43443 14497 43687 14498
tri 43443 14496 43444 14497 ne
rect 43444 14496 43687 14497
tri 43444 14495 43445 14496 ne
rect 43445 14495 43687 14496
tri 43445 14494 43446 14495 ne
rect 43446 14494 43687 14495
tri 43446 14493 43447 14494 ne
rect 43447 14493 43687 14494
tri 43447 14492 43448 14493 ne
rect 43448 14492 43687 14493
tri 43448 14491 43449 14492 ne
rect 43449 14491 43687 14492
tri 43449 14490 43450 14491 ne
rect 43450 14490 43687 14491
tri 43450 14489 43451 14490 ne
rect 43451 14489 43687 14490
tri 43451 14488 43452 14489 ne
rect 43452 14488 43687 14489
tri 43452 14487 43453 14488 ne
rect 43453 14487 43687 14488
tri 43453 14486 43454 14487 ne
rect 43454 14486 43687 14487
tri 43454 14485 43455 14486 ne
rect 43455 14485 43687 14486
tri 43455 14484 43456 14485 ne
rect 43456 14484 43687 14485
tri 43687 14484 43732 14529 sw
tri 43456 14483 43457 14484 ne
rect 43457 14483 43732 14484
tri 43457 14482 43458 14483 ne
rect 43458 14482 43732 14483
tri 43458 14481 43459 14482 ne
rect 43459 14481 43732 14482
tri 43459 14480 43460 14481 ne
rect 43460 14480 43732 14481
tri 43460 14479 43461 14480 ne
rect 43461 14479 43732 14480
tri 43461 14478 43462 14479 ne
rect 43462 14478 43732 14479
tri 43462 14477 43463 14478 ne
rect 43463 14477 43732 14478
tri 43732 14477 43739 14484 sw
tri 43463 14462 43478 14477 ne
rect 43478 14464 43739 14477
rect 43478 14462 43614 14464
tri 43478 14417 43523 14462 ne
rect 43523 14418 43614 14462
rect 43660 14432 43739 14464
tri 43739 14432 43784 14477 sw
rect 70802 14476 71000 14534
rect 43660 14418 43784 14432
rect 43523 14417 43784 14418
tri 43523 14389 43551 14417 ne
rect 43551 14389 43784 14417
tri 43551 14388 43552 14389 ne
rect 43552 14388 43784 14389
tri 43552 14387 43553 14388 ne
rect 43553 14387 43784 14388
tri 43784 14387 43829 14432 sw
rect 70802 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
tri 43553 14386 43554 14387 ne
rect 43554 14386 43829 14387
tri 43554 14385 43555 14386 ne
rect 43555 14385 43829 14386
tri 43555 14384 43556 14385 ne
rect 43556 14384 43829 14385
tri 43556 14383 43557 14384 ne
rect 43557 14383 43829 14384
tri 43557 14382 43558 14383 ne
rect 43558 14382 43829 14383
tri 43558 14381 43559 14382 ne
rect 43559 14381 43829 14382
tri 43559 14380 43560 14381 ne
rect 43560 14380 43829 14381
tri 43560 14379 43561 14380 ne
rect 43561 14379 43829 14380
tri 43561 14378 43562 14379 ne
rect 43562 14378 43829 14379
tri 43562 14377 43563 14378 ne
rect 43563 14377 43829 14378
tri 43563 14376 43564 14377 ne
rect 43564 14376 43829 14377
tri 43564 14375 43565 14376 ne
rect 43565 14375 43829 14376
tri 43565 14374 43566 14375 ne
rect 43566 14374 43829 14375
tri 43566 14373 43567 14374 ne
rect 43567 14373 43829 14374
tri 43567 14372 43568 14373 ne
rect 43568 14372 43829 14373
tri 43568 14371 43569 14372 ne
rect 43569 14371 43829 14372
tri 43569 14370 43570 14371 ne
rect 43570 14370 43829 14371
tri 43570 14369 43571 14370 ne
rect 43571 14369 43829 14370
tri 43571 14368 43572 14369 ne
rect 43572 14368 43829 14369
tri 43572 14367 43573 14368 ne
rect 43573 14367 43829 14368
tri 43573 14366 43574 14367 ne
rect 43574 14366 43829 14367
tri 43574 14365 43575 14366 ne
rect 43575 14365 43829 14366
tri 43575 14364 43576 14365 ne
rect 43576 14364 43829 14365
tri 43576 14363 43577 14364 ne
rect 43577 14363 43829 14364
tri 43577 14362 43578 14363 ne
rect 43578 14362 43829 14363
tri 43578 14361 43579 14362 ne
rect 43579 14361 43829 14362
tri 43579 14360 43580 14361 ne
rect 43580 14360 43829 14361
tri 43580 14359 43581 14360 ne
rect 43581 14359 43829 14360
tri 43581 14358 43582 14359 ne
rect 43582 14358 43829 14359
tri 43582 14357 43583 14358 ne
rect 43583 14357 43829 14358
tri 43583 14356 43584 14357 ne
rect 43584 14356 43829 14357
tri 43584 14355 43585 14356 ne
rect 43585 14355 43829 14356
tri 43585 14354 43586 14355 ne
rect 43586 14354 43829 14355
tri 43586 14353 43587 14354 ne
rect 43587 14353 43829 14354
tri 43587 14352 43588 14353 ne
rect 43588 14352 43829 14353
tri 43588 14351 43589 14352 ne
rect 43589 14351 43829 14352
tri 43589 14350 43590 14351 ne
rect 43590 14350 43829 14351
tri 43590 14349 43591 14350 ne
rect 43591 14349 43829 14350
tri 43591 14348 43592 14349 ne
rect 43592 14348 43829 14349
tri 43592 14347 43593 14348 ne
rect 43593 14347 43829 14348
tri 43593 14346 43594 14347 ne
rect 43594 14346 43829 14347
tri 43594 14345 43595 14346 ne
rect 43595 14345 43829 14346
tri 43595 14344 43596 14345 ne
rect 43596 14344 43829 14345
tri 43596 14343 43597 14344 ne
rect 43597 14343 43829 14344
tri 43597 14342 43598 14343 ne
rect 43598 14342 43829 14343
tri 43829 14342 43874 14387 sw
rect 70802 14372 71000 14430
tri 43598 14341 43599 14342 ne
rect 43599 14341 43874 14342
tri 43599 14340 43600 14341 ne
rect 43600 14340 43874 14341
tri 43600 14339 43601 14340 ne
rect 43601 14339 43874 14340
tri 43601 14338 43602 14339 ne
rect 43602 14338 43874 14339
tri 43602 14337 43603 14338 ne
rect 43603 14337 43874 14338
tri 43603 14336 43604 14337 ne
rect 43604 14336 43874 14337
tri 43874 14336 43880 14342 sw
tri 43604 14335 43605 14336 ne
rect 43605 14335 43880 14336
tri 43605 14334 43606 14335 ne
rect 43606 14334 43880 14335
tri 43606 14333 43607 14334 ne
rect 43607 14333 43880 14334
tri 43607 14332 43608 14333 ne
rect 43608 14332 43880 14333
tri 43608 14331 43609 14332 ne
rect 43609 14331 43746 14332
tri 43609 14330 43610 14331 ne
rect 43610 14330 43746 14331
tri 43610 14329 43611 14330 ne
rect 43611 14329 43746 14330
tri 43611 14328 43612 14329 ne
rect 43612 14328 43746 14329
tri 43612 14327 43613 14328 ne
rect 43613 14327 43746 14328
tri 43613 14326 43614 14327 ne
rect 43614 14326 43746 14327
tri 43614 14325 43615 14326 ne
rect 43615 14325 43746 14326
tri 43615 14324 43616 14325 ne
rect 43616 14324 43746 14325
tri 43616 14323 43617 14324 ne
rect 43617 14323 43746 14324
tri 43617 14322 43618 14323 ne
rect 43618 14322 43746 14323
tri 43618 14321 43619 14322 ne
rect 43619 14321 43746 14322
tri 43619 14320 43620 14321 ne
rect 43620 14320 43746 14321
tri 43620 14319 43621 14320 ne
rect 43621 14319 43746 14320
tri 43621 14318 43622 14319 ne
rect 43622 14318 43746 14319
tri 43622 14317 43623 14318 ne
rect 43623 14317 43746 14318
tri 43623 14316 43624 14317 ne
rect 43624 14316 43746 14317
tri 43624 14315 43625 14316 ne
rect 43625 14315 43746 14316
tri 43625 14314 43626 14315 ne
rect 43626 14314 43746 14315
tri 43626 14313 43627 14314 ne
rect 43627 14313 43746 14314
tri 43627 14312 43628 14313 ne
rect 43628 14312 43746 14313
tri 43628 14311 43629 14312 ne
rect 43629 14311 43746 14312
tri 43629 14310 43630 14311 ne
rect 43630 14310 43746 14311
tri 43630 14309 43631 14310 ne
rect 43631 14309 43746 14310
tri 43631 14308 43632 14309 ne
rect 43632 14308 43746 14309
tri 43632 14307 43633 14308 ne
rect 43633 14307 43746 14308
tri 43633 14306 43634 14307 ne
rect 43634 14306 43746 14307
tri 43634 14305 43635 14306 ne
rect 43635 14305 43746 14306
tri 43635 14304 43636 14305 ne
rect 43636 14304 43746 14305
tri 43636 14303 43637 14304 ne
rect 43637 14303 43746 14304
tri 43637 14302 43638 14303 ne
rect 43638 14302 43746 14303
tri 43638 14301 43639 14302 ne
rect 43639 14301 43746 14302
tri 43639 14300 43640 14301 ne
rect 43640 14300 43746 14301
tri 43640 14299 43641 14300 ne
rect 43641 14299 43746 14300
tri 43641 14298 43642 14299 ne
rect 43642 14298 43746 14299
tri 43642 14297 43643 14298 ne
rect 43643 14297 43746 14298
tri 43643 14296 43644 14297 ne
rect 43644 14296 43746 14297
tri 43644 14295 43645 14296 ne
rect 43645 14295 43746 14296
tri 43645 14294 43646 14295 ne
rect 43646 14294 43746 14295
tri 43646 14293 43647 14294 ne
rect 43647 14293 43746 14294
tri 43647 14292 43648 14293 ne
rect 43648 14292 43746 14293
tri 43648 14291 43649 14292 ne
rect 43649 14291 43746 14292
tri 43649 14290 43650 14291 ne
rect 43650 14290 43746 14291
tri 43650 14289 43651 14290 ne
rect 43651 14289 43746 14290
tri 43651 14288 43652 14289 ne
rect 43652 14288 43746 14289
tri 43652 14287 43653 14288 ne
rect 43653 14287 43746 14288
tri 43653 14286 43654 14287 ne
rect 43654 14286 43746 14287
rect 43792 14291 43880 14332
tri 43880 14291 43925 14336 sw
rect 70802 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43792 14286 43925 14291
tri 43654 14285 43655 14286 ne
rect 43655 14285 43925 14286
tri 43655 14284 43656 14285 ne
rect 43656 14284 43925 14285
tri 43656 14283 43657 14284 ne
rect 43657 14283 43925 14284
tri 43657 14282 43658 14283 ne
rect 43658 14282 43925 14283
tri 43658 14281 43659 14282 ne
rect 43659 14281 43925 14282
tri 43659 14280 43660 14281 ne
rect 43660 14280 43925 14281
tri 43660 14279 43661 14280 ne
rect 43661 14279 43925 14280
tri 43661 14278 43662 14279 ne
rect 43662 14278 43925 14279
tri 43662 14277 43663 14278 ne
rect 43663 14277 43925 14278
tri 43663 14276 43664 14277 ne
rect 43664 14276 43925 14277
tri 43664 14275 43665 14276 ne
rect 43665 14275 43925 14276
tri 43665 14274 43666 14275 ne
rect 43666 14274 43925 14275
tri 43666 14273 43667 14274 ne
rect 43667 14273 43925 14274
tri 43667 14272 43668 14273 ne
rect 43668 14272 43925 14273
tri 43668 14271 43669 14272 ne
rect 43669 14271 43925 14272
tri 43669 14270 43670 14271 ne
rect 43670 14270 43925 14271
tri 43670 14269 43671 14270 ne
rect 43671 14269 43925 14270
tri 43671 14268 43672 14269 ne
rect 43672 14268 43925 14269
tri 43672 14267 43673 14268 ne
rect 43673 14267 43925 14268
tri 43673 14266 43674 14267 ne
rect 43674 14266 43925 14267
tri 43674 14265 43675 14266 ne
rect 43675 14265 43925 14266
tri 43675 14264 43676 14265 ne
rect 43676 14264 43925 14265
tri 43676 14263 43677 14264 ne
rect 43677 14263 43925 14264
tri 43677 14262 43678 14263 ne
rect 43678 14262 43925 14263
tri 43678 14261 43679 14262 ne
rect 43679 14261 43925 14262
tri 43679 14260 43680 14261 ne
rect 43680 14260 43925 14261
tri 43680 14259 43681 14260 ne
rect 43681 14259 43925 14260
tri 43681 14258 43682 14259 ne
rect 43682 14258 43925 14259
tri 43682 14257 43683 14258 ne
rect 43683 14257 43925 14258
tri 43683 14256 43684 14257 ne
rect 43684 14256 43925 14257
tri 43684 14255 43685 14256 ne
rect 43685 14255 43925 14256
tri 43685 14254 43686 14255 ne
rect 43686 14254 43925 14255
tri 43686 14253 43687 14254 ne
rect 43687 14253 43925 14254
tri 43687 14252 43688 14253 ne
rect 43688 14252 43925 14253
tri 43688 14251 43689 14252 ne
rect 43689 14251 43925 14252
tri 43689 14250 43690 14251 ne
rect 43690 14250 43925 14251
tri 43690 14249 43691 14250 ne
rect 43691 14249 43925 14250
tri 43691 14248 43692 14249 ne
rect 43692 14248 43925 14249
tri 43692 14247 43693 14248 ne
rect 43693 14247 43925 14248
tri 43693 14246 43694 14247 ne
rect 43694 14246 43925 14247
tri 43925 14246 43970 14291 sw
rect 70802 14268 71000 14326
tri 43694 14245 43695 14246 ne
rect 43695 14245 43970 14246
tri 43695 14244 43696 14245 ne
rect 43696 14244 43970 14245
tri 43696 14243 43697 14244 ne
rect 43697 14243 43970 14244
tri 43697 14242 43698 14243 ne
rect 43698 14242 43970 14243
tri 43698 14241 43699 14242 ne
rect 43699 14241 43970 14242
tri 43699 14240 43700 14241 ne
rect 43700 14240 43970 14241
tri 43700 14239 43701 14240 ne
rect 43701 14239 43970 14240
tri 43701 14238 43702 14239 ne
rect 43702 14238 43970 14239
tri 43702 14237 43703 14238 ne
rect 43703 14237 43970 14238
tri 43703 14236 43704 14237 ne
rect 43704 14236 43970 14237
tri 43704 14235 43705 14236 ne
rect 43705 14235 43970 14236
tri 43705 14234 43706 14235 ne
rect 43706 14234 43970 14235
tri 43706 14233 43707 14234 ne
rect 43707 14233 43970 14234
tri 43707 14232 43708 14233 ne
rect 43708 14232 43970 14233
tri 43708 14231 43709 14232 ne
rect 43709 14231 43970 14232
tri 43709 14230 43710 14231 ne
rect 43710 14230 43970 14231
tri 43710 14229 43711 14230 ne
rect 43711 14229 43970 14230
tri 43711 14228 43712 14229 ne
rect 43712 14228 43970 14229
tri 43712 14227 43713 14228 ne
rect 43713 14227 43970 14228
tri 43713 14226 43714 14227 ne
rect 43714 14226 43970 14227
tri 43714 14225 43715 14226 ne
rect 43715 14225 43970 14226
tri 43715 14224 43716 14225 ne
rect 43716 14224 43970 14225
tri 43716 14223 43717 14224 ne
rect 43717 14223 43970 14224
tri 43717 14222 43718 14223 ne
rect 43718 14222 43970 14223
tri 43718 14221 43719 14222 ne
rect 43719 14221 43970 14222
tri 43719 14220 43720 14221 ne
rect 43720 14220 43970 14221
tri 43720 14219 43721 14220 ne
rect 43721 14219 43970 14220
tri 43721 14218 43722 14219 ne
rect 43722 14218 43970 14219
tri 43722 14217 43723 14218 ne
rect 43723 14217 43970 14218
tri 43723 14216 43724 14217 ne
rect 43724 14216 43970 14217
tri 43724 14215 43725 14216 ne
rect 43725 14215 43970 14216
tri 43725 14214 43726 14215 ne
rect 43726 14214 43970 14215
tri 43726 14213 43727 14214 ne
rect 43727 14213 43970 14214
tri 43727 14212 43728 14213 ne
rect 43728 14212 43970 14213
tri 43728 14211 43729 14212 ne
rect 43729 14211 43970 14212
tri 43729 14210 43730 14211 ne
rect 43730 14210 43970 14211
tri 43730 14209 43731 14210 ne
rect 43731 14209 43970 14210
tri 43731 14208 43732 14209 ne
rect 43732 14208 43970 14209
tri 43732 14207 43733 14208 ne
rect 43733 14207 43970 14208
tri 43733 14206 43734 14207 ne
rect 43734 14206 43970 14207
tri 43734 14205 43735 14206 ne
rect 43735 14205 43970 14206
tri 43735 14204 43736 14205 ne
rect 43736 14204 43970 14205
tri 43736 14203 43737 14204 ne
rect 43737 14203 43970 14204
tri 43737 14202 43738 14203 ne
rect 43738 14202 43970 14203
tri 43738 14201 43739 14202 ne
rect 43739 14201 43970 14202
tri 43970 14201 44015 14246 sw
rect 70802 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43739 14163 43777 14201 ne
rect 43777 14200 44015 14201
rect 43777 14163 43878 14200
tri 43777 14118 43822 14163 ne
rect 43822 14154 43878 14163
rect 43924 14163 44015 14200
tri 44015 14163 44053 14201 sw
rect 70802 14164 71000 14222
rect 43924 14154 44053 14163
rect 43822 14118 44053 14154
tri 44053 14118 44098 14163 sw
rect 70802 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
tri 43822 14114 43826 14118 ne
rect 43826 14114 44098 14118
tri 43826 14113 43827 14114 ne
rect 43827 14113 44098 14114
tri 43827 14112 43828 14113 ne
rect 43828 14112 44098 14113
tri 43828 14111 43829 14112 ne
rect 43829 14111 44098 14112
tri 43829 14110 43830 14111 ne
rect 43830 14110 44098 14111
tri 43830 14109 43831 14110 ne
rect 43831 14109 44098 14110
tri 43831 14108 43832 14109 ne
rect 43832 14108 44098 14109
tri 43832 14107 43833 14108 ne
rect 43833 14107 44098 14108
tri 43833 14106 43834 14107 ne
rect 43834 14106 44098 14107
tri 43834 14105 43835 14106 ne
rect 43835 14105 44098 14106
tri 43835 14104 43836 14105 ne
rect 43836 14104 44098 14105
tri 43836 14103 43837 14104 ne
rect 43837 14103 44098 14104
tri 43837 14102 43838 14103 ne
rect 43838 14102 44098 14103
tri 43838 14101 43839 14102 ne
rect 43839 14101 44098 14102
tri 43839 14100 43840 14101 ne
rect 43840 14100 44098 14101
tri 43840 14099 43841 14100 ne
rect 43841 14099 44098 14100
tri 43841 14098 43842 14099 ne
rect 43842 14098 44098 14099
tri 43842 14097 43843 14098 ne
rect 43843 14097 44098 14098
tri 43843 14096 43844 14097 ne
rect 43844 14096 44098 14097
tri 43844 14095 43845 14096 ne
rect 43845 14095 44098 14096
tri 43845 14094 43846 14095 ne
rect 43846 14094 44098 14095
tri 43846 14093 43847 14094 ne
rect 43847 14093 44098 14094
tri 43847 14092 43848 14093 ne
rect 43848 14092 44098 14093
tri 43848 14091 43849 14092 ne
rect 43849 14091 44098 14092
tri 43849 14090 43850 14091 ne
rect 43850 14090 44098 14091
tri 43850 14089 43851 14090 ne
rect 43851 14089 44098 14090
tri 43851 14088 43852 14089 ne
rect 43852 14088 44098 14089
tri 43852 14087 43853 14088 ne
rect 43853 14087 44098 14088
tri 43853 14086 43854 14087 ne
rect 43854 14086 44098 14087
tri 43854 14085 43855 14086 ne
rect 43855 14085 44098 14086
tri 43855 14084 43856 14085 ne
rect 43856 14084 44098 14085
tri 43856 14083 43857 14084 ne
rect 43857 14083 44098 14084
tri 43857 14082 43858 14083 ne
rect 43858 14082 44098 14083
tri 43858 14081 43859 14082 ne
rect 43859 14081 44098 14082
tri 43859 14080 43860 14081 ne
rect 43860 14080 44098 14081
tri 43860 14079 43861 14080 ne
rect 43861 14079 44098 14080
tri 43861 14078 43862 14079 ne
rect 43862 14078 44098 14079
tri 43862 14077 43863 14078 ne
rect 43863 14077 44098 14078
tri 43863 14076 43864 14077 ne
rect 43864 14076 44098 14077
tri 43864 14075 43865 14076 ne
rect 43865 14075 44098 14076
tri 43865 14074 43866 14075 ne
rect 43866 14074 44098 14075
tri 43866 14073 43867 14074 ne
rect 43867 14073 44098 14074
tri 44098 14073 44143 14118 sw
tri 43867 14072 43868 14073 ne
rect 43868 14072 44143 14073
tri 43868 14071 43869 14072 ne
rect 43869 14071 44143 14072
tri 43869 14070 43870 14071 ne
rect 43870 14070 44143 14071
tri 43870 14069 43871 14070 ne
rect 43871 14069 44143 14070
tri 43871 14068 43872 14069 ne
rect 43872 14068 44143 14069
tri 43872 14067 43873 14068 ne
rect 43873 14067 44010 14068
tri 43873 14066 43874 14067 ne
rect 43874 14066 44010 14067
tri 43874 14065 43875 14066 ne
rect 43875 14065 44010 14066
tri 43875 14064 43876 14065 ne
rect 43876 14064 44010 14065
tri 43876 14063 43877 14064 ne
rect 43877 14063 44010 14064
tri 43877 14062 43878 14063 ne
rect 43878 14062 44010 14063
tri 43878 14061 43879 14062 ne
rect 43879 14061 44010 14062
tri 43879 14060 43880 14061 ne
rect 43880 14060 44010 14061
tri 43880 14059 43881 14060 ne
rect 43881 14059 44010 14060
tri 43881 14058 43882 14059 ne
rect 43882 14058 44010 14059
tri 43882 14057 43883 14058 ne
rect 43883 14057 44010 14058
tri 43883 14056 43884 14057 ne
rect 43884 14056 44010 14057
tri 43884 14055 43885 14056 ne
rect 43885 14055 44010 14056
tri 43885 14054 43886 14055 ne
rect 43886 14054 44010 14055
tri 43886 14053 43887 14054 ne
rect 43887 14053 44010 14054
tri 43887 14052 43888 14053 ne
rect 43888 14052 44010 14053
tri 43888 14051 43889 14052 ne
rect 43889 14051 44010 14052
tri 43889 14050 43890 14051 ne
rect 43890 14050 44010 14051
tri 43890 14049 43891 14050 ne
rect 43891 14049 44010 14050
tri 43891 14048 43892 14049 ne
rect 43892 14048 44010 14049
tri 43892 14047 43893 14048 ne
rect 43893 14047 44010 14048
tri 43893 14046 43894 14047 ne
rect 43894 14046 44010 14047
tri 43894 14045 43895 14046 ne
rect 43895 14045 44010 14046
tri 43895 14044 43896 14045 ne
rect 43896 14044 44010 14045
tri 43896 14043 43897 14044 ne
rect 43897 14043 44010 14044
tri 43897 14042 43898 14043 ne
rect 43898 14042 44010 14043
tri 43898 14041 43899 14042 ne
rect 43899 14041 44010 14042
tri 43899 14040 43900 14041 ne
rect 43900 14040 44010 14041
tri 43900 14039 43901 14040 ne
rect 43901 14039 44010 14040
tri 43901 14038 43902 14039 ne
rect 43902 14038 44010 14039
tri 43902 14037 43903 14038 ne
rect 43903 14037 44010 14038
tri 43903 14036 43904 14037 ne
rect 43904 14036 44010 14037
tri 43904 14035 43905 14036 ne
rect 43905 14035 44010 14036
tri 43905 14034 43906 14035 ne
rect 43906 14034 44010 14035
tri 43906 14033 43907 14034 ne
rect 43907 14033 44010 14034
tri 43907 14032 43908 14033 ne
rect 43908 14032 44010 14033
tri 43908 14031 43909 14032 ne
rect 43909 14031 44010 14032
tri 43909 14030 43910 14031 ne
rect 43910 14030 44010 14031
tri 43910 14029 43911 14030 ne
rect 43911 14029 44010 14030
tri 43911 14028 43912 14029 ne
rect 43912 14028 44010 14029
tri 43912 14027 43913 14028 ne
rect 43913 14027 44010 14028
tri 43913 14026 43914 14027 ne
rect 43914 14026 44010 14027
tri 43914 14025 43915 14026 ne
rect 43915 14025 44010 14026
tri 43915 14024 43916 14025 ne
rect 43916 14024 44010 14025
tri 43916 14023 43917 14024 ne
rect 43917 14023 44010 14024
tri 43917 14022 43918 14023 ne
rect 43918 14022 44010 14023
rect 44056 14028 44143 14068
tri 44143 14028 44188 14073 sw
rect 70802 14060 71000 14118
rect 44056 14022 44188 14028
tri 43918 14021 43919 14022 ne
rect 43919 14021 44188 14022
tri 43919 14020 43920 14021 ne
rect 43920 14020 44188 14021
tri 43920 14019 43921 14020 ne
rect 43921 14019 44188 14020
tri 43921 14018 43922 14019 ne
rect 43922 14018 44188 14019
tri 43922 14017 43923 14018 ne
rect 43923 14017 44188 14018
tri 43923 14016 43924 14017 ne
rect 43924 14016 44188 14017
tri 43924 14015 43925 14016 ne
rect 43925 14015 44188 14016
tri 44188 14015 44201 14028 sw
tri 43925 14014 43926 14015 ne
rect 43926 14014 44201 14015
tri 43926 14013 43927 14014 ne
rect 43927 14013 44201 14014
tri 43927 14012 43928 14013 ne
rect 43928 14012 44201 14013
tri 43928 14011 43929 14012 ne
rect 43929 14011 44201 14012
tri 43929 14010 43930 14011 ne
rect 43930 14010 44201 14011
tri 43930 14009 43931 14010 ne
rect 43931 14009 44201 14010
tri 43931 14008 43932 14009 ne
rect 43932 14008 44201 14009
tri 43932 14007 43933 14008 ne
rect 43933 14007 44201 14008
tri 43933 14006 43934 14007 ne
rect 43934 14006 44201 14007
tri 43934 14005 43935 14006 ne
rect 43935 14005 44201 14006
tri 43935 14004 43936 14005 ne
rect 43936 14004 44201 14005
tri 43936 14003 43937 14004 ne
rect 43937 14003 44201 14004
tri 43937 14002 43938 14003 ne
rect 43938 14002 44201 14003
tri 43938 14001 43939 14002 ne
rect 43939 14001 44201 14002
tri 43939 14000 43940 14001 ne
rect 43940 14000 44201 14001
tri 43940 13999 43941 14000 ne
rect 43941 13999 44201 14000
tri 43941 13998 43942 13999 ne
rect 43942 13998 44201 13999
tri 43942 13997 43943 13998 ne
rect 43943 13997 44201 13998
tri 43943 13996 43944 13997 ne
rect 43944 13996 44201 13997
tri 43944 13995 43945 13996 ne
rect 43945 13995 44201 13996
tri 43945 13994 43946 13995 ne
rect 43946 13994 44201 13995
tri 43946 13993 43947 13994 ne
rect 43947 13993 44201 13994
tri 43947 13992 43948 13993 ne
rect 43948 13992 44201 13993
tri 43948 13991 43949 13992 ne
rect 43949 13991 44201 13992
tri 43949 13990 43950 13991 ne
rect 43950 13990 44201 13991
tri 43950 13989 43951 13990 ne
rect 43951 13989 44201 13990
tri 43951 13988 43952 13989 ne
rect 43952 13988 44201 13989
tri 43952 13987 43953 13988 ne
rect 43953 13987 44201 13988
tri 43953 13986 43954 13987 ne
rect 43954 13986 44201 13987
tri 43954 13985 43955 13986 ne
rect 43955 13985 44201 13986
tri 43955 13984 43956 13985 ne
rect 43956 13984 44201 13985
tri 43956 13983 43957 13984 ne
rect 43957 13983 44201 13984
tri 43957 13982 43958 13983 ne
rect 43958 13982 44201 13983
tri 43958 13981 43959 13982 ne
rect 43959 13981 44201 13982
tri 43959 13980 43960 13981 ne
rect 43960 13980 44201 13981
tri 43960 13979 43961 13980 ne
rect 43961 13979 44201 13980
tri 43961 13978 43962 13979 ne
rect 43962 13978 44201 13979
tri 43962 13977 43963 13978 ne
rect 43963 13977 44201 13978
tri 43963 13976 43964 13977 ne
rect 43964 13976 44201 13977
tri 43964 13975 43965 13976 ne
rect 43965 13975 44201 13976
tri 43965 13974 43966 13975 ne
rect 43966 13974 44201 13975
tri 43966 13973 43967 13974 ne
rect 43967 13973 44201 13974
tri 43967 13972 43968 13973 ne
rect 43968 13972 44201 13973
tri 43968 13971 43969 13972 ne
rect 43969 13971 44201 13972
tri 43969 13970 43970 13971 ne
rect 43970 13970 44201 13971
tri 44201 13970 44246 14015 sw
rect 70802 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
tri 43970 13969 43971 13970 ne
rect 43971 13969 44246 13970
tri 43971 13968 43972 13969 ne
rect 43972 13968 44246 13969
tri 43972 13967 43973 13968 ne
rect 43973 13967 44246 13968
tri 43973 13966 43974 13967 ne
rect 43974 13966 44246 13967
tri 43974 13965 43975 13966 ne
rect 43975 13965 44246 13966
tri 43975 13964 43976 13965 ne
rect 43976 13964 44246 13965
tri 43976 13963 43977 13964 ne
rect 43977 13963 44246 13964
tri 43977 13962 43978 13963 ne
rect 43978 13962 44246 13963
tri 43978 13961 43979 13962 ne
rect 43979 13961 44246 13962
tri 43979 13960 43980 13961 ne
rect 43980 13960 44246 13961
tri 43980 13959 43981 13960 ne
rect 43981 13959 44246 13960
tri 43981 13958 43982 13959 ne
rect 43982 13958 44246 13959
tri 43982 13957 43983 13958 ne
rect 43983 13957 44246 13958
tri 43983 13956 43984 13957 ne
rect 43984 13956 44246 13957
tri 43984 13955 43985 13956 ne
rect 43985 13955 44246 13956
tri 43985 13954 43986 13955 ne
rect 43986 13954 44246 13955
tri 43986 13953 43987 13954 ne
rect 43987 13953 44246 13954
tri 43987 13952 43988 13953 ne
rect 43988 13952 44246 13953
tri 43988 13951 43989 13952 ne
rect 43989 13951 44246 13952
tri 43989 13950 43990 13951 ne
rect 43990 13950 44246 13951
tri 43990 13949 43991 13950 ne
rect 43991 13949 44246 13950
tri 43991 13948 43992 13949 ne
rect 43992 13948 44246 13949
tri 43992 13947 43993 13948 ne
rect 43993 13947 44246 13948
tri 43993 13946 43994 13947 ne
rect 43994 13946 44246 13947
tri 43994 13945 43995 13946 ne
rect 43995 13945 44246 13946
tri 43995 13944 43996 13945 ne
rect 43996 13944 44246 13945
tri 43996 13943 43997 13944 ne
rect 43997 13943 44246 13944
tri 43997 13942 43998 13943 ne
rect 43998 13942 44246 13943
tri 43998 13941 43999 13942 ne
rect 43999 13941 44246 13942
tri 43999 13940 44000 13941 ne
rect 44000 13940 44246 13941
tri 44000 13939 44001 13940 ne
rect 44001 13939 44246 13940
tri 44001 13938 44002 13939 ne
rect 44002 13938 44246 13939
tri 44002 13937 44003 13938 ne
rect 44003 13937 44246 13938
tri 44003 13936 44004 13937 ne
rect 44004 13936 44246 13937
tri 44004 13935 44005 13936 ne
rect 44005 13935 44142 13936
tri 44005 13934 44006 13935 ne
rect 44006 13934 44142 13935
tri 44006 13933 44007 13934 ne
rect 44007 13933 44142 13934
tri 44007 13932 44008 13933 ne
rect 44008 13932 44142 13933
tri 44008 13931 44009 13932 ne
rect 44009 13931 44142 13932
tri 44009 13930 44010 13931 ne
rect 44010 13930 44142 13931
tri 44010 13929 44011 13930 ne
rect 44011 13929 44142 13930
tri 44011 13928 44012 13929 ne
rect 44012 13928 44142 13929
tri 44012 13927 44013 13928 ne
rect 44013 13927 44142 13928
tri 44013 13926 44014 13927 ne
rect 44014 13926 44142 13927
tri 44014 13925 44015 13926 ne
rect 44015 13925 44142 13926
tri 44015 13880 44060 13925 ne
rect 44060 13890 44142 13925
rect 44188 13925 44246 13936
tri 44246 13925 44291 13970 sw
rect 70802 13956 71000 14014
rect 44188 13890 44291 13925
rect 44060 13880 44291 13890
tri 44291 13880 44336 13925 sw
rect 70802 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
tri 44060 13842 44098 13880 ne
rect 44098 13842 44336 13880
tri 44336 13842 44374 13880 sw
rect 70802 13852 71000 13910
tri 44098 13840 44100 13842 ne
rect 44100 13840 44374 13842
tri 44100 13839 44101 13840 ne
rect 44101 13839 44374 13840
tri 44101 13838 44102 13839 ne
rect 44102 13838 44374 13839
tri 44102 13837 44103 13838 ne
rect 44103 13837 44374 13838
tri 44103 13836 44104 13837 ne
rect 44104 13836 44374 13837
tri 44104 13835 44105 13836 ne
rect 44105 13835 44374 13836
tri 44105 13834 44106 13835 ne
rect 44106 13834 44374 13835
tri 44106 13833 44107 13834 ne
rect 44107 13833 44374 13834
tri 44107 13832 44108 13833 ne
rect 44108 13832 44374 13833
tri 44108 13831 44109 13832 ne
rect 44109 13831 44374 13832
tri 44109 13830 44110 13831 ne
rect 44110 13830 44374 13831
tri 44110 13829 44111 13830 ne
rect 44111 13829 44374 13830
tri 44111 13828 44112 13829 ne
rect 44112 13828 44374 13829
tri 44112 13827 44113 13828 ne
rect 44113 13827 44374 13828
tri 44113 13826 44114 13827 ne
rect 44114 13826 44374 13827
tri 44114 13825 44115 13826 ne
rect 44115 13825 44374 13826
tri 44115 13824 44116 13825 ne
rect 44116 13824 44374 13825
tri 44116 13823 44117 13824 ne
rect 44117 13823 44374 13824
tri 44117 13822 44118 13823 ne
rect 44118 13822 44374 13823
tri 44118 13821 44119 13822 ne
rect 44119 13821 44374 13822
tri 44119 13820 44120 13821 ne
rect 44120 13820 44374 13821
tri 44120 13819 44121 13820 ne
rect 44121 13819 44374 13820
tri 44121 13818 44122 13819 ne
rect 44122 13818 44374 13819
tri 44122 13817 44123 13818 ne
rect 44123 13817 44374 13818
tri 44123 13816 44124 13817 ne
rect 44124 13816 44374 13817
tri 44124 13815 44125 13816 ne
rect 44125 13815 44374 13816
tri 44125 13814 44126 13815 ne
rect 44126 13814 44374 13815
tri 44126 13813 44127 13814 ne
rect 44127 13813 44374 13814
tri 44127 13812 44128 13813 ne
rect 44128 13812 44374 13813
tri 44128 13811 44129 13812 ne
rect 44129 13811 44374 13812
tri 44129 13810 44130 13811 ne
rect 44130 13810 44374 13811
tri 44130 13809 44131 13810 ne
rect 44131 13809 44374 13810
tri 44131 13808 44132 13809 ne
rect 44132 13808 44374 13809
tri 44132 13807 44133 13808 ne
rect 44133 13807 44374 13808
tri 44133 13806 44134 13807 ne
rect 44134 13806 44374 13807
tri 44134 13805 44135 13806 ne
rect 44135 13805 44374 13806
tri 44135 13804 44136 13805 ne
rect 44136 13804 44374 13805
tri 44136 13803 44137 13804 ne
rect 44137 13803 44274 13804
tri 44137 13802 44138 13803 ne
rect 44138 13802 44274 13803
tri 44138 13801 44139 13802 ne
rect 44139 13801 44274 13802
tri 44139 13800 44140 13801 ne
rect 44140 13800 44274 13801
tri 44140 13799 44141 13800 ne
rect 44141 13799 44274 13800
tri 44141 13798 44142 13799 ne
rect 44142 13798 44274 13799
tri 44142 13797 44143 13798 ne
rect 44143 13797 44274 13798
tri 44143 13796 44144 13797 ne
rect 44144 13796 44274 13797
tri 44144 13795 44145 13796 ne
rect 44145 13795 44274 13796
tri 44145 13794 44146 13795 ne
rect 44146 13794 44274 13795
tri 44146 13793 44147 13794 ne
rect 44147 13793 44274 13794
tri 44147 13792 44148 13793 ne
rect 44148 13792 44274 13793
tri 44148 13791 44149 13792 ne
rect 44149 13791 44274 13792
tri 44149 13790 44150 13791 ne
rect 44150 13790 44274 13791
tri 44150 13789 44151 13790 ne
rect 44151 13789 44274 13790
tri 44151 13788 44152 13789 ne
rect 44152 13788 44274 13789
tri 44152 13787 44153 13788 ne
rect 44153 13787 44274 13788
tri 44153 13786 44154 13787 ne
rect 44154 13786 44274 13787
tri 44154 13785 44155 13786 ne
rect 44155 13785 44274 13786
tri 44155 13784 44156 13785 ne
rect 44156 13784 44274 13785
tri 44156 13783 44157 13784 ne
rect 44157 13783 44274 13784
tri 44157 13782 44158 13783 ne
rect 44158 13782 44274 13783
tri 44158 13781 44159 13782 ne
rect 44159 13781 44274 13782
tri 44159 13780 44160 13781 ne
rect 44160 13780 44274 13781
tri 44160 13779 44161 13780 ne
rect 44161 13779 44274 13780
tri 44161 13778 44162 13779 ne
rect 44162 13778 44274 13779
tri 44162 13777 44163 13778 ne
rect 44163 13777 44274 13778
tri 44163 13776 44164 13777 ne
rect 44164 13776 44274 13777
tri 44164 13775 44165 13776 ne
rect 44165 13775 44274 13776
tri 44165 13774 44166 13775 ne
rect 44166 13774 44274 13775
tri 44166 13773 44167 13774 ne
rect 44167 13773 44274 13774
tri 44167 13772 44168 13773 ne
rect 44168 13772 44274 13773
tri 44168 13771 44169 13772 ne
rect 44169 13771 44274 13772
tri 44169 13770 44170 13771 ne
rect 44170 13770 44274 13771
tri 44170 13769 44171 13770 ne
rect 44171 13769 44274 13770
tri 44171 13768 44172 13769 ne
rect 44172 13768 44274 13769
tri 44172 13767 44173 13768 ne
rect 44173 13767 44274 13768
tri 44173 13766 44174 13767 ne
rect 44174 13766 44274 13767
tri 44174 13765 44175 13766 ne
rect 44175 13765 44274 13766
tri 44175 13764 44176 13765 ne
rect 44176 13764 44274 13765
tri 44176 13763 44177 13764 ne
rect 44177 13763 44274 13764
tri 44177 13762 44178 13763 ne
rect 44178 13762 44274 13763
tri 44178 13761 44179 13762 ne
rect 44179 13761 44274 13762
tri 44179 13760 44180 13761 ne
rect 44180 13760 44274 13761
tri 44180 13759 44181 13760 ne
rect 44181 13759 44274 13760
tri 44181 13758 44182 13759 ne
rect 44182 13758 44274 13759
rect 44320 13797 44374 13804
tri 44374 13797 44419 13842 sw
rect 70802 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 44320 13758 44419 13797
tri 44182 13757 44183 13758 ne
rect 44183 13757 44419 13758
tri 44183 13756 44184 13757 ne
rect 44184 13756 44419 13757
tri 44184 13755 44185 13756 ne
rect 44185 13755 44419 13756
tri 44185 13754 44186 13755 ne
rect 44186 13754 44419 13755
tri 44186 13753 44187 13754 ne
rect 44187 13753 44419 13754
tri 44187 13752 44188 13753 ne
rect 44188 13752 44419 13753
tri 44419 13752 44464 13797 sw
tri 44188 13751 44189 13752 ne
rect 44189 13751 44464 13752
tri 44189 13750 44190 13751 ne
rect 44190 13750 44464 13751
tri 44190 13749 44191 13750 ne
rect 44191 13749 44464 13750
tri 44191 13748 44192 13749 ne
rect 44192 13748 44464 13749
tri 44192 13747 44193 13748 ne
rect 44193 13747 44464 13748
tri 44193 13746 44194 13747 ne
rect 44194 13746 44464 13747
tri 44194 13745 44195 13746 ne
rect 44195 13745 44464 13746
tri 44195 13744 44196 13745 ne
rect 44196 13744 44464 13745
tri 44196 13743 44197 13744 ne
rect 44197 13743 44464 13744
tri 44197 13742 44198 13743 ne
rect 44198 13742 44464 13743
tri 44198 13741 44199 13742 ne
rect 44199 13741 44464 13742
tri 44199 13740 44200 13741 ne
rect 44200 13740 44464 13741
tri 44200 13739 44201 13740 ne
rect 44201 13739 44464 13740
tri 44201 13738 44202 13739 ne
rect 44202 13738 44464 13739
tri 44202 13737 44203 13738 ne
rect 44203 13737 44464 13738
tri 44203 13736 44204 13737 ne
rect 44204 13736 44464 13737
tri 44204 13735 44205 13736 ne
rect 44205 13735 44464 13736
tri 44205 13734 44206 13735 ne
rect 44206 13734 44464 13735
tri 44206 13733 44207 13734 ne
rect 44207 13733 44464 13734
tri 44207 13732 44208 13733 ne
rect 44208 13732 44464 13733
tri 44208 13731 44209 13732 ne
rect 44209 13731 44464 13732
tri 44209 13730 44210 13731 ne
rect 44210 13730 44464 13731
tri 44210 13729 44211 13730 ne
rect 44211 13729 44464 13730
tri 44211 13728 44212 13729 ne
rect 44212 13728 44464 13729
tri 44212 13727 44213 13728 ne
rect 44213 13727 44464 13728
tri 44213 13726 44214 13727 ne
rect 44214 13726 44464 13727
tri 44214 13725 44215 13726 ne
rect 44215 13725 44464 13726
tri 44215 13724 44216 13725 ne
rect 44216 13724 44464 13725
tri 44216 13723 44217 13724 ne
rect 44217 13723 44464 13724
tri 44217 13722 44218 13723 ne
rect 44218 13722 44464 13723
tri 44218 13721 44219 13722 ne
rect 44219 13721 44464 13722
tri 44219 13720 44220 13721 ne
rect 44220 13720 44464 13721
tri 44220 13719 44221 13720 ne
rect 44221 13719 44464 13720
tri 44221 13718 44222 13719 ne
rect 44222 13718 44464 13719
tri 44222 13717 44223 13718 ne
rect 44223 13717 44464 13718
tri 44223 13716 44224 13717 ne
rect 44224 13716 44464 13717
tri 44224 13715 44225 13716 ne
rect 44225 13715 44464 13716
tri 44225 13714 44226 13715 ne
rect 44226 13714 44464 13715
tri 44226 13713 44227 13714 ne
rect 44227 13713 44464 13714
tri 44227 13712 44228 13713 ne
rect 44228 13712 44464 13713
tri 44228 13711 44229 13712 ne
rect 44229 13711 44464 13712
tri 44229 13710 44230 13711 ne
rect 44230 13710 44464 13711
tri 44230 13709 44231 13710 ne
rect 44231 13709 44464 13710
tri 44231 13708 44232 13709 ne
rect 44232 13708 44464 13709
tri 44232 13707 44233 13708 ne
rect 44233 13707 44464 13708
tri 44464 13707 44509 13752 sw
rect 70802 13748 71000 13806
tri 44233 13706 44234 13707 ne
rect 44234 13706 44509 13707
tri 44234 13705 44235 13706 ne
rect 44235 13705 44509 13706
tri 44235 13704 44236 13705 ne
rect 44236 13704 44509 13705
tri 44236 13703 44237 13704 ne
rect 44237 13703 44509 13704
tri 44237 13702 44238 13703 ne
rect 44238 13702 44509 13703
tri 44238 13701 44239 13702 ne
rect 44239 13701 44509 13702
tri 44239 13700 44240 13701 ne
rect 44240 13700 44509 13701
tri 44240 13699 44241 13700 ne
rect 44241 13699 44509 13700
tri 44241 13698 44242 13699 ne
rect 44242 13698 44509 13699
tri 44242 13697 44243 13698 ne
rect 44243 13697 44509 13698
tri 44243 13696 44244 13697 ne
rect 44244 13696 44509 13697
tri 44244 13695 44245 13696 ne
rect 44245 13695 44509 13696
tri 44245 13694 44246 13695 ne
rect 44246 13694 44509 13695
tri 44509 13694 44522 13707 sw
rect 70802 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
tri 44246 13693 44247 13694 ne
rect 44247 13693 44522 13694
tri 44247 13692 44248 13693 ne
rect 44248 13692 44522 13693
tri 44248 13691 44249 13692 ne
rect 44249 13691 44522 13692
tri 44249 13690 44250 13691 ne
rect 44250 13690 44522 13691
tri 44250 13689 44251 13690 ne
rect 44251 13689 44522 13690
tri 44251 13688 44252 13689 ne
rect 44252 13688 44522 13689
tri 44252 13687 44253 13688 ne
rect 44253 13687 44522 13688
tri 44253 13686 44254 13687 ne
rect 44254 13686 44522 13687
tri 44254 13685 44255 13686 ne
rect 44255 13685 44522 13686
tri 44255 13684 44256 13685 ne
rect 44256 13684 44522 13685
tri 44256 13683 44257 13684 ne
rect 44257 13683 44522 13684
tri 44257 13682 44258 13683 ne
rect 44258 13682 44522 13683
tri 44258 13681 44259 13682 ne
rect 44259 13681 44522 13682
tri 44259 13680 44260 13681 ne
rect 44260 13680 44522 13681
tri 44260 13679 44261 13680 ne
rect 44261 13679 44522 13680
tri 44261 13678 44262 13679 ne
rect 44262 13678 44522 13679
tri 44262 13677 44263 13678 ne
rect 44263 13677 44522 13678
tri 44263 13676 44264 13677 ne
rect 44264 13676 44522 13677
tri 44264 13675 44265 13676 ne
rect 44265 13675 44522 13676
tri 44265 13674 44266 13675 ne
rect 44266 13674 44522 13675
tri 44266 13673 44267 13674 ne
rect 44267 13673 44522 13674
tri 44267 13672 44268 13673 ne
rect 44268 13672 44522 13673
tri 44268 13671 44269 13672 ne
rect 44269 13671 44406 13672
tri 44269 13670 44270 13671 ne
rect 44270 13670 44406 13671
tri 44270 13669 44271 13670 ne
rect 44271 13669 44406 13670
tri 44271 13668 44272 13669 ne
rect 44272 13668 44406 13669
tri 44272 13667 44273 13668 ne
rect 44273 13667 44406 13668
tri 44273 13666 44274 13667 ne
rect 44274 13666 44406 13667
tri 44274 13665 44275 13666 ne
rect 44275 13665 44406 13666
tri 44275 13664 44276 13665 ne
rect 44276 13664 44406 13665
tri 44276 13663 44277 13664 ne
rect 44277 13663 44406 13664
tri 44277 13662 44278 13663 ne
rect 44278 13662 44406 13663
tri 44278 13661 44279 13662 ne
rect 44279 13661 44406 13662
tri 44279 13660 44280 13661 ne
rect 44280 13660 44406 13661
tri 44280 13659 44281 13660 ne
rect 44281 13659 44406 13660
tri 44281 13658 44282 13659 ne
rect 44282 13658 44406 13659
tri 44282 13657 44283 13658 ne
rect 44283 13657 44406 13658
tri 44283 13656 44284 13657 ne
rect 44284 13656 44406 13657
tri 44284 13655 44285 13656 ne
rect 44285 13655 44406 13656
tri 44285 13654 44286 13655 ne
rect 44286 13654 44406 13655
tri 44286 13653 44287 13654 ne
rect 44287 13653 44406 13654
tri 44287 13652 44288 13653 ne
rect 44288 13652 44406 13653
tri 44288 13651 44289 13652 ne
rect 44289 13651 44406 13652
tri 44289 13650 44290 13651 ne
rect 44290 13650 44406 13651
tri 44290 13649 44291 13650 ne
rect 44291 13649 44406 13650
tri 44291 13604 44336 13649 ne
rect 44336 13626 44406 13649
rect 44452 13649 44522 13672
tri 44522 13649 44567 13694 sw
rect 44452 13626 44567 13649
rect 44336 13604 44567 13626
tri 44567 13604 44612 13649 sw
rect 70802 13644 71000 13702
tri 44336 13565 44375 13604 ne
rect 44375 13565 44612 13604
tri 44375 13564 44376 13565 ne
rect 44376 13564 44612 13565
tri 44376 13563 44377 13564 ne
rect 44377 13563 44612 13564
tri 44377 13562 44378 13563 ne
rect 44378 13562 44612 13563
tri 44378 13561 44379 13562 ne
rect 44379 13561 44612 13562
tri 44379 13560 44380 13561 ne
rect 44380 13560 44612 13561
tri 44380 13559 44381 13560 ne
rect 44381 13559 44612 13560
tri 44612 13559 44657 13604 sw
rect 70802 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
tri 44381 13558 44382 13559 ne
rect 44382 13558 44657 13559
tri 44382 13557 44383 13558 ne
rect 44383 13557 44657 13558
tri 44383 13556 44384 13557 ne
rect 44384 13556 44657 13557
tri 44384 13555 44385 13556 ne
rect 44385 13555 44657 13556
tri 44385 13554 44386 13555 ne
rect 44386 13554 44657 13555
tri 44386 13553 44387 13554 ne
rect 44387 13553 44657 13554
tri 44387 13552 44388 13553 ne
rect 44388 13552 44657 13553
tri 44388 13551 44389 13552 ne
rect 44389 13551 44657 13552
tri 44389 13550 44390 13551 ne
rect 44390 13550 44657 13551
tri 44390 13549 44391 13550 ne
rect 44391 13549 44657 13550
tri 44391 13548 44392 13549 ne
rect 44392 13548 44657 13549
tri 44392 13547 44393 13548 ne
rect 44393 13547 44657 13548
tri 44393 13546 44394 13547 ne
rect 44394 13546 44657 13547
tri 44394 13545 44395 13546 ne
rect 44395 13545 44657 13546
tri 44395 13544 44396 13545 ne
rect 44396 13544 44657 13545
tri 44396 13543 44397 13544 ne
rect 44397 13543 44657 13544
tri 44397 13542 44398 13543 ne
rect 44398 13542 44657 13543
tri 44398 13541 44399 13542 ne
rect 44399 13541 44657 13542
tri 44399 13540 44400 13541 ne
rect 44400 13540 44657 13541
tri 44400 13539 44401 13540 ne
rect 44401 13539 44538 13540
tri 44401 13538 44402 13539 ne
rect 44402 13538 44538 13539
tri 44402 13537 44403 13538 ne
rect 44403 13537 44538 13538
tri 44403 13536 44404 13537 ne
rect 44404 13536 44538 13537
tri 44404 13535 44405 13536 ne
rect 44405 13535 44538 13536
tri 44405 13534 44406 13535 ne
rect 44406 13534 44538 13535
tri 44406 13533 44407 13534 ne
rect 44407 13533 44538 13534
tri 44407 13532 44408 13533 ne
rect 44408 13532 44538 13533
tri 44408 13531 44409 13532 ne
rect 44409 13531 44538 13532
tri 44409 13530 44410 13531 ne
rect 44410 13530 44538 13531
tri 44410 13529 44411 13530 ne
rect 44411 13529 44538 13530
tri 44411 13528 44412 13529 ne
rect 44412 13528 44538 13529
tri 44412 13527 44413 13528 ne
rect 44413 13527 44538 13528
tri 44413 13526 44414 13527 ne
rect 44414 13526 44538 13527
tri 44414 13525 44415 13526 ne
rect 44415 13525 44538 13526
tri 44415 13524 44416 13525 ne
rect 44416 13524 44538 13525
tri 44416 13523 44417 13524 ne
rect 44417 13523 44538 13524
tri 44417 13522 44418 13523 ne
rect 44418 13522 44538 13523
tri 44418 13521 44419 13522 ne
rect 44419 13521 44538 13522
tri 44419 13520 44420 13521 ne
rect 44420 13520 44538 13521
tri 44420 13519 44421 13520 ne
rect 44421 13519 44538 13520
tri 44421 13518 44422 13519 ne
rect 44422 13518 44538 13519
tri 44422 13517 44423 13518 ne
rect 44423 13517 44538 13518
tri 44423 13516 44424 13517 ne
rect 44424 13516 44538 13517
tri 44424 13515 44425 13516 ne
rect 44425 13515 44538 13516
tri 44425 13514 44426 13515 ne
rect 44426 13514 44538 13515
tri 44426 13513 44427 13514 ne
rect 44427 13513 44538 13514
tri 44427 13512 44428 13513 ne
rect 44428 13512 44538 13513
tri 44428 13511 44429 13512 ne
rect 44429 13511 44538 13512
tri 44429 13510 44430 13511 ne
rect 44430 13510 44538 13511
tri 44430 13509 44431 13510 ne
rect 44431 13509 44538 13510
tri 44431 13508 44432 13509 ne
rect 44432 13508 44538 13509
tri 44432 13507 44433 13508 ne
rect 44433 13507 44538 13508
tri 44433 13506 44434 13507 ne
rect 44434 13506 44538 13507
tri 44434 13505 44435 13506 ne
rect 44435 13505 44538 13506
tri 44435 13504 44436 13505 ne
rect 44436 13504 44538 13505
tri 44436 13503 44437 13504 ne
rect 44437 13503 44538 13504
tri 44437 13502 44438 13503 ne
rect 44438 13502 44538 13503
tri 44438 13501 44439 13502 ne
rect 44439 13501 44538 13502
tri 44439 13500 44440 13501 ne
rect 44440 13500 44538 13501
tri 44440 13499 44441 13500 ne
rect 44441 13499 44538 13500
tri 44441 13498 44442 13499 ne
rect 44442 13498 44538 13499
tri 44442 13497 44443 13498 ne
rect 44443 13497 44538 13498
tri 44443 13496 44444 13497 ne
rect 44444 13496 44538 13497
tri 44444 13495 44445 13496 ne
rect 44445 13495 44538 13496
tri 44445 13494 44446 13495 ne
rect 44446 13494 44538 13495
rect 44584 13521 44657 13540
tri 44657 13521 44695 13559 sw
rect 70802 13540 71000 13598
rect 44584 13494 44695 13521
tri 44446 13493 44447 13494 ne
rect 44447 13493 44695 13494
tri 44447 13492 44448 13493 ne
rect 44448 13492 44695 13493
tri 44448 13491 44449 13492 ne
rect 44449 13491 44695 13492
tri 44449 13490 44450 13491 ne
rect 44450 13490 44695 13491
tri 44450 13489 44451 13490 ne
rect 44451 13489 44695 13490
tri 44451 13488 44452 13489 ne
rect 44452 13488 44695 13489
tri 44452 13487 44453 13488 ne
rect 44453 13487 44695 13488
tri 44453 13486 44454 13487 ne
rect 44454 13486 44695 13487
tri 44454 13485 44455 13486 ne
rect 44455 13485 44695 13486
tri 44455 13484 44456 13485 ne
rect 44456 13484 44695 13485
tri 44456 13483 44457 13484 ne
rect 44457 13483 44695 13484
tri 44457 13482 44458 13483 ne
rect 44458 13482 44695 13483
tri 44458 13481 44459 13482 ne
rect 44459 13481 44695 13482
tri 44459 13480 44460 13481 ne
rect 44460 13480 44695 13481
tri 44460 13479 44461 13480 ne
rect 44461 13479 44695 13480
tri 44461 13478 44462 13479 ne
rect 44462 13478 44695 13479
tri 44462 13477 44463 13478 ne
rect 44463 13477 44695 13478
tri 44463 13476 44464 13477 ne
rect 44464 13476 44695 13477
tri 44695 13476 44740 13521 sw
rect 70802 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
tri 44464 13475 44465 13476 ne
rect 44465 13475 44740 13476
tri 44465 13474 44466 13475 ne
rect 44466 13474 44740 13475
tri 44466 13473 44467 13474 ne
rect 44467 13473 44740 13474
tri 44467 13472 44468 13473 ne
rect 44468 13472 44740 13473
tri 44468 13471 44469 13472 ne
rect 44469 13471 44740 13472
tri 44469 13470 44470 13471 ne
rect 44470 13470 44740 13471
tri 44470 13469 44471 13470 ne
rect 44471 13469 44740 13470
tri 44471 13468 44472 13469 ne
rect 44472 13468 44740 13469
tri 44472 13467 44473 13468 ne
rect 44473 13467 44740 13468
tri 44473 13466 44474 13467 ne
rect 44474 13466 44740 13467
tri 44474 13465 44475 13466 ne
rect 44475 13465 44740 13466
tri 44475 13464 44476 13465 ne
rect 44476 13464 44740 13465
tri 44476 13463 44477 13464 ne
rect 44477 13463 44740 13464
tri 44477 13462 44478 13463 ne
rect 44478 13462 44740 13463
tri 44478 13461 44479 13462 ne
rect 44479 13461 44740 13462
tri 44479 13460 44480 13461 ne
rect 44480 13460 44740 13461
tri 44480 13459 44481 13460 ne
rect 44481 13459 44740 13460
tri 44481 13458 44482 13459 ne
rect 44482 13458 44740 13459
tri 44482 13457 44483 13458 ne
rect 44483 13457 44740 13458
tri 44483 13456 44484 13457 ne
rect 44484 13456 44740 13457
tri 44484 13455 44485 13456 ne
rect 44485 13455 44740 13456
tri 44485 13454 44486 13455 ne
rect 44486 13454 44740 13455
tri 44486 13453 44487 13454 ne
rect 44487 13453 44740 13454
tri 44487 13452 44488 13453 ne
rect 44488 13452 44740 13453
tri 44488 13451 44489 13452 ne
rect 44489 13451 44740 13452
tri 44489 13450 44490 13451 ne
rect 44490 13450 44740 13451
tri 44490 13449 44491 13450 ne
rect 44491 13449 44740 13450
tri 44491 13448 44492 13449 ne
rect 44492 13448 44740 13449
tri 44492 13447 44493 13448 ne
rect 44493 13447 44740 13448
tri 44493 13446 44494 13447 ne
rect 44494 13446 44740 13447
tri 44494 13445 44495 13446 ne
rect 44495 13445 44740 13446
tri 44495 13444 44496 13445 ne
rect 44496 13444 44740 13445
tri 44496 13443 44497 13444 ne
rect 44497 13443 44740 13444
tri 44497 13442 44498 13443 ne
rect 44498 13442 44740 13443
tri 44498 13441 44499 13442 ne
rect 44499 13441 44740 13442
tri 44499 13440 44500 13441 ne
rect 44500 13440 44740 13441
tri 44500 13439 44501 13440 ne
rect 44501 13439 44740 13440
tri 44501 13438 44502 13439 ne
rect 44502 13438 44740 13439
tri 44502 13437 44503 13438 ne
rect 44503 13437 44740 13438
tri 44503 13436 44504 13437 ne
rect 44504 13436 44740 13437
tri 44504 13435 44505 13436 ne
rect 44505 13435 44740 13436
tri 44505 13434 44506 13435 ne
rect 44506 13434 44740 13435
tri 44506 13433 44507 13434 ne
rect 44507 13433 44740 13434
tri 44507 13432 44508 13433 ne
rect 44508 13432 44740 13433
tri 44508 13431 44509 13432 ne
rect 44509 13431 44740 13432
tri 44740 13431 44785 13476 sw
rect 70802 13436 71000 13494
tri 44509 13430 44510 13431 ne
rect 44510 13430 44785 13431
tri 44510 13429 44511 13430 ne
rect 44511 13429 44785 13430
tri 44511 13428 44512 13429 ne
rect 44512 13428 44785 13429
tri 44512 13427 44513 13428 ne
rect 44513 13427 44785 13428
tri 44513 13426 44514 13427 ne
rect 44514 13426 44785 13427
tri 44514 13425 44515 13426 ne
rect 44515 13425 44785 13426
tri 44515 13424 44516 13425 ne
rect 44516 13424 44785 13425
tri 44516 13423 44517 13424 ne
rect 44517 13423 44785 13424
tri 44517 13422 44518 13423 ne
rect 44518 13422 44785 13423
tri 44518 13421 44519 13422 ne
rect 44519 13421 44785 13422
tri 44519 13420 44520 13421 ne
rect 44520 13420 44785 13421
tri 44520 13419 44521 13420 ne
rect 44521 13419 44785 13420
tri 44521 13418 44522 13419 ne
rect 44522 13418 44785 13419
tri 44522 13417 44523 13418 ne
rect 44523 13417 44785 13418
tri 44523 13416 44524 13417 ne
rect 44524 13416 44785 13417
tri 44524 13415 44525 13416 ne
rect 44525 13415 44785 13416
tri 44525 13414 44526 13415 ne
rect 44526 13414 44785 13415
tri 44526 13413 44527 13414 ne
rect 44527 13413 44785 13414
tri 44527 13412 44528 13413 ne
rect 44528 13412 44785 13413
tri 44528 13411 44529 13412 ne
rect 44529 13411 44785 13412
tri 44529 13410 44530 13411 ne
rect 44530 13410 44785 13411
tri 44530 13409 44531 13410 ne
rect 44531 13409 44785 13410
tri 44531 13408 44532 13409 ne
rect 44532 13408 44785 13409
tri 44532 13407 44533 13408 ne
rect 44533 13407 44670 13408
tri 44533 13406 44534 13407 ne
rect 44534 13406 44670 13407
tri 44534 13405 44535 13406 ne
rect 44535 13405 44670 13406
tri 44535 13404 44536 13405 ne
rect 44536 13404 44670 13405
tri 44536 13403 44537 13404 ne
rect 44537 13403 44670 13404
tri 44537 13402 44538 13403 ne
rect 44538 13402 44670 13403
tri 44538 13401 44539 13402 ne
rect 44539 13401 44670 13402
tri 44539 13400 44540 13401 ne
rect 44540 13400 44670 13401
tri 44540 13399 44541 13400 ne
rect 44541 13399 44670 13400
tri 44541 13398 44542 13399 ne
rect 44542 13398 44670 13399
tri 44542 13397 44543 13398 ne
rect 44543 13397 44670 13398
tri 44543 13396 44544 13397 ne
rect 44544 13396 44670 13397
tri 44544 13395 44545 13396 ne
rect 44545 13395 44670 13396
tri 44545 13394 44546 13395 ne
rect 44546 13394 44670 13395
tri 44546 13393 44547 13394 ne
rect 44547 13393 44670 13394
tri 44547 13392 44548 13393 ne
rect 44548 13392 44670 13393
tri 44548 13391 44549 13392 ne
rect 44549 13391 44670 13392
tri 44549 13390 44550 13391 ne
rect 44550 13390 44670 13391
tri 44550 13389 44551 13390 ne
rect 44551 13389 44670 13390
tri 44551 13388 44552 13389 ne
rect 44552 13388 44670 13389
tri 44552 13387 44553 13388 ne
rect 44553 13387 44670 13388
tri 44553 13386 44554 13387 ne
rect 44554 13386 44670 13387
tri 44554 13385 44555 13386 ne
rect 44555 13385 44670 13386
tri 44555 13384 44556 13385 ne
rect 44556 13384 44670 13385
tri 44556 13383 44557 13384 ne
rect 44557 13383 44670 13384
tri 44557 13382 44558 13383 ne
rect 44558 13382 44670 13383
tri 44558 13381 44559 13382 ne
rect 44559 13381 44670 13382
tri 44559 13380 44560 13381 ne
rect 44560 13380 44670 13381
tri 44560 13379 44561 13380 ne
rect 44561 13379 44670 13380
tri 44561 13378 44562 13379 ne
rect 44562 13378 44670 13379
tri 44562 13377 44563 13378 ne
rect 44563 13377 44670 13378
tri 44563 13376 44564 13377 ne
rect 44564 13376 44670 13377
tri 44564 13375 44565 13376 ne
rect 44565 13375 44670 13376
tri 44565 13374 44566 13375 ne
rect 44566 13374 44670 13375
tri 44566 13373 44567 13374 ne
rect 44567 13373 44670 13374
tri 44567 13368 44572 13373 ne
rect 44572 13368 44670 13373
tri 44572 13323 44617 13368 ne
rect 44617 13362 44670 13368
rect 44716 13386 44785 13408
tri 44785 13386 44830 13431 sw
rect 70802 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13373 44830 13386
tri 44830 13373 44843 13386 sw
rect 44716 13368 44843 13373
tri 44843 13368 44848 13373 sw
rect 44716 13362 44848 13368
rect 44617 13323 44848 13362
tri 44848 13323 44893 13368 sw
tri 44617 13291 44649 13323 ne
rect 44649 13291 44893 13323
tri 44893 13291 44925 13323 sw
rect 70802 13291 71000 13390
tri 44649 13246 44694 13291 ne
rect 44694 13269 71000 13291
rect 44694 13256 45088 13269
rect 44694 13246 44850 13256
tri 44694 13201 44739 13246 ne
rect 44739 13210 44850 13246
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44739 13201 71000 13210
tri 44739 13200 44740 13201 ne
rect 44740 13200 71000 13201
tri 44740 13155 44785 13200 ne
rect 44785 13165 71000 13200
rect 44785 13155 45088 13165
tri 44785 13110 44830 13155 ne
rect 44830 13119 45088 13155
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44830 13110 71000 13119
tri 44830 13097 44843 13110 ne
rect 44843 13097 71000 13110
<< psubdiffcont >>
rect 13119 70929 13165 70975
rect 13223 70929 13269 70975
rect 13377 70929 13423 70975
rect 13481 70929 13527 70975
rect 13585 70929 13631 70975
rect 13689 70929 13735 70975
rect 13793 70929 13839 70975
rect 13897 70929 13943 70975
rect 14001 70929 14047 70975
rect 14105 70929 14151 70975
rect 14209 70929 14255 70975
rect 14313 70929 14359 70975
rect 14417 70929 14463 70975
rect 14521 70929 14567 70975
rect 14625 70929 14671 70975
rect 14729 70929 14775 70975
rect 14833 70929 14879 70975
rect 14937 70929 14983 70975
rect 15041 70929 15087 70975
rect 15145 70929 15191 70975
rect 15249 70929 15295 70975
rect 15353 70929 15399 70975
rect 15457 70929 15503 70975
rect 15561 70929 15607 70975
rect 15665 70929 15711 70975
rect 15769 70929 15815 70975
rect 15873 70929 15919 70975
rect 15977 70929 16023 70975
rect 16081 70929 16127 70975
rect 16185 70929 16231 70975
rect 16289 70929 16335 70975
rect 16393 70929 16439 70975
rect 16497 70929 16543 70975
rect 16601 70929 16647 70975
rect 16705 70929 16751 70975
rect 16809 70929 16855 70975
rect 16913 70929 16959 70975
rect 17017 70929 17063 70975
rect 17121 70929 17167 70975
rect 17225 70929 17271 70975
rect 17329 70929 17375 70975
rect 17433 70929 17479 70975
rect 17537 70929 17583 70975
rect 17641 70929 17687 70975
rect 17745 70929 17791 70975
rect 17849 70929 17895 70975
rect 17953 70929 17999 70975
rect 18057 70929 18103 70975
rect 18161 70929 18207 70975
rect 18265 70929 18311 70975
rect 18369 70929 18415 70975
rect 18473 70929 18519 70975
rect 18577 70929 18623 70975
rect 18681 70929 18727 70975
rect 18785 70929 18831 70975
rect 18889 70929 18935 70975
rect 18993 70929 19039 70975
rect 19097 70929 19143 70975
rect 19201 70929 19247 70975
rect 19305 70929 19351 70975
rect 19409 70929 19455 70975
rect 19513 70929 19559 70975
rect 19617 70929 19663 70975
rect 19721 70929 19767 70975
rect 19825 70929 19871 70975
rect 19929 70929 19975 70975
rect 20033 70929 20079 70975
rect 20137 70929 20183 70975
rect 20241 70929 20287 70975
rect 20345 70929 20391 70975
rect 20449 70929 20495 70975
rect 20553 70929 20599 70975
rect 20657 70929 20703 70975
rect 20761 70929 20807 70975
rect 20865 70929 20911 70975
rect 20969 70929 21015 70975
rect 21073 70929 21119 70975
rect 21177 70929 21223 70975
rect 21281 70929 21327 70975
rect 21385 70929 21431 70975
rect 21489 70929 21535 70975
rect 21593 70929 21639 70975
rect 21697 70929 21743 70975
rect 21801 70929 21847 70975
rect 21905 70929 21951 70975
rect 22009 70929 22055 70975
rect 22113 70929 22159 70975
rect 22217 70929 22263 70975
rect 22321 70929 22367 70975
rect 22425 70929 22471 70975
rect 22529 70929 22575 70975
rect 22633 70929 22679 70975
rect 22737 70929 22783 70975
rect 22841 70929 22887 70975
rect 22945 70929 22991 70975
rect 23049 70929 23095 70975
rect 23153 70929 23199 70975
rect 23257 70929 23303 70975
rect 23361 70929 23407 70975
rect 23465 70929 23511 70975
rect 23569 70929 23615 70975
rect 23673 70929 23719 70975
rect 23777 70929 23823 70975
rect 23881 70929 23927 70975
rect 23985 70929 24031 70975
rect 24089 70929 24135 70975
rect 24193 70929 24239 70975
rect 24297 70929 24343 70975
rect 24401 70929 24447 70975
rect 24505 70929 24551 70975
rect 24609 70929 24655 70975
rect 24713 70929 24759 70975
rect 24817 70929 24863 70975
rect 24921 70929 24967 70975
rect 25025 70929 25071 70975
rect 25129 70929 25175 70975
rect 25233 70929 25279 70975
rect 25337 70929 25383 70975
rect 25441 70929 25487 70975
rect 25545 70929 25591 70975
rect 25649 70929 25695 70975
rect 25753 70929 25799 70975
rect 25857 70929 25903 70975
rect 25961 70929 26007 70975
rect 26065 70929 26111 70975
rect 26169 70929 26215 70975
rect 26273 70929 26319 70975
rect 26377 70929 26423 70975
rect 26481 70929 26527 70975
rect 26585 70929 26631 70975
rect 26689 70929 26735 70975
rect 26793 70929 26839 70975
rect 26897 70929 26943 70975
rect 27001 70929 27047 70975
rect 27105 70929 27151 70975
rect 27209 70929 27255 70975
rect 27313 70929 27359 70975
rect 27417 70929 27463 70975
rect 27521 70929 27567 70975
rect 27625 70929 27671 70975
rect 27729 70929 27775 70975
rect 27833 70929 27879 70975
rect 27937 70929 27983 70975
rect 28041 70929 28087 70975
rect 28145 70929 28191 70975
rect 28249 70929 28295 70975
rect 28353 70929 28399 70975
rect 28457 70929 28503 70975
rect 28561 70929 28607 70975
rect 28665 70929 28711 70975
rect 28769 70929 28815 70975
rect 28873 70929 28919 70975
rect 28977 70929 29023 70975
rect 29081 70929 29127 70975
rect 29185 70929 29231 70975
rect 29289 70929 29335 70975
rect 29393 70929 29439 70975
rect 29497 70929 29543 70975
rect 29601 70929 29647 70975
rect 29705 70929 29751 70975
rect 29809 70929 29855 70975
rect 29913 70929 29959 70975
rect 30017 70929 30063 70975
rect 30121 70929 30167 70975
rect 30225 70929 30271 70975
rect 30329 70929 30375 70975
rect 30433 70929 30479 70975
rect 30537 70929 30583 70975
rect 30641 70929 30687 70975
rect 30745 70929 30791 70975
rect 30849 70929 30895 70975
rect 30953 70929 30999 70975
rect 31057 70929 31103 70975
rect 31161 70929 31207 70975
rect 31265 70929 31311 70975
rect 31369 70929 31415 70975
rect 31473 70929 31519 70975
rect 31577 70929 31623 70975
rect 31681 70929 31727 70975
rect 31785 70929 31831 70975
rect 31889 70929 31935 70975
rect 31993 70929 32039 70975
rect 32097 70929 32143 70975
rect 32201 70929 32247 70975
rect 32305 70929 32351 70975
rect 32409 70929 32455 70975
rect 32513 70929 32559 70975
rect 32617 70929 32663 70975
rect 32721 70929 32767 70975
rect 32825 70929 32871 70975
rect 32929 70929 32975 70975
rect 33033 70929 33079 70975
rect 33137 70929 33183 70975
rect 33241 70929 33287 70975
rect 33345 70929 33391 70975
rect 33449 70929 33495 70975
rect 33553 70929 33599 70975
rect 33657 70929 33703 70975
rect 33761 70929 33807 70975
rect 33865 70929 33911 70975
rect 33969 70929 34015 70975
rect 34073 70929 34119 70975
rect 34177 70929 34223 70975
rect 34281 70929 34327 70975
rect 34385 70929 34431 70975
rect 34489 70929 34535 70975
rect 34593 70929 34639 70975
rect 34697 70929 34743 70975
rect 34801 70929 34847 70975
rect 34905 70929 34951 70975
rect 35009 70929 35055 70975
rect 35113 70929 35159 70975
rect 35217 70929 35263 70975
rect 35321 70929 35367 70975
rect 35425 70929 35471 70975
rect 35529 70929 35575 70975
rect 35633 70929 35679 70975
rect 35737 70929 35783 70975
rect 35841 70929 35887 70975
rect 35945 70929 35991 70975
rect 36049 70929 36095 70975
rect 36153 70929 36199 70975
rect 36257 70929 36303 70975
rect 36361 70929 36407 70975
rect 36465 70929 36511 70975
rect 36569 70929 36615 70975
rect 36673 70929 36719 70975
rect 36777 70929 36823 70975
rect 36881 70929 36927 70975
rect 36985 70929 37031 70975
rect 37089 70929 37135 70975
rect 37193 70929 37239 70975
rect 37297 70929 37343 70975
rect 37401 70929 37447 70975
rect 37505 70929 37551 70975
rect 37609 70929 37655 70975
rect 37713 70929 37759 70975
rect 37817 70929 37863 70975
rect 37921 70929 37967 70975
rect 38025 70929 38071 70975
rect 38129 70929 38175 70975
rect 38233 70929 38279 70975
rect 38337 70929 38383 70975
rect 38441 70929 38487 70975
rect 38545 70929 38591 70975
rect 38649 70929 38695 70975
rect 38753 70929 38799 70975
rect 38857 70929 38903 70975
rect 38961 70929 39007 70975
rect 39065 70929 39111 70975
rect 39169 70929 39215 70975
rect 39273 70929 39319 70975
rect 39377 70929 39423 70975
rect 39481 70929 39527 70975
rect 39585 70929 39631 70975
rect 39689 70929 39735 70975
rect 39793 70929 39839 70975
rect 39897 70929 39943 70975
rect 40001 70929 40047 70975
rect 40105 70929 40151 70975
rect 40209 70929 40255 70975
rect 40313 70929 40359 70975
rect 40417 70929 40463 70975
rect 40521 70929 40567 70975
rect 40625 70929 40671 70975
rect 40729 70929 40775 70975
rect 40833 70929 40879 70975
rect 40937 70929 40983 70975
rect 41041 70929 41087 70975
rect 41145 70929 41191 70975
rect 41249 70929 41295 70975
rect 41353 70929 41399 70975
rect 41457 70929 41503 70975
rect 41561 70929 41607 70975
rect 41665 70929 41711 70975
rect 41769 70929 41815 70975
rect 41873 70929 41919 70975
rect 41977 70929 42023 70975
rect 42081 70929 42127 70975
rect 42185 70929 42231 70975
rect 42289 70929 42335 70975
rect 42393 70929 42439 70975
rect 42497 70929 42543 70975
rect 42601 70929 42647 70975
rect 42705 70929 42751 70975
rect 42809 70929 42855 70975
rect 42913 70929 42959 70975
rect 43017 70929 43063 70975
rect 43121 70929 43167 70975
rect 43225 70929 43271 70975
rect 43329 70929 43375 70975
rect 43433 70929 43479 70975
rect 43537 70929 43583 70975
rect 43641 70929 43687 70975
rect 43745 70929 43791 70975
rect 43849 70929 43895 70975
rect 43953 70929 43999 70975
rect 44057 70929 44103 70975
rect 44161 70929 44207 70975
rect 44265 70929 44311 70975
rect 44369 70929 44415 70975
rect 44473 70929 44519 70975
rect 44577 70929 44623 70975
rect 44681 70929 44727 70975
rect 44785 70929 44831 70975
rect 44889 70929 44935 70975
rect 44993 70929 45039 70975
rect 45097 70929 45143 70975
rect 45201 70929 45247 70975
rect 45305 70929 45351 70975
rect 45409 70929 45455 70975
rect 45513 70929 45559 70975
rect 45617 70929 45663 70975
rect 45721 70929 45767 70975
rect 45825 70929 45871 70975
rect 45929 70929 45975 70975
rect 46033 70929 46079 70975
rect 46137 70929 46183 70975
rect 46241 70929 46287 70975
rect 46345 70929 46391 70975
rect 46449 70929 46495 70975
rect 46553 70929 46599 70975
rect 46657 70929 46703 70975
rect 46761 70929 46807 70975
rect 46865 70929 46911 70975
rect 46969 70929 47015 70975
rect 47073 70929 47119 70975
rect 47177 70929 47223 70975
rect 47281 70929 47327 70975
rect 47385 70929 47431 70975
rect 47489 70929 47535 70975
rect 47593 70929 47639 70975
rect 47697 70929 47743 70975
rect 47801 70929 47847 70975
rect 47905 70929 47951 70975
rect 48009 70929 48055 70975
rect 48113 70929 48159 70975
rect 48217 70929 48263 70975
rect 48321 70929 48367 70975
rect 48425 70929 48471 70975
rect 48529 70929 48575 70975
rect 48633 70929 48679 70975
rect 48737 70929 48783 70975
rect 48841 70929 48887 70975
rect 48945 70929 48991 70975
rect 49049 70929 49095 70975
rect 49153 70929 49199 70975
rect 49257 70929 49303 70975
rect 49361 70929 49407 70975
rect 49465 70929 49511 70975
rect 49569 70929 49615 70975
rect 49673 70929 49719 70975
rect 49777 70929 49823 70975
rect 49881 70929 49927 70975
rect 49985 70929 50031 70975
rect 50089 70929 50135 70975
rect 50193 70929 50239 70975
rect 50297 70929 50343 70975
rect 50401 70929 50447 70975
rect 50505 70929 50551 70975
rect 50609 70929 50655 70975
rect 50713 70929 50759 70975
rect 50817 70929 50863 70975
rect 50921 70929 50967 70975
rect 51025 70929 51071 70975
rect 51129 70929 51175 70975
rect 51233 70929 51279 70975
rect 51337 70929 51383 70975
rect 51441 70929 51487 70975
rect 51545 70929 51591 70975
rect 51649 70929 51695 70975
rect 51753 70929 51799 70975
rect 51857 70929 51903 70975
rect 51961 70929 52007 70975
rect 52065 70929 52111 70975
rect 52169 70929 52215 70975
rect 52273 70929 52319 70975
rect 52377 70929 52423 70975
rect 52481 70929 52527 70975
rect 52585 70929 52631 70975
rect 52689 70929 52735 70975
rect 52793 70929 52839 70975
rect 52897 70929 52943 70975
rect 53001 70929 53047 70975
rect 53105 70929 53151 70975
rect 53209 70929 53255 70975
rect 53313 70929 53359 70975
rect 53417 70929 53463 70975
rect 53521 70929 53567 70975
rect 53625 70929 53671 70975
rect 53729 70929 53775 70975
rect 53833 70929 53879 70975
rect 53937 70929 53983 70975
rect 54041 70929 54087 70975
rect 54145 70929 54191 70975
rect 54249 70929 54295 70975
rect 54353 70929 54399 70975
rect 54457 70929 54503 70975
rect 54561 70929 54607 70975
rect 54665 70929 54711 70975
rect 54769 70929 54815 70975
rect 54873 70929 54919 70975
rect 54977 70929 55023 70975
rect 55081 70929 55127 70975
rect 55185 70929 55231 70975
rect 55289 70929 55335 70975
rect 55393 70929 55439 70975
rect 55497 70929 55543 70975
rect 55601 70929 55647 70975
rect 55705 70929 55751 70975
rect 55809 70929 55855 70975
rect 55913 70929 55959 70975
rect 56017 70929 56063 70975
rect 56121 70929 56167 70975
rect 56225 70929 56271 70975
rect 56329 70929 56375 70975
rect 56433 70929 56479 70975
rect 56537 70929 56583 70975
rect 56641 70929 56687 70975
rect 56745 70929 56791 70975
rect 56849 70929 56895 70975
rect 56953 70929 56999 70975
rect 57057 70929 57103 70975
rect 57161 70929 57207 70975
rect 57265 70929 57311 70975
rect 57369 70929 57415 70975
rect 57473 70929 57519 70975
rect 57577 70929 57623 70975
rect 57681 70929 57727 70975
rect 57785 70929 57831 70975
rect 57889 70929 57935 70975
rect 57993 70929 58039 70975
rect 58097 70929 58143 70975
rect 58201 70929 58247 70975
rect 58305 70929 58351 70975
rect 58409 70929 58455 70975
rect 58513 70929 58559 70975
rect 58617 70929 58663 70975
rect 58721 70929 58767 70975
rect 58825 70929 58871 70975
rect 58929 70929 58975 70975
rect 59033 70929 59079 70975
rect 59137 70929 59183 70975
rect 59241 70929 59287 70975
rect 59345 70929 59391 70975
rect 59449 70929 59495 70975
rect 59553 70929 59599 70975
rect 59657 70929 59703 70975
rect 59761 70929 59807 70975
rect 59865 70929 59911 70975
rect 59969 70929 60015 70975
rect 60073 70929 60119 70975
rect 60177 70929 60223 70975
rect 60281 70929 60327 70975
rect 60385 70929 60431 70975
rect 60489 70929 60535 70975
rect 60593 70929 60639 70975
rect 60697 70929 60743 70975
rect 60801 70929 60847 70975
rect 60905 70929 60951 70975
rect 61009 70929 61055 70975
rect 61113 70929 61159 70975
rect 61217 70929 61263 70975
rect 61321 70929 61367 70975
rect 61425 70929 61471 70975
rect 61529 70929 61575 70975
rect 61633 70929 61679 70975
rect 61737 70929 61783 70975
rect 61841 70929 61887 70975
rect 61945 70929 61991 70975
rect 62049 70929 62095 70975
rect 62153 70929 62199 70975
rect 62257 70929 62303 70975
rect 62361 70929 62407 70975
rect 62465 70929 62511 70975
rect 62569 70929 62615 70975
rect 62673 70929 62719 70975
rect 62777 70929 62823 70975
rect 62881 70929 62927 70975
rect 62985 70929 63031 70975
rect 63089 70929 63135 70975
rect 63193 70929 63239 70975
rect 63297 70929 63343 70975
rect 63401 70929 63447 70975
rect 63505 70929 63551 70975
rect 63609 70929 63655 70975
rect 63713 70929 63759 70975
rect 63817 70929 63863 70975
rect 63921 70929 63967 70975
rect 64025 70929 64071 70975
rect 64129 70929 64175 70975
rect 64233 70929 64279 70975
rect 64337 70929 64383 70975
rect 64441 70929 64487 70975
rect 64545 70929 64591 70975
rect 64649 70929 64695 70975
rect 64753 70929 64799 70975
rect 64857 70929 64903 70975
rect 64961 70929 65007 70975
rect 65065 70929 65111 70975
rect 65169 70929 65215 70975
rect 65273 70929 65319 70975
rect 65377 70929 65423 70975
rect 65481 70929 65527 70975
rect 65585 70929 65631 70975
rect 65689 70929 65735 70975
rect 65793 70929 65839 70975
rect 65897 70929 65943 70975
rect 66001 70929 66047 70975
rect 66105 70929 66151 70975
rect 66209 70929 66255 70975
rect 66313 70929 66359 70975
rect 66417 70929 66463 70975
rect 66521 70929 66567 70975
rect 66625 70929 66671 70975
rect 66729 70929 66775 70975
rect 66833 70929 66879 70975
rect 66937 70929 66983 70975
rect 67041 70929 67087 70975
rect 67145 70929 67191 70975
rect 67249 70929 67295 70975
rect 67353 70929 67399 70975
rect 67457 70929 67503 70975
rect 67561 70929 67607 70975
rect 67665 70929 67711 70975
rect 67769 70929 67815 70975
rect 67873 70929 67919 70975
rect 67977 70929 68023 70975
rect 68081 70929 68127 70975
rect 68185 70929 68231 70975
rect 68289 70929 68335 70975
rect 68393 70929 68439 70975
rect 68497 70929 68543 70975
rect 68601 70929 68647 70975
rect 68705 70929 68751 70975
rect 68809 70929 68855 70975
rect 68913 70929 68959 70975
rect 69017 70929 69063 70975
rect 69121 70929 69167 70975
rect 69225 70929 69271 70975
rect 69329 70929 69375 70975
rect 69433 70929 69479 70975
rect 69537 70929 69583 70975
rect 69641 70929 69687 70975
rect 69745 70929 69791 70975
rect 69849 70929 69895 70975
rect 13119 70825 13165 70871
rect 13223 70825 13269 70871
rect 13377 70825 13423 70871
rect 13481 70825 13527 70871
rect 13585 70825 13631 70871
rect 13689 70825 13735 70871
rect 13793 70825 13839 70871
rect 13897 70825 13943 70871
rect 14001 70825 14047 70871
rect 14105 70825 14151 70871
rect 14209 70825 14255 70871
rect 14313 70825 14359 70871
rect 14417 70825 14463 70871
rect 14521 70825 14567 70871
rect 14625 70825 14671 70871
rect 14729 70825 14775 70871
rect 14833 70825 14879 70871
rect 14937 70825 14983 70871
rect 15041 70825 15087 70871
rect 15145 70825 15191 70871
rect 15249 70825 15295 70871
rect 15353 70825 15399 70871
rect 15457 70825 15503 70871
rect 15561 70825 15607 70871
rect 15665 70825 15711 70871
rect 15769 70825 15815 70871
rect 15873 70825 15919 70871
rect 15977 70825 16023 70871
rect 16081 70825 16127 70871
rect 16185 70825 16231 70871
rect 16289 70825 16335 70871
rect 16393 70825 16439 70871
rect 16497 70825 16543 70871
rect 16601 70825 16647 70871
rect 16705 70825 16751 70871
rect 16809 70825 16855 70871
rect 16913 70825 16959 70871
rect 17017 70825 17063 70871
rect 17121 70825 17167 70871
rect 17225 70825 17271 70871
rect 17329 70825 17375 70871
rect 17433 70825 17479 70871
rect 17537 70825 17583 70871
rect 17641 70825 17687 70871
rect 17745 70825 17791 70871
rect 17849 70825 17895 70871
rect 17953 70825 17999 70871
rect 18057 70825 18103 70871
rect 18161 70825 18207 70871
rect 18265 70825 18311 70871
rect 18369 70825 18415 70871
rect 18473 70825 18519 70871
rect 18577 70825 18623 70871
rect 18681 70825 18727 70871
rect 18785 70825 18831 70871
rect 18889 70825 18935 70871
rect 18993 70825 19039 70871
rect 19097 70825 19143 70871
rect 19201 70825 19247 70871
rect 19305 70825 19351 70871
rect 19409 70825 19455 70871
rect 19513 70825 19559 70871
rect 19617 70825 19663 70871
rect 19721 70825 19767 70871
rect 19825 70825 19871 70871
rect 19929 70825 19975 70871
rect 20033 70825 20079 70871
rect 20137 70825 20183 70871
rect 20241 70825 20287 70871
rect 20345 70825 20391 70871
rect 20449 70825 20495 70871
rect 20553 70825 20599 70871
rect 20657 70825 20703 70871
rect 20761 70825 20807 70871
rect 20865 70825 20911 70871
rect 20969 70825 21015 70871
rect 21073 70825 21119 70871
rect 21177 70825 21223 70871
rect 21281 70825 21327 70871
rect 21385 70825 21431 70871
rect 21489 70825 21535 70871
rect 21593 70825 21639 70871
rect 21697 70825 21743 70871
rect 21801 70825 21847 70871
rect 21905 70825 21951 70871
rect 22009 70825 22055 70871
rect 22113 70825 22159 70871
rect 22217 70825 22263 70871
rect 22321 70825 22367 70871
rect 22425 70825 22471 70871
rect 22529 70825 22575 70871
rect 22633 70825 22679 70871
rect 22737 70825 22783 70871
rect 22841 70825 22887 70871
rect 22945 70825 22991 70871
rect 23049 70825 23095 70871
rect 23153 70825 23199 70871
rect 23257 70825 23303 70871
rect 23361 70825 23407 70871
rect 23465 70825 23511 70871
rect 23569 70825 23615 70871
rect 23673 70825 23719 70871
rect 23777 70825 23823 70871
rect 23881 70825 23927 70871
rect 23985 70825 24031 70871
rect 24089 70825 24135 70871
rect 24193 70825 24239 70871
rect 24297 70825 24343 70871
rect 24401 70825 24447 70871
rect 24505 70825 24551 70871
rect 24609 70825 24655 70871
rect 24713 70825 24759 70871
rect 24817 70825 24863 70871
rect 24921 70825 24967 70871
rect 25025 70825 25071 70871
rect 25129 70825 25175 70871
rect 25233 70825 25279 70871
rect 25337 70825 25383 70871
rect 25441 70825 25487 70871
rect 25545 70825 25591 70871
rect 25649 70825 25695 70871
rect 25753 70825 25799 70871
rect 25857 70825 25903 70871
rect 25961 70825 26007 70871
rect 26065 70825 26111 70871
rect 26169 70825 26215 70871
rect 26273 70825 26319 70871
rect 26377 70825 26423 70871
rect 26481 70825 26527 70871
rect 26585 70825 26631 70871
rect 26689 70825 26735 70871
rect 26793 70825 26839 70871
rect 26897 70825 26943 70871
rect 27001 70825 27047 70871
rect 27105 70825 27151 70871
rect 27209 70825 27255 70871
rect 27313 70825 27359 70871
rect 27417 70825 27463 70871
rect 27521 70825 27567 70871
rect 27625 70825 27671 70871
rect 27729 70825 27775 70871
rect 27833 70825 27879 70871
rect 27937 70825 27983 70871
rect 28041 70825 28087 70871
rect 28145 70825 28191 70871
rect 28249 70825 28295 70871
rect 28353 70825 28399 70871
rect 28457 70825 28503 70871
rect 28561 70825 28607 70871
rect 28665 70825 28711 70871
rect 28769 70825 28815 70871
rect 28873 70825 28919 70871
rect 28977 70825 29023 70871
rect 29081 70825 29127 70871
rect 29185 70825 29231 70871
rect 29289 70825 29335 70871
rect 29393 70825 29439 70871
rect 29497 70825 29543 70871
rect 29601 70825 29647 70871
rect 29705 70825 29751 70871
rect 29809 70825 29855 70871
rect 29913 70825 29959 70871
rect 30017 70825 30063 70871
rect 30121 70825 30167 70871
rect 30225 70825 30271 70871
rect 30329 70825 30375 70871
rect 30433 70825 30479 70871
rect 30537 70825 30583 70871
rect 30641 70825 30687 70871
rect 30745 70825 30791 70871
rect 30849 70825 30895 70871
rect 30953 70825 30999 70871
rect 31057 70825 31103 70871
rect 31161 70825 31207 70871
rect 31265 70825 31311 70871
rect 31369 70825 31415 70871
rect 31473 70825 31519 70871
rect 31577 70825 31623 70871
rect 31681 70825 31727 70871
rect 31785 70825 31831 70871
rect 31889 70825 31935 70871
rect 31993 70825 32039 70871
rect 32097 70825 32143 70871
rect 32201 70825 32247 70871
rect 32305 70825 32351 70871
rect 32409 70825 32455 70871
rect 32513 70825 32559 70871
rect 32617 70825 32663 70871
rect 32721 70825 32767 70871
rect 32825 70825 32871 70871
rect 32929 70825 32975 70871
rect 33033 70825 33079 70871
rect 33137 70825 33183 70871
rect 33241 70825 33287 70871
rect 33345 70825 33391 70871
rect 33449 70825 33495 70871
rect 33553 70825 33599 70871
rect 33657 70825 33703 70871
rect 33761 70825 33807 70871
rect 33865 70825 33911 70871
rect 33969 70825 34015 70871
rect 34073 70825 34119 70871
rect 34177 70825 34223 70871
rect 34281 70825 34327 70871
rect 34385 70825 34431 70871
rect 34489 70825 34535 70871
rect 34593 70825 34639 70871
rect 34697 70825 34743 70871
rect 34801 70825 34847 70871
rect 34905 70825 34951 70871
rect 35009 70825 35055 70871
rect 35113 70825 35159 70871
rect 35217 70825 35263 70871
rect 35321 70825 35367 70871
rect 35425 70825 35471 70871
rect 35529 70825 35575 70871
rect 35633 70825 35679 70871
rect 35737 70825 35783 70871
rect 35841 70825 35887 70871
rect 35945 70825 35991 70871
rect 36049 70825 36095 70871
rect 36153 70825 36199 70871
rect 36257 70825 36303 70871
rect 36361 70825 36407 70871
rect 36465 70825 36511 70871
rect 36569 70825 36615 70871
rect 36673 70825 36719 70871
rect 36777 70825 36823 70871
rect 36881 70825 36927 70871
rect 36985 70825 37031 70871
rect 37089 70825 37135 70871
rect 37193 70825 37239 70871
rect 37297 70825 37343 70871
rect 37401 70825 37447 70871
rect 37505 70825 37551 70871
rect 37609 70825 37655 70871
rect 37713 70825 37759 70871
rect 37817 70825 37863 70871
rect 37921 70825 37967 70871
rect 38025 70825 38071 70871
rect 38129 70825 38175 70871
rect 38233 70825 38279 70871
rect 38337 70825 38383 70871
rect 38441 70825 38487 70871
rect 38545 70825 38591 70871
rect 38649 70825 38695 70871
rect 38753 70825 38799 70871
rect 38857 70825 38903 70871
rect 38961 70825 39007 70871
rect 39065 70825 39111 70871
rect 39169 70825 39215 70871
rect 39273 70825 39319 70871
rect 39377 70825 39423 70871
rect 39481 70825 39527 70871
rect 39585 70825 39631 70871
rect 39689 70825 39735 70871
rect 39793 70825 39839 70871
rect 39897 70825 39943 70871
rect 40001 70825 40047 70871
rect 40105 70825 40151 70871
rect 40209 70825 40255 70871
rect 40313 70825 40359 70871
rect 40417 70825 40463 70871
rect 40521 70825 40567 70871
rect 40625 70825 40671 70871
rect 40729 70825 40775 70871
rect 40833 70825 40879 70871
rect 40937 70825 40983 70871
rect 41041 70825 41087 70871
rect 41145 70825 41191 70871
rect 41249 70825 41295 70871
rect 41353 70825 41399 70871
rect 41457 70825 41503 70871
rect 41561 70825 41607 70871
rect 41665 70825 41711 70871
rect 41769 70825 41815 70871
rect 41873 70825 41919 70871
rect 41977 70825 42023 70871
rect 42081 70825 42127 70871
rect 42185 70825 42231 70871
rect 42289 70825 42335 70871
rect 42393 70825 42439 70871
rect 42497 70825 42543 70871
rect 42601 70825 42647 70871
rect 42705 70825 42751 70871
rect 42809 70825 42855 70871
rect 42913 70825 42959 70871
rect 43017 70825 43063 70871
rect 43121 70825 43167 70871
rect 43225 70825 43271 70871
rect 43329 70825 43375 70871
rect 43433 70825 43479 70871
rect 43537 70825 43583 70871
rect 43641 70825 43687 70871
rect 43745 70825 43791 70871
rect 43849 70825 43895 70871
rect 43953 70825 43999 70871
rect 44057 70825 44103 70871
rect 44161 70825 44207 70871
rect 44265 70825 44311 70871
rect 44369 70825 44415 70871
rect 44473 70825 44519 70871
rect 44577 70825 44623 70871
rect 44681 70825 44727 70871
rect 44785 70825 44831 70871
rect 44889 70825 44935 70871
rect 44993 70825 45039 70871
rect 45097 70825 45143 70871
rect 45201 70825 45247 70871
rect 45305 70825 45351 70871
rect 45409 70825 45455 70871
rect 45513 70825 45559 70871
rect 45617 70825 45663 70871
rect 45721 70825 45767 70871
rect 45825 70825 45871 70871
rect 45929 70825 45975 70871
rect 46033 70825 46079 70871
rect 46137 70825 46183 70871
rect 46241 70825 46287 70871
rect 46345 70825 46391 70871
rect 46449 70825 46495 70871
rect 46553 70825 46599 70871
rect 46657 70825 46703 70871
rect 46761 70825 46807 70871
rect 46865 70825 46911 70871
rect 46969 70825 47015 70871
rect 47073 70825 47119 70871
rect 47177 70825 47223 70871
rect 47281 70825 47327 70871
rect 47385 70825 47431 70871
rect 47489 70825 47535 70871
rect 47593 70825 47639 70871
rect 47697 70825 47743 70871
rect 47801 70825 47847 70871
rect 47905 70825 47951 70871
rect 48009 70825 48055 70871
rect 48113 70825 48159 70871
rect 48217 70825 48263 70871
rect 48321 70825 48367 70871
rect 48425 70825 48471 70871
rect 48529 70825 48575 70871
rect 48633 70825 48679 70871
rect 48737 70825 48783 70871
rect 48841 70825 48887 70871
rect 48945 70825 48991 70871
rect 49049 70825 49095 70871
rect 49153 70825 49199 70871
rect 49257 70825 49303 70871
rect 49361 70825 49407 70871
rect 49465 70825 49511 70871
rect 49569 70825 49615 70871
rect 49673 70825 49719 70871
rect 49777 70825 49823 70871
rect 49881 70825 49927 70871
rect 49985 70825 50031 70871
rect 50089 70825 50135 70871
rect 50193 70825 50239 70871
rect 50297 70825 50343 70871
rect 50401 70825 50447 70871
rect 50505 70825 50551 70871
rect 50609 70825 50655 70871
rect 50713 70825 50759 70871
rect 50817 70825 50863 70871
rect 50921 70825 50967 70871
rect 51025 70825 51071 70871
rect 51129 70825 51175 70871
rect 51233 70825 51279 70871
rect 51337 70825 51383 70871
rect 51441 70825 51487 70871
rect 51545 70825 51591 70871
rect 51649 70825 51695 70871
rect 51753 70825 51799 70871
rect 51857 70825 51903 70871
rect 51961 70825 52007 70871
rect 52065 70825 52111 70871
rect 52169 70825 52215 70871
rect 52273 70825 52319 70871
rect 52377 70825 52423 70871
rect 52481 70825 52527 70871
rect 52585 70825 52631 70871
rect 52689 70825 52735 70871
rect 52793 70825 52839 70871
rect 52897 70825 52943 70871
rect 53001 70825 53047 70871
rect 53105 70825 53151 70871
rect 53209 70825 53255 70871
rect 53313 70825 53359 70871
rect 53417 70825 53463 70871
rect 53521 70825 53567 70871
rect 53625 70825 53671 70871
rect 53729 70825 53775 70871
rect 53833 70825 53879 70871
rect 53937 70825 53983 70871
rect 54041 70825 54087 70871
rect 54145 70825 54191 70871
rect 54249 70825 54295 70871
rect 54353 70825 54399 70871
rect 54457 70825 54503 70871
rect 54561 70825 54607 70871
rect 54665 70825 54711 70871
rect 54769 70825 54815 70871
rect 54873 70825 54919 70871
rect 54977 70825 55023 70871
rect 55081 70825 55127 70871
rect 55185 70825 55231 70871
rect 55289 70825 55335 70871
rect 55393 70825 55439 70871
rect 55497 70825 55543 70871
rect 55601 70825 55647 70871
rect 55705 70825 55751 70871
rect 55809 70825 55855 70871
rect 55913 70825 55959 70871
rect 56017 70825 56063 70871
rect 56121 70825 56167 70871
rect 56225 70825 56271 70871
rect 56329 70825 56375 70871
rect 56433 70825 56479 70871
rect 56537 70825 56583 70871
rect 56641 70825 56687 70871
rect 56745 70825 56791 70871
rect 56849 70825 56895 70871
rect 56953 70825 56999 70871
rect 57057 70825 57103 70871
rect 57161 70825 57207 70871
rect 57265 70825 57311 70871
rect 57369 70825 57415 70871
rect 57473 70825 57519 70871
rect 57577 70825 57623 70871
rect 57681 70825 57727 70871
rect 57785 70825 57831 70871
rect 57889 70825 57935 70871
rect 57993 70825 58039 70871
rect 58097 70825 58143 70871
rect 58201 70825 58247 70871
rect 58305 70825 58351 70871
rect 58409 70825 58455 70871
rect 58513 70825 58559 70871
rect 58617 70825 58663 70871
rect 58721 70825 58767 70871
rect 58825 70825 58871 70871
rect 58929 70825 58975 70871
rect 59033 70825 59079 70871
rect 59137 70825 59183 70871
rect 59241 70825 59287 70871
rect 59345 70825 59391 70871
rect 59449 70825 59495 70871
rect 59553 70825 59599 70871
rect 59657 70825 59703 70871
rect 59761 70825 59807 70871
rect 59865 70825 59911 70871
rect 59969 70825 60015 70871
rect 60073 70825 60119 70871
rect 60177 70825 60223 70871
rect 60281 70825 60327 70871
rect 60385 70825 60431 70871
rect 60489 70825 60535 70871
rect 60593 70825 60639 70871
rect 60697 70825 60743 70871
rect 60801 70825 60847 70871
rect 60905 70825 60951 70871
rect 61009 70825 61055 70871
rect 61113 70825 61159 70871
rect 61217 70825 61263 70871
rect 61321 70825 61367 70871
rect 61425 70825 61471 70871
rect 61529 70825 61575 70871
rect 61633 70825 61679 70871
rect 61737 70825 61783 70871
rect 61841 70825 61887 70871
rect 61945 70825 61991 70871
rect 62049 70825 62095 70871
rect 62153 70825 62199 70871
rect 62257 70825 62303 70871
rect 62361 70825 62407 70871
rect 62465 70825 62511 70871
rect 62569 70825 62615 70871
rect 62673 70825 62719 70871
rect 62777 70825 62823 70871
rect 62881 70825 62927 70871
rect 62985 70825 63031 70871
rect 63089 70825 63135 70871
rect 63193 70825 63239 70871
rect 63297 70825 63343 70871
rect 63401 70825 63447 70871
rect 63505 70825 63551 70871
rect 63609 70825 63655 70871
rect 63713 70825 63759 70871
rect 63817 70825 63863 70871
rect 63921 70825 63967 70871
rect 64025 70825 64071 70871
rect 64129 70825 64175 70871
rect 64233 70825 64279 70871
rect 64337 70825 64383 70871
rect 64441 70825 64487 70871
rect 64545 70825 64591 70871
rect 64649 70825 64695 70871
rect 64753 70825 64799 70871
rect 64857 70825 64903 70871
rect 64961 70825 65007 70871
rect 65065 70825 65111 70871
rect 65169 70825 65215 70871
rect 65273 70825 65319 70871
rect 65377 70825 65423 70871
rect 65481 70825 65527 70871
rect 65585 70825 65631 70871
rect 65689 70825 65735 70871
rect 65793 70825 65839 70871
rect 65897 70825 65943 70871
rect 66001 70825 66047 70871
rect 66105 70825 66151 70871
rect 66209 70825 66255 70871
rect 66313 70825 66359 70871
rect 66417 70825 66463 70871
rect 66521 70825 66567 70871
rect 66625 70825 66671 70871
rect 66729 70825 66775 70871
rect 66833 70825 66879 70871
rect 66937 70825 66983 70871
rect 67041 70825 67087 70871
rect 67145 70825 67191 70871
rect 67249 70825 67295 70871
rect 67353 70825 67399 70871
rect 67457 70825 67503 70871
rect 67561 70825 67607 70871
rect 67665 70825 67711 70871
rect 67769 70825 67815 70871
rect 67873 70825 67919 70871
rect 67977 70825 68023 70871
rect 68081 70825 68127 70871
rect 68185 70825 68231 70871
rect 68289 70825 68335 70871
rect 68393 70825 68439 70871
rect 68497 70825 68543 70871
rect 68601 70825 68647 70871
rect 68705 70825 68751 70871
rect 68809 70825 68855 70871
rect 68913 70825 68959 70871
rect 69017 70825 69063 70871
rect 69121 70825 69167 70871
rect 69225 70825 69271 70871
rect 69329 70825 69375 70871
rect 69433 70825 69479 70871
rect 69537 70825 69583 70871
rect 69641 70825 69687 70871
rect 69745 70825 69791 70871
rect 69849 70825 69895 70871
rect 13119 70721 13165 70767
rect 13223 70721 13269 70767
rect 13119 70617 13165 70663
rect 13223 70617 13269 70663
rect 13119 70513 13165 70559
rect 13223 70513 13269 70559
rect 13119 70409 13165 70455
rect 13223 70409 13269 70455
rect 13119 70305 13165 70351
rect 13223 70305 13269 70351
rect 13119 70201 13165 70247
rect 13223 70201 13269 70247
rect 13119 70097 13165 70143
rect 13223 70097 13269 70143
rect 13119 69993 13165 70039
rect 13223 69993 13269 70039
rect 13119 69889 13165 69935
rect 13223 69889 13269 69935
rect 13119 69785 13165 69831
rect 13223 69785 13269 69831
rect 69796 70674 69842 70720
rect 69900 70674 69946 70720
rect 69796 70570 69842 70616
rect 69900 70570 69946 70616
rect 69796 70466 69842 70512
rect 69900 70466 69946 70512
rect 69796 70362 69842 70408
rect 69900 70362 69946 70408
rect 69796 70258 69842 70304
rect 69900 70258 69946 70304
rect 69796 70154 69842 70200
rect 69900 70154 69946 70200
rect 69796 70050 69842 70096
rect 69900 70050 69946 70096
rect 69796 69900 69842 69946
rect 69900 69900 69946 69946
rect 70004 69900 70050 69946
rect 70108 69900 70154 69946
rect 70212 69900 70258 69946
rect 70316 69900 70362 69946
rect 70420 69900 70466 69946
rect 70524 69900 70570 69946
rect 70628 69900 70674 69946
rect 70824 69862 70870 69908
rect 70928 69862 70974 69908
rect 69796 69796 69842 69842
rect 69900 69796 69946 69842
rect 70004 69796 70050 69842
rect 70108 69796 70154 69842
rect 70212 69796 70258 69842
rect 70316 69796 70362 69842
rect 70420 69796 70466 69842
rect 70524 69796 70570 69842
rect 70628 69796 70674 69842
rect 13119 69681 13165 69727
rect 13223 69681 13269 69727
rect 13119 69577 13165 69623
rect 13223 69577 13269 69623
rect 13119 69473 13165 69519
rect 13223 69473 13269 69519
rect 13119 69369 13165 69415
rect 13223 69369 13269 69415
rect 13119 69265 13165 69311
rect 13223 69265 13269 69311
rect 13119 69161 13165 69207
rect 13223 69161 13269 69207
rect 13119 69057 13165 69103
rect 13223 69057 13269 69103
rect 13119 68953 13165 68999
rect 13223 68953 13269 68999
rect 13119 68849 13165 68895
rect 13223 68849 13269 68895
rect 13119 68745 13165 68791
rect 13223 68745 13269 68791
rect 13119 68641 13165 68687
rect 13223 68641 13269 68687
rect 13119 68537 13165 68583
rect 13223 68537 13269 68583
rect 13119 68433 13165 68479
rect 13223 68433 13269 68479
rect 13119 68329 13165 68375
rect 13223 68329 13269 68375
rect 13119 68225 13165 68271
rect 13223 68225 13269 68271
rect 13119 68121 13165 68167
rect 13223 68121 13269 68167
rect 13119 68017 13165 68063
rect 13223 68017 13269 68063
rect 13119 67913 13165 67959
rect 13223 67913 13269 67959
rect 13119 67809 13165 67855
rect 13223 67809 13269 67855
rect 13119 67705 13165 67751
rect 13223 67705 13269 67751
rect 13119 67601 13165 67647
rect 13223 67601 13269 67647
rect 13119 67497 13165 67543
rect 13223 67497 13269 67543
rect 13119 67393 13165 67439
rect 13223 67393 13269 67439
rect 13119 67289 13165 67335
rect 13223 67289 13269 67335
rect 13119 67185 13165 67231
rect 13223 67185 13269 67231
rect 13119 67081 13165 67127
rect 13223 67081 13269 67127
rect 13119 66977 13165 67023
rect 13223 66977 13269 67023
rect 13119 66873 13165 66919
rect 13223 66873 13269 66919
rect 13119 66769 13165 66815
rect 13223 66769 13269 66815
rect 13119 66665 13165 66711
rect 13223 66665 13269 66711
rect 13119 66561 13165 66607
rect 13223 66561 13269 66607
rect 13119 66457 13165 66503
rect 13223 66457 13269 66503
rect 13119 66353 13165 66399
rect 13223 66353 13269 66399
rect 13119 66249 13165 66295
rect 13223 66249 13269 66295
rect 13119 66145 13165 66191
rect 13223 66145 13269 66191
rect 13119 66041 13165 66087
rect 13223 66041 13269 66087
rect 13119 65937 13165 65983
rect 13223 65937 13269 65983
rect 13119 65833 13165 65879
rect 13223 65833 13269 65879
rect 13119 65729 13165 65775
rect 13223 65729 13269 65775
rect 13119 65625 13165 65671
rect 13223 65625 13269 65671
rect 13119 65521 13165 65567
rect 13223 65521 13269 65567
rect 13119 65417 13165 65463
rect 13223 65417 13269 65463
rect 13119 65313 13165 65359
rect 13223 65313 13269 65359
rect 13119 65209 13165 65255
rect 13223 65209 13269 65255
rect 13119 65105 13165 65151
rect 13223 65105 13269 65151
rect 13119 65001 13165 65047
rect 13223 65001 13269 65047
rect 13119 64897 13165 64943
rect 13223 64897 13269 64943
rect 13119 64793 13165 64839
rect 13223 64793 13269 64839
rect 13119 64689 13165 64735
rect 13223 64689 13269 64735
rect 13119 64585 13165 64631
rect 13223 64585 13269 64631
rect 13119 64481 13165 64527
rect 13223 64481 13269 64527
rect 13119 64377 13165 64423
rect 13223 64377 13269 64423
rect 13119 64273 13165 64319
rect 13223 64273 13269 64319
rect 13119 64169 13165 64215
rect 13223 64169 13269 64215
rect 13119 64065 13165 64111
rect 13223 64065 13269 64111
rect 13119 63961 13165 64007
rect 13223 63961 13269 64007
rect 13119 63857 13165 63903
rect 13223 63857 13269 63903
rect 13119 63753 13165 63799
rect 13223 63753 13269 63799
rect 13119 63649 13165 63695
rect 13223 63649 13269 63695
rect 13119 63545 13165 63591
rect 13223 63545 13269 63591
rect 13119 63441 13165 63487
rect 13223 63441 13269 63487
rect 13119 63337 13165 63383
rect 13223 63337 13269 63383
rect 13119 63233 13165 63279
rect 13223 63233 13269 63279
rect 13119 63129 13165 63175
rect 13223 63129 13269 63175
rect 13119 63025 13165 63071
rect 13223 63025 13269 63071
rect 13119 62921 13165 62967
rect 13223 62921 13269 62967
rect 13119 62817 13165 62863
rect 13223 62817 13269 62863
rect 13119 62713 13165 62759
rect 13223 62713 13269 62759
rect 13119 62609 13165 62655
rect 13223 62609 13269 62655
rect 13119 62505 13165 62551
rect 13223 62505 13269 62551
rect 13119 62401 13165 62447
rect 13223 62401 13269 62447
rect 13119 62297 13165 62343
rect 13223 62297 13269 62343
rect 13119 62193 13165 62239
rect 13223 62193 13269 62239
rect 13119 62089 13165 62135
rect 13223 62089 13269 62135
rect 13119 61985 13165 62031
rect 13223 61985 13269 62031
rect 13119 61881 13165 61927
rect 13223 61881 13269 61927
rect 13119 61777 13165 61823
rect 13223 61777 13269 61823
rect 13119 61673 13165 61719
rect 13223 61673 13269 61719
rect 13119 61569 13165 61615
rect 13223 61569 13269 61615
rect 13119 61465 13165 61511
rect 13223 61465 13269 61511
rect 13119 61361 13165 61407
rect 13223 61361 13269 61407
rect 13119 61257 13165 61303
rect 13223 61257 13269 61303
rect 13119 61153 13165 61199
rect 13223 61153 13269 61199
rect 13119 61049 13165 61095
rect 13223 61049 13269 61095
rect 13119 60945 13165 60991
rect 13223 60945 13269 60991
rect 13119 60841 13165 60887
rect 13223 60841 13269 60887
rect 13119 60737 13165 60783
rect 13223 60737 13269 60783
rect 13119 60633 13165 60679
rect 13223 60633 13269 60679
rect 13119 60529 13165 60575
rect 13223 60529 13269 60575
rect 13119 60425 13165 60471
rect 13223 60425 13269 60471
rect 13119 60321 13165 60367
rect 13223 60321 13269 60367
rect 13119 60217 13165 60263
rect 13223 60217 13269 60263
rect 13119 60113 13165 60159
rect 13223 60113 13269 60159
rect 13119 60009 13165 60055
rect 13223 60009 13269 60055
rect 13119 59905 13165 59951
rect 13223 59905 13269 59951
rect 13119 59801 13165 59847
rect 13223 59801 13269 59847
rect 13119 59697 13165 59743
rect 13223 59697 13269 59743
rect 13119 59593 13165 59639
rect 13223 59593 13269 59639
rect 13119 59489 13165 59535
rect 13223 59489 13269 59535
rect 13119 59385 13165 59431
rect 13223 59385 13269 59431
rect 13119 59281 13165 59327
rect 13223 59281 13269 59327
rect 13119 59177 13165 59223
rect 13223 59177 13269 59223
rect 13119 59073 13165 59119
rect 13223 59073 13269 59119
rect 13119 58969 13165 59015
rect 13223 58969 13269 59015
rect 13119 58865 13165 58911
rect 13223 58865 13269 58911
rect 13119 58761 13165 58807
rect 13223 58761 13269 58807
rect 13119 58657 13165 58703
rect 13223 58657 13269 58703
rect 13119 58553 13165 58599
rect 13223 58553 13269 58599
rect 13119 58449 13165 58495
rect 13223 58449 13269 58495
rect 13119 58345 13165 58391
rect 13223 58345 13269 58391
rect 13119 58241 13165 58287
rect 13223 58241 13269 58287
rect 13119 58137 13165 58183
rect 13223 58137 13269 58183
rect 13119 58033 13165 58079
rect 13223 58033 13269 58079
rect 13119 57929 13165 57975
rect 13223 57929 13269 57975
rect 13119 57825 13165 57871
rect 13223 57825 13269 57871
rect 13119 57721 13165 57767
rect 13223 57721 13269 57767
rect 13119 57617 13165 57663
rect 13223 57617 13269 57663
rect 13119 57513 13165 57559
rect 13223 57513 13269 57559
rect 13119 57409 13165 57455
rect 13223 57409 13269 57455
rect 13119 57305 13165 57351
rect 13223 57305 13269 57351
rect 13119 57201 13165 57247
rect 13223 57201 13269 57247
rect 13119 57097 13165 57143
rect 13223 57097 13269 57143
rect 13119 56993 13165 57039
rect 13223 56993 13269 57039
rect 13119 56889 13165 56935
rect 13223 56889 13269 56935
rect 13119 56785 13165 56831
rect 13223 56785 13269 56831
rect 13119 56681 13165 56727
rect 13223 56681 13269 56727
rect 13119 56577 13165 56623
rect 13223 56577 13269 56623
rect 13119 56473 13165 56519
rect 13223 56473 13269 56519
rect 13119 56369 13165 56415
rect 13223 56369 13269 56415
rect 13119 56265 13165 56311
rect 13223 56265 13269 56311
rect 13119 56161 13165 56207
rect 13223 56161 13269 56207
rect 13119 56057 13165 56103
rect 13223 56057 13269 56103
rect 13119 55953 13165 55999
rect 13223 55953 13269 55999
rect 13119 55849 13165 55895
rect 13223 55849 13269 55895
rect 13119 55745 13165 55791
rect 13223 55745 13269 55791
rect 13119 55641 13165 55687
rect 13223 55641 13269 55687
rect 13119 55537 13165 55583
rect 13223 55537 13269 55583
rect 13119 55433 13165 55479
rect 13223 55433 13269 55479
rect 13119 55329 13165 55375
rect 13223 55329 13269 55375
rect 13119 55225 13165 55271
rect 13223 55225 13269 55271
rect 13119 55121 13165 55167
rect 13223 55121 13269 55167
rect 13119 55017 13165 55063
rect 13223 55017 13269 55063
rect 13119 54913 13165 54959
rect 13223 54913 13269 54959
rect 13119 54809 13165 54855
rect 13223 54809 13269 54855
rect 13119 54705 13165 54751
rect 13223 54705 13269 54751
rect 13119 54601 13165 54647
rect 13223 54601 13269 54647
rect 13119 54497 13165 54543
rect 13223 54497 13269 54543
rect 13119 54393 13165 54439
rect 13223 54393 13269 54439
rect 13119 54289 13165 54335
rect 13223 54289 13269 54335
rect 13119 54185 13165 54231
rect 13223 54185 13269 54231
rect 13119 54081 13165 54127
rect 13223 54081 13269 54127
rect 13119 53977 13165 54023
rect 13223 53977 13269 54023
rect 13119 53873 13165 53919
rect 13223 53873 13269 53919
rect 13119 53769 13165 53815
rect 13223 53769 13269 53815
rect 13119 53665 13165 53711
rect 13223 53665 13269 53711
rect 13119 53561 13165 53607
rect 13223 53561 13269 53607
rect 13119 53457 13165 53503
rect 13223 53457 13269 53503
rect 13119 53353 13165 53399
rect 13223 53353 13269 53399
rect 13119 53249 13165 53295
rect 13223 53249 13269 53295
rect 13119 53145 13165 53191
rect 13223 53145 13269 53191
rect 13119 53041 13165 53087
rect 13223 53041 13269 53087
rect 13119 52937 13165 52983
rect 13223 52937 13269 52983
rect 13119 52833 13165 52879
rect 13223 52833 13269 52879
rect 13119 52729 13165 52775
rect 13223 52729 13269 52775
rect 13119 52625 13165 52671
rect 13223 52625 13269 52671
rect 13119 52521 13165 52567
rect 13223 52521 13269 52567
rect 13119 52417 13165 52463
rect 13223 52417 13269 52463
rect 13119 52313 13165 52359
rect 13223 52313 13269 52359
rect 13119 52209 13165 52255
rect 13223 52209 13269 52255
rect 13119 52105 13165 52151
rect 13223 52105 13269 52151
rect 13119 52001 13165 52047
rect 13223 52001 13269 52047
rect 13119 51897 13165 51943
rect 13223 51897 13269 51943
rect 13119 51793 13165 51839
rect 13223 51793 13269 51839
rect 13119 51689 13165 51735
rect 13223 51689 13269 51735
rect 13119 51585 13165 51631
rect 13223 51585 13269 51631
rect 13119 51481 13165 51527
rect 13223 51481 13269 51527
rect 13119 51377 13165 51423
rect 13223 51377 13269 51423
rect 13119 51273 13165 51319
rect 13223 51273 13269 51319
rect 13119 51169 13165 51215
rect 13223 51169 13269 51215
rect 13119 51065 13165 51111
rect 13223 51065 13269 51111
rect 13119 50961 13165 51007
rect 13223 50961 13269 51007
rect 13119 50857 13165 50903
rect 13223 50857 13269 50903
rect 13119 50753 13165 50799
rect 13223 50753 13269 50799
rect 13119 50649 13165 50695
rect 13223 50649 13269 50695
rect 13119 50545 13165 50591
rect 13223 50545 13269 50591
rect 13119 50441 13165 50487
rect 13223 50441 13269 50487
rect 13119 50337 13165 50383
rect 13223 50337 13269 50383
rect 13119 50233 13165 50279
rect 13223 50233 13269 50279
rect 13119 50129 13165 50175
rect 13223 50129 13269 50175
rect 13119 50025 13165 50071
rect 13223 50025 13269 50071
rect 13119 49921 13165 49967
rect 13223 49921 13269 49967
rect 13119 49817 13165 49863
rect 13223 49817 13269 49863
rect 13119 49713 13165 49759
rect 13223 49713 13269 49759
rect 13119 49609 13165 49655
rect 13223 49609 13269 49655
rect 13119 49505 13165 49551
rect 13223 49505 13269 49551
rect 13119 49401 13165 49447
rect 13223 49401 13269 49447
rect 13119 49297 13165 49343
rect 13223 49297 13269 49343
rect 13119 49193 13165 49239
rect 13223 49193 13269 49239
rect 13119 49089 13165 49135
rect 13223 49089 13269 49135
rect 13119 48985 13165 49031
rect 13223 48985 13269 49031
rect 13119 48881 13165 48927
rect 13223 48881 13269 48927
rect 13119 48777 13165 48823
rect 13223 48777 13269 48823
rect 13119 48673 13165 48719
rect 13223 48673 13269 48719
rect 13119 48569 13165 48615
rect 13223 48569 13269 48615
rect 13119 48465 13165 48511
rect 13223 48465 13269 48511
rect 13119 48361 13165 48407
rect 13223 48361 13269 48407
rect 13119 48257 13165 48303
rect 13223 48257 13269 48303
rect 13119 48153 13165 48199
rect 13223 48153 13269 48199
rect 13119 48049 13165 48095
rect 13223 48049 13269 48095
rect 13119 47945 13165 47991
rect 13223 47945 13269 47991
rect 13119 47841 13165 47887
rect 13223 47841 13269 47887
rect 13119 47737 13165 47783
rect 13223 47737 13269 47783
rect 13119 47633 13165 47679
rect 13223 47633 13269 47679
rect 13119 47529 13165 47575
rect 13223 47529 13269 47575
rect 13119 47425 13165 47471
rect 13223 47425 13269 47471
rect 13119 47321 13165 47367
rect 13223 47321 13269 47367
rect 13119 47217 13165 47263
rect 13223 47217 13269 47263
rect 13119 47113 13165 47159
rect 13223 47113 13269 47159
rect 13119 47009 13165 47055
rect 13223 47009 13269 47055
rect 13119 46905 13165 46951
rect 13223 46905 13269 46951
rect 13119 46801 13165 46847
rect 13223 46801 13269 46847
rect 13119 46697 13165 46743
rect 13223 46697 13269 46743
rect 13119 46593 13165 46639
rect 13223 46593 13269 46639
rect 13119 46489 13165 46535
rect 13223 46489 13269 46535
rect 13119 46385 13165 46431
rect 13223 46385 13269 46431
rect 13119 46281 13165 46327
rect 13223 46281 13269 46327
rect 13119 46177 13165 46223
rect 13223 46177 13269 46223
rect 13119 46073 13165 46119
rect 13223 46073 13269 46119
rect 13119 45969 13165 46015
rect 13223 45969 13269 46015
rect 13119 45865 13165 45911
rect 13223 45865 13269 45911
rect 13119 45761 13165 45807
rect 13223 45761 13269 45807
rect 13119 45657 13165 45703
rect 13223 45657 13269 45703
rect 13119 45553 13165 45599
rect 13223 45553 13269 45599
rect 13119 45449 13165 45495
rect 13223 45449 13269 45495
rect 13119 45345 13165 45391
rect 13223 45345 13269 45391
rect 13119 45241 13165 45287
rect 13223 45241 13269 45287
rect 13119 45137 13165 45183
rect 13223 45137 13269 45183
rect 13119 45033 13165 45079
rect 13223 45033 13269 45079
rect 70824 69758 70870 69804
rect 70928 69758 70974 69804
rect 70824 69654 70870 69700
rect 70928 69654 70974 69700
rect 70824 69550 70870 69596
rect 70928 69550 70974 69596
rect 70824 69446 70870 69492
rect 70928 69446 70974 69492
rect 70824 69342 70870 69388
rect 70928 69342 70974 69388
rect 70824 69238 70870 69284
rect 70928 69238 70974 69284
rect 70824 69134 70870 69180
rect 70928 69134 70974 69180
rect 70824 69030 70870 69076
rect 70928 69030 70974 69076
rect 70824 68926 70870 68972
rect 70928 68926 70974 68972
rect 70824 68822 70870 68868
rect 70928 68822 70974 68868
rect 70824 68718 70870 68764
rect 70928 68718 70974 68764
rect 70824 68614 70870 68660
rect 70928 68614 70974 68660
rect 70824 68510 70870 68556
rect 70928 68510 70974 68556
rect 70824 68406 70870 68452
rect 70928 68406 70974 68452
rect 70824 68302 70870 68348
rect 70928 68302 70974 68348
rect 70824 68198 70870 68244
rect 70928 68198 70974 68244
rect 70824 68094 70870 68140
rect 70928 68094 70974 68140
rect 70824 67990 70870 68036
rect 70928 67990 70974 68036
rect 70824 67886 70870 67932
rect 70928 67886 70974 67932
rect 70824 67782 70870 67828
rect 70928 67782 70974 67828
rect 70824 67678 70870 67724
rect 70928 67678 70974 67724
rect 70824 67574 70870 67620
rect 70928 67574 70974 67620
rect 70824 67470 70870 67516
rect 70928 67470 70974 67516
rect 70824 67366 70870 67412
rect 70928 67366 70974 67412
rect 70824 67262 70870 67308
rect 70928 67262 70974 67308
rect 70824 67158 70870 67204
rect 70928 67158 70974 67204
rect 70824 67054 70870 67100
rect 70928 67054 70974 67100
rect 70824 66950 70870 66996
rect 70928 66950 70974 66996
rect 70824 66846 70870 66892
rect 70928 66846 70974 66892
rect 70824 66742 70870 66788
rect 70928 66742 70974 66788
rect 70824 66638 70870 66684
rect 70928 66638 70974 66684
rect 70824 66534 70870 66580
rect 70928 66534 70974 66580
rect 70824 66430 70870 66476
rect 70928 66430 70974 66476
rect 70824 66326 70870 66372
rect 70928 66326 70974 66372
rect 70824 66222 70870 66268
rect 70928 66222 70974 66268
rect 70824 66118 70870 66164
rect 70928 66118 70974 66164
rect 70824 66014 70870 66060
rect 70928 66014 70974 66060
rect 70824 65910 70870 65956
rect 70928 65910 70974 65956
rect 70824 65806 70870 65852
rect 70928 65806 70974 65852
rect 70824 65702 70870 65748
rect 70928 65702 70974 65748
rect 70824 65598 70870 65644
rect 70928 65598 70974 65644
rect 70824 65494 70870 65540
rect 70928 65494 70974 65540
rect 70824 65390 70870 65436
rect 70928 65390 70974 65436
rect 70824 65286 70870 65332
rect 70928 65286 70974 65332
rect 70824 65182 70870 65228
rect 70928 65182 70974 65228
rect 70824 65078 70870 65124
rect 70928 65078 70974 65124
rect 70824 64974 70870 65020
rect 70928 64974 70974 65020
rect 70824 64870 70870 64916
rect 70928 64870 70974 64916
rect 70824 64766 70870 64812
rect 70928 64766 70974 64812
rect 70824 64662 70870 64708
rect 70928 64662 70974 64708
rect 70824 64558 70870 64604
rect 70928 64558 70974 64604
rect 70824 64454 70870 64500
rect 70928 64454 70974 64500
rect 70824 64350 70870 64396
rect 70928 64350 70974 64396
rect 70824 64246 70870 64292
rect 70928 64246 70974 64292
rect 70824 64142 70870 64188
rect 70928 64142 70974 64188
rect 70824 64038 70870 64084
rect 70928 64038 70974 64084
rect 70824 63934 70870 63980
rect 70928 63934 70974 63980
rect 70824 63830 70870 63876
rect 70928 63830 70974 63876
rect 70824 63726 70870 63772
rect 70928 63726 70974 63772
rect 70824 63622 70870 63668
rect 70928 63622 70974 63668
rect 70824 63518 70870 63564
rect 70928 63518 70974 63564
rect 70824 63414 70870 63460
rect 70928 63414 70974 63460
rect 70824 63310 70870 63356
rect 70928 63310 70974 63356
rect 70824 63206 70870 63252
rect 70928 63206 70974 63252
rect 70824 63102 70870 63148
rect 70928 63102 70974 63148
rect 70824 62998 70870 63044
rect 70928 62998 70974 63044
rect 70824 62894 70870 62940
rect 70928 62894 70974 62940
rect 70824 62790 70870 62836
rect 70928 62790 70974 62836
rect 70824 62686 70870 62732
rect 70928 62686 70974 62732
rect 70824 62582 70870 62628
rect 70928 62582 70974 62628
rect 70824 62478 70870 62524
rect 70928 62478 70974 62524
rect 70824 62374 70870 62420
rect 70928 62374 70974 62420
rect 70824 62270 70870 62316
rect 70928 62270 70974 62316
rect 70824 62166 70870 62212
rect 70928 62166 70974 62212
rect 70824 62062 70870 62108
rect 70928 62062 70974 62108
rect 70824 61958 70870 62004
rect 70928 61958 70974 62004
rect 70824 61854 70870 61900
rect 70928 61854 70974 61900
rect 70824 61750 70870 61796
rect 70928 61750 70974 61796
rect 70824 61646 70870 61692
rect 70928 61646 70974 61692
rect 70824 61542 70870 61588
rect 70928 61542 70974 61588
rect 70824 61438 70870 61484
rect 70928 61438 70974 61484
rect 70824 61334 70870 61380
rect 70928 61334 70974 61380
rect 70824 61230 70870 61276
rect 70928 61230 70974 61276
rect 70824 61126 70870 61172
rect 70928 61126 70974 61172
rect 70824 61022 70870 61068
rect 70928 61022 70974 61068
rect 70824 60918 70870 60964
rect 70928 60918 70974 60964
rect 70824 60814 70870 60860
rect 70928 60814 70974 60860
rect 70824 60710 70870 60756
rect 70928 60710 70974 60756
rect 70824 60606 70870 60652
rect 70928 60606 70974 60652
rect 70824 60502 70870 60548
rect 70928 60502 70974 60548
rect 70824 60398 70870 60444
rect 70928 60398 70974 60444
rect 70824 60294 70870 60340
rect 70928 60294 70974 60340
rect 70824 60190 70870 60236
rect 70928 60190 70974 60236
rect 70824 60086 70870 60132
rect 70928 60086 70974 60132
rect 70824 59982 70870 60028
rect 70928 59982 70974 60028
rect 70824 59878 70870 59924
rect 70928 59878 70974 59924
rect 70824 59774 70870 59820
rect 70928 59774 70974 59820
rect 70824 59670 70870 59716
rect 70928 59670 70974 59716
rect 70824 59566 70870 59612
rect 70928 59566 70974 59612
rect 70824 59462 70870 59508
rect 70928 59462 70974 59508
rect 70824 59358 70870 59404
rect 70928 59358 70974 59404
rect 70824 59254 70870 59300
rect 70928 59254 70974 59300
rect 70824 59150 70870 59196
rect 70928 59150 70974 59196
rect 70824 59046 70870 59092
rect 70928 59046 70974 59092
rect 70824 58942 70870 58988
rect 70928 58942 70974 58988
rect 70824 58838 70870 58884
rect 70928 58838 70974 58884
rect 70824 58734 70870 58780
rect 70928 58734 70974 58780
rect 70824 58630 70870 58676
rect 70928 58630 70974 58676
rect 70824 58526 70870 58572
rect 70928 58526 70974 58572
rect 70824 58422 70870 58468
rect 70928 58422 70974 58468
rect 70824 58318 70870 58364
rect 70928 58318 70974 58364
rect 70824 58214 70870 58260
rect 70928 58214 70974 58260
rect 70824 58110 70870 58156
rect 70928 58110 70974 58156
rect 70824 58006 70870 58052
rect 70928 58006 70974 58052
rect 70824 57902 70870 57948
rect 70928 57902 70974 57948
rect 70824 57798 70870 57844
rect 70928 57798 70974 57844
rect 70824 57694 70870 57740
rect 70928 57694 70974 57740
rect 70824 57590 70870 57636
rect 70928 57590 70974 57636
rect 70824 57486 70870 57532
rect 70928 57486 70974 57532
rect 70824 57382 70870 57428
rect 70928 57382 70974 57428
rect 70824 57278 70870 57324
rect 70928 57278 70974 57324
rect 70824 57174 70870 57220
rect 70928 57174 70974 57220
rect 70824 57070 70870 57116
rect 70928 57070 70974 57116
rect 70824 56966 70870 57012
rect 70928 56966 70974 57012
rect 70824 56862 70870 56908
rect 70928 56862 70974 56908
rect 70824 56758 70870 56804
rect 70928 56758 70974 56804
rect 70824 56654 70870 56700
rect 70928 56654 70974 56700
rect 70824 56550 70870 56596
rect 70928 56550 70974 56596
rect 70824 56446 70870 56492
rect 70928 56446 70974 56492
rect 70824 56342 70870 56388
rect 70928 56342 70974 56388
rect 70824 56238 70870 56284
rect 70928 56238 70974 56284
rect 70824 56134 70870 56180
rect 70928 56134 70974 56180
rect 70824 56030 70870 56076
rect 70928 56030 70974 56076
rect 70824 55926 70870 55972
rect 70928 55926 70974 55972
rect 70824 55822 70870 55868
rect 70928 55822 70974 55868
rect 70824 55718 70870 55764
rect 70928 55718 70974 55764
rect 70824 55614 70870 55660
rect 70928 55614 70974 55660
rect 70824 55510 70870 55556
rect 70928 55510 70974 55556
rect 70824 55406 70870 55452
rect 70928 55406 70974 55452
rect 70824 55302 70870 55348
rect 70928 55302 70974 55348
rect 70824 55198 70870 55244
rect 70928 55198 70974 55244
rect 70824 55094 70870 55140
rect 70928 55094 70974 55140
rect 70824 54990 70870 55036
rect 70928 54990 70974 55036
rect 70824 54886 70870 54932
rect 70928 54886 70974 54932
rect 70824 54782 70870 54828
rect 70928 54782 70974 54828
rect 70824 54678 70870 54724
rect 70928 54678 70974 54724
rect 70824 54574 70870 54620
rect 70928 54574 70974 54620
rect 70824 54470 70870 54516
rect 70928 54470 70974 54516
rect 70824 54366 70870 54412
rect 70928 54366 70974 54412
rect 70824 54262 70870 54308
rect 70928 54262 70974 54308
rect 70824 54158 70870 54204
rect 70928 54158 70974 54204
rect 70824 54054 70870 54100
rect 70928 54054 70974 54100
rect 70824 53950 70870 53996
rect 70928 53950 70974 53996
rect 70824 53846 70870 53892
rect 70928 53846 70974 53892
rect 70824 53742 70870 53788
rect 70928 53742 70974 53788
rect 70824 53638 70870 53684
rect 70928 53638 70974 53684
rect 70824 53534 70870 53580
rect 70928 53534 70974 53580
rect 70824 53430 70870 53476
rect 70928 53430 70974 53476
rect 70824 53326 70870 53372
rect 70928 53326 70974 53372
rect 70824 53222 70870 53268
rect 70928 53222 70974 53268
rect 70824 53118 70870 53164
rect 70928 53118 70974 53164
rect 70824 53014 70870 53060
rect 70928 53014 70974 53060
rect 70824 52910 70870 52956
rect 70928 52910 70974 52956
rect 70824 52806 70870 52852
rect 70928 52806 70974 52852
rect 70824 52702 70870 52748
rect 70928 52702 70974 52748
rect 70824 52598 70870 52644
rect 70928 52598 70974 52644
rect 70824 52494 70870 52540
rect 70928 52494 70974 52540
rect 70824 52390 70870 52436
rect 70928 52390 70974 52436
rect 70824 52286 70870 52332
rect 70928 52286 70974 52332
rect 70824 52182 70870 52228
rect 70928 52182 70974 52228
rect 70824 52078 70870 52124
rect 70928 52078 70974 52124
rect 70824 51974 70870 52020
rect 70928 51974 70974 52020
rect 70824 51870 70870 51916
rect 70928 51870 70974 51916
rect 70824 51766 70870 51812
rect 70928 51766 70974 51812
rect 70824 51662 70870 51708
rect 70928 51662 70974 51708
rect 70824 51558 70870 51604
rect 70928 51558 70974 51604
rect 70824 51454 70870 51500
rect 70928 51454 70974 51500
rect 70824 51350 70870 51396
rect 70928 51350 70974 51396
rect 70824 51246 70870 51292
rect 70928 51246 70974 51292
rect 70824 51142 70870 51188
rect 70928 51142 70974 51188
rect 70824 51038 70870 51084
rect 70928 51038 70974 51084
rect 70824 50934 70870 50980
rect 70928 50934 70974 50980
rect 70824 50830 70870 50876
rect 70928 50830 70974 50876
rect 70824 50726 70870 50772
rect 70928 50726 70974 50772
rect 70824 50622 70870 50668
rect 70928 50622 70974 50668
rect 70824 50518 70870 50564
rect 70928 50518 70974 50564
rect 70824 50414 70870 50460
rect 70928 50414 70974 50460
rect 70824 50310 70870 50356
rect 70928 50310 70974 50356
rect 70824 50206 70870 50252
rect 70928 50206 70974 50252
rect 70824 50102 70870 50148
rect 70928 50102 70974 50148
rect 70824 49998 70870 50044
rect 70928 49998 70974 50044
rect 70824 49894 70870 49940
rect 70928 49894 70974 49940
rect 70824 49790 70870 49836
rect 70928 49790 70974 49836
rect 70824 49686 70870 49732
rect 70928 49686 70974 49732
rect 70824 49582 70870 49628
rect 70928 49582 70974 49628
rect 70824 49478 70870 49524
rect 70928 49478 70974 49524
rect 70824 49374 70870 49420
rect 70928 49374 70974 49420
rect 70824 49270 70870 49316
rect 70928 49270 70974 49316
rect 70824 49166 70870 49212
rect 70928 49166 70974 49212
rect 70824 49062 70870 49108
rect 70928 49062 70974 49108
rect 70824 48958 70870 49004
rect 70928 48958 70974 49004
rect 70824 48854 70870 48900
rect 70928 48854 70974 48900
rect 70824 48750 70870 48796
rect 70928 48750 70974 48796
rect 70824 48646 70870 48692
rect 70928 48646 70974 48692
rect 70824 48542 70870 48588
rect 70928 48542 70974 48588
rect 70824 48438 70870 48484
rect 70928 48438 70974 48484
rect 70824 48334 70870 48380
rect 70928 48334 70974 48380
rect 70824 48230 70870 48276
rect 70928 48230 70974 48276
rect 70824 48126 70870 48172
rect 70928 48126 70974 48172
rect 70824 48022 70870 48068
rect 70928 48022 70974 48068
rect 70824 47918 70870 47964
rect 70928 47918 70974 47964
rect 70824 47814 70870 47860
rect 70928 47814 70974 47860
rect 70824 47710 70870 47756
rect 70928 47710 70974 47756
rect 70824 47606 70870 47652
rect 70928 47606 70974 47652
rect 70824 47502 70870 47548
rect 70928 47502 70974 47548
rect 70824 47398 70870 47444
rect 70928 47398 70974 47444
rect 70824 47294 70870 47340
rect 70928 47294 70974 47340
rect 70824 47190 70870 47236
rect 70928 47190 70974 47236
rect 70824 47086 70870 47132
rect 70928 47086 70974 47132
rect 70824 46982 70870 47028
rect 70928 46982 70974 47028
rect 70824 46878 70870 46924
rect 70928 46878 70974 46924
rect 70824 46774 70870 46820
rect 70928 46774 70974 46820
rect 70824 46670 70870 46716
rect 70928 46670 70974 46716
rect 70824 46566 70870 46612
rect 70928 46566 70974 46612
rect 70824 46462 70870 46508
rect 70928 46462 70974 46508
rect 70824 46358 70870 46404
rect 70928 46358 70974 46404
rect 70824 46254 70870 46300
rect 70928 46254 70974 46300
rect 70824 46150 70870 46196
rect 70928 46150 70974 46196
rect 70824 46046 70870 46092
rect 70928 46046 70974 46092
rect 70824 45942 70870 45988
rect 70928 45942 70974 45988
rect 70824 45838 70870 45884
rect 70928 45838 70974 45884
rect 70824 45734 70870 45780
rect 70928 45734 70974 45780
rect 70824 45630 70870 45676
rect 70928 45630 70974 45676
rect 70824 45526 70870 45572
rect 70928 45526 70974 45572
rect 70824 45422 70870 45468
rect 70928 45422 70974 45468
rect 70824 45318 70870 45364
rect 70928 45318 70974 45364
rect 70824 45214 70870 45260
rect 70928 45214 70974 45260
rect 70824 45110 70870 45156
rect 70928 45110 70974 45156
rect 70824 45006 70870 45052
rect 70928 45006 70974 45052
rect 70824 44902 70870 44948
rect 70928 44902 70974 44948
rect 13254 44778 13300 44824
rect 70824 44798 70870 44844
rect 70928 44798 70974 44844
rect 13386 44646 13432 44692
rect 70824 44694 70870 44740
rect 70928 44694 70974 44740
rect 70824 44590 70870 44636
rect 70928 44590 70974 44636
rect 13518 44514 13564 44560
rect 70824 44486 70870 44532
rect 70928 44486 70974 44532
rect 13650 44382 13696 44428
rect 70824 44382 70870 44428
rect 70928 44382 70974 44428
rect 13782 44250 13828 44296
rect 70824 44278 70870 44324
rect 70928 44278 70974 44324
rect 13914 44118 13960 44164
rect 70824 44174 70870 44220
rect 70928 44174 70974 44220
rect 70824 44070 70870 44116
rect 70928 44070 70974 44116
rect 14046 43986 14092 44032
rect 70824 43966 70870 44012
rect 70928 43966 70974 44012
rect 14178 43854 14224 43900
rect 70824 43862 70870 43908
rect 70928 43862 70974 43908
rect 14310 43722 14356 43768
rect 70824 43758 70870 43804
rect 70928 43758 70974 43804
rect 70824 43654 70870 43700
rect 70928 43654 70974 43700
rect 14442 43590 14488 43636
rect 70824 43550 70870 43596
rect 70928 43550 70974 43596
rect 14574 43458 14620 43504
rect 70824 43446 70870 43492
rect 70928 43446 70974 43492
rect 14706 43326 14752 43372
rect 70824 43342 70870 43388
rect 70928 43342 70974 43388
rect 14838 43194 14884 43240
rect 70824 43238 70870 43284
rect 70928 43238 70974 43284
rect 70824 43134 70870 43180
rect 70928 43134 70974 43180
rect 14970 43062 15016 43108
rect 70824 43030 70870 43076
rect 70928 43030 70974 43076
rect 15102 42930 15148 42976
rect 70824 42926 70870 42972
rect 70928 42926 70974 42972
rect 15234 42798 15280 42844
rect 70824 42822 70870 42868
rect 70928 42822 70974 42868
rect 15366 42666 15412 42712
rect 70824 42718 70870 42764
rect 70928 42718 70974 42764
rect 70824 42614 70870 42660
rect 70928 42614 70974 42660
rect 15498 42534 15544 42580
rect 70824 42510 70870 42556
rect 70928 42510 70974 42556
rect 15630 42402 15676 42448
rect 70824 42406 70870 42452
rect 70928 42406 70974 42452
rect 15762 42270 15808 42316
rect 70824 42302 70870 42348
rect 70928 42302 70974 42348
rect 15894 42138 15940 42184
rect 70824 42198 70870 42244
rect 70928 42198 70974 42244
rect 70824 42094 70870 42140
rect 70928 42094 70974 42140
rect 16026 42006 16072 42052
rect 70824 41990 70870 42036
rect 70928 41990 70974 42036
rect 16158 41874 16204 41920
rect 70824 41886 70870 41932
rect 70928 41886 70974 41932
rect 16290 41742 16336 41788
rect 70824 41782 70870 41828
rect 70928 41782 70974 41828
rect 70824 41678 70870 41724
rect 70928 41678 70974 41724
rect 16422 41610 16468 41656
rect 70824 41574 70870 41620
rect 70928 41574 70974 41620
rect 16554 41478 16600 41524
rect 70824 41470 70870 41516
rect 70928 41470 70974 41516
rect 16686 41346 16732 41392
rect 70824 41366 70870 41412
rect 70928 41366 70974 41412
rect 16818 41214 16864 41260
rect 70824 41262 70870 41308
rect 70928 41262 70974 41308
rect 70824 41158 70870 41204
rect 70928 41158 70974 41204
rect 16950 41082 16996 41128
rect 70824 41054 70870 41100
rect 70928 41054 70974 41100
rect 17082 40950 17128 40996
rect 70824 40950 70870 40996
rect 70928 40950 70974 40996
rect 17214 40818 17260 40864
rect 70824 40846 70870 40892
rect 70928 40846 70974 40892
rect 70824 40742 70870 40788
rect 70928 40742 70974 40788
rect 17346 40686 17392 40732
rect 70824 40638 70870 40684
rect 70928 40638 70974 40684
rect 17478 40554 17524 40600
rect 70824 40534 70870 40580
rect 70928 40534 70974 40580
rect 17610 40422 17656 40468
rect 70824 40430 70870 40476
rect 70928 40430 70974 40476
rect 17742 40290 17788 40336
rect 70824 40326 70870 40372
rect 70928 40326 70974 40372
rect 17874 40158 17920 40204
rect 70824 40222 70870 40268
rect 70928 40222 70974 40268
rect 70824 40118 70870 40164
rect 70928 40118 70974 40164
rect 18006 40026 18052 40072
rect 70824 40014 70870 40060
rect 70928 40014 70974 40060
rect 18138 39894 18184 39940
rect 70824 39910 70870 39956
rect 70928 39910 70974 39956
rect 18270 39762 18316 39808
rect 70824 39806 70870 39852
rect 70928 39806 70974 39852
rect 70824 39702 70870 39748
rect 70928 39702 70974 39748
rect 18402 39630 18448 39676
rect 70824 39598 70870 39644
rect 70928 39598 70974 39644
rect 18534 39498 18580 39544
rect 70824 39494 70870 39540
rect 70928 39494 70974 39540
rect 18666 39366 18712 39412
rect 70824 39390 70870 39436
rect 70928 39390 70974 39436
rect 18798 39234 18844 39280
rect 70824 39286 70870 39332
rect 70928 39286 70974 39332
rect 18930 39102 18976 39148
rect 70824 39182 70870 39228
rect 70928 39182 70974 39228
rect 70824 39078 70870 39124
rect 70928 39078 70974 39124
rect 19062 38970 19108 39016
rect 70824 38974 70870 39020
rect 70928 38974 70974 39020
rect 19194 38838 19240 38884
rect 70824 38870 70870 38916
rect 70928 38870 70974 38916
rect 70824 38766 70870 38812
rect 70928 38766 70974 38812
rect 19326 38706 19372 38752
rect 70824 38662 70870 38708
rect 70928 38662 70974 38708
rect 19458 38574 19504 38620
rect 70824 38558 70870 38604
rect 70928 38558 70974 38604
rect 19590 38442 19636 38488
rect 70824 38454 70870 38500
rect 70928 38454 70974 38500
rect 19722 38310 19768 38356
rect 70824 38350 70870 38396
rect 70928 38350 70974 38396
rect 19854 38178 19900 38224
rect 70824 38246 70870 38292
rect 70928 38246 70974 38292
rect 70824 38142 70870 38188
rect 70928 38142 70974 38188
rect 19986 38046 20032 38092
rect 70824 38038 70870 38084
rect 70928 38038 70974 38084
rect 20118 37914 20164 37960
rect 70824 37934 70870 37980
rect 70928 37934 70974 37980
rect 20250 37782 20296 37828
rect 70824 37830 70870 37876
rect 70928 37830 70974 37876
rect 70824 37726 70870 37772
rect 70928 37726 70974 37772
rect 20382 37650 20428 37696
rect 70824 37622 70870 37668
rect 70928 37622 70974 37668
rect 20514 37518 20560 37564
rect 70824 37518 70870 37564
rect 70928 37518 70974 37564
rect 20646 37386 20692 37432
rect 70824 37414 70870 37460
rect 70928 37414 70974 37460
rect 20778 37254 20824 37300
rect 70824 37310 70870 37356
rect 70928 37310 70974 37356
rect 70824 37206 70870 37252
rect 70928 37206 70974 37252
rect 20910 37122 20956 37168
rect 70824 37102 70870 37148
rect 70928 37102 70974 37148
rect 21042 36990 21088 37036
rect 70824 36998 70870 37044
rect 70928 36998 70974 37044
rect 21174 36858 21220 36904
rect 70824 36894 70870 36940
rect 70928 36894 70974 36940
rect 21306 36726 21352 36772
rect 70824 36790 70870 36836
rect 70928 36790 70974 36836
rect 70824 36686 70870 36732
rect 70928 36686 70974 36732
rect 21438 36594 21484 36640
rect 70824 36582 70870 36628
rect 70928 36582 70974 36628
rect 21570 36462 21616 36508
rect 70824 36478 70870 36524
rect 70928 36478 70974 36524
rect 21702 36330 21748 36376
rect 70824 36374 70870 36420
rect 70928 36374 70974 36420
rect 21834 36198 21880 36244
rect 70824 36270 70870 36316
rect 70928 36270 70974 36316
rect 70824 36166 70870 36212
rect 70928 36166 70974 36212
rect 21966 36066 22012 36112
rect 70824 36062 70870 36108
rect 70928 36062 70974 36108
rect 22098 35934 22144 35980
rect 70824 35958 70870 36004
rect 70928 35958 70974 36004
rect 22230 35802 22276 35848
rect 70824 35854 70870 35900
rect 70928 35854 70974 35900
rect 70824 35750 70870 35796
rect 70928 35750 70974 35796
rect 22362 35670 22408 35716
rect 70824 35646 70870 35692
rect 70928 35646 70974 35692
rect 22494 35538 22540 35584
rect 70824 35542 70870 35588
rect 70928 35542 70974 35588
rect 22626 35406 22672 35452
rect 70824 35438 70870 35484
rect 70928 35438 70974 35484
rect 22758 35274 22804 35320
rect 70824 35334 70870 35380
rect 70928 35334 70974 35380
rect 70824 35230 70870 35276
rect 70928 35230 70974 35276
rect 22890 35142 22936 35188
rect 70824 35126 70870 35172
rect 70928 35126 70974 35172
rect 23022 35010 23068 35056
rect 70824 35022 70870 35068
rect 70928 35022 70974 35068
rect 23154 34878 23200 34924
rect 70824 34918 70870 34964
rect 70928 34918 70974 34964
rect 70824 34814 70870 34860
rect 70928 34814 70974 34860
rect 23286 34746 23332 34792
rect 70824 34710 70870 34756
rect 70928 34710 70974 34756
rect 23418 34614 23464 34660
rect 70824 34606 70870 34652
rect 70928 34606 70974 34652
rect 23550 34482 23596 34528
rect 70824 34502 70870 34548
rect 70928 34502 70974 34548
rect 23682 34350 23728 34396
rect 70824 34398 70870 34444
rect 70928 34398 70974 34444
rect 70824 34294 70870 34340
rect 70928 34294 70974 34340
rect 23814 34218 23860 34264
rect 70824 34190 70870 34236
rect 70928 34190 70974 34236
rect 23946 34086 23992 34132
rect 70824 34086 70870 34132
rect 70928 34086 70974 34132
rect 24078 33954 24124 34000
rect 70824 33982 70870 34028
rect 70928 33982 70974 34028
rect 24210 33822 24256 33868
rect 70824 33878 70870 33924
rect 70928 33878 70974 33924
rect 70824 33774 70870 33820
rect 70928 33774 70974 33820
rect 24342 33690 24388 33736
rect 70824 33670 70870 33716
rect 70928 33670 70974 33716
rect 24474 33558 24520 33604
rect 70824 33566 70870 33612
rect 70928 33566 70974 33612
rect 24606 33426 24652 33472
rect 70824 33462 70870 33508
rect 70928 33462 70974 33508
rect 24738 33294 24784 33340
rect 70824 33358 70870 33404
rect 70928 33358 70974 33404
rect 70824 33254 70870 33300
rect 70928 33254 70974 33300
rect 24870 33162 24916 33208
rect 70824 33150 70870 33196
rect 70928 33150 70974 33196
rect 25002 33030 25048 33076
rect 70824 33046 70870 33092
rect 70928 33046 70974 33092
rect 25134 32898 25180 32944
rect 70824 32942 70870 32988
rect 70928 32942 70974 32988
rect 70824 32838 70870 32884
rect 70928 32838 70974 32884
rect 25266 32766 25312 32812
rect 70824 32734 70870 32780
rect 70928 32734 70974 32780
rect 25398 32634 25444 32680
rect 70824 32630 70870 32676
rect 70928 32630 70974 32676
rect 25530 32502 25576 32548
rect 70824 32526 70870 32572
rect 70928 32526 70974 32572
rect 70824 32422 70870 32468
rect 70928 32422 70974 32468
rect 25662 32370 25708 32416
rect 25794 32238 25840 32284
rect 70824 32318 70870 32364
rect 70928 32318 70974 32364
rect 70824 32214 70870 32260
rect 70928 32214 70974 32260
rect 25926 32106 25972 32152
rect 70824 32110 70870 32156
rect 70928 32110 70974 32156
rect 26058 31974 26104 32020
rect 70824 32006 70870 32052
rect 70928 32006 70974 32052
rect 26190 31842 26236 31888
rect 70824 31902 70870 31948
rect 70928 31902 70974 31948
rect 70824 31798 70870 31844
rect 70928 31798 70974 31844
rect 26322 31710 26368 31756
rect 70824 31694 70870 31740
rect 70928 31694 70974 31740
rect 26454 31578 26500 31624
rect 70824 31590 70870 31636
rect 70928 31590 70974 31636
rect 26586 31446 26632 31492
rect 70824 31486 70870 31532
rect 70928 31486 70974 31532
rect 70824 31382 70870 31428
rect 70928 31382 70974 31428
rect 26718 31314 26764 31360
rect 70824 31278 70870 31324
rect 70928 31278 70974 31324
rect 26850 31182 26896 31228
rect 70824 31174 70870 31220
rect 70928 31174 70974 31220
rect 26982 31050 27028 31096
rect 70824 31070 70870 31116
rect 70928 31070 70974 31116
rect 27114 30918 27160 30964
rect 70824 30966 70870 31012
rect 70928 30966 70974 31012
rect 70824 30862 70870 30908
rect 70928 30862 70974 30908
rect 27246 30786 27292 30832
rect 70824 30758 70870 30804
rect 70928 30758 70974 30804
rect 27378 30654 27424 30700
rect 70824 30654 70870 30700
rect 70928 30654 70974 30700
rect 27510 30522 27556 30568
rect 70824 30550 70870 30596
rect 70928 30550 70974 30596
rect 70824 30446 70870 30492
rect 70928 30446 70974 30492
rect 27642 30390 27688 30436
rect 70824 30342 70870 30388
rect 70928 30342 70974 30388
rect 27774 30258 27820 30304
rect 70824 30238 70870 30284
rect 70928 30238 70974 30284
rect 27906 30126 27952 30172
rect 70824 30134 70870 30180
rect 70928 30134 70974 30180
rect 28038 29994 28084 30040
rect 70824 30030 70870 30076
rect 70928 30030 70974 30076
rect 28170 29862 28216 29908
rect 70824 29926 70870 29972
rect 70928 29926 70974 29972
rect 70824 29822 70870 29868
rect 70928 29822 70974 29868
rect 28302 29730 28348 29776
rect 70824 29718 70870 29764
rect 70928 29718 70974 29764
rect 28434 29598 28480 29644
rect 70824 29614 70870 29660
rect 70928 29614 70974 29660
rect 28566 29466 28612 29512
rect 70824 29510 70870 29556
rect 70928 29510 70974 29556
rect 70824 29406 70870 29452
rect 70928 29406 70974 29452
rect 28698 29334 28744 29380
rect 70824 29302 70870 29348
rect 70928 29302 70974 29348
rect 28830 29202 28876 29248
rect 70824 29198 70870 29244
rect 70928 29198 70974 29244
rect 28962 29070 29008 29116
rect 70824 29094 70870 29140
rect 70928 29094 70974 29140
rect 29094 28938 29140 28984
rect 70824 28990 70870 29036
rect 70928 28990 70974 29036
rect 70824 28886 70870 28932
rect 70928 28886 70974 28932
rect 29226 28806 29272 28852
rect 70824 28782 70870 28828
rect 70928 28782 70974 28828
rect 29358 28674 29404 28720
rect 70824 28678 70870 28724
rect 70928 28678 70974 28724
rect 29490 28542 29536 28588
rect 70824 28574 70870 28620
rect 70928 28574 70974 28620
rect 29622 28410 29668 28456
rect 70824 28470 70870 28516
rect 70928 28470 70974 28516
rect 70824 28366 70870 28412
rect 70928 28366 70974 28412
rect 29754 28278 29800 28324
rect 70824 28262 70870 28308
rect 70928 28262 70974 28308
rect 29886 28146 29932 28192
rect 70824 28158 70870 28204
rect 70928 28158 70974 28204
rect 30018 28014 30064 28060
rect 70824 28054 70870 28100
rect 70928 28054 70974 28100
rect 30150 27882 30196 27928
rect 70824 27950 70870 27996
rect 70928 27950 70974 27996
rect 70824 27846 70870 27892
rect 70928 27846 70974 27892
rect 30282 27750 30328 27796
rect 70824 27742 70870 27788
rect 70928 27742 70974 27788
rect 30414 27618 30460 27664
rect 70824 27638 70870 27684
rect 70928 27638 70974 27684
rect 30546 27486 30592 27532
rect 70824 27534 70870 27580
rect 70928 27534 70974 27580
rect 70824 27430 70870 27476
rect 70928 27430 70974 27476
rect 30678 27354 30724 27400
rect 70824 27326 70870 27372
rect 70928 27326 70974 27372
rect 30810 27222 30856 27268
rect 70824 27222 70870 27268
rect 70928 27222 70974 27268
rect 30942 27090 30988 27136
rect 70824 27118 70870 27164
rect 70928 27118 70974 27164
rect 31074 26958 31120 27004
rect 70824 27014 70870 27060
rect 70928 27014 70974 27060
rect 70824 26910 70870 26956
rect 70928 26910 70974 26956
rect 31206 26826 31252 26872
rect 70824 26806 70870 26852
rect 70928 26806 70974 26852
rect 31338 26694 31384 26740
rect 70824 26702 70870 26748
rect 70928 26702 70974 26748
rect 31470 26562 31516 26608
rect 70824 26598 70870 26644
rect 70928 26598 70974 26644
rect 31602 26430 31648 26476
rect 70824 26494 70870 26540
rect 70928 26494 70974 26540
rect 70824 26390 70870 26436
rect 70928 26390 70974 26436
rect 31734 26298 31780 26344
rect 70824 26286 70870 26332
rect 70928 26286 70974 26332
rect 31866 26166 31912 26212
rect 70824 26182 70870 26228
rect 70928 26182 70974 26228
rect 31998 26034 32044 26080
rect 70824 26078 70870 26124
rect 70928 26078 70974 26124
rect 70824 25974 70870 26020
rect 70928 25974 70974 26020
rect 32130 25902 32176 25948
rect 70824 25870 70870 25916
rect 70928 25870 70974 25916
rect 32262 25770 32308 25816
rect 70824 25766 70870 25812
rect 70928 25766 70974 25812
rect 32394 25638 32440 25684
rect 70824 25662 70870 25708
rect 70928 25662 70974 25708
rect 32526 25506 32572 25552
rect 70824 25558 70870 25604
rect 70928 25558 70974 25604
rect 32658 25374 32704 25420
rect 70824 25454 70870 25500
rect 70928 25454 70974 25500
rect 70824 25350 70870 25396
rect 70928 25350 70974 25396
rect 32790 25242 32836 25288
rect 70824 25246 70870 25292
rect 70928 25246 70974 25292
rect 32922 25110 32968 25156
rect 70824 25142 70870 25188
rect 70928 25142 70974 25188
rect 33054 24978 33100 25024
rect 70824 25038 70870 25084
rect 70928 25038 70974 25084
rect 70824 24934 70870 24980
rect 70928 24934 70974 24980
rect 33186 24846 33232 24892
rect 70824 24830 70870 24876
rect 70928 24830 70974 24876
rect 33318 24714 33364 24760
rect 70824 24726 70870 24772
rect 70928 24726 70974 24772
rect 33450 24582 33496 24628
rect 70824 24622 70870 24668
rect 70928 24622 70974 24668
rect 70824 24518 70870 24564
rect 70928 24518 70974 24564
rect 33582 24450 33628 24496
rect 70824 24414 70870 24460
rect 70928 24414 70974 24460
rect 33714 24318 33760 24364
rect 70824 24310 70870 24356
rect 70928 24310 70974 24356
rect 33846 24186 33892 24232
rect 70824 24206 70870 24252
rect 70928 24206 70974 24252
rect 33978 24054 34024 24100
rect 70824 24102 70870 24148
rect 70928 24102 70974 24148
rect 34110 23922 34156 23968
rect 70824 23998 70870 24044
rect 70928 23998 70974 24044
rect 70824 23894 70870 23940
rect 70928 23894 70974 23940
rect 34242 23790 34288 23836
rect 70824 23790 70870 23836
rect 70928 23790 70974 23836
rect 34374 23658 34420 23704
rect 70824 23686 70870 23732
rect 70928 23686 70974 23732
rect 34506 23526 34552 23572
rect 70824 23582 70870 23628
rect 70928 23582 70974 23628
rect 70824 23478 70870 23524
rect 70928 23478 70974 23524
rect 34638 23394 34684 23440
rect 70824 23374 70870 23420
rect 70928 23374 70974 23420
rect 34770 23262 34816 23308
rect 70824 23270 70870 23316
rect 70928 23270 70974 23316
rect 34902 23130 34948 23176
rect 70824 23166 70870 23212
rect 70928 23166 70974 23212
rect 35034 22998 35080 23044
rect 70824 23062 70870 23108
rect 70928 23062 70974 23108
rect 70824 22958 70870 23004
rect 70928 22958 70974 23004
rect 35166 22866 35212 22912
rect 70824 22854 70870 22900
rect 70928 22854 70974 22900
rect 35298 22734 35344 22780
rect 70824 22750 70870 22796
rect 70928 22750 70974 22796
rect 35430 22602 35476 22648
rect 70824 22646 70870 22692
rect 70928 22646 70974 22692
rect 70824 22542 70870 22588
rect 70928 22542 70974 22588
rect 35562 22470 35608 22516
rect 70824 22438 70870 22484
rect 70928 22438 70974 22484
rect 35694 22338 35740 22384
rect 70824 22334 70870 22380
rect 70928 22334 70974 22380
rect 35826 22206 35872 22252
rect 70824 22230 70870 22276
rect 70928 22230 70974 22276
rect 70824 22126 70870 22172
rect 70928 22126 70974 22172
rect 35958 22074 36004 22120
rect 70824 22022 70870 22068
rect 70928 22022 70974 22068
rect 36090 21942 36136 21988
rect 70824 21918 70870 21964
rect 70928 21918 70974 21964
rect 36222 21810 36268 21856
rect 70824 21814 70870 21860
rect 70928 21814 70974 21860
rect 36354 21678 36400 21724
rect 70824 21710 70870 21756
rect 70928 21710 70974 21756
rect 36486 21546 36532 21592
rect 70824 21606 70870 21652
rect 70928 21606 70974 21652
rect 70824 21502 70870 21548
rect 70928 21502 70974 21548
rect 36618 21414 36664 21460
rect 70824 21398 70870 21444
rect 70928 21398 70974 21444
rect 36750 21282 36796 21328
rect 70824 21294 70870 21340
rect 70928 21294 70974 21340
rect 36882 21150 36928 21196
rect 70824 21190 70870 21236
rect 70928 21190 70974 21236
rect 70824 21086 70870 21132
rect 70928 21086 70974 21132
rect 37014 21018 37060 21064
rect 70824 20982 70870 21028
rect 70928 20982 70974 21028
rect 37146 20886 37192 20932
rect 70824 20878 70870 20924
rect 70928 20878 70974 20924
rect 37278 20754 37324 20800
rect 70824 20774 70870 20820
rect 70928 20774 70974 20820
rect 37410 20622 37456 20668
rect 70824 20670 70870 20716
rect 70928 20670 70974 20716
rect 70824 20566 70870 20612
rect 70928 20566 70974 20612
rect 37542 20490 37588 20536
rect 70824 20462 70870 20508
rect 70928 20462 70974 20508
rect 37674 20358 37720 20404
rect 70824 20358 70870 20404
rect 70928 20358 70974 20404
rect 37806 20226 37852 20272
rect 70824 20254 70870 20300
rect 70928 20254 70974 20300
rect 37938 20094 37984 20140
rect 70824 20150 70870 20196
rect 70928 20150 70974 20196
rect 70824 20046 70870 20092
rect 70928 20046 70974 20092
rect 38070 19962 38116 20008
rect 70824 19942 70870 19988
rect 70928 19942 70974 19988
rect 38202 19830 38248 19876
rect 70824 19838 70870 19884
rect 70928 19838 70974 19884
rect 38334 19698 38380 19744
rect 70824 19734 70870 19780
rect 70928 19734 70974 19780
rect 38466 19566 38512 19612
rect 70824 19630 70870 19676
rect 70928 19630 70974 19676
rect 70824 19526 70870 19572
rect 70928 19526 70974 19572
rect 38598 19434 38644 19480
rect 70824 19422 70870 19468
rect 70928 19422 70974 19468
rect 38730 19302 38776 19348
rect 70824 19318 70870 19364
rect 70928 19318 70974 19364
rect 38862 19170 38908 19216
rect 70824 19214 70870 19260
rect 70928 19214 70974 19260
rect 38994 19038 39040 19084
rect 70824 19110 70870 19156
rect 70928 19110 70974 19156
rect 70824 19006 70870 19052
rect 70928 19006 70974 19052
rect 39126 18906 39172 18952
rect 70824 18902 70870 18948
rect 70928 18902 70974 18948
rect 39258 18774 39304 18820
rect 70824 18798 70870 18844
rect 70928 18798 70974 18844
rect 39390 18642 39436 18688
rect 70824 18694 70870 18740
rect 70928 18694 70974 18740
rect 39522 18510 39568 18556
rect 70824 18590 70870 18636
rect 70928 18590 70974 18636
rect 70824 18486 70870 18532
rect 70928 18486 70974 18532
rect 39654 18378 39700 18424
rect 70824 18382 70870 18428
rect 70928 18382 70974 18428
rect 39786 18246 39832 18292
rect 70824 18278 70870 18324
rect 70928 18278 70974 18324
rect 39918 18114 39964 18160
rect 70824 18174 70870 18220
rect 70928 18174 70974 18220
rect 70824 18070 70870 18116
rect 70928 18070 70974 18116
rect 40050 17982 40096 18028
rect 70824 17966 70870 18012
rect 70928 17966 70974 18012
rect 40182 17850 40228 17896
rect 70824 17862 70870 17908
rect 70928 17862 70974 17908
rect 40314 17718 40360 17764
rect 70824 17758 70870 17804
rect 70928 17758 70974 17804
rect 70824 17654 70870 17700
rect 70928 17654 70974 17700
rect 40446 17586 40492 17632
rect 70824 17550 70870 17596
rect 70928 17550 70974 17596
rect 40578 17454 40624 17500
rect 70824 17446 70870 17492
rect 70928 17446 70974 17492
rect 40710 17322 40756 17368
rect 70824 17342 70870 17388
rect 70928 17342 70974 17388
rect 70824 17238 70870 17284
rect 70928 17238 70974 17284
rect 40842 17190 40888 17236
rect 40974 17058 41020 17104
rect 70824 17134 70870 17180
rect 70928 17134 70974 17180
rect 70824 17030 70870 17076
rect 70928 17030 70974 17076
rect 41106 16926 41152 16972
rect 70824 16926 70870 16972
rect 70928 16926 70974 16972
rect 41238 16794 41284 16840
rect 70824 16822 70870 16868
rect 70928 16822 70974 16868
rect 41370 16662 41416 16708
rect 70824 16718 70870 16764
rect 70928 16718 70974 16764
rect 70824 16614 70870 16660
rect 70928 16614 70974 16660
rect 41502 16530 41548 16576
rect 70824 16510 70870 16556
rect 70928 16510 70974 16556
rect 41634 16398 41680 16444
rect 70824 16406 70870 16452
rect 70928 16406 70974 16452
rect 41766 16266 41812 16312
rect 70824 16302 70870 16348
rect 70928 16302 70974 16348
rect 41898 16134 41944 16180
rect 70824 16198 70870 16244
rect 70928 16198 70974 16244
rect 70824 16094 70870 16140
rect 70928 16094 70974 16140
rect 42030 16002 42076 16048
rect 70824 15990 70870 16036
rect 70928 15990 70974 16036
rect 42162 15870 42208 15916
rect 70824 15886 70870 15932
rect 70928 15886 70974 15932
rect 42294 15738 42340 15784
rect 70824 15782 70870 15828
rect 70928 15782 70974 15828
rect 70824 15678 70870 15724
rect 70928 15678 70974 15724
rect 42426 15606 42472 15652
rect 70824 15574 70870 15620
rect 70928 15574 70974 15620
rect 42558 15474 42604 15520
rect 70824 15470 70870 15516
rect 70928 15470 70974 15516
rect 42690 15342 42736 15388
rect 70824 15366 70870 15412
rect 70928 15366 70974 15412
rect 70824 15262 70870 15308
rect 70928 15262 70974 15308
rect 42822 15210 42868 15256
rect 70824 15158 70870 15204
rect 70928 15158 70974 15204
rect 42954 15078 43000 15124
rect 70824 15054 70870 15100
rect 70928 15054 70974 15100
rect 43086 14946 43132 14992
rect 70824 14950 70870 14996
rect 70928 14950 70974 14996
rect 43218 14814 43264 14860
rect 70824 14846 70870 14892
rect 70928 14846 70974 14892
rect 43350 14682 43396 14728
rect 70824 14742 70870 14788
rect 70928 14742 70974 14788
rect 70824 14638 70870 14684
rect 70928 14638 70974 14684
rect 43482 14550 43528 14596
rect 70824 14534 70870 14580
rect 70928 14534 70974 14580
rect 43614 14418 43660 14464
rect 70824 14430 70870 14476
rect 70928 14430 70974 14476
rect 43746 14286 43792 14332
rect 70824 14326 70870 14372
rect 70928 14326 70974 14372
rect 70824 14222 70870 14268
rect 70928 14222 70974 14268
rect 43878 14154 43924 14200
rect 70824 14118 70870 14164
rect 70928 14118 70974 14164
rect 44010 14022 44056 14068
rect 70824 14014 70870 14060
rect 70928 14014 70974 14060
rect 44142 13890 44188 13936
rect 70824 13910 70870 13956
rect 70928 13910 70974 13956
rect 44274 13758 44320 13804
rect 70824 13806 70870 13852
rect 70928 13806 70974 13852
rect 70824 13702 70870 13748
rect 70928 13702 70974 13748
rect 44406 13626 44452 13672
rect 70824 13598 70870 13644
rect 70928 13598 70974 13644
rect 44538 13494 44584 13540
rect 70824 13494 70870 13540
rect 70928 13494 70974 13540
rect 44670 13362 44716 13408
rect 70824 13390 70870 13436
rect 70928 13390 70974 13436
rect 44850 13210 44896 13256
rect 45088 13223 45134 13269
rect 45192 13223 45238 13269
rect 45296 13223 45342 13269
rect 45400 13223 45446 13269
rect 45504 13223 45550 13269
rect 45608 13223 45654 13269
rect 45712 13223 45758 13269
rect 45816 13223 45862 13269
rect 45920 13223 45966 13269
rect 46024 13223 46070 13269
rect 46128 13223 46174 13269
rect 46232 13223 46278 13269
rect 46336 13223 46382 13269
rect 46440 13223 46486 13269
rect 46544 13223 46590 13269
rect 46648 13223 46694 13269
rect 46752 13223 46798 13269
rect 46856 13223 46902 13269
rect 46960 13223 47006 13269
rect 47064 13223 47110 13269
rect 47168 13223 47214 13269
rect 47272 13223 47318 13269
rect 47376 13223 47422 13269
rect 47480 13223 47526 13269
rect 47584 13223 47630 13269
rect 47688 13223 47734 13269
rect 47792 13223 47838 13269
rect 47896 13223 47942 13269
rect 48000 13223 48046 13269
rect 48104 13223 48150 13269
rect 48208 13223 48254 13269
rect 48312 13223 48358 13269
rect 48416 13223 48462 13269
rect 48520 13223 48566 13269
rect 48624 13223 48670 13269
rect 48728 13223 48774 13269
rect 48832 13223 48878 13269
rect 48936 13223 48982 13269
rect 49040 13223 49086 13269
rect 49144 13223 49190 13269
rect 49248 13223 49294 13269
rect 49352 13223 49398 13269
rect 49456 13223 49502 13269
rect 49560 13223 49606 13269
rect 49664 13223 49710 13269
rect 49768 13223 49814 13269
rect 49872 13223 49918 13269
rect 49976 13223 50022 13269
rect 50080 13223 50126 13269
rect 50184 13223 50230 13269
rect 50288 13223 50334 13269
rect 50392 13223 50438 13269
rect 50496 13223 50542 13269
rect 50600 13223 50646 13269
rect 50704 13223 50750 13269
rect 50808 13223 50854 13269
rect 50912 13223 50958 13269
rect 51016 13223 51062 13269
rect 51120 13223 51166 13269
rect 51224 13223 51270 13269
rect 51328 13223 51374 13269
rect 51432 13223 51478 13269
rect 51536 13223 51582 13269
rect 51640 13223 51686 13269
rect 51744 13223 51790 13269
rect 51848 13223 51894 13269
rect 51952 13223 51998 13269
rect 52056 13223 52102 13269
rect 52160 13223 52206 13269
rect 52264 13223 52310 13269
rect 52368 13223 52414 13269
rect 52472 13223 52518 13269
rect 52576 13223 52622 13269
rect 52680 13223 52726 13269
rect 52784 13223 52830 13269
rect 52888 13223 52934 13269
rect 52992 13223 53038 13269
rect 53096 13223 53142 13269
rect 53200 13223 53246 13269
rect 53304 13223 53350 13269
rect 53408 13223 53454 13269
rect 53512 13223 53558 13269
rect 53616 13223 53662 13269
rect 53720 13223 53766 13269
rect 53824 13223 53870 13269
rect 53928 13223 53974 13269
rect 54032 13223 54078 13269
rect 54136 13223 54182 13269
rect 54240 13223 54286 13269
rect 54344 13223 54390 13269
rect 54448 13223 54494 13269
rect 54552 13223 54598 13269
rect 54656 13223 54702 13269
rect 54760 13223 54806 13269
rect 54864 13223 54910 13269
rect 54968 13223 55014 13269
rect 55072 13223 55118 13269
rect 55176 13223 55222 13269
rect 55280 13223 55326 13269
rect 55384 13223 55430 13269
rect 55488 13223 55534 13269
rect 55592 13223 55638 13269
rect 55696 13223 55742 13269
rect 55800 13223 55846 13269
rect 55904 13223 55950 13269
rect 56008 13223 56054 13269
rect 56112 13223 56158 13269
rect 56216 13223 56262 13269
rect 56320 13223 56366 13269
rect 56424 13223 56470 13269
rect 56528 13223 56574 13269
rect 56632 13223 56678 13269
rect 56736 13223 56782 13269
rect 56840 13223 56886 13269
rect 56944 13223 56990 13269
rect 57048 13223 57094 13269
rect 57152 13223 57198 13269
rect 57256 13223 57302 13269
rect 57360 13223 57406 13269
rect 57464 13223 57510 13269
rect 57568 13223 57614 13269
rect 57672 13223 57718 13269
rect 57776 13223 57822 13269
rect 57880 13223 57926 13269
rect 57984 13223 58030 13269
rect 58088 13223 58134 13269
rect 58192 13223 58238 13269
rect 58296 13223 58342 13269
rect 58400 13223 58446 13269
rect 58504 13223 58550 13269
rect 58608 13223 58654 13269
rect 58712 13223 58758 13269
rect 58816 13223 58862 13269
rect 58920 13223 58966 13269
rect 59024 13223 59070 13269
rect 59128 13223 59174 13269
rect 59232 13223 59278 13269
rect 59336 13223 59382 13269
rect 59440 13223 59486 13269
rect 59544 13223 59590 13269
rect 59648 13223 59694 13269
rect 59752 13223 59798 13269
rect 59856 13223 59902 13269
rect 59960 13223 60006 13269
rect 60064 13223 60110 13269
rect 60168 13223 60214 13269
rect 60272 13223 60318 13269
rect 60376 13223 60422 13269
rect 60480 13223 60526 13269
rect 60584 13223 60630 13269
rect 60688 13223 60734 13269
rect 60792 13223 60838 13269
rect 60896 13223 60942 13269
rect 61000 13223 61046 13269
rect 61104 13223 61150 13269
rect 61208 13223 61254 13269
rect 61312 13223 61358 13269
rect 61416 13223 61462 13269
rect 61520 13223 61566 13269
rect 61624 13223 61670 13269
rect 61728 13223 61774 13269
rect 61832 13223 61878 13269
rect 61936 13223 61982 13269
rect 62040 13223 62086 13269
rect 62144 13223 62190 13269
rect 62248 13223 62294 13269
rect 62352 13223 62398 13269
rect 62456 13223 62502 13269
rect 62560 13223 62606 13269
rect 62664 13223 62710 13269
rect 62768 13223 62814 13269
rect 62872 13223 62918 13269
rect 62976 13223 63022 13269
rect 63080 13223 63126 13269
rect 63184 13223 63230 13269
rect 63288 13223 63334 13269
rect 63392 13223 63438 13269
rect 63496 13223 63542 13269
rect 63600 13223 63646 13269
rect 63704 13223 63750 13269
rect 63808 13223 63854 13269
rect 63912 13223 63958 13269
rect 64016 13223 64062 13269
rect 64120 13223 64166 13269
rect 64224 13223 64270 13269
rect 64328 13223 64374 13269
rect 64432 13223 64478 13269
rect 64536 13223 64582 13269
rect 64640 13223 64686 13269
rect 64744 13223 64790 13269
rect 64848 13223 64894 13269
rect 64952 13223 64998 13269
rect 65056 13223 65102 13269
rect 65160 13223 65206 13269
rect 65264 13223 65310 13269
rect 65368 13223 65414 13269
rect 65472 13223 65518 13269
rect 65576 13223 65622 13269
rect 65680 13223 65726 13269
rect 65784 13223 65830 13269
rect 65888 13223 65934 13269
rect 65992 13223 66038 13269
rect 66096 13223 66142 13269
rect 66200 13223 66246 13269
rect 66304 13223 66350 13269
rect 66408 13223 66454 13269
rect 66512 13223 66558 13269
rect 66616 13223 66662 13269
rect 66720 13223 66766 13269
rect 66824 13223 66870 13269
rect 66928 13223 66974 13269
rect 67032 13223 67078 13269
rect 67136 13223 67182 13269
rect 67240 13223 67286 13269
rect 67344 13223 67390 13269
rect 67448 13223 67494 13269
rect 67552 13223 67598 13269
rect 67656 13223 67702 13269
rect 67760 13223 67806 13269
rect 67864 13223 67910 13269
rect 67968 13223 68014 13269
rect 68072 13223 68118 13269
rect 68176 13223 68222 13269
rect 68280 13223 68326 13269
rect 68384 13223 68430 13269
rect 68488 13223 68534 13269
rect 68592 13223 68638 13269
rect 68696 13223 68742 13269
rect 68800 13223 68846 13269
rect 68904 13223 68950 13269
rect 69008 13223 69054 13269
rect 69112 13223 69158 13269
rect 69216 13223 69262 13269
rect 69320 13223 69366 13269
rect 69424 13223 69470 13269
rect 69528 13223 69574 13269
rect 69632 13223 69678 13269
rect 69736 13223 69782 13269
rect 69840 13223 69886 13269
rect 69944 13223 69990 13269
rect 70048 13223 70094 13269
rect 70152 13223 70198 13269
rect 70256 13223 70302 13269
rect 70360 13223 70406 13269
rect 70464 13223 70510 13269
rect 70568 13223 70614 13269
rect 70672 13223 70718 13269
rect 70776 13223 70822 13269
rect 70880 13223 70926 13269
rect 45088 13119 45134 13165
rect 45192 13119 45238 13165
rect 45296 13119 45342 13165
rect 45400 13119 45446 13165
rect 45504 13119 45550 13165
rect 45608 13119 45654 13165
rect 45712 13119 45758 13165
rect 45816 13119 45862 13165
rect 45920 13119 45966 13165
rect 46024 13119 46070 13165
rect 46128 13119 46174 13165
rect 46232 13119 46278 13165
rect 46336 13119 46382 13165
rect 46440 13119 46486 13165
rect 46544 13119 46590 13165
rect 46648 13119 46694 13165
rect 46752 13119 46798 13165
rect 46856 13119 46902 13165
rect 46960 13119 47006 13165
rect 47064 13119 47110 13165
rect 47168 13119 47214 13165
rect 47272 13119 47318 13165
rect 47376 13119 47422 13165
rect 47480 13119 47526 13165
rect 47584 13119 47630 13165
rect 47688 13119 47734 13165
rect 47792 13119 47838 13165
rect 47896 13119 47942 13165
rect 48000 13119 48046 13165
rect 48104 13119 48150 13165
rect 48208 13119 48254 13165
rect 48312 13119 48358 13165
rect 48416 13119 48462 13165
rect 48520 13119 48566 13165
rect 48624 13119 48670 13165
rect 48728 13119 48774 13165
rect 48832 13119 48878 13165
rect 48936 13119 48982 13165
rect 49040 13119 49086 13165
rect 49144 13119 49190 13165
rect 49248 13119 49294 13165
rect 49352 13119 49398 13165
rect 49456 13119 49502 13165
rect 49560 13119 49606 13165
rect 49664 13119 49710 13165
rect 49768 13119 49814 13165
rect 49872 13119 49918 13165
rect 49976 13119 50022 13165
rect 50080 13119 50126 13165
rect 50184 13119 50230 13165
rect 50288 13119 50334 13165
rect 50392 13119 50438 13165
rect 50496 13119 50542 13165
rect 50600 13119 50646 13165
rect 50704 13119 50750 13165
rect 50808 13119 50854 13165
rect 50912 13119 50958 13165
rect 51016 13119 51062 13165
rect 51120 13119 51166 13165
rect 51224 13119 51270 13165
rect 51328 13119 51374 13165
rect 51432 13119 51478 13165
rect 51536 13119 51582 13165
rect 51640 13119 51686 13165
rect 51744 13119 51790 13165
rect 51848 13119 51894 13165
rect 51952 13119 51998 13165
rect 52056 13119 52102 13165
rect 52160 13119 52206 13165
rect 52264 13119 52310 13165
rect 52368 13119 52414 13165
rect 52472 13119 52518 13165
rect 52576 13119 52622 13165
rect 52680 13119 52726 13165
rect 52784 13119 52830 13165
rect 52888 13119 52934 13165
rect 52992 13119 53038 13165
rect 53096 13119 53142 13165
rect 53200 13119 53246 13165
rect 53304 13119 53350 13165
rect 53408 13119 53454 13165
rect 53512 13119 53558 13165
rect 53616 13119 53662 13165
rect 53720 13119 53766 13165
rect 53824 13119 53870 13165
rect 53928 13119 53974 13165
rect 54032 13119 54078 13165
rect 54136 13119 54182 13165
rect 54240 13119 54286 13165
rect 54344 13119 54390 13165
rect 54448 13119 54494 13165
rect 54552 13119 54598 13165
rect 54656 13119 54702 13165
rect 54760 13119 54806 13165
rect 54864 13119 54910 13165
rect 54968 13119 55014 13165
rect 55072 13119 55118 13165
rect 55176 13119 55222 13165
rect 55280 13119 55326 13165
rect 55384 13119 55430 13165
rect 55488 13119 55534 13165
rect 55592 13119 55638 13165
rect 55696 13119 55742 13165
rect 55800 13119 55846 13165
rect 55904 13119 55950 13165
rect 56008 13119 56054 13165
rect 56112 13119 56158 13165
rect 56216 13119 56262 13165
rect 56320 13119 56366 13165
rect 56424 13119 56470 13165
rect 56528 13119 56574 13165
rect 56632 13119 56678 13165
rect 56736 13119 56782 13165
rect 56840 13119 56886 13165
rect 56944 13119 56990 13165
rect 57048 13119 57094 13165
rect 57152 13119 57198 13165
rect 57256 13119 57302 13165
rect 57360 13119 57406 13165
rect 57464 13119 57510 13165
rect 57568 13119 57614 13165
rect 57672 13119 57718 13165
rect 57776 13119 57822 13165
rect 57880 13119 57926 13165
rect 57984 13119 58030 13165
rect 58088 13119 58134 13165
rect 58192 13119 58238 13165
rect 58296 13119 58342 13165
rect 58400 13119 58446 13165
rect 58504 13119 58550 13165
rect 58608 13119 58654 13165
rect 58712 13119 58758 13165
rect 58816 13119 58862 13165
rect 58920 13119 58966 13165
rect 59024 13119 59070 13165
rect 59128 13119 59174 13165
rect 59232 13119 59278 13165
rect 59336 13119 59382 13165
rect 59440 13119 59486 13165
rect 59544 13119 59590 13165
rect 59648 13119 59694 13165
rect 59752 13119 59798 13165
rect 59856 13119 59902 13165
rect 59960 13119 60006 13165
rect 60064 13119 60110 13165
rect 60168 13119 60214 13165
rect 60272 13119 60318 13165
rect 60376 13119 60422 13165
rect 60480 13119 60526 13165
rect 60584 13119 60630 13165
rect 60688 13119 60734 13165
rect 60792 13119 60838 13165
rect 60896 13119 60942 13165
rect 61000 13119 61046 13165
rect 61104 13119 61150 13165
rect 61208 13119 61254 13165
rect 61312 13119 61358 13165
rect 61416 13119 61462 13165
rect 61520 13119 61566 13165
rect 61624 13119 61670 13165
rect 61728 13119 61774 13165
rect 61832 13119 61878 13165
rect 61936 13119 61982 13165
rect 62040 13119 62086 13165
rect 62144 13119 62190 13165
rect 62248 13119 62294 13165
rect 62352 13119 62398 13165
rect 62456 13119 62502 13165
rect 62560 13119 62606 13165
rect 62664 13119 62710 13165
rect 62768 13119 62814 13165
rect 62872 13119 62918 13165
rect 62976 13119 63022 13165
rect 63080 13119 63126 13165
rect 63184 13119 63230 13165
rect 63288 13119 63334 13165
rect 63392 13119 63438 13165
rect 63496 13119 63542 13165
rect 63600 13119 63646 13165
rect 63704 13119 63750 13165
rect 63808 13119 63854 13165
rect 63912 13119 63958 13165
rect 64016 13119 64062 13165
rect 64120 13119 64166 13165
rect 64224 13119 64270 13165
rect 64328 13119 64374 13165
rect 64432 13119 64478 13165
rect 64536 13119 64582 13165
rect 64640 13119 64686 13165
rect 64744 13119 64790 13165
rect 64848 13119 64894 13165
rect 64952 13119 64998 13165
rect 65056 13119 65102 13165
rect 65160 13119 65206 13165
rect 65264 13119 65310 13165
rect 65368 13119 65414 13165
rect 65472 13119 65518 13165
rect 65576 13119 65622 13165
rect 65680 13119 65726 13165
rect 65784 13119 65830 13165
rect 65888 13119 65934 13165
rect 65992 13119 66038 13165
rect 66096 13119 66142 13165
rect 66200 13119 66246 13165
rect 66304 13119 66350 13165
rect 66408 13119 66454 13165
rect 66512 13119 66558 13165
rect 66616 13119 66662 13165
rect 66720 13119 66766 13165
rect 66824 13119 66870 13165
rect 66928 13119 66974 13165
rect 67032 13119 67078 13165
rect 67136 13119 67182 13165
rect 67240 13119 67286 13165
rect 67344 13119 67390 13165
rect 67448 13119 67494 13165
rect 67552 13119 67598 13165
rect 67656 13119 67702 13165
rect 67760 13119 67806 13165
rect 67864 13119 67910 13165
rect 67968 13119 68014 13165
rect 68072 13119 68118 13165
rect 68176 13119 68222 13165
rect 68280 13119 68326 13165
rect 68384 13119 68430 13165
rect 68488 13119 68534 13165
rect 68592 13119 68638 13165
rect 68696 13119 68742 13165
rect 68800 13119 68846 13165
rect 68904 13119 68950 13165
rect 69008 13119 69054 13165
rect 69112 13119 69158 13165
rect 69216 13119 69262 13165
rect 69320 13119 69366 13165
rect 69424 13119 69470 13165
rect 69528 13119 69574 13165
rect 69632 13119 69678 13165
rect 69736 13119 69782 13165
rect 69840 13119 69886 13165
rect 69944 13119 69990 13165
rect 70048 13119 70094 13165
rect 70152 13119 70198 13165
rect 70256 13119 70302 13165
rect 70360 13119 70406 13165
rect 70464 13119 70510 13165
rect 70568 13119 70614 13165
rect 70672 13119 70718 13165
rect 70776 13119 70822 13165
rect 70880 13119 70926 13165
<< metal1 >>
rect 13108 70975 69957 71000
rect 13108 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69957 70975
rect 13108 70871 69957 70929
rect 13108 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69957 70871
rect 13108 70814 69957 70825
rect 13108 70767 13280 70814
rect 13108 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13280 70767
rect 13108 70663 13280 70721
rect 13108 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13280 70663
rect 13108 70559 13280 70617
rect 13108 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13280 70559
rect 13108 70455 13280 70513
rect 13108 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13280 70455
rect 13108 70351 13280 70409
rect 13108 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13280 70351
rect 13108 70247 13280 70305
rect 13108 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13280 70247
rect 13108 70143 13280 70201
rect 13108 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13280 70143
rect 13108 70039 13280 70097
rect 13108 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13280 70039
rect 13108 69935 13280 69993
rect 13108 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13280 69935
rect 13108 69831 13280 69889
rect 13108 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13280 69831
rect 69785 70720 69957 70814
rect 69785 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69957 70720
rect 69785 70616 69957 70674
rect 69785 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69957 70616
rect 69785 70512 69957 70570
rect 69785 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69957 70512
rect 69785 70408 69957 70466
rect 69785 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69957 70408
rect 69785 70304 69957 70362
rect 69785 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69957 70304
rect 69785 70200 69957 70258
rect 69785 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69957 70200
rect 69785 70096 69957 70154
rect 69785 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69957 70096
rect 69785 69957 69957 70050
rect 69785 69946 71000 69957
rect 69785 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69785 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69785 69842 71000 69862
rect 69785 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69785 69785 70824 69796
rect 13108 69727 13280 69785
rect 13108 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13280 69727
rect 13108 69623 13280 69681
rect 13108 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13280 69623
rect 13108 69519 13280 69577
rect 13108 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13280 69519
rect 13108 69415 13280 69473
rect 13108 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13280 69415
rect 13108 69311 13280 69369
rect 13108 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13280 69311
rect 13108 69207 13280 69265
rect 13108 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13280 69207
rect 13108 69103 13280 69161
rect 13108 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13280 69103
rect 13108 68999 13280 69057
rect 13108 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13280 68999
rect 13108 68895 13280 68953
rect 13108 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13280 68895
rect 13108 68791 13280 68849
rect 13108 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13280 68791
rect 13108 68687 13280 68745
rect 13108 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13280 68687
rect 13108 68583 13280 68641
rect 13108 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13280 68583
rect 13108 68479 13280 68537
rect 13108 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13280 68479
rect 13108 68375 13280 68433
rect 13108 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13280 68375
rect 13108 68271 13280 68329
rect 13108 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13280 68271
rect 13108 68167 13280 68225
rect 13108 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13280 68167
rect 13108 68063 13280 68121
rect 13108 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13280 68063
rect 13108 67959 13280 68017
rect 13108 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13280 67959
rect 13108 67855 13280 67913
rect 13108 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13280 67855
rect 13108 67751 13280 67809
rect 13108 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13280 67751
rect 13108 67647 13280 67705
rect 13108 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13280 67647
rect 13108 67543 13280 67601
rect 13108 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13280 67543
rect 13108 67439 13280 67497
rect 13108 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13280 67439
rect 13108 67335 13280 67393
rect 13108 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13280 67335
rect 13108 67231 13280 67289
rect 13108 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13280 67231
rect 13108 67127 13280 67185
rect 13108 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13280 67127
rect 13108 67023 13280 67081
rect 13108 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13280 67023
rect 13108 66919 13280 66977
rect 13108 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13280 66919
rect 13108 66815 13280 66873
rect 13108 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13280 66815
rect 13108 66711 13280 66769
rect 13108 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13280 66711
rect 13108 66607 13280 66665
rect 13108 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13280 66607
rect 13108 66503 13280 66561
rect 13108 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13280 66503
rect 13108 66399 13280 66457
rect 13108 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13280 66399
rect 13108 66295 13280 66353
rect 13108 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13280 66295
rect 13108 66191 13280 66249
rect 13108 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13280 66191
rect 13108 66087 13280 66145
rect 13108 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13280 66087
rect 13108 65983 13280 66041
rect 13108 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13280 65983
rect 13108 65879 13280 65937
rect 13108 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13280 65879
rect 13108 65775 13280 65833
rect 13108 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13280 65775
rect 13108 65671 13280 65729
rect 13108 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13280 65671
rect 13108 65567 13280 65625
rect 13108 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13280 65567
rect 13108 65463 13280 65521
rect 13108 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13280 65463
rect 13108 65359 13280 65417
rect 13108 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13280 65359
rect 13108 65255 13280 65313
rect 13108 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13280 65255
rect 13108 65151 13280 65209
rect 13108 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13280 65151
rect 13108 65047 13280 65105
rect 13108 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13280 65047
rect 13108 64943 13280 65001
rect 13108 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13280 64943
rect 13108 64839 13280 64897
rect 13108 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13280 64839
rect 13108 64735 13280 64793
rect 13108 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13280 64735
rect 13108 64631 13280 64689
rect 13108 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13280 64631
rect 13108 64527 13280 64585
rect 13108 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13280 64527
rect 13108 64423 13280 64481
rect 13108 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13280 64423
rect 13108 64319 13280 64377
rect 13108 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13280 64319
rect 13108 64215 13280 64273
rect 13108 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13280 64215
rect 13108 64111 13280 64169
rect 13108 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13280 64111
rect 13108 64007 13280 64065
rect 13108 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13280 64007
rect 13108 63903 13280 63961
rect 13108 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13280 63903
rect 13108 63799 13280 63857
rect 13108 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13280 63799
rect 13108 63695 13280 63753
rect 13108 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13280 63695
rect 13108 63591 13280 63649
rect 13108 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13280 63591
rect 13108 63487 13280 63545
rect 13108 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13280 63487
rect 13108 63383 13280 63441
rect 13108 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13280 63383
rect 13108 63279 13280 63337
rect 13108 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13280 63279
rect 13108 63175 13280 63233
rect 13108 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13280 63175
rect 13108 63071 13280 63129
rect 13108 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13280 63071
rect 13108 62967 13280 63025
rect 13108 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13280 62967
rect 13108 62863 13280 62921
rect 13108 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13280 62863
rect 13108 62759 13280 62817
rect 13108 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13280 62759
rect 13108 62655 13280 62713
rect 13108 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13280 62655
rect 13108 62551 13280 62609
rect 13108 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13280 62551
rect 13108 62447 13280 62505
rect 13108 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13280 62447
rect 13108 62343 13280 62401
rect 13108 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13280 62343
rect 13108 62239 13280 62297
rect 13108 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13280 62239
rect 13108 62135 13280 62193
rect 13108 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13280 62135
rect 13108 62031 13280 62089
rect 13108 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13280 62031
rect 13108 61927 13280 61985
rect 13108 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13280 61927
rect 13108 61823 13280 61881
rect 13108 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13280 61823
rect 13108 61719 13280 61777
rect 13108 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13280 61719
rect 13108 61615 13280 61673
rect 13108 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13280 61615
rect 13108 61511 13280 61569
rect 13108 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13280 61511
rect 13108 61407 13280 61465
rect 13108 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13280 61407
rect 13108 61303 13280 61361
rect 13108 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13280 61303
rect 13108 61199 13280 61257
rect 13108 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13280 61199
rect 13108 61095 13280 61153
rect 13108 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13280 61095
rect 13108 60991 13280 61049
rect 13108 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13280 60991
rect 13108 60887 13280 60945
rect 13108 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13280 60887
rect 13108 60783 13280 60841
rect 13108 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13280 60783
rect 13108 60679 13280 60737
rect 13108 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13280 60679
rect 13108 60575 13280 60633
rect 13108 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13280 60575
rect 13108 60471 13280 60529
rect 13108 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13280 60471
rect 13108 60367 13280 60425
rect 13108 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13280 60367
rect 13108 60263 13280 60321
rect 13108 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13280 60263
rect 13108 60159 13280 60217
rect 13108 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13280 60159
rect 13108 60055 13280 60113
rect 13108 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13280 60055
rect 13108 59951 13280 60009
rect 13108 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13280 59951
rect 13108 59847 13280 59905
rect 13108 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13280 59847
rect 13108 59743 13280 59801
rect 13108 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13280 59743
rect 13108 59639 13280 59697
rect 13108 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13280 59639
rect 13108 59535 13280 59593
rect 13108 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13280 59535
rect 13108 59431 13280 59489
rect 13108 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13280 59431
rect 13108 59327 13280 59385
rect 13108 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13280 59327
rect 13108 59223 13280 59281
rect 13108 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13280 59223
rect 13108 59119 13280 59177
rect 13108 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13280 59119
rect 13108 59015 13280 59073
rect 13108 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13280 59015
rect 13108 58911 13280 58969
rect 13108 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13280 58911
rect 13108 58807 13280 58865
rect 13108 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13280 58807
rect 13108 58703 13280 58761
rect 13108 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13280 58703
rect 13108 58599 13280 58657
rect 13108 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13280 58599
rect 13108 58495 13280 58553
rect 13108 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13280 58495
rect 13108 58391 13280 58449
rect 13108 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13280 58391
rect 13108 58287 13280 58345
rect 13108 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13280 58287
rect 13108 58183 13280 58241
rect 13108 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13280 58183
rect 13108 58079 13280 58137
rect 13108 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13280 58079
rect 13108 57975 13280 58033
rect 13108 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13280 57975
rect 13108 57871 13280 57929
rect 13108 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13280 57871
rect 13108 57767 13280 57825
rect 13108 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13280 57767
rect 13108 57663 13280 57721
rect 13108 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13280 57663
rect 13108 57559 13280 57617
rect 13108 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13280 57559
rect 13108 57455 13280 57513
rect 13108 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13280 57455
rect 13108 57351 13280 57409
rect 13108 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13280 57351
rect 13108 57247 13280 57305
rect 13108 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13280 57247
rect 13108 57143 13280 57201
rect 13108 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13280 57143
rect 13108 57039 13280 57097
rect 13108 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13280 57039
rect 13108 56935 13280 56993
rect 13108 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13280 56935
rect 13108 56831 13280 56889
rect 13108 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13280 56831
rect 13108 56727 13280 56785
rect 13108 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13280 56727
rect 13108 56623 13280 56681
rect 13108 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13280 56623
rect 13108 56519 13280 56577
rect 13108 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13280 56519
rect 13108 56415 13280 56473
rect 13108 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13280 56415
rect 13108 56311 13280 56369
rect 13108 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13280 56311
rect 13108 56207 13280 56265
rect 13108 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13280 56207
rect 13108 56103 13280 56161
rect 13108 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13280 56103
rect 13108 55999 13280 56057
rect 13108 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13280 55999
rect 13108 55895 13280 55953
rect 13108 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13280 55895
rect 13108 55791 13280 55849
rect 13108 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13280 55791
rect 13108 55687 13280 55745
rect 13108 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13280 55687
rect 13108 55583 13280 55641
rect 13108 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13280 55583
rect 13108 55479 13280 55537
rect 13108 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13280 55479
rect 13108 55375 13280 55433
rect 13108 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13280 55375
rect 13108 55271 13280 55329
rect 13108 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13280 55271
rect 13108 55167 13280 55225
rect 13108 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13280 55167
rect 13108 55063 13280 55121
rect 13108 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13280 55063
rect 13108 54959 13280 55017
rect 13108 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13280 54959
rect 13108 54855 13280 54913
rect 13108 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13280 54855
rect 13108 54751 13280 54809
rect 13108 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13280 54751
rect 13108 54647 13280 54705
rect 13108 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13280 54647
rect 13108 54543 13280 54601
rect 13108 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13280 54543
rect 13108 54439 13280 54497
rect 13108 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13280 54439
rect 13108 54335 13280 54393
rect 13108 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13280 54335
rect 13108 54231 13280 54289
rect 13108 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13280 54231
rect 13108 54127 13280 54185
rect 13108 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13280 54127
rect 13108 54023 13280 54081
rect 13108 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13280 54023
rect 13108 53919 13280 53977
rect 13108 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13280 53919
rect 13108 53815 13280 53873
rect 13108 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13280 53815
rect 13108 53711 13280 53769
rect 13108 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13280 53711
rect 13108 53607 13280 53665
rect 13108 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13280 53607
rect 13108 53503 13280 53561
rect 13108 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13280 53503
rect 13108 53399 13280 53457
rect 13108 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13280 53399
rect 13108 53295 13280 53353
rect 13108 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13280 53295
rect 13108 53191 13280 53249
rect 13108 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13280 53191
rect 13108 53087 13280 53145
rect 13108 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13280 53087
rect 13108 52983 13280 53041
rect 13108 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13280 52983
rect 13108 52879 13280 52937
rect 13108 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13280 52879
rect 13108 52775 13280 52833
rect 13108 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13280 52775
rect 13108 52671 13280 52729
rect 13108 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13280 52671
rect 13108 52567 13280 52625
rect 13108 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13280 52567
rect 13108 52463 13280 52521
rect 13108 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13280 52463
rect 13108 52359 13280 52417
rect 13108 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13280 52359
rect 13108 52255 13280 52313
rect 13108 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13280 52255
rect 13108 52151 13280 52209
rect 13108 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13280 52151
rect 13108 52047 13280 52105
rect 13108 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13280 52047
rect 13108 51943 13280 52001
rect 13108 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13280 51943
rect 13108 51839 13280 51897
rect 13108 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13280 51839
rect 13108 51735 13280 51793
rect 13108 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13280 51735
rect 13108 51631 13280 51689
rect 13108 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13280 51631
rect 13108 51527 13280 51585
rect 13108 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13280 51527
rect 13108 51423 13280 51481
rect 13108 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13280 51423
rect 13108 51319 13280 51377
rect 13108 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13280 51319
rect 13108 51215 13280 51273
rect 13108 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13280 51215
rect 13108 51111 13280 51169
rect 13108 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13280 51111
rect 13108 51007 13280 51065
rect 13108 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13280 51007
rect 13108 50903 13280 50961
rect 13108 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13280 50903
rect 13108 50799 13280 50857
rect 13108 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13280 50799
rect 13108 50695 13280 50753
rect 13108 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13280 50695
rect 13108 50591 13280 50649
rect 13108 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13280 50591
rect 13108 50487 13280 50545
rect 13108 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13280 50487
rect 13108 50383 13280 50441
rect 13108 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13280 50383
rect 13108 50279 13280 50337
rect 13108 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13280 50279
rect 13108 50175 13280 50233
rect 13108 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13280 50175
rect 13108 50071 13280 50129
rect 13108 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13280 50071
rect 13108 49967 13280 50025
rect 13108 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13280 49967
rect 13108 49863 13280 49921
rect 13108 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13280 49863
rect 13108 49759 13280 49817
rect 13108 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13280 49759
rect 13108 49655 13280 49713
rect 13108 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13280 49655
rect 13108 49551 13280 49609
rect 13108 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13280 49551
rect 13108 49447 13280 49505
rect 13108 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13280 49447
rect 13108 49343 13280 49401
rect 13108 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13280 49343
rect 13108 49239 13280 49297
rect 13108 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13280 49239
rect 13108 49135 13280 49193
rect 13108 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13280 49135
rect 13108 49031 13280 49089
rect 13108 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13280 49031
rect 13108 48927 13280 48985
rect 13108 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13280 48927
rect 13108 48823 13280 48881
rect 13108 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13280 48823
rect 13108 48719 13280 48777
rect 13108 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13280 48719
rect 13108 48615 13280 48673
rect 13108 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13280 48615
rect 13108 48511 13280 48569
rect 13108 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13280 48511
rect 13108 48407 13280 48465
rect 13108 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13280 48407
rect 13108 48303 13280 48361
rect 13108 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13280 48303
rect 13108 48199 13280 48257
rect 13108 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13280 48199
rect 13108 48095 13280 48153
rect 13108 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13280 48095
rect 13108 47991 13280 48049
rect 13108 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13280 47991
rect 13108 47887 13280 47945
rect 13108 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13280 47887
rect 13108 47783 13280 47841
rect 13108 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13280 47783
rect 13108 47679 13280 47737
rect 13108 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13280 47679
rect 13108 47575 13280 47633
rect 13108 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13280 47575
rect 13108 47471 13280 47529
rect 13108 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13280 47471
rect 13108 47367 13280 47425
rect 13108 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13280 47367
rect 13108 47263 13280 47321
rect 13108 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13280 47263
rect 13108 47159 13280 47217
rect 13108 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13280 47159
rect 13108 47055 13280 47113
rect 13108 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13280 47055
rect 13108 46951 13280 47009
rect 13108 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13280 46951
rect 13108 46847 13280 46905
rect 13108 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13280 46847
rect 13108 46743 13280 46801
rect 13108 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13280 46743
rect 13108 46639 13280 46697
rect 13108 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13280 46639
rect 13108 46535 13280 46593
rect 13108 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13280 46535
rect 13108 46431 13280 46489
rect 13108 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13280 46431
rect 13108 46327 13280 46385
rect 13108 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13280 46327
rect 13108 46223 13280 46281
rect 13108 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13280 46223
rect 13108 46119 13280 46177
rect 13108 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13280 46119
rect 13108 46015 13280 46073
rect 13108 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13280 46015
rect 13108 45911 13280 45969
rect 13108 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13280 45911
rect 13108 45807 13280 45865
rect 13108 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13280 45807
rect 13108 45703 13280 45761
rect 13108 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13280 45703
rect 13108 45599 13280 45657
rect 13108 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13280 45599
rect 13108 45495 13280 45553
rect 13108 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13280 45495
rect 13108 45391 13280 45449
rect 13108 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13280 45391
rect 13108 45287 13280 45345
rect 13108 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13280 45287
rect 13108 45183 13280 45241
rect 13108 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13280 45183
rect 13108 45079 13280 45137
rect 13108 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13280 45079
rect 13108 44902 13280 45033
rect 70813 69758 70824 69785
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70813 69700 71000 69758
rect 70813 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70813 69596 71000 69654
rect 70813 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70813 69492 71000 69550
rect 70813 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70813 69388 71000 69446
rect 70813 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70813 69284 71000 69342
rect 70813 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70813 69180 71000 69238
rect 70813 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70813 69076 71000 69134
rect 70813 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70813 68972 71000 69030
rect 70813 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70813 68868 71000 68926
rect 70813 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70813 68764 71000 68822
rect 70813 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70813 68660 71000 68718
rect 70813 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70813 68556 71000 68614
rect 70813 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70813 68452 71000 68510
rect 70813 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70813 68348 71000 68406
rect 70813 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70813 68244 71000 68302
rect 70813 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70813 68140 71000 68198
rect 70813 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70813 68036 71000 68094
rect 70813 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70813 67932 71000 67990
rect 70813 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70813 67828 71000 67886
rect 70813 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70813 67724 71000 67782
rect 70813 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70813 67620 71000 67678
rect 70813 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70813 67516 71000 67574
rect 70813 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70813 67412 71000 67470
rect 70813 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70813 67308 71000 67366
rect 70813 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70813 67204 71000 67262
rect 70813 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70813 67100 71000 67158
rect 70813 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70813 66996 71000 67054
rect 70813 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70813 66892 71000 66950
rect 70813 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70813 66788 71000 66846
rect 70813 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70813 66684 71000 66742
rect 70813 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70813 66580 71000 66638
rect 70813 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70813 66476 71000 66534
rect 70813 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70813 66372 71000 66430
rect 70813 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70813 66268 71000 66326
rect 70813 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70813 66164 71000 66222
rect 70813 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70813 66060 71000 66118
rect 70813 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70813 65956 71000 66014
rect 70813 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70813 65852 71000 65910
rect 70813 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70813 65748 71000 65806
rect 70813 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70813 65644 71000 65702
rect 70813 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70813 65540 71000 65598
rect 70813 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70813 65436 71000 65494
rect 70813 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70813 65332 71000 65390
rect 70813 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70813 65228 71000 65286
rect 70813 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70813 65124 71000 65182
rect 70813 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70813 65020 71000 65078
rect 70813 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70813 64916 71000 64974
rect 70813 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70813 64812 71000 64870
rect 70813 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70813 64708 71000 64766
rect 70813 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70813 64604 71000 64662
rect 70813 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70813 64500 71000 64558
rect 70813 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70813 64396 71000 64454
rect 70813 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70813 64292 71000 64350
rect 70813 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70813 64188 71000 64246
rect 70813 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70813 64084 71000 64142
rect 70813 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70813 63980 71000 64038
rect 70813 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70813 63876 71000 63934
rect 70813 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70813 63772 71000 63830
rect 70813 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70813 63668 71000 63726
rect 70813 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70813 63564 71000 63622
rect 70813 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70813 63460 71000 63518
rect 70813 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70813 63356 71000 63414
rect 70813 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70813 63252 71000 63310
rect 70813 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70813 63148 71000 63206
rect 70813 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70813 63044 71000 63102
rect 70813 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70813 62940 71000 62998
rect 70813 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70813 62836 71000 62894
rect 70813 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70813 62732 71000 62790
rect 70813 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70813 62628 71000 62686
rect 70813 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70813 62524 71000 62582
rect 70813 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70813 62420 71000 62478
rect 70813 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70813 62316 71000 62374
rect 70813 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70813 62212 71000 62270
rect 70813 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70813 62108 71000 62166
rect 70813 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70813 62004 71000 62062
rect 70813 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70813 61900 71000 61958
rect 70813 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70813 61796 71000 61854
rect 70813 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70813 61692 71000 61750
rect 70813 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70813 61588 71000 61646
rect 70813 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70813 61484 71000 61542
rect 70813 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70813 61380 71000 61438
rect 70813 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70813 61276 71000 61334
rect 70813 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70813 61172 71000 61230
rect 70813 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70813 61068 71000 61126
rect 70813 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70813 60964 71000 61022
rect 70813 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70813 60860 71000 60918
rect 70813 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70813 60756 71000 60814
rect 70813 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70813 60652 71000 60710
rect 70813 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70813 60548 71000 60606
rect 70813 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70813 60444 71000 60502
rect 70813 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70813 60340 71000 60398
rect 70813 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70813 60236 71000 60294
rect 70813 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70813 60132 71000 60190
rect 70813 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70813 60028 71000 60086
rect 70813 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70813 59924 71000 59982
rect 70813 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70813 59820 71000 59878
rect 70813 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70813 59716 71000 59774
rect 70813 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70813 59612 71000 59670
rect 70813 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70813 59508 71000 59566
rect 70813 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70813 59404 71000 59462
rect 70813 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70813 59300 71000 59358
rect 70813 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70813 59196 71000 59254
rect 70813 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70813 59092 71000 59150
rect 70813 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70813 58988 71000 59046
rect 70813 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70813 58884 71000 58942
rect 70813 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70813 58780 71000 58838
rect 70813 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70813 58676 71000 58734
rect 70813 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70813 58572 71000 58630
rect 70813 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70813 58468 71000 58526
rect 70813 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70813 58364 71000 58422
rect 70813 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70813 58260 71000 58318
rect 70813 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70813 58156 71000 58214
rect 70813 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70813 58052 71000 58110
rect 70813 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70813 57948 71000 58006
rect 70813 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70813 57844 71000 57902
rect 70813 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70813 57740 71000 57798
rect 70813 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70813 57636 71000 57694
rect 70813 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70813 57532 71000 57590
rect 70813 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70813 57428 71000 57486
rect 70813 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70813 57324 71000 57382
rect 70813 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70813 57220 71000 57278
rect 70813 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70813 57116 71000 57174
rect 70813 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70813 57012 71000 57070
rect 70813 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70813 56908 71000 56966
rect 70813 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70813 56804 71000 56862
rect 70813 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70813 56700 71000 56758
rect 70813 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70813 56596 71000 56654
rect 70813 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70813 56492 71000 56550
rect 70813 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70813 56388 71000 56446
rect 70813 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70813 56284 71000 56342
rect 70813 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70813 56180 71000 56238
rect 70813 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70813 56076 71000 56134
rect 70813 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70813 55972 71000 56030
rect 70813 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70813 55868 71000 55926
rect 70813 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70813 55764 71000 55822
rect 70813 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70813 55660 71000 55718
rect 70813 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70813 55556 71000 55614
rect 70813 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70813 55452 71000 55510
rect 70813 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70813 55348 71000 55406
rect 70813 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70813 55244 71000 55302
rect 70813 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70813 55140 71000 55198
rect 70813 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70813 55036 71000 55094
rect 70813 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70813 54932 71000 54990
rect 70813 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70813 54828 71000 54886
rect 70813 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70813 54724 71000 54782
rect 70813 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70813 54620 71000 54678
rect 70813 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70813 54516 71000 54574
rect 70813 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70813 54412 71000 54470
rect 70813 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70813 54308 71000 54366
rect 70813 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70813 54204 71000 54262
rect 70813 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70813 54100 71000 54158
rect 70813 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70813 53996 71000 54054
rect 70813 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70813 53892 71000 53950
rect 70813 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70813 53788 71000 53846
rect 70813 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70813 53684 71000 53742
rect 70813 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70813 53580 71000 53638
rect 70813 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70813 53476 71000 53534
rect 70813 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70813 53372 71000 53430
rect 70813 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70813 53268 71000 53326
rect 70813 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70813 53164 71000 53222
rect 70813 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70813 53060 71000 53118
rect 70813 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70813 52956 71000 53014
rect 70813 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70813 52852 71000 52910
rect 70813 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70813 52748 71000 52806
rect 70813 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70813 52644 71000 52702
rect 70813 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70813 52540 71000 52598
rect 70813 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70813 52436 71000 52494
rect 70813 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70813 52332 71000 52390
rect 70813 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70813 52228 71000 52286
rect 70813 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70813 52124 71000 52182
rect 70813 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70813 52020 71000 52078
rect 70813 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70813 51916 71000 51974
rect 70813 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70813 51812 71000 51870
rect 70813 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70813 51708 71000 51766
rect 70813 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70813 51604 71000 51662
rect 70813 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70813 51500 71000 51558
rect 70813 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70813 51396 71000 51454
rect 70813 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70813 51292 71000 51350
rect 70813 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70813 51188 71000 51246
rect 70813 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70813 51084 71000 51142
rect 70813 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70813 50980 71000 51038
rect 70813 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70813 50876 71000 50934
rect 70813 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70813 50772 71000 50830
rect 70813 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70813 50668 71000 50726
rect 70813 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70813 50564 71000 50622
rect 70813 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70813 50460 71000 50518
rect 70813 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70813 50356 71000 50414
rect 70813 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70813 50252 71000 50310
rect 70813 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70813 50148 71000 50206
rect 70813 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70813 50044 71000 50102
rect 70813 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70813 49940 71000 49998
rect 70813 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70813 49836 71000 49894
rect 70813 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70813 49732 71000 49790
rect 70813 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70813 49628 71000 49686
rect 70813 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70813 49524 71000 49582
rect 70813 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70813 49420 71000 49478
rect 70813 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70813 49316 71000 49374
rect 70813 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70813 49212 71000 49270
rect 70813 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70813 49108 71000 49166
rect 70813 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70813 49004 71000 49062
rect 70813 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70813 48900 71000 48958
rect 70813 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70813 48796 71000 48854
rect 70813 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70813 48692 71000 48750
rect 70813 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70813 48588 71000 48646
rect 70813 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70813 48484 71000 48542
rect 70813 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70813 48380 71000 48438
rect 70813 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70813 48276 71000 48334
rect 70813 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70813 48172 71000 48230
rect 70813 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70813 48068 71000 48126
rect 70813 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70813 47964 71000 48022
rect 70813 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70813 47860 71000 47918
rect 70813 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70813 47756 71000 47814
rect 70813 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70813 47652 71000 47710
rect 70813 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70813 47548 71000 47606
rect 70813 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70813 47444 71000 47502
rect 70813 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70813 47340 71000 47398
rect 70813 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70813 47236 71000 47294
rect 70813 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70813 47132 71000 47190
rect 70813 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70813 47028 71000 47086
rect 70813 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70813 46924 71000 46982
rect 70813 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70813 46820 71000 46878
rect 70813 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70813 46716 71000 46774
rect 70813 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70813 46612 71000 46670
rect 70813 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70813 46508 71000 46566
rect 70813 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70813 46404 71000 46462
rect 70813 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70813 46300 71000 46358
rect 70813 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70813 46196 71000 46254
rect 70813 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70813 46092 71000 46150
rect 70813 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70813 45988 71000 46046
rect 70813 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70813 45884 71000 45942
rect 70813 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70813 45780 71000 45838
rect 70813 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70813 45676 71000 45734
rect 70813 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70813 45572 71000 45630
rect 70813 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70813 45468 71000 45526
rect 70813 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70813 45364 71000 45422
rect 70813 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70813 45260 71000 45318
rect 70813 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70813 45156 71000 45214
rect 70813 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70813 45052 71000 45110
rect 70813 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70813 44948 71000 45006
tri 13280 44902 13298 44920 sw
rect 70813 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13108 44848 13298 44902
tri 13108 44844 13112 44848 ne
rect 13112 44844 13298 44848
tri 13298 44844 13356 44902 sw
rect 70813 44844 71000 44902
tri 13112 44828 13128 44844 ne
rect 13128 44828 13356 44844
tri 13356 44828 13372 44844 sw
tri 13128 44824 13132 44828 ne
rect 13132 44824 13372 44828
tri 13132 44778 13178 44824 ne
rect 13178 44778 13254 44824
rect 13300 44798 13372 44824
tri 13372 44798 13402 44828 sw
rect 70813 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 13300 44778 13402 44798
tri 13178 44740 13216 44778 ne
rect 13216 44740 13402 44778
tri 13402 44740 13460 44798 sw
rect 70813 44740 71000 44798
tri 13216 44694 13262 44740 ne
rect 13262 44694 13460 44740
tri 13460 44694 13506 44740 sw
rect 70813 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
tri 13262 44692 13264 44694 ne
rect 13264 44692 13506 44694
tri 13506 44692 13508 44694 sw
tri 13264 44646 13310 44692 ne
rect 13310 44646 13386 44692
rect 13432 44646 13508 44692
tri 13508 44646 13554 44692 sw
tri 13310 44636 13320 44646 ne
rect 13320 44636 13554 44646
tri 13554 44636 13564 44646 sw
rect 70813 44636 71000 44694
tri 13320 44590 13366 44636 ne
rect 13366 44590 13564 44636
tri 13564 44590 13610 44636 sw
rect 70813 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13366 44584 13372 44590 ne
rect 13372 44584 13610 44590
tri 13610 44584 13616 44590 sw
tri 13372 44560 13396 44584 ne
rect 13396 44560 13616 44584
tri 13396 44514 13442 44560 ne
rect 13442 44514 13518 44560
rect 13564 44532 13616 44560
tri 13616 44532 13668 44584 sw
rect 70813 44532 71000 44590
rect 13564 44514 13668 44532
tri 13442 44486 13470 44514 ne
rect 13470 44486 13668 44514
tri 13668 44486 13714 44532 sw
rect 70813 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
tri 13470 44428 13528 44486 ne
rect 13528 44428 13714 44486
tri 13714 44428 13772 44486 sw
rect 70813 44428 71000 44486
tri 13528 44382 13574 44428 ne
rect 13574 44382 13650 44428
rect 13696 44382 13772 44428
tri 13772 44382 13818 44428 sw
rect 70813 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
tri 13574 44340 13616 44382 ne
rect 13616 44340 13818 44382
tri 13818 44340 13860 44382 sw
tri 13616 44324 13632 44340 ne
rect 13632 44324 13860 44340
tri 13860 44324 13876 44340 sw
rect 70813 44324 71000 44382
tri 13632 44296 13660 44324 ne
rect 13660 44296 13876 44324
tri 13660 44250 13706 44296 ne
rect 13706 44250 13782 44296
rect 13828 44278 13876 44296
tri 13876 44278 13922 44324 sw
rect 70813 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 13828 44250 13922 44278
tri 13706 44220 13736 44250 ne
rect 13736 44220 13922 44250
tri 13922 44220 13980 44278 sw
rect 70813 44220 71000 44278
tri 13736 44174 13782 44220 ne
rect 13782 44174 13980 44220
tri 13980 44174 14026 44220 sw
rect 70813 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
tri 13782 44164 13792 44174 ne
rect 13792 44164 14026 44174
tri 14026 44164 14036 44174 sw
tri 13792 44118 13838 44164 ne
rect 13838 44118 13914 44164
rect 13960 44118 14036 44164
tri 14036 44118 14082 44164 sw
tri 13838 44116 13840 44118 ne
rect 13840 44116 14082 44118
tri 14082 44116 14084 44118 sw
rect 70813 44116 71000 44174
tri 13840 44096 13860 44116 ne
rect 13860 44096 14084 44116
tri 14084 44096 14104 44116 sw
tri 13860 44070 13886 44096 ne
rect 13886 44070 14104 44096
tri 14104 44070 14130 44096 sw
rect 70813 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
tri 13886 44032 13924 44070 ne
rect 13924 44032 14130 44070
tri 13924 43986 13970 44032 ne
rect 13970 43986 14046 44032
rect 14092 44012 14130 44032
tri 14130 44012 14188 44070 sw
rect 70813 44012 71000 44070
rect 14092 43986 14188 44012
tri 13970 43966 13990 43986 ne
rect 13990 43966 14188 43986
tri 14188 43966 14234 44012 sw
rect 70813 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13990 43908 14048 43966 ne
rect 14048 43908 14234 43966
tri 14234 43908 14292 43966 sw
rect 70813 43908 71000 43966
tri 14048 43900 14056 43908 ne
rect 14056 43900 14292 43908
tri 14292 43900 14300 43908 sw
tri 14056 43854 14102 43900 ne
rect 14102 43854 14178 43900
rect 14224 43862 14300 43900
tri 14300 43862 14338 43900 sw
rect 70813 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 14224 43854 14338 43862
tri 14338 43854 14346 43862 sw
tri 14102 43852 14104 43854 ne
rect 14104 43852 14346 43854
tri 14346 43852 14348 43854 sw
tri 14104 43804 14152 43852 ne
rect 14152 43804 14348 43852
tri 14348 43804 14396 43852 sw
rect 70813 43804 71000 43862
tri 14152 43768 14188 43804 ne
rect 14188 43768 14396 43804
tri 14396 43768 14432 43804 sw
tri 14188 43722 14234 43768 ne
rect 14234 43722 14310 43768
rect 14356 43758 14432 43768
tri 14432 43758 14442 43768 sw
rect 70813 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43722 14442 43758
tri 14442 43722 14478 43758 sw
tri 14234 43700 14256 43722 ne
rect 14256 43700 14478 43722
tri 14478 43700 14500 43722 sw
rect 70813 43700 71000 43758
tri 14256 43654 14302 43700 ne
rect 14302 43654 14500 43700
tri 14500 43654 14546 43700 sw
rect 70813 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
tri 14302 43636 14320 43654 ne
rect 14320 43636 14546 43654
tri 14546 43636 14564 43654 sw
tri 14320 43608 14348 43636 ne
rect 14348 43608 14442 43636
tri 14348 43590 14366 43608 ne
rect 14366 43590 14442 43608
rect 14488 43608 14564 43636
tri 14564 43608 14592 43636 sw
rect 14488 43596 14592 43608
tri 14592 43596 14604 43608 sw
rect 70813 43596 71000 43654
rect 14488 43590 14604 43596
tri 14366 43550 14406 43590 ne
rect 14406 43550 14604 43590
tri 14604 43550 14650 43596 sw
rect 70813 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
tri 14406 43504 14452 43550 ne
rect 14452 43504 14650 43550
tri 14650 43504 14696 43550 sw
tri 14452 43458 14498 43504 ne
rect 14498 43458 14574 43504
rect 14620 43492 14696 43504
tri 14696 43492 14708 43504 sw
rect 70813 43492 71000 43550
rect 14620 43458 14708 43492
tri 14708 43458 14742 43492 sw
tri 14498 43446 14510 43458 ne
rect 14510 43446 14742 43458
tri 14742 43446 14754 43458 sw
rect 70813 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14510 43388 14568 43446 ne
rect 14568 43388 14754 43446
tri 14754 43388 14812 43446 sw
rect 70813 43388 71000 43446
tri 14568 43372 14584 43388 ne
rect 14584 43372 14812 43388
tri 14812 43372 14828 43388 sw
tri 14584 43364 14592 43372 ne
rect 14592 43364 14706 43372
tri 14592 43326 14630 43364 ne
rect 14630 43326 14706 43364
rect 14752 43364 14828 43372
tri 14828 43364 14836 43372 sw
rect 14752 43342 14836 43364
tri 14836 43342 14858 43364 sw
rect 70813 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 14752 43326 14858 43342
tri 14630 43284 14672 43326 ne
rect 14672 43284 14858 43326
tri 14858 43284 14916 43342 sw
rect 70813 43284 71000 43342
tri 14672 43240 14716 43284 ne
rect 14716 43240 14916 43284
tri 14916 43240 14960 43284 sw
tri 14716 43194 14762 43240 ne
rect 14762 43194 14838 43240
rect 14884 43238 14960 43240
tri 14960 43238 14962 43240 sw
rect 70813 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43194 14962 43238
tri 14962 43194 15006 43238 sw
tri 14762 43180 14776 43194 ne
rect 14776 43180 15006 43194
tri 15006 43180 15020 43194 sw
rect 70813 43180 71000 43238
tri 14776 43134 14822 43180 ne
rect 14822 43134 15020 43180
tri 15020 43134 15066 43180 sw
rect 70813 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14822 43120 14836 43134 ne
rect 14836 43120 15066 43134
tri 15066 43120 15080 43134 sw
tri 14836 43108 14848 43120 ne
rect 14848 43108 15080 43120
tri 14848 43062 14894 43108 ne
rect 14894 43062 14970 43108
rect 15016 43076 15080 43108
tri 15080 43076 15124 43120 sw
rect 70813 43076 71000 43134
rect 15016 43062 15124 43076
tri 14894 43030 14926 43062 ne
rect 14926 43030 15124 43062
tri 15124 43030 15170 43076 sw
rect 70813 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14926 42976 14980 43030 ne
rect 14980 42976 15170 43030
tri 15170 42976 15224 43030 sw
tri 14980 42930 15026 42976 ne
rect 15026 42930 15102 42976
rect 15148 42972 15224 42976
tri 15224 42972 15228 42976 sw
rect 70813 42972 71000 43030
rect 15148 42930 15228 42972
tri 15228 42930 15270 42972 sw
tri 15026 42926 15030 42930 ne
rect 15030 42926 15270 42930
tri 15270 42926 15274 42930 sw
rect 70813 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15030 42876 15080 42926 ne
rect 15080 42876 15274 42926
tri 15274 42876 15324 42926 sw
tri 15080 42868 15088 42876 ne
rect 15088 42868 15324 42876
tri 15324 42868 15332 42876 sw
rect 70813 42868 71000 42926
tri 15088 42844 15112 42868 ne
rect 15112 42844 15332 42868
tri 15112 42798 15158 42844 ne
rect 15158 42798 15234 42844
rect 15280 42822 15332 42844
tri 15332 42822 15378 42868 sw
rect 70813 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 15280 42798 15378 42822
tri 15158 42764 15192 42798 ne
rect 15192 42764 15378 42798
tri 15378 42764 15436 42822 sw
rect 70813 42764 71000 42822
tri 15192 42718 15238 42764 ne
rect 15238 42718 15436 42764
tri 15436 42718 15482 42764 sw
rect 70813 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
tri 15238 42712 15244 42718 ne
rect 15244 42712 15482 42718
tri 15482 42712 15488 42718 sw
tri 15244 42666 15290 42712 ne
rect 15290 42666 15366 42712
rect 15412 42666 15488 42712
tri 15488 42666 15534 42712 sw
tri 15290 42660 15296 42666 ne
rect 15296 42660 15534 42666
tri 15534 42660 15540 42666 sw
rect 70813 42660 71000 42718
tri 15296 42632 15324 42660 ne
rect 15324 42632 15540 42660
tri 15540 42632 15568 42660 sw
tri 15324 42614 15342 42632 ne
rect 15342 42614 15568 42632
tri 15568 42614 15586 42632 sw
rect 70813 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15342 42580 15376 42614 ne
rect 15376 42580 15586 42614
tri 15376 42534 15422 42580 ne
rect 15422 42534 15498 42580
rect 15544 42556 15586 42580
tri 15586 42556 15644 42614 sw
rect 70813 42556 71000 42614
rect 15544 42534 15644 42556
tri 15422 42510 15446 42534 ne
rect 15446 42510 15644 42534
tri 15644 42510 15690 42556 sw
rect 70813 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
tri 15446 42452 15504 42510 ne
rect 15504 42452 15690 42510
tri 15690 42452 15748 42510 sw
rect 70813 42452 71000 42510
tri 15504 42448 15508 42452 ne
rect 15508 42448 15748 42452
tri 15748 42448 15752 42452 sw
tri 15508 42402 15554 42448 ne
rect 15554 42402 15630 42448
rect 15676 42406 15752 42448
tri 15752 42406 15794 42448 sw
rect 70813 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 15676 42402 15794 42406
tri 15794 42402 15798 42406 sw
tri 15554 42388 15568 42402 ne
rect 15568 42388 15798 42402
tri 15798 42388 15812 42402 sw
tri 15568 42348 15608 42388 ne
rect 15608 42348 15812 42388
tri 15812 42348 15852 42388 sw
rect 70813 42348 71000 42406
tri 15608 42316 15640 42348 ne
rect 15640 42316 15852 42348
tri 15640 42270 15686 42316 ne
rect 15686 42270 15762 42316
rect 15808 42302 15852 42316
tri 15852 42302 15898 42348 sw
rect 70813 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42270 15898 42302
tri 15686 42244 15712 42270 ne
rect 15712 42244 15898 42270
tri 15898 42244 15956 42302 sw
rect 70813 42244 71000 42302
tri 15712 42198 15758 42244 ne
rect 15758 42198 15956 42244
tri 15956 42198 16002 42244 sw
rect 70813 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
tri 15758 42184 15772 42198 ne
rect 15772 42184 16002 42198
tri 16002 42184 16016 42198 sw
tri 15772 42144 15812 42184 ne
rect 15812 42144 15894 42184
tri 15812 42138 15818 42144 ne
rect 15818 42138 15894 42144
rect 15940 42144 16016 42184
tri 16016 42144 16056 42184 sw
rect 15940 42140 16056 42144
tri 16056 42140 16060 42144 sw
rect 70813 42140 71000 42198
rect 15940 42138 16060 42140
tri 15818 42094 15862 42138 ne
rect 15862 42094 16060 42138
tri 16060 42094 16106 42140 sw
rect 70813 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15862 42052 15904 42094 ne
rect 15904 42052 16106 42094
tri 16106 42052 16148 42094 sw
tri 15904 42006 15950 42052 ne
rect 15950 42006 16026 42052
rect 16072 42036 16148 42052
tri 16148 42036 16164 42052 sw
rect 70813 42036 71000 42094
rect 16072 42006 16164 42036
tri 16164 42006 16194 42036 sw
tri 15950 41990 15966 42006 ne
rect 15966 41990 16194 42006
tri 16194 41990 16210 42006 sw
rect 70813 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15966 41932 16024 41990 ne
rect 16024 41932 16210 41990
tri 16210 41932 16268 41990 sw
rect 70813 41932 71000 41990
tri 16024 41920 16036 41932 ne
rect 16036 41920 16268 41932
tri 16268 41920 16280 41932 sw
tri 16036 41900 16056 41920 ne
rect 16056 41900 16158 41920
tri 16056 41874 16082 41900 ne
rect 16082 41874 16158 41900
rect 16204 41900 16280 41920
tri 16280 41900 16300 41920 sw
rect 16204 41886 16300 41900
tri 16300 41886 16314 41900 sw
rect 70813 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 16204 41874 16314 41886
tri 16082 41828 16128 41874 ne
rect 16128 41828 16314 41874
tri 16314 41828 16372 41886 sw
rect 70813 41828 71000 41886
tri 16128 41788 16168 41828 ne
rect 16168 41788 16372 41828
tri 16372 41788 16412 41828 sw
tri 16168 41742 16214 41788 ne
rect 16214 41742 16290 41788
rect 16336 41782 16412 41788
tri 16412 41782 16418 41788 sw
rect 70813 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41742 16418 41782
tri 16418 41742 16458 41782 sw
tri 16214 41724 16232 41742 ne
rect 16232 41724 16458 41742
tri 16458 41724 16476 41742 sw
rect 70813 41724 71000 41782
tri 16232 41678 16278 41724 ne
rect 16278 41678 16476 41724
tri 16476 41678 16522 41724 sw
rect 70813 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
tri 16278 41656 16300 41678 ne
rect 16300 41656 16522 41678
tri 16522 41656 16544 41678 sw
tri 16300 41610 16346 41656 ne
rect 16346 41610 16422 41656
rect 16468 41620 16544 41656
tri 16544 41620 16580 41656 sw
rect 70813 41620 71000 41678
rect 16468 41610 16580 41620
tri 16346 41574 16382 41610 ne
rect 16382 41574 16580 41610
tri 16580 41574 16626 41620 sw
rect 70813 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16382 41524 16432 41574 ne
rect 16432 41524 16626 41574
tri 16626 41524 16676 41574 sw
tri 16432 41478 16478 41524 ne
rect 16478 41478 16554 41524
rect 16600 41516 16676 41524
tri 16676 41516 16684 41524 sw
rect 70813 41516 71000 41574
rect 16600 41478 16684 41516
tri 16684 41478 16722 41516 sw
tri 16478 41470 16486 41478 ne
rect 16486 41470 16722 41478
tri 16722 41470 16730 41478 sw
rect 70813 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
tri 16486 41412 16544 41470 ne
rect 16544 41412 16730 41470
tri 16730 41412 16788 41470 sw
rect 70813 41412 71000 41470
tri 16544 41392 16564 41412 ne
rect 16564 41392 16788 41412
tri 16564 41346 16610 41392 ne
rect 16610 41346 16686 41392
rect 16732 41366 16788 41392
tri 16788 41366 16834 41412 sw
rect 70813 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 16732 41346 16834 41366
tri 16610 41308 16648 41346 ne
rect 16648 41308 16834 41346
tri 16834 41308 16892 41366 sw
rect 70813 41308 71000 41366
tri 16648 41262 16694 41308 ne
rect 16694 41262 16892 41308
tri 16892 41262 16938 41308 sw
rect 70813 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
tri 16694 41260 16696 41262 ne
rect 16696 41260 16938 41262
tri 16938 41260 16940 41262 sw
tri 16696 41214 16742 41260 ne
rect 16742 41214 16818 41260
rect 16864 41214 16940 41260
tri 16940 41214 16986 41260 sw
tri 16742 41204 16752 41214 ne
rect 16752 41204 16986 41214
tri 16986 41204 16996 41214 sw
rect 70813 41204 71000 41262
tri 16752 41168 16788 41204 ne
rect 16788 41168 16996 41204
tri 16996 41168 17032 41204 sw
tri 16788 41158 16798 41168 ne
rect 16798 41158 17032 41168
tri 17032 41158 17042 41168 sw
rect 70813 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
tri 16798 41128 16828 41158 ne
rect 16828 41128 17042 41158
tri 16828 41082 16874 41128 ne
rect 16874 41082 16950 41128
rect 16996 41100 17042 41128
tri 17042 41100 17100 41158 sw
rect 70813 41100 71000 41158
rect 16996 41082 17100 41100
tri 16874 41054 16902 41082 ne
rect 16902 41054 17100 41082
tri 17100 41054 17146 41100 sw
rect 70813 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
tri 16902 40996 16960 41054 ne
rect 16960 40996 17146 41054
tri 17146 40996 17204 41054 sw
rect 70813 40996 71000 41054
tri 16960 40950 17006 40996 ne
rect 17006 40950 17082 40996
rect 17128 40950 17204 40996
tri 17204 40950 17250 40996 sw
rect 70813 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
tri 17006 40924 17032 40950 ne
rect 17032 40924 17250 40950
tri 17250 40924 17276 40950 sw
tri 17032 40892 17064 40924 ne
rect 17064 40892 17276 40924
tri 17276 40892 17308 40924 sw
rect 70813 40892 71000 40950
tri 17064 40864 17092 40892 ne
rect 17092 40864 17308 40892
tri 17092 40818 17138 40864 ne
rect 17138 40818 17214 40864
rect 17260 40846 17308 40864
tri 17308 40846 17354 40892 sw
rect 70813 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40818 17354 40846
tri 17138 40788 17168 40818 ne
rect 17168 40788 17354 40818
tri 17354 40788 17412 40846 sw
rect 70813 40788 71000 40846
tri 17168 40742 17214 40788 ne
rect 17214 40742 17412 40788
tri 17412 40742 17458 40788 sw
rect 70813 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
tri 17214 40732 17224 40742 ne
rect 17224 40732 17458 40742
tri 17458 40732 17468 40742 sw
tri 17224 40686 17270 40732 ne
rect 17270 40686 17346 40732
rect 17392 40686 17468 40732
tri 17468 40686 17514 40732 sw
tri 17270 40684 17272 40686 ne
rect 17272 40684 17514 40686
tri 17514 40684 17516 40686 sw
rect 70813 40684 71000 40742
tri 17272 40680 17276 40684 ne
rect 17276 40680 17516 40684
tri 17516 40680 17520 40684 sw
tri 17276 40638 17318 40680 ne
rect 17318 40638 17520 40680
tri 17520 40638 17562 40680 sw
rect 70813 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17318 40600 17356 40638 ne
rect 17356 40600 17562 40638
tri 17562 40600 17600 40638 sw
tri 17356 40554 17402 40600 ne
rect 17402 40554 17478 40600
rect 17524 40580 17600 40600
tri 17600 40580 17620 40600 sw
rect 70813 40580 71000 40638
rect 17524 40554 17620 40580
tri 17620 40554 17646 40580 sw
tri 17402 40534 17422 40554 ne
rect 17422 40534 17646 40554
tri 17646 40534 17666 40554 sw
rect 70813 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17422 40476 17480 40534 ne
rect 17480 40476 17666 40534
tri 17666 40476 17724 40534 sw
rect 70813 40476 71000 40534
tri 17480 40468 17488 40476 ne
rect 17488 40468 17724 40476
tri 17724 40468 17732 40476 sw
tri 17488 40436 17520 40468 ne
rect 17520 40436 17610 40468
tri 17520 40422 17534 40436 ne
rect 17534 40422 17610 40436
rect 17656 40436 17732 40468
tri 17732 40436 17764 40468 sw
rect 17656 40430 17764 40436
tri 17764 40430 17770 40436 sw
rect 70813 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 17656 40422 17770 40430
tri 17534 40372 17584 40422 ne
rect 17584 40372 17770 40422
tri 17770 40372 17828 40430 sw
rect 70813 40372 71000 40430
tri 17584 40336 17620 40372 ne
rect 17620 40336 17828 40372
tri 17828 40336 17864 40372 sw
tri 17620 40290 17666 40336 ne
rect 17666 40290 17742 40336
rect 17788 40326 17864 40336
tri 17864 40326 17874 40336 sw
rect 70813 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17788 40290 17874 40326
tri 17874 40290 17910 40326 sw
tri 17666 40268 17688 40290 ne
rect 17688 40268 17910 40290
tri 17910 40268 17932 40290 sw
rect 70813 40268 71000 40326
tri 17688 40222 17734 40268 ne
rect 17734 40222 17932 40268
tri 17932 40222 17978 40268 sw
rect 70813 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
tri 17734 40204 17752 40222 ne
rect 17752 40204 17978 40222
tri 17978 40204 17996 40222 sw
tri 17752 40192 17764 40204 ne
rect 17764 40192 17874 40204
tri 17764 40158 17798 40192 ne
rect 17798 40158 17874 40192
rect 17920 40192 17996 40204
tri 17996 40192 18008 40204 sw
rect 17920 40164 18008 40192
tri 18008 40164 18036 40192 sw
rect 70813 40164 71000 40222
rect 17920 40158 18036 40164
tri 17798 40118 17838 40158 ne
rect 17838 40118 18036 40158
tri 18036 40118 18082 40164 sw
rect 70813 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17838 40072 17884 40118 ne
rect 17884 40072 18082 40118
tri 18082 40072 18128 40118 sw
tri 17884 40026 17930 40072 ne
rect 17930 40026 18006 40072
rect 18052 40060 18128 40072
tri 18128 40060 18140 40072 sw
rect 70813 40060 71000 40118
rect 18052 40026 18140 40060
tri 18140 40026 18174 40060 sw
tri 17930 40014 17942 40026 ne
rect 17942 40014 18174 40026
tri 18174 40014 18186 40026 sw
rect 70813 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
tri 17942 39956 18000 40014 ne
rect 18000 39956 18186 40014
tri 18186 39956 18244 40014 sw
rect 70813 39956 71000 40014
tri 18000 39948 18008 39956 ne
rect 18008 39948 18244 39956
tri 18244 39948 18252 39956 sw
tri 18008 39940 18016 39948 ne
rect 18016 39940 18252 39948
tri 18016 39894 18062 39940 ne
rect 18062 39894 18138 39940
rect 18184 39910 18252 39940
tri 18252 39910 18290 39948 sw
rect 70813 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 18184 39894 18290 39910
tri 18062 39852 18104 39894 ne
rect 18104 39852 18290 39894
tri 18290 39852 18348 39910 sw
rect 70813 39852 71000 39910
tri 18104 39808 18148 39852 ne
rect 18148 39808 18348 39852
tri 18348 39808 18392 39852 sw
tri 18148 39762 18194 39808 ne
rect 18194 39762 18270 39808
rect 18316 39806 18392 39808
tri 18392 39806 18394 39808 sw
rect 70813 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39762 18394 39806
tri 18394 39762 18438 39806 sw
tri 18194 39748 18208 39762 ne
rect 18208 39748 18438 39762
tri 18438 39748 18452 39762 sw
rect 70813 39748 71000 39806
tri 18208 39704 18252 39748 ne
rect 18252 39704 18452 39748
tri 18452 39704 18496 39748 sw
tri 18252 39702 18254 39704 ne
rect 18254 39702 18496 39704
tri 18496 39702 18498 39704 sw
rect 70813 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
tri 18254 39676 18280 39702 ne
rect 18280 39676 18498 39702
tri 18280 39630 18326 39676 ne
rect 18326 39630 18402 39676
rect 18448 39644 18498 39676
tri 18498 39644 18556 39702 sw
rect 70813 39644 71000 39702
rect 18448 39630 18556 39644
tri 18326 39598 18358 39630 ne
rect 18358 39598 18556 39630
tri 18556 39598 18602 39644 sw
rect 70813 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18358 39544 18412 39598 ne
rect 18412 39544 18602 39598
tri 18602 39544 18656 39598 sw
tri 18412 39498 18458 39544 ne
rect 18458 39498 18534 39544
rect 18580 39540 18656 39544
tri 18656 39540 18660 39544 sw
rect 70813 39540 71000 39598
rect 18580 39498 18660 39540
tri 18660 39498 18702 39540 sw
tri 18458 39494 18462 39498 ne
rect 18462 39494 18702 39498
tri 18702 39494 18706 39498 sw
rect 70813 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18462 39460 18496 39494 ne
rect 18496 39460 18706 39494
tri 18706 39460 18740 39494 sw
tri 18496 39436 18520 39460 ne
rect 18520 39436 18740 39460
tri 18740 39436 18764 39460 sw
rect 70813 39436 71000 39494
tri 18520 39412 18544 39436 ne
rect 18544 39412 18764 39436
tri 18544 39366 18590 39412 ne
rect 18590 39366 18666 39412
rect 18712 39390 18764 39412
tri 18764 39390 18810 39436 sw
rect 70813 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 18712 39366 18810 39390
tri 18590 39332 18624 39366 ne
rect 18624 39332 18810 39366
tri 18810 39332 18868 39390 sw
rect 70813 39332 71000 39390
tri 18624 39286 18670 39332 ne
rect 18670 39286 18868 39332
tri 18868 39286 18914 39332 sw
rect 70813 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
tri 18670 39280 18676 39286 ne
rect 18676 39280 18914 39286
tri 18914 39280 18920 39286 sw
tri 18676 39234 18722 39280 ne
rect 18722 39234 18798 39280
rect 18844 39234 18920 39280
tri 18920 39234 18966 39280 sw
tri 18722 39228 18728 39234 ne
rect 18728 39228 18966 39234
tri 18966 39228 18972 39234 sw
rect 70813 39228 71000 39286
tri 18728 39216 18740 39228 ne
rect 18740 39216 18972 39228
tri 18972 39216 18984 39228 sw
tri 18740 39182 18774 39216 ne
rect 18774 39182 18984 39216
tri 18984 39182 19018 39216 sw
rect 70813 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
tri 18774 39148 18808 39182 ne
rect 18808 39148 19018 39182
tri 18808 39102 18854 39148 ne
rect 18854 39102 18930 39148
rect 18976 39124 19018 39148
tri 19018 39124 19076 39182 sw
rect 70813 39124 71000 39182
rect 18976 39102 19076 39124
tri 18854 39078 18878 39102 ne
rect 18878 39078 19076 39102
tri 19076 39078 19122 39124 sw
rect 70813 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18878 39020 18936 39078 ne
rect 18936 39020 19122 39078
tri 19122 39020 19180 39078 sw
rect 70813 39020 71000 39078
tri 18936 39016 18940 39020 ne
rect 18940 39016 19180 39020
tri 19180 39016 19184 39020 sw
tri 18940 38972 18984 39016 ne
rect 18984 38972 19062 39016
tri 18984 38970 18986 38972 ne
rect 18986 38970 19062 38972
rect 19108 38974 19184 39016
tri 19184 38974 19226 39016 sw
rect 70813 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 19108 38972 19226 38974
tri 19226 38972 19228 38974 sw
rect 19108 38970 19228 38972
tri 18986 38916 19040 38970 ne
rect 19040 38916 19228 38970
tri 19228 38916 19284 38972 sw
rect 70813 38916 71000 38974
tri 19040 38884 19072 38916 ne
rect 19072 38884 19284 38916
tri 19284 38884 19316 38916 sw
tri 19072 38838 19118 38884 ne
rect 19118 38838 19194 38884
rect 19240 38870 19316 38884
tri 19316 38870 19330 38884 sw
rect 70813 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38838 19330 38870
tri 19330 38838 19362 38870 sw
tri 19118 38812 19144 38838 ne
rect 19144 38812 19362 38838
tri 19362 38812 19388 38838 sw
rect 70813 38812 71000 38870
tri 19144 38766 19190 38812 ne
rect 19190 38766 19388 38812
tri 19388 38766 19434 38812 sw
rect 70813 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19190 38752 19204 38766 ne
rect 19204 38752 19434 38766
tri 19434 38752 19448 38766 sw
tri 19204 38728 19228 38752 ne
rect 19228 38728 19326 38752
tri 19228 38706 19250 38728 ne
rect 19250 38706 19326 38728
rect 19372 38728 19448 38752
tri 19448 38728 19472 38752 sw
rect 19372 38708 19472 38728
tri 19472 38708 19492 38728 sw
rect 70813 38708 71000 38766
rect 19372 38706 19492 38708
tri 19250 38662 19294 38706 ne
rect 19294 38662 19492 38706
tri 19492 38662 19538 38708 sw
rect 70813 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19294 38620 19336 38662 ne
rect 19336 38620 19538 38662
tri 19538 38620 19580 38662 sw
tri 19336 38574 19382 38620 ne
rect 19382 38574 19458 38620
rect 19504 38604 19580 38620
tri 19580 38604 19596 38620 sw
rect 70813 38604 71000 38662
rect 19504 38574 19596 38604
tri 19596 38574 19626 38604 sw
tri 19382 38558 19398 38574 ne
rect 19398 38558 19626 38574
tri 19626 38558 19642 38574 sw
rect 70813 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
tri 19398 38500 19456 38558 ne
rect 19456 38500 19642 38558
tri 19642 38500 19700 38558 sw
rect 70813 38500 71000 38558
tri 19456 38488 19468 38500 ne
rect 19468 38488 19700 38500
tri 19700 38488 19712 38500 sw
tri 19468 38484 19472 38488 ne
rect 19472 38484 19590 38488
tri 19472 38442 19514 38484 ne
rect 19514 38442 19590 38484
rect 19636 38484 19712 38488
tri 19712 38484 19716 38488 sw
rect 19636 38454 19716 38484
tri 19716 38454 19746 38484 sw
rect 70813 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19746 38454
tri 19514 38396 19560 38442 ne
rect 19560 38396 19746 38442
tri 19746 38396 19804 38454 sw
rect 70813 38396 71000 38454
tri 19560 38356 19600 38396 ne
rect 19600 38356 19804 38396
tri 19804 38356 19844 38396 sw
tri 19600 38310 19646 38356 ne
rect 19646 38310 19722 38356
rect 19768 38350 19844 38356
tri 19844 38350 19850 38356 sw
rect 70813 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 19768 38310 19850 38350
tri 19850 38310 19890 38350 sw
tri 19646 38292 19664 38310 ne
rect 19664 38292 19890 38310
tri 19890 38292 19908 38310 sw
rect 70813 38292 71000 38350
tri 19664 38246 19710 38292 ne
rect 19710 38246 19908 38292
tri 19908 38246 19954 38292 sw
rect 70813 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
tri 19710 38240 19716 38246 ne
rect 19716 38240 19954 38246
tri 19954 38240 19960 38246 sw
tri 19716 38224 19732 38240 ne
rect 19732 38224 19960 38240
tri 19732 38178 19778 38224 ne
rect 19778 38178 19854 38224
rect 19900 38188 19960 38224
tri 19960 38188 20012 38240 sw
rect 70813 38188 71000 38246
rect 19900 38178 20012 38188
tri 19778 38142 19814 38178 ne
rect 19814 38142 20012 38178
tri 20012 38142 20058 38188 sw
rect 70813 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
tri 19814 38092 19864 38142 ne
rect 19864 38092 20058 38142
tri 20058 38092 20108 38142 sw
tri 19864 38046 19910 38092 ne
rect 19910 38046 19986 38092
rect 20032 38084 20108 38092
tri 20108 38084 20116 38092 sw
rect 70813 38084 71000 38142
rect 20032 38046 20116 38084
tri 20116 38046 20154 38084 sw
tri 19910 38038 19918 38046 ne
rect 19918 38038 20154 38046
tri 20154 38038 20162 38046 sw
rect 70813 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
tri 19918 37996 19960 38038 ne
rect 19960 37996 20162 38038
tri 20162 37996 20204 38038 sw
tri 19960 37980 19976 37996 ne
rect 19976 37980 20204 37996
tri 20204 37980 20220 37996 sw
rect 70813 37980 71000 38038
tri 19976 37960 19996 37980 ne
rect 19996 37960 20220 37980
tri 19996 37914 20042 37960 ne
rect 20042 37914 20118 37960
rect 20164 37934 20220 37960
tri 20220 37934 20266 37980 sw
rect 70813 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 20164 37914 20266 37934
tri 20042 37876 20080 37914 ne
rect 20080 37876 20266 37914
tri 20266 37876 20324 37934 sw
rect 70813 37876 71000 37934
tri 20080 37830 20126 37876 ne
rect 20126 37830 20324 37876
tri 20324 37830 20370 37876 sw
rect 70813 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
tri 20126 37828 20128 37830 ne
rect 20128 37828 20370 37830
tri 20370 37828 20372 37830 sw
tri 20128 37782 20174 37828 ne
rect 20174 37782 20250 37828
rect 20296 37782 20372 37828
tri 20372 37782 20418 37828 sw
tri 20174 37772 20184 37782 ne
rect 20184 37772 20418 37782
tri 20418 37772 20428 37782 sw
rect 70813 37772 71000 37830
tri 20184 37752 20204 37772 ne
rect 20204 37752 20428 37772
tri 20428 37752 20448 37772 sw
tri 20204 37726 20230 37752 ne
rect 20230 37726 20448 37752
tri 20448 37726 20474 37752 sw
rect 70813 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
tri 20230 37696 20260 37726 ne
rect 20260 37696 20474 37726
tri 20260 37650 20306 37696 ne
rect 20306 37650 20382 37696
rect 20428 37668 20474 37696
tri 20474 37668 20532 37726 sw
rect 70813 37668 71000 37726
rect 20428 37650 20532 37668
tri 20306 37622 20334 37650 ne
rect 20334 37622 20532 37650
tri 20532 37622 20578 37668 sw
rect 70813 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20334 37564 20392 37622 ne
rect 20392 37564 20578 37622
tri 20578 37564 20636 37622 sw
rect 70813 37564 71000 37622
tri 20392 37518 20438 37564 ne
rect 20438 37518 20514 37564
rect 20560 37518 20636 37564
tri 20636 37518 20682 37564 sw
rect 70813 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
tri 20438 37508 20448 37518 ne
rect 20448 37508 20682 37518
tri 20682 37508 20692 37518 sw
tri 20448 37460 20496 37508 ne
rect 20496 37460 20692 37508
tri 20692 37460 20740 37508 sw
rect 70813 37460 71000 37518
tri 20496 37432 20524 37460 ne
rect 20524 37432 20740 37460
tri 20524 37386 20570 37432 ne
rect 20570 37386 20646 37432
rect 20692 37414 20740 37432
tri 20740 37414 20786 37460 sw
rect 70813 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 20692 37386 20786 37414
tri 20570 37356 20600 37386 ne
rect 20600 37356 20786 37386
tri 20786 37356 20844 37414 sw
rect 70813 37356 71000 37414
tri 20600 37310 20646 37356 ne
rect 20646 37310 20844 37356
tri 20844 37310 20890 37356 sw
rect 70813 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
tri 20646 37300 20656 37310 ne
rect 20656 37300 20890 37310
tri 20890 37300 20900 37310 sw
tri 20656 37264 20692 37300 ne
rect 20692 37264 20778 37300
tri 20692 37254 20702 37264 ne
rect 20702 37254 20778 37264
rect 20824 37264 20900 37300
tri 20900 37264 20936 37300 sw
rect 20824 37254 20936 37264
tri 20702 37252 20704 37254 ne
rect 20704 37252 20936 37254
tri 20936 37252 20948 37264 sw
rect 70813 37252 71000 37310
tri 20704 37206 20750 37252 ne
rect 20750 37206 20948 37252
tri 20948 37206 20994 37252 sw
rect 70813 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
tri 20750 37168 20788 37206 ne
rect 20788 37168 20994 37206
tri 20994 37168 21032 37206 sw
tri 20788 37122 20834 37168 ne
rect 20834 37122 20910 37168
rect 20956 37148 21032 37168
tri 21032 37148 21052 37168 sw
rect 70813 37148 71000 37206
rect 20956 37122 21052 37148
tri 21052 37122 21078 37148 sw
tri 20834 37102 20854 37122 ne
rect 20854 37102 21078 37122
tri 21078 37102 21098 37122 sw
rect 70813 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20854 37044 20912 37102 ne
rect 20912 37044 21098 37102
tri 21098 37044 21156 37102 sw
rect 70813 37044 71000 37102
tri 20912 37036 20920 37044 ne
rect 20920 37036 21156 37044
tri 21156 37036 21164 37044 sw
tri 20920 37020 20936 37036 ne
rect 20936 37020 21042 37036
tri 20936 36990 20966 37020 ne
rect 20966 36990 21042 37020
rect 21088 37020 21164 37036
tri 21164 37020 21180 37036 sw
rect 21088 36998 21180 37020
tri 21180 36998 21202 37020 sw
rect 70813 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 21088 36990 21202 36998
tri 20966 36940 21016 36990 ne
rect 21016 36940 21202 36990
tri 21202 36940 21260 36998 sw
rect 70813 36940 71000 36998
tri 21016 36904 21052 36940 ne
rect 21052 36904 21260 36940
tri 21260 36904 21296 36940 sw
tri 21052 36858 21098 36904 ne
rect 21098 36858 21174 36904
rect 21220 36894 21296 36904
tri 21296 36894 21306 36904 sw
rect 70813 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 21220 36858 21306 36894
tri 21306 36858 21342 36894 sw
tri 21098 36836 21120 36858 ne
rect 21120 36836 21342 36858
tri 21342 36836 21364 36858 sw
rect 70813 36836 71000 36894
tri 21120 36790 21166 36836 ne
rect 21166 36790 21364 36836
tri 21364 36790 21410 36836 sw
rect 70813 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
tri 21166 36776 21180 36790 ne
rect 21180 36776 21410 36790
tri 21410 36776 21424 36790 sw
tri 21180 36772 21184 36776 ne
rect 21184 36772 21424 36776
tri 21184 36726 21230 36772 ne
rect 21230 36726 21306 36772
rect 21352 36732 21424 36772
tri 21424 36732 21468 36776 sw
rect 70813 36732 71000 36790
rect 21352 36726 21468 36732
tri 21230 36686 21270 36726 ne
rect 21270 36686 21468 36726
tri 21468 36686 21514 36732 sw
rect 70813 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
tri 21270 36640 21316 36686 ne
rect 21316 36640 21514 36686
tri 21514 36640 21560 36686 sw
tri 21316 36594 21362 36640 ne
rect 21362 36594 21438 36640
rect 21484 36628 21560 36640
tri 21560 36628 21572 36640 sw
rect 70813 36628 71000 36686
rect 21484 36594 21572 36628
tri 21572 36594 21606 36628 sw
tri 21362 36582 21374 36594 ne
rect 21374 36582 21606 36594
tri 21606 36582 21618 36594 sw
rect 70813 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21374 36532 21424 36582 ne
rect 21424 36532 21618 36582
tri 21618 36532 21668 36582 sw
tri 21424 36524 21432 36532 ne
rect 21432 36524 21668 36532
tri 21668 36524 21676 36532 sw
rect 70813 36524 71000 36582
tri 21432 36508 21448 36524 ne
rect 21448 36508 21676 36524
tri 21448 36462 21494 36508 ne
rect 21494 36462 21570 36508
rect 21616 36478 21676 36508
tri 21676 36478 21722 36524 sw
rect 70813 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 21616 36462 21722 36478
tri 21494 36420 21536 36462 ne
rect 21536 36420 21722 36462
tri 21722 36420 21780 36478 sw
rect 70813 36420 71000 36478
tri 21536 36376 21580 36420 ne
rect 21580 36376 21780 36420
tri 21780 36376 21824 36420 sw
tri 21580 36330 21626 36376 ne
rect 21626 36330 21702 36376
rect 21748 36374 21824 36376
tri 21824 36374 21826 36376 sw
rect 70813 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36330 21826 36374
tri 21826 36330 21870 36374 sw
tri 21626 36316 21640 36330 ne
rect 21640 36316 21870 36330
tri 21870 36316 21884 36330 sw
rect 70813 36316 71000 36374
tri 21640 36288 21668 36316 ne
rect 21668 36288 21884 36316
tri 21884 36288 21912 36316 sw
tri 21668 36270 21686 36288 ne
rect 21686 36270 21912 36288
tri 21912 36270 21930 36288 sw
rect 70813 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
tri 21686 36244 21712 36270 ne
rect 21712 36244 21930 36270
tri 21712 36198 21758 36244 ne
rect 21758 36198 21834 36244
rect 21880 36212 21930 36244
tri 21930 36212 21988 36270 sw
rect 70813 36212 71000 36270
rect 21880 36198 21988 36212
tri 21758 36166 21790 36198 ne
rect 21790 36166 21988 36198
tri 21988 36166 22034 36212 sw
rect 70813 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21790 36112 21844 36166 ne
rect 21844 36112 22034 36166
tri 22034 36112 22088 36166 sw
tri 21844 36066 21890 36112 ne
rect 21890 36066 21966 36112
rect 22012 36108 22088 36112
tri 22088 36108 22092 36112 sw
rect 70813 36108 71000 36166
rect 22012 36066 22092 36108
tri 22092 36066 22134 36108 sw
tri 21890 36062 21894 36066 ne
rect 21894 36062 22134 36066
tri 22134 36062 22138 36066 sw
rect 70813 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
tri 21894 36044 21912 36062 ne
rect 21912 36044 22138 36062
tri 22138 36044 22156 36062 sw
tri 21912 36004 21952 36044 ne
rect 21952 36004 22156 36044
tri 22156 36004 22196 36044 sw
rect 70813 36004 71000 36062
tri 21952 35980 21976 36004 ne
rect 21976 35980 22196 36004
tri 21976 35934 22022 35980 ne
rect 22022 35934 22098 35980
rect 22144 35958 22196 35980
tri 22196 35958 22242 36004 sw
rect 70813 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22144 35934 22242 35958
tri 22022 35900 22056 35934 ne
rect 22056 35900 22242 35934
tri 22242 35900 22300 35958 sw
rect 70813 35900 71000 35958
tri 22056 35854 22102 35900 ne
rect 22102 35854 22300 35900
tri 22300 35854 22346 35900 sw
rect 70813 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
tri 22102 35848 22108 35854 ne
rect 22108 35848 22346 35854
tri 22346 35848 22352 35854 sw
tri 22108 35802 22154 35848 ne
rect 22154 35802 22230 35848
rect 22276 35802 22352 35848
tri 22352 35802 22398 35848 sw
tri 22154 35800 22156 35802 ne
rect 22156 35800 22398 35802
tri 22398 35800 22400 35802 sw
tri 22156 35796 22160 35800 ne
rect 22160 35796 22400 35800
tri 22400 35796 22404 35800 sw
rect 70813 35796 71000 35854
tri 22160 35750 22206 35796 ne
rect 22206 35750 22404 35796
tri 22404 35750 22450 35796 sw
rect 70813 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22206 35716 22240 35750 ne
rect 22240 35716 22450 35750
tri 22450 35716 22484 35750 sw
tri 22240 35670 22286 35716 ne
rect 22286 35670 22362 35716
rect 22408 35692 22484 35716
tri 22484 35692 22508 35716 sw
rect 70813 35692 71000 35750
rect 22408 35670 22508 35692
tri 22508 35670 22530 35692 sw
tri 22286 35646 22310 35670 ne
rect 22310 35646 22530 35670
tri 22530 35646 22554 35670 sw
rect 70813 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
tri 22310 35588 22368 35646 ne
rect 22368 35588 22554 35646
tri 22554 35588 22612 35646 sw
rect 70813 35588 71000 35646
tri 22368 35584 22372 35588 ne
rect 22372 35584 22612 35588
tri 22612 35584 22616 35588 sw
tri 22372 35556 22400 35584 ne
rect 22400 35556 22494 35584
tri 22400 35538 22418 35556 ne
rect 22418 35538 22494 35556
rect 22540 35556 22616 35584
tri 22616 35556 22644 35584 sw
rect 22540 35542 22644 35556
tri 22644 35542 22658 35556 sw
rect 70813 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 22540 35538 22658 35542
tri 22418 35484 22472 35538 ne
rect 22472 35484 22658 35538
tri 22658 35484 22716 35542 sw
rect 70813 35484 71000 35542
tri 22472 35452 22504 35484 ne
rect 22504 35452 22716 35484
tri 22716 35452 22748 35484 sw
tri 22504 35406 22550 35452 ne
rect 22550 35406 22626 35452
rect 22672 35438 22748 35452
tri 22748 35438 22762 35452 sw
rect 70813 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35406 22762 35438
tri 22762 35406 22794 35438 sw
tri 22550 35380 22576 35406 ne
rect 22576 35380 22794 35406
tri 22794 35380 22820 35406 sw
rect 70813 35380 71000 35438
tri 22576 35334 22622 35380 ne
rect 22622 35334 22820 35380
tri 22820 35334 22866 35380 sw
rect 70813 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
tri 22622 35320 22636 35334 ne
rect 22636 35320 22866 35334
tri 22866 35320 22880 35334 sw
tri 22636 35312 22644 35320 ne
rect 22644 35312 22758 35320
tri 22644 35274 22682 35312 ne
rect 22682 35274 22758 35312
rect 22804 35312 22880 35320
tri 22880 35312 22888 35320 sw
rect 22804 35276 22888 35312
tri 22888 35276 22924 35312 sw
rect 70813 35276 71000 35334
rect 22804 35274 22924 35276
tri 22682 35230 22726 35274 ne
rect 22726 35230 22924 35274
tri 22924 35230 22970 35276 sw
rect 70813 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22726 35188 22768 35230 ne
rect 22768 35188 22970 35230
tri 22970 35188 23012 35230 sw
tri 22768 35142 22814 35188 ne
rect 22814 35142 22890 35188
rect 22936 35172 23012 35188
tri 23012 35172 23028 35188 sw
rect 70813 35172 71000 35230
rect 22936 35142 23028 35172
tri 23028 35142 23058 35172 sw
tri 22814 35126 22830 35142 ne
rect 22830 35126 23058 35142
tri 23058 35126 23074 35142 sw
rect 70813 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
tri 22830 35068 22888 35126 ne
rect 22888 35068 23074 35126
tri 23074 35068 23132 35126 sw
rect 70813 35068 71000 35126
tri 22888 35056 22900 35068 ne
rect 22900 35056 23132 35068
tri 22900 35010 22946 35056 ne
rect 22946 35010 23022 35056
rect 23068 35022 23132 35056
tri 23132 35022 23178 35068 sw
rect 70813 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 23068 35010 23178 35022
tri 22946 34964 22992 35010 ne
rect 22992 34964 23178 35010
tri 23178 34964 23236 35022 sw
rect 70813 34964 71000 35022
tri 22992 34924 23032 34964 ne
rect 23032 34924 23236 34964
tri 23236 34924 23276 34964 sw
tri 23032 34878 23078 34924 ne
rect 23078 34878 23154 34924
rect 23200 34918 23276 34924
tri 23276 34918 23282 34924 sw
rect 70813 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34878 23282 34918
tri 23282 34878 23322 34918 sw
tri 23078 34860 23096 34878 ne
rect 23096 34860 23322 34878
tri 23322 34860 23340 34878 sw
rect 70813 34860 71000 34918
tri 23096 34824 23132 34860 ne
rect 23132 34824 23340 34860
tri 23340 34824 23376 34860 sw
tri 23132 34814 23142 34824 ne
rect 23142 34814 23376 34824
tri 23376 34814 23386 34824 sw
rect 70813 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
tri 23142 34792 23164 34814 ne
rect 23164 34792 23386 34814
tri 23164 34746 23210 34792 ne
rect 23210 34746 23286 34792
rect 23332 34756 23386 34792
tri 23386 34756 23444 34814 sw
rect 70813 34756 71000 34814
rect 23332 34746 23444 34756
tri 23210 34710 23246 34746 ne
rect 23246 34710 23444 34746
tri 23444 34710 23490 34756 sw
rect 70813 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23246 34660 23296 34710 ne
rect 23296 34660 23490 34710
tri 23490 34660 23540 34710 sw
tri 23296 34614 23342 34660 ne
rect 23342 34614 23418 34660
rect 23464 34652 23540 34660
tri 23540 34652 23548 34660 sw
rect 70813 34652 71000 34710
rect 23464 34614 23548 34652
tri 23548 34614 23586 34652 sw
tri 23342 34606 23350 34614 ne
rect 23350 34606 23586 34614
tri 23586 34606 23594 34614 sw
rect 70813 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
tri 23350 34580 23376 34606 ne
rect 23376 34580 23594 34606
tri 23594 34580 23620 34606 sw
tri 23376 34548 23408 34580 ne
rect 23408 34548 23620 34580
tri 23620 34548 23652 34580 sw
rect 70813 34548 71000 34606
tri 23408 34528 23428 34548 ne
rect 23428 34528 23652 34548
tri 23428 34482 23474 34528 ne
rect 23474 34482 23550 34528
rect 23596 34502 23652 34528
tri 23652 34502 23698 34548 sw
rect 70813 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 23596 34482 23698 34502
tri 23474 34444 23512 34482 ne
rect 23512 34444 23698 34482
tri 23698 34444 23756 34502 sw
rect 70813 34444 71000 34502
tri 23512 34398 23558 34444 ne
rect 23558 34398 23756 34444
tri 23756 34398 23802 34444 sw
rect 70813 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
tri 23558 34396 23560 34398 ne
rect 23560 34396 23802 34398
tri 23802 34396 23804 34398 sw
tri 23560 34350 23606 34396 ne
rect 23606 34350 23682 34396
rect 23728 34350 23804 34396
tri 23804 34350 23850 34396 sw
tri 23606 34340 23616 34350 ne
rect 23616 34340 23850 34350
tri 23850 34340 23860 34350 sw
rect 70813 34340 71000 34398
tri 23616 34336 23620 34340 ne
rect 23620 34336 23860 34340
tri 23860 34336 23864 34340 sw
tri 23620 34294 23662 34336 ne
rect 23662 34294 23864 34336
tri 23864 34294 23906 34336 sw
rect 70813 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23662 34264 23692 34294 ne
rect 23692 34264 23906 34294
tri 23692 34218 23738 34264 ne
rect 23738 34218 23814 34264
rect 23860 34236 23906 34264
tri 23906 34236 23964 34294 sw
rect 70813 34236 71000 34294
rect 23860 34218 23964 34236
tri 23738 34190 23766 34218 ne
rect 23766 34190 23964 34218
tri 23964 34190 24010 34236 sw
rect 70813 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
tri 23766 34132 23824 34190 ne
rect 23824 34132 24010 34190
tri 24010 34132 24068 34190 sw
rect 70813 34132 71000 34190
tri 23824 34092 23864 34132 ne
rect 23864 34092 23946 34132
tri 23864 34086 23870 34092 ne
rect 23870 34086 23946 34092
rect 23992 34092 24068 34132
tri 24068 34092 24108 34132 sw
rect 23992 34086 24108 34092
tri 24108 34086 24114 34092 sw
rect 70813 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
tri 23870 34028 23928 34086 ne
rect 23928 34028 24114 34086
tri 24114 34028 24172 34086 sw
rect 70813 34028 71000 34086
tri 23928 34000 23956 34028 ne
rect 23956 34000 24172 34028
tri 24172 34000 24200 34028 sw
tri 23956 33954 24002 34000 ne
rect 24002 33954 24078 34000
rect 24124 33982 24200 34000
tri 24200 33982 24218 34000 sw
rect 70813 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33954 24218 33982
tri 24218 33954 24246 33982 sw
tri 24002 33924 24032 33954 ne
rect 24032 33924 24246 33954
tri 24246 33924 24276 33954 sw
rect 70813 33924 71000 33982
tri 24032 33878 24078 33924 ne
rect 24078 33878 24276 33924
tri 24276 33878 24322 33924 sw
rect 70813 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
tri 24078 33868 24088 33878 ne
rect 24088 33868 24322 33878
tri 24322 33868 24332 33878 sw
tri 24088 33848 24108 33868 ne
rect 24108 33848 24210 33868
tri 24108 33822 24134 33848 ne
rect 24134 33822 24210 33848
rect 24256 33848 24332 33868
tri 24332 33848 24352 33868 sw
rect 24256 33822 24352 33848
tri 24134 33820 24136 33822 ne
rect 24136 33820 24352 33822
tri 24352 33820 24380 33848 sw
rect 70813 33820 71000 33878
tri 24136 33774 24182 33820 ne
rect 24182 33774 24380 33820
tri 24380 33774 24426 33820 sw
rect 70813 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24182 33736 24220 33774 ne
rect 24220 33736 24426 33774
tri 24426 33736 24464 33774 sw
tri 24220 33690 24266 33736 ne
rect 24266 33690 24342 33736
rect 24388 33716 24464 33736
tri 24464 33716 24484 33736 sw
rect 70813 33716 71000 33774
rect 24388 33690 24484 33716
tri 24484 33690 24510 33716 sw
tri 24266 33670 24286 33690 ne
rect 24286 33670 24510 33690
tri 24510 33670 24530 33690 sw
rect 70813 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
tri 24286 33612 24344 33670 ne
rect 24344 33612 24530 33670
tri 24530 33612 24588 33670 sw
rect 70813 33612 71000 33670
tri 24344 33604 24352 33612 ne
rect 24352 33604 24588 33612
tri 24588 33604 24596 33612 sw
tri 24352 33558 24398 33604 ne
rect 24398 33558 24474 33604
rect 24520 33566 24596 33604
tri 24596 33566 24634 33604 sw
rect 70813 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 24520 33558 24634 33566
tri 24398 33508 24448 33558 ne
rect 24448 33508 24634 33558
tri 24634 33508 24692 33566 sw
rect 70813 33508 71000 33566
tri 24448 33472 24484 33508 ne
rect 24484 33472 24692 33508
tri 24692 33472 24728 33508 sw
tri 24484 33426 24530 33472 ne
rect 24530 33426 24606 33472
rect 24652 33462 24728 33472
tri 24728 33462 24738 33472 sw
rect 70813 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24652 33426 24738 33462
tri 24738 33426 24774 33462 sw
tri 24530 33404 24552 33426 ne
rect 24552 33404 24774 33426
tri 24774 33404 24796 33426 sw
rect 70813 33404 71000 33462
tri 24552 33360 24596 33404 ne
rect 24596 33360 24796 33404
tri 24796 33360 24840 33404 sw
tri 24596 33358 24598 33360 ne
rect 24598 33358 24840 33360
tri 24840 33358 24842 33360 sw
rect 70813 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
tri 24598 33340 24616 33358 ne
rect 24616 33340 24842 33358
tri 24616 33294 24662 33340 ne
rect 24662 33294 24738 33340
rect 24784 33300 24842 33340
tri 24842 33300 24900 33358 sw
rect 70813 33300 71000 33358
rect 24784 33294 24900 33300
tri 24662 33254 24702 33294 ne
rect 24702 33254 24900 33294
tri 24900 33254 24946 33300 sw
rect 70813 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24702 33208 24748 33254 ne
rect 24748 33208 24946 33254
tri 24946 33208 24992 33254 sw
tri 24748 33162 24794 33208 ne
rect 24794 33162 24870 33208
rect 24916 33196 24992 33208
tri 24992 33196 25004 33208 sw
rect 70813 33196 71000 33254
rect 24916 33162 25004 33196
tri 25004 33162 25038 33196 sw
tri 24794 33150 24806 33162 ne
rect 24806 33150 25038 33162
tri 25038 33150 25050 33162 sw
rect 70813 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
tri 24806 33116 24840 33150 ne
rect 24840 33116 25050 33150
tri 25050 33116 25084 33150 sw
tri 24840 33092 24864 33116 ne
rect 24864 33092 25084 33116
tri 25084 33092 25108 33116 sw
rect 70813 33092 71000 33150
tri 24864 33076 24880 33092 ne
rect 24880 33076 25108 33092
tri 24880 33030 24926 33076 ne
rect 24926 33030 25002 33076
rect 25048 33046 25108 33076
tri 25108 33046 25154 33092 sw
rect 70813 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 25048 33030 25154 33046
tri 24926 32988 24968 33030 ne
rect 24968 32988 25154 33030
tri 25154 32988 25212 33046 sw
rect 70813 32988 71000 33046
tri 24968 32944 25012 32988 ne
rect 25012 32944 25212 32988
tri 25212 32944 25256 32988 sw
tri 25012 32898 25058 32944 ne
rect 25058 32898 25134 32944
rect 25180 32942 25256 32944
tri 25256 32942 25258 32944 sw
rect 70813 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32898 25258 32942
tri 25258 32898 25302 32942 sw
tri 25058 32884 25072 32898 ne
rect 25072 32884 25302 32898
tri 25302 32884 25316 32898 sw
rect 70813 32884 71000 32942
tri 25072 32872 25084 32884 ne
rect 25084 32872 25316 32884
tri 25316 32872 25328 32884 sw
tri 25084 32838 25118 32872 ne
rect 25118 32838 25328 32872
tri 25328 32838 25362 32872 sw
rect 70813 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
tri 25118 32812 25144 32838 ne
rect 25144 32812 25362 32838
tri 25144 32766 25190 32812 ne
rect 25190 32766 25266 32812
rect 25312 32780 25362 32812
tri 25362 32780 25420 32838 sw
rect 70813 32780 71000 32838
rect 25312 32766 25420 32780
tri 25190 32734 25222 32766 ne
rect 25222 32734 25420 32766
tri 25420 32734 25466 32780 sw
rect 70813 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25222 32680 25276 32734 ne
rect 25276 32680 25466 32734
tri 25466 32680 25520 32734 sw
tri 25276 32634 25322 32680 ne
rect 25322 32634 25398 32680
rect 25444 32676 25520 32680
tri 25520 32676 25524 32680 sw
rect 70813 32676 71000 32734
rect 25444 32634 25524 32676
tri 25524 32634 25566 32676 sw
tri 25322 32630 25326 32634 ne
rect 25326 32630 25566 32634
tri 25566 32630 25570 32634 sw
rect 70813 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25326 32628 25328 32630 ne
rect 25328 32628 25570 32630
tri 25570 32628 25572 32630 sw
tri 25328 32572 25384 32628 ne
rect 25384 32572 25572 32628
tri 25572 32572 25628 32628 sw
rect 70813 32572 71000 32630
tri 25384 32548 25408 32572 ne
rect 25408 32548 25628 32572
tri 25628 32548 25652 32572 sw
tri 25408 32502 25454 32548 ne
rect 25454 32502 25530 32548
rect 25576 32526 25652 32548
tri 25652 32526 25674 32548 sw
rect 70813 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 25576 32502 25674 32526
tri 25674 32502 25698 32526 sw
tri 25454 32468 25488 32502 ne
rect 25488 32468 25698 32502
tri 25698 32468 25732 32502 sw
rect 70813 32468 71000 32526
tri 25488 32422 25534 32468 ne
rect 25534 32422 25732 32468
tri 25732 32422 25778 32468 sw
rect 70813 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
tri 25534 32416 25540 32422 ne
rect 25540 32416 25778 32422
tri 25778 32416 25784 32422 sw
tri 25540 32384 25572 32416 ne
rect 25572 32384 25662 32416
tri 25572 32370 25586 32384 ne
rect 25586 32370 25662 32384
rect 25708 32384 25784 32416
tri 25784 32384 25816 32416 sw
rect 25708 32370 25816 32384
tri 25586 32364 25592 32370 ne
rect 25592 32364 25816 32370
tri 25816 32364 25836 32384 sw
rect 70813 32364 71000 32422
tri 25592 32318 25638 32364 ne
rect 25638 32318 25836 32364
tri 25836 32318 25882 32364 sw
rect 70813 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
tri 25638 32284 25672 32318 ne
rect 25672 32284 25882 32318
tri 25882 32284 25916 32318 sw
tri 25672 32238 25718 32284 ne
rect 25718 32238 25794 32284
rect 25840 32260 25916 32284
tri 25916 32260 25940 32284 sw
rect 70813 32260 71000 32318
rect 25840 32238 25940 32260
tri 25940 32238 25962 32260 sw
tri 25718 32214 25742 32238 ne
rect 25742 32214 25962 32238
tri 25962 32214 25986 32238 sw
rect 70813 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25742 32156 25800 32214 ne
rect 25800 32156 25986 32214
tri 25986 32156 26044 32214 sw
rect 70813 32156 71000 32214
tri 25800 32152 25804 32156 ne
rect 25804 32152 26044 32156
tri 26044 32152 26048 32156 sw
tri 25804 32140 25816 32152 ne
rect 25816 32140 25926 32152
tri 25816 32106 25850 32140 ne
rect 25850 32106 25926 32140
rect 25972 32140 26048 32152
tri 26048 32140 26060 32152 sw
rect 25972 32110 26060 32140
tri 26060 32110 26090 32140 sw
rect 70813 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 25972 32106 26090 32110
tri 25850 32052 25904 32106 ne
rect 25904 32052 26090 32106
tri 26090 32052 26148 32110 sw
rect 70813 32052 71000 32110
tri 25904 32020 25936 32052 ne
rect 25936 32020 26148 32052
tri 26148 32020 26180 32052 sw
tri 25936 31974 25982 32020 ne
rect 25982 31974 26058 32020
rect 26104 32006 26180 32020
tri 26180 32006 26194 32020 sw
rect 70813 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 26104 31974 26194 32006
tri 26194 31974 26226 32006 sw
tri 25982 31948 26008 31974 ne
rect 26008 31948 26226 31974
tri 26226 31948 26252 31974 sw
rect 70813 31948 71000 32006
tri 26008 31902 26054 31948 ne
rect 26054 31902 26252 31948
tri 26252 31902 26298 31948 sw
rect 70813 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
tri 26054 31896 26060 31902 ne
rect 26060 31896 26298 31902
tri 26298 31896 26304 31902 sw
tri 26060 31888 26068 31896 ne
rect 26068 31888 26304 31896
tri 26068 31842 26114 31888 ne
rect 26114 31842 26190 31888
rect 26236 31844 26304 31888
tri 26304 31844 26356 31896 sw
rect 70813 31844 71000 31902
rect 26236 31842 26356 31844
tri 26114 31798 26158 31842 ne
rect 26158 31798 26356 31842
tri 26356 31798 26402 31844 sw
rect 70813 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
tri 26158 31756 26200 31798 ne
rect 26200 31756 26402 31798
tri 26402 31756 26444 31798 sw
tri 26200 31710 26246 31756 ne
rect 26246 31710 26322 31756
rect 26368 31740 26444 31756
tri 26444 31740 26460 31756 sw
rect 70813 31740 71000 31798
rect 26368 31710 26460 31740
tri 26460 31710 26490 31740 sw
tri 26246 31694 26262 31710 ne
rect 26262 31694 26490 31710
tri 26490 31694 26506 31710 sw
rect 70813 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
tri 26262 31652 26304 31694 ne
rect 26304 31652 26506 31694
tri 26506 31652 26548 31694 sw
tri 26304 31636 26320 31652 ne
rect 26320 31636 26548 31652
tri 26548 31636 26564 31652 sw
rect 70813 31636 71000 31694
tri 26320 31624 26332 31636 ne
rect 26332 31624 26564 31636
tri 26332 31578 26378 31624 ne
rect 26378 31578 26454 31624
rect 26500 31590 26564 31624
tri 26564 31590 26610 31636 sw
rect 70813 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 26500 31578 26610 31590
tri 26378 31532 26424 31578 ne
rect 26424 31532 26610 31578
tri 26610 31532 26668 31590 sw
rect 70813 31532 71000 31590
tri 26424 31492 26464 31532 ne
rect 26464 31492 26668 31532
tri 26668 31492 26708 31532 sw
tri 26464 31446 26510 31492 ne
rect 26510 31446 26586 31492
rect 26632 31486 26708 31492
tri 26708 31486 26714 31492 sw
rect 70813 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31446 26714 31486
tri 26714 31446 26754 31486 sw
tri 26510 31428 26528 31446 ne
rect 26528 31428 26754 31446
tri 26754 31428 26772 31446 sw
rect 70813 31428 71000 31486
tri 26528 31408 26548 31428 ne
rect 26548 31408 26772 31428
tri 26772 31408 26792 31428 sw
tri 26548 31382 26574 31408 ne
rect 26574 31382 26792 31408
tri 26792 31382 26818 31408 sw
rect 70813 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
tri 26574 31360 26596 31382 ne
rect 26596 31360 26818 31382
tri 26596 31314 26642 31360 ne
rect 26642 31314 26718 31360
rect 26764 31324 26818 31360
tri 26818 31324 26876 31382 sw
rect 70813 31324 71000 31382
rect 26764 31314 26876 31324
tri 26642 31278 26678 31314 ne
rect 26678 31278 26876 31314
tri 26876 31278 26922 31324 sw
rect 70813 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
tri 26678 31228 26728 31278 ne
rect 26728 31228 26922 31278
tri 26922 31228 26972 31278 sw
tri 26728 31182 26774 31228 ne
rect 26774 31182 26850 31228
rect 26896 31220 26972 31228
tri 26972 31220 26980 31228 sw
rect 70813 31220 71000 31278
rect 26896 31182 26980 31220
tri 26980 31182 27018 31220 sw
tri 26774 31174 26782 31182 ne
rect 26782 31174 27018 31182
tri 27018 31174 27026 31182 sw
rect 70813 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
tri 26782 31164 26792 31174 ne
rect 26792 31164 27026 31174
tri 27026 31164 27036 31174 sw
tri 26792 31116 26840 31164 ne
rect 26840 31116 27036 31164
tri 27036 31116 27084 31164 sw
rect 70813 31116 71000 31174
tri 26840 31096 26860 31116 ne
rect 26860 31096 27084 31116
tri 26860 31050 26906 31096 ne
rect 26906 31050 26982 31096
rect 27028 31070 27084 31096
tri 27084 31070 27130 31116 sw
rect 70813 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 27028 31050 27130 31070
tri 26906 31012 26944 31050 ne
rect 26944 31012 27130 31050
tri 27130 31012 27188 31070 sw
rect 70813 31012 71000 31070
tri 26944 30966 26990 31012 ne
rect 26990 30966 27188 31012
tri 27188 30966 27234 31012 sw
rect 70813 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
tri 26990 30964 26992 30966 ne
rect 26992 30964 27234 30966
tri 27234 30964 27236 30966 sw
tri 26992 30920 27036 30964 ne
rect 27036 30920 27114 30964
tri 27036 30918 27038 30920 ne
rect 27038 30918 27114 30920
rect 27160 30920 27236 30964
tri 27236 30920 27280 30964 sw
rect 27160 30918 27280 30920
tri 27038 30908 27048 30918 ne
rect 27048 30908 27280 30918
tri 27280 30908 27292 30920 sw
rect 70813 30908 71000 30966
tri 27048 30862 27094 30908 ne
rect 27094 30862 27292 30908
tri 27292 30862 27338 30908 sw
rect 70813 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
tri 27094 30832 27124 30862 ne
rect 27124 30832 27338 30862
tri 27338 30832 27368 30862 sw
tri 27124 30786 27170 30832 ne
rect 27170 30786 27246 30832
rect 27292 30804 27368 30832
tri 27368 30804 27396 30832 sw
rect 70813 30804 71000 30862
rect 27292 30786 27396 30804
tri 27396 30786 27414 30804 sw
tri 27170 30758 27198 30786 ne
rect 27198 30758 27414 30786
tri 27414 30758 27442 30786 sw
rect 70813 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27198 30700 27256 30758 ne
rect 27256 30700 27442 30758
tri 27442 30700 27500 30758 sw
rect 70813 30700 71000 30758
tri 27256 30676 27280 30700 ne
rect 27280 30676 27378 30700
tri 27280 30654 27302 30676 ne
rect 27302 30654 27378 30676
rect 27424 30676 27500 30700
tri 27500 30676 27524 30700 sw
rect 27424 30654 27524 30676
tri 27524 30654 27546 30676 sw
rect 70813 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
tri 27302 30596 27360 30654 ne
rect 27360 30596 27546 30654
tri 27546 30596 27604 30654 sw
rect 70813 30596 71000 30654
tri 27360 30568 27388 30596 ne
rect 27388 30568 27604 30596
tri 27604 30568 27632 30596 sw
tri 27388 30522 27434 30568 ne
rect 27434 30522 27510 30568
rect 27556 30550 27632 30568
tri 27632 30550 27650 30568 sw
rect 70813 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30522 27650 30550
tri 27650 30522 27678 30550 sw
tri 27434 30492 27464 30522 ne
rect 27464 30492 27678 30522
tri 27678 30492 27708 30522 sw
rect 70813 30492 71000 30550
tri 27464 30446 27510 30492 ne
rect 27510 30446 27708 30492
tri 27708 30446 27754 30492 sw
rect 70813 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
tri 27510 30436 27520 30446 ne
rect 27520 30436 27754 30446
tri 27754 30436 27764 30446 sw
tri 27520 30432 27524 30436 ne
rect 27524 30432 27642 30436
tri 27524 30390 27566 30432 ne
rect 27566 30390 27642 30432
rect 27688 30432 27764 30436
tri 27764 30432 27768 30436 sw
rect 27688 30390 27768 30432
tri 27566 30388 27568 30390 ne
rect 27568 30388 27768 30390
tri 27768 30388 27812 30432 sw
rect 70813 30388 71000 30446
tri 27568 30342 27614 30388 ne
rect 27614 30342 27812 30388
tri 27812 30342 27858 30388 sw
rect 70813 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27614 30304 27652 30342 ne
rect 27652 30304 27858 30342
tri 27858 30304 27896 30342 sw
tri 27652 30258 27698 30304 ne
rect 27698 30258 27774 30304
rect 27820 30284 27896 30304
tri 27896 30284 27916 30304 sw
rect 70813 30284 71000 30342
rect 27820 30258 27916 30284
tri 27916 30258 27942 30284 sw
tri 27698 30238 27718 30258 ne
rect 27718 30238 27942 30258
tri 27942 30238 27962 30258 sw
rect 70813 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27718 30188 27768 30238 ne
rect 27768 30188 27962 30238
tri 27962 30188 28012 30238 sw
tri 27768 30180 27776 30188 ne
rect 27776 30180 28012 30188
tri 28012 30180 28020 30188 sw
rect 70813 30180 71000 30238
tri 27776 30172 27784 30180 ne
rect 27784 30172 28020 30180
tri 27784 30126 27830 30172 ne
rect 27830 30126 27906 30172
rect 27952 30134 28020 30172
tri 28020 30134 28066 30180 sw
rect 70813 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 27952 30126 28066 30134
tri 27830 30076 27880 30126 ne
rect 27880 30076 28066 30126
tri 28066 30076 28124 30134 sw
rect 70813 30076 71000 30134
tri 27880 30040 27916 30076 ne
rect 27916 30040 28124 30076
tri 28124 30040 28160 30076 sw
tri 27916 29994 27962 30040 ne
rect 27962 29994 28038 30040
rect 28084 30030 28160 30040
tri 28160 30030 28170 30040 sw
rect 70813 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 29994 28170 30030
tri 28170 29994 28206 30030 sw
tri 27962 29972 27984 29994 ne
rect 27984 29972 28206 29994
tri 28206 29972 28228 29994 sw
rect 70813 29972 71000 30030
tri 27984 29944 28012 29972 ne
rect 28012 29944 28228 29972
tri 28228 29944 28256 29972 sw
tri 28012 29926 28030 29944 ne
rect 28030 29926 28256 29944
tri 28256 29926 28274 29944 sw
rect 70813 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
tri 28030 29908 28048 29926 ne
rect 28048 29908 28274 29926
tri 28048 29862 28094 29908 ne
rect 28094 29862 28170 29908
rect 28216 29868 28274 29908
tri 28274 29868 28332 29926 sw
rect 70813 29868 71000 29926
rect 28216 29862 28332 29868
tri 28094 29822 28134 29862 ne
rect 28134 29822 28332 29862
tri 28332 29822 28378 29868 sw
rect 70813 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
tri 28134 29776 28180 29822 ne
rect 28180 29776 28378 29822
tri 28378 29776 28424 29822 sw
tri 28180 29730 28226 29776 ne
rect 28226 29730 28302 29776
rect 28348 29764 28424 29776
tri 28424 29764 28436 29776 sw
rect 70813 29764 71000 29822
rect 28348 29730 28436 29764
tri 28436 29730 28470 29764 sw
tri 28226 29718 28238 29730 ne
rect 28238 29718 28470 29730
tri 28470 29718 28482 29730 sw
rect 70813 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
tri 28238 29700 28256 29718 ne
rect 28256 29700 28482 29718
tri 28482 29700 28500 29718 sw
tri 28256 29660 28296 29700 ne
rect 28296 29660 28500 29700
tri 28500 29660 28540 29700 sw
rect 70813 29660 71000 29718
tri 28296 29644 28312 29660 ne
rect 28312 29644 28540 29660
tri 28312 29598 28358 29644 ne
rect 28358 29598 28434 29644
rect 28480 29614 28540 29644
tri 28540 29614 28586 29660 sw
rect 70813 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 28480 29598 28586 29614
tri 28358 29556 28400 29598 ne
rect 28400 29556 28586 29598
tri 28586 29556 28644 29614 sw
rect 70813 29556 71000 29614
tri 28400 29512 28444 29556 ne
rect 28444 29512 28644 29556
tri 28644 29512 28688 29556 sw
tri 28444 29466 28490 29512 ne
rect 28490 29466 28566 29512
rect 28612 29510 28688 29512
tri 28688 29510 28690 29512 sw
rect 70813 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29466 28690 29510
tri 28690 29466 28734 29510 sw
tri 28490 29456 28500 29466 ne
rect 28500 29456 28734 29466
tri 28734 29456 28744 29466 sw
tri 28500 29452 28504 29456 ne
rect 28504 29452 28744 29456
tri 28744 29452 28748 29456 sw
rect 70813 29452 71000 29510
tri 28504 29406 28550 29452 ne
rect 28550 29406 28748 29452
tri 28748 29406 28794 29452 sw
rect 70813 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28550 29380 28576 29406 ne
rect 28576 29380 28794 29406
tri 28576 29334 28622 29380 ne
rect 28622 29334 28698 29380
rect 28744 29348 28794 29380
tri 28794 29348 28852 29406 sw
rect 70813 29348 71000 29406
rect 28744 29334 28852 29348
tri 28622 29302 28654 29334 ne
rect 28654 29302 28852 29334
tri 28852 29302 28898 29348 sw
rect 70813 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28654 29248 28708 29302 ne
rect 28708 29248 28898 29302
tri 28898 29248 28952 29302 sw
tri 28708 29212 28744 29248 ne
rect 28744 29212 28830 29248
tri 28744 29202 28754 29212 ne
rect 28754 29202 28830 29212
rect 28876 29244 28952 29248
tri 28952 29244 28956 29248 sw
rect 70813 29244 71000 29302
rect 28876 29212 28956 29244
tri 28956 29212 28988 29244 sw
rect 28876 29202 28988 29212
tri 28754 29198 28758 29202 ne
rect 28758 29198 28988 29202
tri 28988 29198 29002 29212 sw
rect 70813 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
tri 28758 29140 28816 29198 ne
rect 28816 29140 29002 29198
tri 29002 29140 29060 29198 sw
rect 70813 29140 71000 29198
tri 28816 29116 28840 29140 ne
rect 28840 29116 29060 29140
tri 29060 29116 29084 29140 sw
tri 28840 29070 28886 29116 ne
rect 28886 29070 28962 29116
rect 29008 29094 29084 29116
tri 29084 29094 29106 29116 sw
rect 70813 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 29008 29070 29106 29094
tri 29106 29070 29130 29094 sw
tri 28886 29036 28920 29070 ne
rect 28920 29036 29130 29070
tri 29130 29036 29164 29070 sw
rect 70813 29036 71000 29094
tri 28920 28990 28966 29036 ne
rect 28966 28990 29164 29036
tri 29164 28990 29210 29036 sw
rect 70813 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
tri 28966 28984 28972 28990 ne
rect 28972 28984 29210 28990
tri 29210 28984 29216 28990 sw
tri 28972 28968 28988 28984 ne
rect 28988 28968 29094 28984
tri 28988 28938 29018 28968 ne
rect 29018 28938 29094 28968
rect 29140 28968 29216 28984
tri 29216 28968 29232 28984 sw
rect 29140 28938 29232 28968
tri 29018 28932 29024 28938 ne
rect 29024 28932 29232 28938
tri 29232 28932 29268 28968 sw
rect 70813 28932 71000 28990
tri 29024 28886 29070 28932 ne
rect 29070 28886 29268 28932
tri 29268 28886 29314 28932 sw
rect 70813 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29070 28852 29104 28886 ne
rect 29104 28852 29314 28886
tri 29314 28852 29348 28886 sw
tri 29104 28806 29150 28852 ne
rect 29150 28806 29226 28852
rect 29272 28828 29348 28852
tri 29348 28828 29372 28852 sw
rect 70813 28828 71000 28886
rect 29272 28806 29372 28828
tri 29372 28806 29394 28828 sw
tri 29150 28782 29174 28806 ne
rect 29174 28782 29394 28806
tri 29394 28782 29418 28806 sw
rect 70813 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
tri 29174 28724 29232 28782 ne
rect 29232 28724 29418 28782
tri 29418 28724 29476 28782 sw
rect 70813 28724 71000 28782
tri 29232 28720 29236 28724 ne
rect 29236 28720 29476 28724
tri 29236 28674 29282 28720 ne
rect 29282 28674 29358 28720
rect 29404 28678 29476 28720
tri 29476 28678 29522 28724 sw
rect 70813 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 29404 28674 29522 28678
tri 29282 28620 29336 28674 ne
rect 29336 28620 29522 28674
tri 29522 28620 29580 28678 sw
rect 70813 28620 71000 28678
tri 29336 28588 29368 28620 ne
rect 29368 28588 29580 28620
tri 29580 28588 29612 28620 sw
tri 29368 28542 29414 28588 ne
rect 29414 28542 29490 28588
rect 29536 28574 29612 28588
tri 29612 28574 29626 28588 sw
rect 70813 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28542 29626 28574
tri 29626 28542 29658 28574 sw
tri 29414 28516 29440 28542 ne
rect 29440 28516 29658 28542
tri 29658 28516 29684 28542 sw
rect 70813 28516 71000 28574
tri 29440 28480 29476 28516 ne
rect 29476 28480 29684 28516
tri 29684 28480 29720 28516 sw
tri 29476 28470 29486 28480 ne
rect 29486 28470 29720 28480
tri 29720 28470 29730 28480 sw
rect 70813 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
tri 29486 28456 29500 28470 ne
rect 29500 28456 29730 28470
tri 29500 28410 29546 28456 ne
rect 29546 28410 29622 28456
rect 29668 28412 29730 28456
tri 29730 28412 29788 28470 sw
rect 70813 28412 71000 28470
rect 29668 28410 29788 28412
tri 29546 28366 29590 28410 ne
rect 29590 28366 29788 28410
tri 29788 28366 29834 28412 sw
rect 70813 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29590 28324 29632 28366 ne
rect 29632 28324 29834 28366
tri 29834 28324 29876 28366 sw
tri 29632 28278 29678 28324 ne
rect 29678 28278 29754 28324
rect 29800 28308 29876 28324
tri 29876 28308 29892 28324 sw
rect 70813 28308 71000 28366
rect 29800 28278 29892 28308
tri 29892 28278 29922 28308 sw
tri 29678 28262 29694 28278 ne
rect 29694 28262 29922 28278
tri 29922 28262 29938 28278 sw
rect 70813 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
tri 29694 28236 29720 28262 ne
rect 29720 28236 29938 28262
tri 29938 28236 29964 28262 sw
tri 29720 28204 29752 28236 ne
rect 29752 28204 29964 28236
tri 29964 28204 29996 28236 sw
rect 70813 28204 71000 28262
tri 29752 28192 29764 28204 ne
rect 29764 28192 29996 28204
tri 29764 28146 29810 28192 ne
rect 29810 28146 29886 28192
rect 29932 28158 29996 28192
tri 29996 28158 30042 28204 sw
rect 70813 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 29932 28146 30042 28158
tri 29810 28100 29856 28146 ne
rect 29856 28100 30042 28146
tri 30042 28100 30100 28158 sw
rect 70813 28100 71000 28158
tri 29856 28060 29896 28100 ne
rect 29896 28060 30100 28100
tri 30100 28060 30140 28100 sw
tri 29896 28014 29942 28060 ne
rect 29942 28014 30018 28060
rect 30064 28054 30140 28060
tri 30140 28054 30146 28060 sw
rect 70813 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28014 30146 28054
tri 30146 28014 30186 28054 sw
tri 29942 27996 29960 28014 ne
rect 29960 27996 30186 28014
tri 30186 27996 30204 28014 sw
rect 70813 27996 71000 28054
tri 29960 27992 29964 27996 ne
rect 29964 27992 30204 27996
tri 30204 27992 30208 27996 sw
tri 29964 27950 30006 27992 ne
rect 30006 27950 30208 27992
tri 30208 27950 30250 27992 sw
rect 70813 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
tri 30006 27928 30028 27950 ne
rect 30028 27928 30250 27950
tri 30028 27882 30074 27928 ne
rect 30074 27882 30150 27928
rect 30196 27892 30250 27928
tri 30250 27892 30308 27950 sw
rect 70813 27892 71000 27950
rect 30196 27882 30308 27892
tri 30074 27846 30110 27882 ne
rect 30110 27846 30308 27882
tri 30308 27846 30354 27892 sw
rect 70813 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30110 27796 30160 27846 ne
rect 30160 27796 30354 27846
tri 30354 27796 30404 27846 sw
tri 30160 27750 30206 27796 ne
rect 30206 27750 30282 27796
rect 30328 27788 30404 27796
tri 30404 27788 30412 27796 sw
rect 70813 27788 71000 27846
rect 30328 27750 30412 27788
tri 30412 27750 30450 27788 sw
tri 30206 27748 30208 27750 ne
rect 30208 27748 30450 27750
tri 30450 27748 30452 27750 sw
tri 30208 27742 30214 27748 ne
rect 30214 27742 30452 27748
tri 30452 27742 30458 27748 sw
rect 70813 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
tri 30214 27684 30272 27742 ne
rect 30272 27684 30458 27742
tri 30458 27684 30516 27742 sw
rect 70813 27684 71000 27742
tri 30272 27664 30292 27684 ne
rect 30292 27664 30516 27684
tri 30516 27664 30536 27684 sw
tri 30292 27618 30338 27664 ne
rect 30338 27618 30414 27664
rect 30460 27638 30536 27664
tri 30536 27638 30562 27664 sw
rect 70813 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30460 27618 30562 27638
tri 30562 27618 30582 27638 sw
tri 30338 27580 30376 27618 ne
rect 30376 27580 30582 27618
tri 30582 27580 30620 27618 sw
rect 70813 27580 71000 27638
tri 30376 27534 30422 27580 ne
rect 30422 27534 30620 27580
tri 30620 27534 30666 27580 sw
rect 70813 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
tri 30422 27532 30424 27534 ne
rect 30424 27532 30666 27534
tri 30666 27532 30668 27534 sw
tri 30424 27504 30452 27532 ne
rect 30452 27504 30546 27532
tri 30452 27486 30470 27504 ne
rect 30470 27486 30546 27504
rect 30592 27504 30668 27532
tri 30668 27504 30696 27532 sw
rect 30592 27486 30696 27504
tri 30470 27476 30480 27486 ne
rect 30480 27476 30696 27486
tri 30696 27476 30724 27504 sw
rect 70813 27476 71000 27534
tri 30480 27430 30526 27476 ne
rect 30526 27430 30724 27476
tri 30724 27430 30770 27476 sw
rect 70813 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30526 27400 30556 27430 ne
rect 30556 27400 30770 27430
tri 30770 27400 30800 27430 sw
tri 30556 27354 30602 27400 ne
rect 30602 27354 30678 27400
rect 30724 27372 30800 27400
tri 30800 27372 30828 27400 sw
rect 70813 27372 71000 27430
rect 30724 27354 30828 27372
tri 30828 27354 30846 27372 sw
tri 30602 27326 30630 27354 ne
rect 30630 27326 30846 27354
tri 30846 27326 30874 27354 sw
rect 70813 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
tri 30630 27268 30688 27326 ne
rect 30688 27268 30874 27326
tri 30874 27268 30932 27326 sw
rect 70813 27268 71000 27326
tri 30688 27260 30696 27268 ne
rect 30696 27260 30810 27268
tri 30696 27222 30734 27260 ne
rect 30734 27222 30810 27260
rect 30856 27260 30932 27268
tri 30932 27260 30940 27268 sw
rect 30856 27222 30940 27260
tri 30940 27222 30978 27260 sw
rect 70813 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30734 27164 30792 27222 ne
rect 30792 27164 30978 27222
tri 30978 27164 31036 27222 sw
rect 70813 27164 71000 27222
tri 30792 27136 30820 27164 ne
rect 30820 27136 31036 27164
tri 31036 27136 31064 27164 sw
tri 30820 27090 30866 27136 ne
rect 30866 27090 30942 27136
rect 30988 27118 31064 27136
tri 31064 27118 31082 27136 sw
rect 70813 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 30988 27090 31082 27118
tri 31082 27090 31110 27118 sw
tri 30866 27060 30896 27090 ne
rect 30896 27060 31110 27090
tri 31110 27060 31140 27090 sw
rect 70813 27060 71000 27118
tri 30896 27016 30940 27060 ne
rect 30940 27016 31140 27060
tri 31140 27016 31184 27060 sw
tri 30940 27014 30942 27016 ne
rect 30942 27014 31184 27016
tri 31184 27014 31186 27016 sw
rect 70813 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
tri 30942 27004 30952 27014 ne
rect 30952 27004 31186 27014
tri 30952 26958 30998 27004 ne
rect 30998 26958 31074 27004
rect 31120 26958 31186 27004
tri 30998 26956 31000 26958 ne
rect 31000 26956 31186 26958
tri 31186 26956 31244 27014 sw
rect 70813 26956 71000 27014
tri 31000 26910 31046 26956 ne
rect 31046 26910 31244 26956
tri 31244 26910 31290 26956 sw
rect 70813 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31046 26872 31084 26910 ne
rect 31084 26872 31290 26910
tri 31290 26872 31328 26910 sw
tri 31084 26826 31130 26872 ne
rect 31130 26826 31206 26872
rect 31252 26852 31328 26872
tri 31328 26852 31348 26872 sw
rect 70813 26852 71000 26910
rect 31252 26826 31348 26852
tri 31348 26826 31374 26852 sw
tri 31130 26806 31150 26826 ne
rect 31150 26806 31374 26826
tri 31374 26806 31394 26826 sw
rect 70813 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
tri 31150 26772 31184 26806 ne
rect 31184 26772 31394 26806
tri 31394 26772 31428 26806 sw
tri 31184 26748 31208 26772 ne
rect 31208 26748 31428 26772
tri 31428 26748 31452 26772 sw
rect 70813 26748 71000 26806
tri 31208 26740 31216 26748 ne
rect 31216 26740 31452 26748
tri 31216 26694 31262 26740 ne
rect 31262 26694 31338 26740
rect 31384 26702 31452 26740
tri 31452 26702 31498 26748 sw
rect 70813 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 31384 26694 31498 26702
tri 31262 26644 31312 26694 ne
rect 31312 26644 31498 26694
tri 31498 26644 31556 26702 sw
rect 70813 26644 71000 26702
tri 31312 26608 31348 26644 ne
rect 31348 26608 31556 26644
tri 31556 26608 31592 26644 sw
tri 31348 26562 31394 26608 ne
rect 31394 26562 31470 26608
rect 31516 26598 31592 26608
tri 31592 26598 31602 26608 sw
rect 70813 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 31516 26562 31602 26598
tri 31602 26562 31638 26598 sw
tri 31394 26540 31416 26562 ne
rect 31416 26540 31638 26562
tri 31638 26540 31660 26562 sw
rect 70813 26540 71000 26598
tri 31416 26528 31428 26540 ne
rect 31428 26528 31660 26540
tri 31660 26528 31672 26540 sw
tri 31428 26494 31462 26528 ne
rect 31462 26494 31672 26528
tri 31672 26494 31706 26528 sw
rect 70813 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
tri 31462 26476 31480 26494 ne
rect 31480 26476 31706 26494
tri 31480 26430 31526 26476 ne
rect 31526 26430 31602 26476
rect 31648 26436 31706 26476
tri 31706 26436 31764 26494 sw
rect 70813 26436 71000 26494
rect 31648 26430 31764 26436
tri 31526 26390 31566 26430 ne
rect 31566 26390 31764 26430
tri 31764 26390 31810 26436 sw
rect 70813 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31566 26344 31612 26390 ne
rect 31612 26344 31810 26390
tri 31810 26344 31856 26390 sw
tri 31612 26298 31658 26344 ne
rect 31658 26298 31734 26344
rect 31780 26332 31856 26344
tri 31856 26332 31868 26344 sw
rect 70813 26332 71000 26390
rect 31780 26298 31868 26332
tri 31868 26298 31902 26332 sw
tri 31658 26286 31670 26298 ne
rect 31670 26286 31902 26298
tri 31902 26286 31914 26298 sw
rect 70813 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31670 26284 31672 26286 ne
rect 31672 26284 31914 26286
tri 31914 26284 31916 26286 sw
tri 31672 26228 31728 26284 ne
rect 31728 26228 31916 26284
tri 31916 26228 31972 26284 sw
rect 70813 26228 71000 26286
tri 31728 26212 31744 26228 ne
rect 31744 26212 31972 26228
tri 31744 26166 31790 26212 ne
rect 31790 26166 31866 26212
rect 31912 26182 31972 26212
tri 31972 26182 32018 26228 sw
rect 70813 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 31912 26166 32018 26182
tri 31790 26124 31832 26166 ne
rect 31832 26124 32018 26166
tri 32018 26124 32076 26182 sw
rect 70813 26124 71000 26182
tri 31832 26080 31876 26124 ne
rect 31876 26080 32076 26124
tri 32076 26080 32120 26124 sw
tri 31876 26040 31916 26080 ne
rect 31916 26040 31998 26080
tri 31916 26034 31922 26040 ne
rect 31922 26034 31998 26040
rect 32044 26078 32120 26080
tri 32120 26078 32122 26080 sw
rect 70813 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26040 32122 26078
tri 32122 26040 32160 26078 sw
rect 32044 26034 32160 26040
tri 31922 26020 31936 26034 ne
rect 31936 26020 32160 26034
tri 32160 26020 32180 26040 sw
rect 70813 26020 71000 26078
tri 31936 25974 31982 26020 ne
rect 31982 25974 32180 26020
tri 32180 25974 32226 26020 sw
rect 70813 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
tri 31982 25948 32008 25974 ne
rect 32008 25948 32226 25974
tri 32226 25948 32252 25974 sw
tri 32008 25902 32054 25948 ne
rect 32054 25902 32130 25948
rect 32176 25916 32252 25948
tri 32252 25916 32284 25948 sw
rect 70813 25916 71000 25974
rect 32176 25902 32284 25916
tri 32284 25902 32298 25916 sw
tri 32054 25870 32086 25902 ne
rect 32086 25870 32298 25902
tri 32298 25870 32330 25902 sw
rect 70813 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32086 25816 32140 25870 ne
rect 32140 25816 32330 25870
tri 32330 25816 32384 25870 sw
tri 32140 25796 32160 25816 ne
rect 32160 25796 32262 25816
tri 32160 25770 32186 25796 ne
rect 32186 25770 32262 25796
rect 32308 25812 32384 25816
tri 32384 25812 32388 25816 sw
rect 70813 25812 71000 25870
rect 32308 25796 32388 25812
tri 32388 25796 32404 25812 sw
rect 32308 25770 32404 25796
tri 32186 25766 32190 25770 ne
rect 32190 25766 32404 25770
tri 32404 25766 32434 25796 sw
rect 70813 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
tri 32190 25708 32248 25766 ne
rect 32248 25708 32434 25766
tri 32434 25708 32492 25766 sw
rect 70813 25708 71000 25766
tri 32248 25684 32272 25708 ne
rect 32272 25684 32492 25708
tri 32492 25684 32516 25708 sw
tri 32272 25638 32318 25684 ne
rect 32318 25638 32394 25684
rect 32440 25662 32516 25684
tri 32516 25662 32538 25684 sw
rect 70813 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25638 32538 25662
tri 32538 25638 32562 25662 sw
tri 32318 25604 32352 25638 ne
rect 32352 25604 32562 25638
tri 32562 25604 32596 25638 sw
rect 70813 25604 71000 25662
tri 32352 25558 32398 25604 ne
rect 32398 25558 32596 25604
tri 32596 25558 32642 25604 sw
rect 70813 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
tri 32398 25552 32404 25558 ne
rect 32404 25552 32642 25558
tri 32642 25552 32648 25558 sw
tri 32404 25506 32450 25552 ne
rect 32450 25506 32526 25552
rect 32572 25506 32648 25552
tri 32450 25500 32456 25506 ne
rect 32456 25500 32648 25506
tri 32648 25500 32700 25552 sw
rect 70813 25500 71000 25558
tri 32456 25454 32502 25500 ne
rect 32502 25454 32700 25500
tri 32700 25454 32746 25500 sw
rect 70813 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
tri 32502 25420 32536 25454 ne
rect 32536 25420 32746 25454
tri 32746 25420 32780 25454 sw
tri 32536 25374 32582 25420 ne
rect 32582 25374 32658 25420
rect 32704 25396 32780 25420
tri 32780 25396 32804 25420 sw
rect 70813 25396 71000 25454
rect 32704 25374 32804 25396
tri 32804 25374 32826 25396 sw
tri 32582 25350 32606 25374 ne
rect 32606 25350 32826 25374
tri 32826 25350 32850 25374 sw
rect 70813 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
tri 32606 25308 32648 25350 ne
rect 32648 25308 32850 25350
tri 32850 25308 32892 25350 sw
tri 32648 25292 32664 25308 ne
rect 32664 25292 32892 25308
tri 32892 25292 32908 25308 sw
rect 70813 25292 71000 25350
tri 32664 25288 32668 25292 ne
rect 32668 25288 32908 25292
tri 32668 25242 32714 25288 ne
rect 32714 25242 32790 25288
rect 32836 25246 32908 25288
tri 32908 25246 32954 25292 sw
rect 70813 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 32836 25242 32954 25246
tri 32714 25188 32768 25242 ne
rect 32768 25188 32954 25242
tri 32954 25188 33012 25246 sw
rect 70813 25188 71000 25246
tri 32768 25156 32800 25188 ne
rect 32800 25156 33012 25188
tri 33012 25156 33044 25188 sw
tri 32800 25110 32846 25156 ne
rect 32846 25110 32922 25156
rect 32968 25142 33044 25156
tri 33044 25142 33058 25156 sw
rect 70813 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 32968 25110 33058 25142
tri 33058 25110 33090 25142 sw
tri 32846 25084 32872 25110 ne
rect 32872 25084 33090 25110
tri 33090 25084 33116 25110 sw
rect 70813 25084 71000 25142
tri 32872 25064 32892 25084 ne
rect 32892 25064 33116 25084
tri 33116 25064 33136 25084 sw
tri 32892 25038 32918 25064 ne
rect 32918 25038 33136 25064
tri 33136 25038 33162 25064 sw
rect 70813 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
tri 32918 25024 32932 25038 ne
rect 32932 25024 33162 25038
tri 32932 24978 32978 25024 ne
rect 32978 24978 33054 25024
rect 33100 24980 33162 25024
tri 33162 24980 33220 25038 sw
rect 70813 24980 71000 25038
rect 33100 24978 33220 24980
tri 32978 24934 33022 24978 ne
rect 33022 24934 33220 24978
tri 33220 24934 33266 24980 sw
rect 70813 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33022 24892 33064 24934 ne
rect 33064 24892 33266 24934
tri 33266 24892 33308 24934 sw
tri 33064 24846 33110 24892 ne
rect 33110 24846 33186 24892
rect 33232 24876 33308 24892
tri 33308 24876 33324 24892 sw
rect 70813 24876 71000 24934
rect 33232 24846 33324 24876
tri 33324 24846 33354 24876 sw
tri 33110 24830 33126 24846 ne
rect 33126 24830 33354 24846
tri 33354 24830 33370 24846 sw
rect 70813 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
tri 33126 24820 33136 24830 ne
rect 33136 24820 33370 24830
tri 33370 24820 33380 24830 sw
tri 33136 24772 33184 24820 ne
rect 33184 24772 33380 24820
tri 33380 24772 33428 24820 sw
rect 70813 24772 71000 24830
tri 33184 24760 33196 24772 ne
rect 33196 24760 33428 24772
tri 33196 24714 33242 24760 ne
rect 33242 24714 33318 24760
rect 33364 24726 33428 24760
tri 33428 24726 33474 24772 sw
rect 70813 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 33364 24714 33474 24726
tri 33242 24668 33288 24714 ne
rect 33288 24668 33474 24714
tri 33474 24668 33532 24726 sw
rect 70813 24668 71000 24726
tri 33288 24628 33328 24668 ne
rect 33328 24628 33532 24668
tri 33532 24628 33572 24668 sw
tri 33328 24582 33374 24628 ne
rect 33374 24582 33450 24628
rect 33496 24622 33572 24628
tri 33572 24622 33578 24628 sw
rect 70813 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24582 33578 24622
tri 33578 24582 33618 24622 sw
tri 33374 24576 33380 24582 ne
rect 33380 24576 33618 24582
tri 33618 24576 33624 24582 sw
tri 33380 24564 33392 24576 ne
rect 33392 24564 33624 24576
tri 33624 24564 33636 24576 sw
rect 70813 24564 71000 24622
tri 33392 24518 33438 24564 ne
rect 33438 24518 33636 24564
tri 33636 24518 33682 24564 sw
rect 70813 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33438 24496 33460 24518 ne
rect 33460 24496 33682 24518
tri 33682 24496 33704 24518 sw
tri 33460 24450 33506 24496 ne
rect 33506 24450 33582 24496
rect 33628 24460 33704 24496
tri 33704 24460 33740 24496 sw
rect 70813 24460 71000 24518
rect 33628 24450 33740 24460
tri 33740 24450 33750 24460 sw
tri 33506 24414 33542 24450 ne
rect 33542 24414 33750 24450
tri 33750 24414 33786 24450 sw
rect 70813 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33542 24364 33592 24414 ne
rect 33592 24364 33786 24414
tri 33786 24364 33836 24414 sw
tri 33592 24332 33624 24364 ne
rect 33624 24332 33714 24364
tri 33624 24318 33638 24332 ne
rect 33638 24318 33714 24332
rect 33760 24356 33836 24364
tri 33836 24356 33844 24364 sw
rect 70813 24356 71000 24414
rect 33760 24332 33844 24356
tri 33844 24332 33868 24356 sw
rect 33760 24318 33868 24332
tri 33638 24310 33646 24318 ne
rect 33646 24310 33868 24318
tri 33868 24310 33890 24332 sw
rect 70813 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
tri 33646 24252 33704 24310 ne
rect 33704 24252 33890 24310
tri 33890 24252 33948 24310 sw
rect 70813 24252 71000 24310
tri 33704 24232 33724 24252 ne
rect 33724 24232 33948 24252
tri 33948 24232 33968 24252 sw
tri 33724 24186 33770 24232 ne
rect 33770 24186 33846 24232
rect 33892 24206 33968 24232
tri 33968 24206 33994 24232 sw
rect 70813 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 33892 24186 33994 24206
tri 33994 24186 34014 24206 sw
tri 33770 24148 33808 24186 ne
rect 33808 24148 34014 24186
tri 34014 24148 34052 24186 sw
rect 70813 24148 71000 24206
tri 33808 24102 33854 24148 ne
rect 33854 24102 34052 24148
tri 34052 24102 34098 24148 sw
rect 70813 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
tri 33854 24100 33856 24102 ne
rect 33856 24100 34098 24102
tri 34098 24100 34100 24102 sw
tri 33856 24088 33868 24100 ne
rect 33868 24088 33978 24100
tri 33868 24054 33902 24088 ne
rect 33902 24054 33978 24088
rect 34024 24088 34100 24100
tri 34100 24088 34112 24100 sw
rect 34024 24054 34112 24088
tri 33902 24044 33912 24054 ne
rect 33912 24044 34112 24054
tri 34112 24044 34156 24088 sw
rect 70813 24044 71000 24102
tri 33912 23998 33958 24044 ne
rect 33958 23998 34156 24044
tri 34156 23998 34202 24044 sw
rect 70813 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33958 23968 33988 23998 ne
rect 33988 23968 34202 23998
tri 34202 23968 34232 23998 sw
tri 33988 23922 34034 23968 ne
rect 34034 23922 34110 23968
rect 34156 23940 34232 23968
tri 34232 23940 34260 23968 sw
rect 70813 23940 71000 23998
rect 34156 23922 34260 23940
tri 34260 23922 34278 23940 sw
tri 34034 23894 34062 23922 ne
rect 34062 23894 34278 23922
tri 34278 23894 34306 23922 sw
rect 70813 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34062 23844 34112 23894 ne
rect 34112 23844 34306 23894
tri 34306 23844 34356 23894 sw
tri 34112 23836 34120 23844 ne
rect 34120 23836 34356 23844
tri 34356 23836 34364 23844 sw
rect 70813 23836 71000 23894
tri 34120 23790 34166 23836 ne
rect 34166 23790 34242 23836
rect 34288 23790 34364 23836
tri 34364 23790 34410 23836 sw
rect 70813 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
tri 34166 23732 34224 23790 ne
rect 34224 23732 34410 23790
tri 34410 23732 34468 23790 sw
rect 70813 23732 71000 23790
tri 34224 23704 34252 23732 ne
rect 34252 23704 34468 23732
tri 34468 23704 34496 23732 sw
tri 34252 23658 34298 23704 ne
rect 34298 23658 34374 23704
rect 34420 23686 34496 23704
tri 34496 23686 34514 23704 sw
rect 70813 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23658 34514 23686
tri 34514 23658 34542 23686 sw
tri 34298 23628 34328 23658 ne
rect 34328 23628 34542 23658
tri 34542 23628 34572 23658 sw
rect 70813 23628 71000 23686
tri 34328 23600 34356 23628 ne
rect 34356 23600 34572 23628
tri 34572 23600 34600 23628 sw
tri 34356 23582 34374 23600 ne
rect 34374 23582 34600 23600
tri 34600 23582 34618 23600 sw
rect 70813 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
tri 34374 23572 34384 23582 ne
rect 34384 23572 34618 23582
tri 34384 23526 34430 23572 ne
rect 34430 23526 34506 23572
rect 34552 23526 34618 23572
tri 34430 23524 34432 23526 ne
rect 34432 23524 34618 23526
tri 34618 23524 34676 23582 sw
rect 70813 23524 71000 23582
tri 34432 23478 34478 23524 ne
rect 34478 23478 34676 23524
tri 34676 23478 34722 23524 sw
rect 70813 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
tri 34478 23440 34516 23478 ne
rect 34516 23440 34722 23478
tri 34722 23440 34760 23478 sw
tri 34516 23394 34562 23440 ne
rect 34562 23394 34638 23440
rect 34684 23420 34760 23440
tri 34760 23420 34780 23440 sw
rect 70813 23420 71000 23478
rect 34684 23394 34780 23420
tri 34780 23394 34806 23420 sw
tri 34562 23374 34582 23394 ne
rect 34582 23374 34806 23394
tri 34806 23374 34826 23394 sw
rect 70813 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34582 23356 34600 23374 ne
rect 34600 23356 34826 23374
tri 34826 23356 34844 23374 sw
tri 34600 23316 34640 23356 ne
rect 34640 23316 34844 23356
tri 34844 23316 34884 23356 sw
rect 70813 23316 71000 23374
tri 34640 23308 34648 23316 ne
rect 34648 23308 34884 23316
tri 34648 23262 34694 23308 ne
rect 34694 23262 34770 23308
rect 34816 23270 34884 23308
tri 34884 23270 34930 23316 sw
rect 70813 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 34816 23262 34930 23270
tri 34694 23212 34744 23262 ne
rect 34744 23212 34930 23262
tri 34930 23212 34988 23270 sw
rect 70813 23212 71000 23270
tri 34744 23176 34780 23212 ne
rect 34780 23176 34988 23212
tri 34988 23176 35024 23212 sw
tri 34780 23130 34826 23176 ne
rect 34826 23130 34902 23176
rect 34948 23166 35024 23176
tri 35024 23166 35034 23176 sw
rect 70813 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 34948 23130 35034 23166
tri 35034 23130 35070 23166 sw
tri 34826 23112 34844 23130 ne
rect 34844 23112 35070 23130
tri 35070 23112 35088 23130 sw
tri 34844 23108 34848 23112 ne
rect 34848 23108 35088 23112
tri 35088 23108 35092 23112 sw
rect 70813 23108 71000 23166
tri 34848 23062 34894 23108 ne
rect 34894 23062 35092 23108
tri 35092 23062 35138 23108 sw
rect 70813 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
tri 34894 23044 34912 23062 ne
rect 34912 23044 35138 23062
tri 34912 22998 34958 23044 ne
rect 34958 22998 35034 23044
rect 35080 23004 35138 23044
tri 35138 23004 35196 23062 sw
rect 70813 23004 71000 23062
rect 35080 22998 35196 23004
tri 34958 22958 34998 22998 ne
rect 34998 22958 35196 22998
tri 35196 22958 35242 23004 sw
rect 70813 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 34998 22912 35044 22958 ne
rect 35044 22912 35242 22958
tri 35242 22912 35288 22958 sw
tri 35044 22868 35088 22912 ne
rect 35088 22868 35166 22912
tri 35088 22866 35090 22868 ne
rect 35090 22866 35166 22868
rect 35212 22900 35288 22912
tri 35288 22900 35300 22912 sw
rect 70813 22900 71000 22958
rect 35212 22868 35300 22900
tri 35300 22868 35332 22900 sw
rect 35212 22866 35332 22868
tri 35090 22854 35102 22866 ne
rect 35102 22854 35332 22866
tri 35332 22854 35346 22868 sw
rect 70813 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
tri 35102 22796 35160 22854 ne
rect 35160 22796 35346 22854
tri 35346 22796 35404 22854 sw
rect 70813 22796 71000 22854
tri 35160 22780 35176 22796 ne
rect 35176 22780 35404 22796
tri 35404 22780 35420 22796 sw
tri 35176 22734 35222 22780 ne
rect 35222 22734 35298 22780
rect 35344 22750 35420 22780
tri 35420 22750 35450 22780 sw
rect 70813 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 35344 22734 35450 22750
tri 35450 22734 35466 22750 sw
tri 35222 22692 35264 22734 ne
rect 35264 22692 35466 22734
tri 35466 22692 35508 22734 sw
rect 70813 22692 71000 22750
tri 35264 22648 35308 22692 ne
rect 35308 22648 35508 22692
tri 35508 22648 35552 22692 sw
tri 35308 22624 35332 22648 ne
rect 35332 22624 35430 22648
tri 35332 22602 35354 22624 ne
rect 35354 22602 35430 22624
rect 35476 22646 35552 22648
tri 35552 22646 35554 22648 sw
rect 70813 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22624 35554 22646
tri 35554 22624 35576 22646 sw
rect 35476 22602 35576 22624
tri 35354 22588 35368 22602 ne
rect 35368 22588 35576 22602
tri 35576 22588 35612 22624 sw
rect 70813 22588 71000 22646
tri 35368 22542 35414 22588 ne
rect 35414 22542 35612 22588
tri 35612 22542 35658 22588 sw
rect 70813 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35414 22516 35440 22542 ne
rect 35440 22516 35658 22542
tri 35658 22516 35684 22542 sw
tri 35440 22470 35486 22516 ne
rect 35486 22470 35562 22516
rect 35608 22484 35684 22516
tri 35684 22484 35716 22516 sw
rect 70813 22484 71000 22542
rect 35608 22470 35716 22484
tri 35716 22470 35730 22484 sw
tri 35486 22438 35518 22470 ne
rect 35518 22438 35730 22470
tri 35730 22438 35762 22470 sw
rect 70813 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35518 22384 35572 22438 ne
rect 35572 22384 35762 22438
tri 35762 22384 35816 22438 sw
tri 35572 22380 35576 22384 ne
rect 35576 22380 35694 22384
tri 35576 22338 35618 22380 ne
rect 35618 22338 35694 22380
rect 35740 22380 35816 22384
tri 35816 22380 35820 22384 sw
rect 70813 22380 71000 22438
rect 35740 22338 35820 22380
tri 35618 22334 35622 22338 ne
rect 35622 22334 35820 22338
tri 35820 22334 35866 22380 sw
rect 70813 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35622 22276 35680 22334 ne
rect 35680 22276 35866 22334
tri 35866 22276 35924 22334 sw
rect 70813 22276 71000 22334
tri 35680 22252 35704 22276 ne
rect 35704 22252 35924 22276
tri 35924 22252 35948 22276 sw
tri 35704 22206 35750 22252 ne
rect 35750 22206 35826 22252
rect 35872 22230 35948 22252
tri 35948 22230 35970 22252 sw
rect 70813 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22206 35970 22230
tri 35970 22206 35994 22230 sw
tri 35750 22172 35784 22206 ne
rect 35784 22172 35994 22206
tri 35994 22172 36028 22206 sw
rect 70813 22172 71000 22230
tri 35784 22136 35820 22172 ne
rect 35820 22136 36028 22172
tri 36028 22136 36064 22172 sw
tri 35820 22126 35830 22136 ne
rect 35830 22126 36064 22136
tri 36064 22126 36074 22136 sw
rect 70813 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
tri 35830 22120 35836 22126 ne
rect 35836 22120 36074 22126
tri 35836 22074 35882 22120 ne
rect 35882 22074 35958 22120
rect 36004 22074 36074 22120
tri 35882 22068 35888 22074 ne
rect 35888 22068 36074 22074
tri 36074 22068 36132 22126 sw
rect 70813 22068 71000 22126
tri 35888 22022 35934 22068 ne
rect 35934 22022 36132 22068
tri 36132 22022 36178 22068 sw
rect 70813 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35934 21988 35968 22022 ne
rect 35968 21988 36178 22022
tri 36178 21988 36212 22022 sw
tri 35968 21942 36014 21988 ne
rect 36014 21942 36090 21988
rect 36136 21964 36212 21988
tri 36212 21964 36236 21988 sw
rect 70813 21964 71000 22022
rect 36136 21942 36236 21964
tri 36236 21942 36258 21964 sw
tri 36014 21918 36038 21942 ne
rect 36038 21918 36258 21942
tri 36258 21918 36282 21942 sw
rect 70813 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
tri 36038 21892 36064 21918 ne
rect 36064 21892 36282 21918
tri 36282 21892 36308 21918 sw
tri 36064 21860 36096 21892 ne
rect 36096 21860 36308 21892
tri 36308 21860 36340 21892 sw
rect 70813 21860 71000 21918
tri 36096 21856 36100 21860 ne
rect 36100 21856 36340 21860
tri 36100 21810 36146 21856 ne
rect 36146 21810 36222 21856
rect 36268 21814 36340 21856
tri 36340 21814 36386 21860 sw
rect 70813 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 36268 21810 36386 21814
tri 36146 21756 36200 21810 ne
rect 36200 21756 36386 21810
tri 36386 21756 36444 21814 sw
rect 70813 21756 71000 21814
tri 36200 21724 36232 21756 ne
rect 36232 21724 36444 21756
tri 36444 21724 36476 21756 sw
tri 36232 21678 36278 21724 ne
rect 36278 21678 36354 21724
rect 36400 21710 36476 21724
tri 36476 21710 36490 21724 sw
rect 70813 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 36400 21678 36490 21710
tri 36490 21678 36522 21710 sw
tri 36278 21652 36304 21678 ne
rect 36304 21652 36522 21678
tri 36522 21652 36548 21678 sw
rect 70813 21652 71000 21710
tri 36304 21648 36308 21652 ne
rect 36308 21648 36548 21652
tri 36548 21648 36552 21652 sw
tri 36308 21606 36350 21648 ne
rect 36350 21606 36552 21648
tri 36552 21606 36594 21648 sw
rect 70813 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
tri 36350 21592 36364 21606 ne
rect 36364 21592 36594 21606
tri 36364 21546 36410 21592 ne
rect 36410 21546 36486 21592
rect 36532 21548 36594 21592
tri 36594 21548 36652 21606 sw
rect 70813 21548 71000 21606
rect 36532 21546 36652 21548
tri 36410 21502 36454 21546 ne
rect 36454 21502 36652 21546
tri 36652 21502 36698 21548 sw
rect 70813 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36454 21460 36496 21502 ne
rect 36496 21460 36698 21502
tri 36698 21460 36740 21502 sw
tri 36496 21414 36542 21460 ne
rect 36542 21414 36618 21460
rect 36664 21444 36740 21460
tri 36740 21444 36756 21460 sw
rect 70813 21444 71000 21502
rect 36664 21414 36756 21444
tri 36756 21414 36786 21444 sw
tri 36542 21404 36552 21414 ne
rect 36552 21404 36786 21414
tri 36786 21404 36796 21414 sw
tri 36552 21398 36558 21404 ne
rect 36558 21398 36796 21404
tri 36796 21398 36802 21404 sw
rect 70813 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36558 21340 36616 21398 ne
rect 36616 21340 36802 21398
tri 36802 21340 36860 21398 sw
rect 70813 21340 71000 21398
tri 36616 21328 36628 21340 ne
rect 36628 21328 36860 21340
tri 36628 21282 36674 21328 ne
rect 36674 21282 36750 21328
rect 36796 21294 36860 21328
tri 36860 21294 36906 21340 sw
rect 70813 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36796 21282 36906 21294
tri 36674 21236 36720 21282 ne
rect 36720 21236 36906 21282
tri 36906 21236 36964 21294 sw
rect 70813 21236 71000 21294
tri 36720 21196 36760 21236 ne
rect 36760 21196 36964 21236
tri 36964 21196 37004 21236 sw
tri 36760 21160 36796 21196 ne
rect 36796 21160 36882 21196
tri 36796 21150 36806 21160 ne
rect 36806 21150 36882 21160
rect 36928 21190 37004 21196
tri 37004 21190 37010 21196 sw
rect 70813 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21160 37010 21190
tri 37010 21160 37040 21190 sw
rect 36928 21150 37040 21160
tri 36806 21132 36824 21150 ne
rect 36824 21132 37040 21150
tri 37040 21132 37068 21160 sw
rect 70813 21132 71000 21190
tri 36824 21086 36870 21132 ne
rect 36870 21086 37068 21132
tri 37068 21086 37114 21132 sw
rect 70813 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
tri 36870 21064 36892 21086 ne
rect 36892 21064 37114 21086
tri 37114 21064 37136 21086 sw
tri 36892 21018 36938 21064 ne
rect 36938 21018 37014 21064
rect 37060 21028 37136 21064
tri 37136 21028 37172 21064 sw
rect 70813 21028 71000 21086
rect 37060 21018 37172 21028
tri 37172 21018 37182 21028 sw
tri 36938 20982 36974 21018 ne
rect 36974 20982 37182 21018
tri 37182 20982 37218 21018 sw
rect 70813 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 36974 20932 37024 20982 ne
rect 37024 20932 37218 20982
tri 37218 20932 37268 20982 sw
tri 37024 20916 37040 20932 ne
rect 37040 20916 37146 20932
tri 37040 20886 37070 20916 ne
rect 37070 20886 37146 20916
rect 37192 20924 37268 20932
tri 37268 20924 37276 20932 sw
rect 70813 20924 71000 20982
rect 37192 20916 37276 20924
tri 37276 20916 37284 20924 sw
rect 37192 20886 37284 20916
tri 37070 20878 37078 20886 ne
rect 37078 20878 37284 20886
tri 37284 20878 37322 20916 sw
rect 70813 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
tri 37078 20820 37136 20878 ne
rect 37136 20820 37322 20878
tri 37322 20820 37380 20878 sw
rect 70813 20820 71000 20878
tri 37136 20800 37156 20820 ne
rect 37156 20800 37380 20820
tri 37380 20800 37400 20820 sw
tri 37156 20754 37202 20800 ne
rect 37202 20754 37278 20800
rect 37324 20774 37400 20800
tri 37400 20774 37426 20800 sw
rect 70813 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 37324 20754 37426 20774
tri 37426 20754 37446 20774 sw
tri 37202 20716 37240 20754 ne
rect 37240 20716 37446 20754
tri 37446 20716 37484 20754 sw
rect 70813 20716 71000 20774
tri 37240 20672 37284 20716 ne
rect 37284 20672 37484 20716
tri 37484 20672 37528 20716 sw
tri 37284 20670 37286 20672 ne
rect 37286 20670 37528 20672
tri 37528 20670 37530 20672 sw
rect 70813 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
tri 37286 20668 37288 20670 ne
rect 37288 20668 37530 20670
tri 37288 20622 37334 20668 ne
rect 37334 20622 37410 20668
rect 37456 20622 37530 20668
tri 37334 20612 37344 20622 ne
rect 37344 20612 37530 20622
tri 37530 20612 37588 20670 sw
rect 70813 20612 71000 20670
tri 37344 20566 37390 20612 ne
rect 37390 20566 37588 20612
tri 37588 20566 37634 20612 sw
rect 70813 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
tri 37390 20536 37420 20566 ne
rect 37420 20536 37634 20566
tri 37634 20536 37664 20566 sw
tri 37420 20490 37466 20536 ne
rect 37466 20490 37542 20536
rect 37588 20508 37664 20536
tri 37664 20508 37692 20536 sw
rect 70813 20508 71000 20566
rect 37588 20490 37692 20508
tri 37692 20490 37710 20508 sw
tri 37466 20462 37494 20490 ne
rect 37494 20462 37710 20490
tri 37710 20462 37738 20490 sw
rect 70813 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
tri 37494 20428 37528 20462 ne
rect 37528 20428 37738 20462
tri 37738 20428 37772 20462 sw
tri 37528 20404 37552 20428 ne
rect 37552 20404 37772 20428
tri 37772 20404 37796 20428 sw
rect 70813 20404 71000 20462
tri 37552 20358 37598 20404 ne
rect 37598 20358 37674 20404
rect 37720 20358 37796 20404
tri 37796 20358 37842 20404 sw
rect 70813 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37598 20300 37656 20358 ne
rect 37656 20300 37842 20358
tri 37842 20300 37900 20358 sw
rect 70813 20300 71000 20358
tri 37656 20272 37684 20300 ne
rect 37684 20272 37900 20300
tri 37900 20272 37928 20300 sw
tri 37684 20226 37730 20272 ne
rect 37730 20226 37806 20272
rect 37852 20254 37928 20272
tri 37928 20254 37946 20272 sw
rect 70813 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20226 37946 20254
tri 37946 20226 37974 20254 sw
tri 37730 20196 37760 20226 ne
rect 37760 20196 37974 20226
tri 37974 20196 38004 20226 sw
rect 70813 20196 71000 20254
tri 37760 20184 37772 20196 ne
rect 37772 20184 38004 20196
tri 38004 20184 38016 20196 sw
tri 37772 20150 37806 20184 ne
rect 37806 20150 38016 20184
tri 38016 20150 38050 20184 sw
rect 70813 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
tri 37806 20140 37816 20150 ne
rect 37816 20140 38050 20150
tri 37816 20094 37862 20140 ne
rect 37862 20094 37938 20140
rect 37984 20094 38050 20140
tri 37862 20092 37864 20094 ne
rect 37864 20092 38050 20094
tri 38050 20092 38108 20150 sw
rect 70813 20092 71000 20150
tri 37864 20046 37910 20092 ne
rect 37910 20046 38108 20092
tri 38108 20046 38154 20092 sw
rect 70813 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37910 20008 37948 20046 ne
rect 37948 20008 38154 20046
tri 38154 20008 38192 20046 sw
tri 37948 19962 37994 20008 ne
rect 37994 19962 38070 20008
rect 38116 19988 38192 20008
tri 38192 19988 38212 20008 sw
rect 70813 19988 71000 20046
rect 38116 19962 38212 19988
tri 38212 19962 38238 19988 sw
tri 37994 19942 38014 19962 ne
rect 38014 19942 38238 19962
tri 38238 19942 38258 19962 sw
rect 70813 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
tri 38014 19940 38016 19942 ne
rect 38016 19940 38258 19942
tri 38258 19940 38260 19942 sw
tri 38016 19884 38072 19940 ne
rect 38072 19884 38260 19940
tri 38260 19884 38316 19940 sw
rect 70813 19884 71000 19942
tri 38072 19876 38080 19884 ne
rect 38080 19876 38316 19884
tri 38080 19830 38126 19876 ne
rect 38126 19830 38202 19876
rect 38248 19838 38316 19876
tri 38316 19838 38362 19884 sw
rect 70813 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 38248 19830 38362 19838
tri 38126 19780 38176 19830 ne
rect 38176 19780 38362 19830
tri 38362 19780 38420 19838 sw
rect 70813 19780 71000 19838
tri 38176 19744 38212 19780 ne
rect 38212 19744 38420 19780
tri 38420 19744 38456 19780 sw
tri 38212 19698 38258 19744 ne
rect 38258 19698 38334 19744
rect 38380 19734 38456 19744
tri 38456 19734 38466 19744 sw
rect 70813 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 38380 19698 38466 19734
tri 38466 19698 38502 19734 sw
tri 38258 19696 38260 19698 ne
rect 38260 19696 38502 19698
tri 38502 19696 38504 19698 sw
tri 38260 19676 38280 19696 ne
rect 38280 19676 38504 19696
tri 38504 19676 38524 19696 sw
rect 70813 19676 71000 19734
tri 38280 19630 38326 19676 ne
rect 38326 19630 38524 19676
tri 38524 19630 38570 19676 sw
rect 70813 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
tri 38326 19612 38344 19630 ne
rect 38344 19612 38570 19630
tri 38570 19612 38588 19630 sw
tri 38344 19566 38390 19612 ne
rect 38390 19566 38466 19612
rect 38512 19572 38588 19612
tri 38588 19572 38628 19612 sw
rect 70813 19572 71000 19630
rect 38512 19566 38628 19572
tri 38628 19566 38634 19572 sw
tri 38390 19526 38430 19566 ne
rect 38430 19526 38634 19566
tri 38634 19526 38674 19566 sw
rect 70813 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38430 19480 38476 19526 ne
rect 38476 19480 38674 19526
tri 38674 19480 38720 19526 sw
tri 38476 19452 38504 19480 ne
rect 38504 19452 38598 19480
tri 38504 19434 38522 19452 ne
rect 38522 19434 38598 19452
rect 38644 19468 38720 19480
tri 38720 19468 38732 19480 sw
rect 70813 19468 71000 19526
rect 38644 19452 38732 19468
tri 38732 19452 38748 19468 sw
rect 38644 19434 38748 19452
tri 38522 19422 38534 19434 ne
rect 38534 19422 38748 19434
tri 38748 19422 38778 19452 sw
rect 70813 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
tri 38534 19364 38592 19422 ne
rect 38592 19364 38778 19422
tri 38778 19364 38836 19422 sw
rect 70813 19364 71000 19422
tri 38592 19348 38608 19364 ne
rect 38608 19348 38836 19364
tri 38836 19348 38852 19364 sw
tri 38608 19302 38654 19348 ne
rect 38654 19302 38730 19348
rect 38776 19318 38852 19348
tri 38852 19318 38882 19348 sw
rect 70813 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 38776 19302 38882 19318
tri 38882 19302 38898 19318 sw
tri 38654 19260 38696 19302 ne
rect 38696 19260 38898 19302
tri 38898 19260 38940 19302 sw
rect 70813 19260 71000 19318
tri 38696 19216 38740 19260 ne
rect 38740 19216 38940 19260
tri 38940 19216 38984 19260 sw
tri 38740 19208 38748 19216 ne
rect 38748 19208 38862 19216
tri 38748 19170 38786 19208 ne
rect 38786 19170 38862 19208
rect 38908 19214 38984 19216
tri 38984 19214 38986 19216 sw
rect 70813 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19208 38986 19214
tri 38986 19208 38992 19214 sw
rect 38908 19170 38992 19208
tri 38786 19156 38800 19170 ne
rect 38800 19156 38992 19170
tri 38992 19156 39044 19208 sw
rect 70813 19156 71000 19214
tri 38800 19110 38846 19156 ne
rect 38846 19110 39044 19156
tri 39044 19110 39090 19156 sw
rect 70813 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
tri 38846 19084 38872 19110 ne
rect 38872 19084 39090 19110
tri 39090 19084 39116 19110 sw
tri 38872 19038 38918 19084 ne
rect 38918 19038 38994 19084
rect 39040 19052 39116 19084
tri 39116 19052 39148 19084 sw
rect 70813 19052 71000 19110
rect 39040 19038 39148 19052
tri 39148 19038 39162 19052 sw
tri 38918 19006 38950 19038 ne
rect 38950 19006 39162 19038
tri 39162 19006 39194 19038 sw
rect 70813 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
tri 38950 18964 38992 19006 ne
rect 38992 18964 39194 19006
tri 39194 18964 39236 19006 sw
tri 38992 18952 39004 18964 ne
rect 39004 18952 39236 18964
tri 39004 18906 39050 18952 ne
rect 39050 18906 39126 18952
rect 39172 18948 39236 18952
tri 39236 18948 39252 18964 sw
rect 70813 18948 71000 19006
rect 39172 18906 39252 18948
tri 39050 18902 39054 18906 ne
rect 39054 18902 39252 18906
tri 39252 18902 39298 18948 sw
rect 70813 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
tri 39054 18844 39112 18902 ne
rect 39112 18844 39298 18902
tri 39298 18844 39356 18902 sw
rect 70813 18844 71000 18902
tri 39112 18820 39136 18844 ne
rect 39136 18820 39356 18844
tri 39356 18820 39380 18844 sw
tri 39136 18774 39182 18820 ne
rect 39182 18774 39258 18820
rect 39304 18798 39380 18820
tri 39380 18798 39402 18820 sw
rect 70813 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18774 39402 18798
tri 39402 18774 39426 18798 sw
tri 39182 18740 39216 18774 ne
rect 39216 18740 39426 18774
tri 39426 18740 39460 18774 sw
rect 70813 18740 71000 18798
tri 39216 18720 39236 18740 ne
rect 39236 18720 39460 18740
tri 39460 18720 39480 18740 sw
tri 39236 18694 39262 18720 ne
rect 39262 18694 39480 18720
tri 39480 18694 39506 18720 sw
rect 70813 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
tri 39262 18688 39268 18694 ne
rect 39268 18688 39506 18694
tri 39268 18642 39314 18688 ne
rect 39314 18642 39390 18688
rect 39436 18642 39506 18688
tri 39314 18636 39320 18642 ne
rect 39320 18636 39506 18642
tri 39506 18636 39564 18694 sw
rect 70813 18636 71000 18694
tri 39320 18590 39366 18636 ne
rect 39366 18590 39564 18636
tri 39564 18590 39610 18636 sw
rect 70813 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
tri 39366 18556 39400 18590 ne
rect 39400 18556 39610 18590
tri 39610 18556 39644 18590 sw
tri 39400 18510 39446 18556 ne
rect 39446 18510 39522 18556
rect 39568 18532 39644 18556
tri 39644 18532 39668 18556 sw
rect 70813 18532 71000 18590
rect 39568 18510 39668 18532
tri 39668 18510 39690 18532 sw
tri 39446 18486 39470 18510 ne
rect 39470 18486 39690 18510
tri 39690 18486 39714 18510 sw
rect 70813 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
tri 39470 18476 39480 18486 ne
rect 39480 18476 39714 18486
tri 39714 18476 39724 18486 sw
tri 39480 18428 39528 18476 ne
rect 39528 18428 39724 18476
tri 39724 18428 39772 18476 sw
rect 70813 18428 71000 18486
tri 39528 18424 39532 18428 ne
rect 39532 18424 39772 18428
tri 39532 18378 39578 18424 ne
rect 39578 18378 39654 18424
rect 39700 18382 39772 18424
tri 39772 18382 39818 18428 sw
rect 70813 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 39700 18378 39818 18382
tri 39578 18324 39632 18378 ne
rect 39632 18324 39818 18378
tri 39818 18324 39876 18382 sw
rect 70813 18324 71000 18382
tri 39632 18292 39664 18324 ne
rect 39664 18292 39876 18324
tri 39876 18292 39908 18324 sw
tri 39664 18246 39710 18292 ne
rect 39710 18246 39786 18292
rect 39832 18278 39908 18292
tri 39908 18278 39922 18292 sw
rect 70813 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 39832 18246 39922 18278
tri 39922 18246 39954 18278 sw
tri 39710 18232 39724 18246 ne
rect 39724 18232 39954 18246
tri 39954 18232 39968 18246 sw
tri 39724 18220 39736 18232 ne
rect 39736 18220 39968 18232
tri 39968 18220 39980 18232 sw
rect 70813 18220 71000 18278
tri 39736 18174 39782 18220 ne
rect 39782 18174 39980 18220
tri 39980 18174 40026 18220 sw
rect 70813 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
tri 39782 18160 39796 18174 ne
rect 39796 18160 40026 18174
tri 39796 18114 39842 18160 ne
rect 39842 18114 39918 18160
rect 39964 18116 40026 18160
tri 40026 18116 40084 18174 sw
rect 70813 18116 71000 18174
rect 39964 18114 40084 18116
tri 39842 18070 39886 18114 ne
rect 39886 18070 40084 18114
tri 40084 18070 40130 18116 sw
rect 70813 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39886 18028 39928 18070 ne
rect 39928 18028 40130 18070
tri 40130 18028 40172 18070 sw
tri 39928 17988 39968 18028 ne
rect 39968 17988 40050 18028
tri 39968 17982 39974 17988 ne
rect 39974 17982 40050 17988
rect 40096 18012 40172 18028
tri 40172 18012 40188 18028 sw
rect 70813 18012 71000 18070
rect 40096 17988 40188 18012
tri 40188 17988 40212 18012 sw
rect 40096 17982 40212 17988
tri 39974 17966 39990 17982 ne
rect 39990 17966 40212 17982
tri 40212 17966 40234 17988 sw
rect 70813 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
tri 39990 17908 40048 17966 ne
rect 40048 17908 40234 17966
tri 40234 17908 40292 17966 sw
rect 70813 17908 71000 17966
tri 40048 17896 40060 17908 ne
rect 40060 17896 40292 17908
tri 40292 17896 40304 17908 sw
tri 40060 17850 40106 17896 ne
rect 40106 17850 40182 17896
rect 40228 17862 40304 17896
tri 40304 17862 40338 17896 sw
rect 70813 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 40228 17850 40338 17862
tri 40338 17850 40350 17862 sw
tri 40106 17804 40152 17850 ne
rect 40152 17804 40350 17850
tri 40350 17804 40396 17850 sw
rect 70813 17804 71000 17862
tri 40152 17764 40192 17804 ne
rect 40192 17764 40396 17804
tri 40396 17764 40436 17804 sw
tri 40192 17744 40212 17764 ne
rect 40212 17744 40314 17764
tri 40212 17718 40238 17744 ne
rect 40238 17718 40314 17744
rect 40360 17758 40436 17764
tri 40436 17758 40442 17764 sw
rect 70813 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17744 40442 17758
tri 40442 17744 40456 17758 sw
rect 40360 17718 40456 17744
tri 40238 17700 40256 17718 ne
rect 40256 17700 40456 17718
tri 40456 17700 40500 17744 sw
rect 70813 17700 71000 17758
tri 40256 17654 40302 17700 ne
rect 40302 17654 40500 17700
tri 40500 17654 40546 17700 sw
rect 70813 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40302 17632 40324 17654 ne
rect 40324 17632 40546 17654
tri 40546 17632 40568 17654 sw
tri 40324 17586 40370 17632 ne
rect 40370 17586 40446 17632
rect 40492 17596 40568 17632
tri 40568 17596 40604 17632 sw
rect 70813 17596 71000 17654
rect 40492 17586 40604 17596
tri 40604 17586 40614 17596 sw
tri 40370 17550 40406 17586 ne
rect 40406 17550 40614 17586
tri 40614 17550 40650 17586 sw
rect 70813 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
tri 40406 17500 40456 17550 ne
rect 40456 17500 40650 17550
tri 40650 17500 40700 17550 sw
tri 40456 17454 40502 17500 ne
rect 40502 17454 40578 17500
rect 40624 17492 40700 17500
tri 40700 17492 40708 17500 sw
rect 70813 17492 71000 17550
rect 40624 17454 40708 17492
tri 40502 17446 40510 17454 ne
rect 40510 17446 40708 17454
tri 40708 17446 40754 17492 sw
rect 70813 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
tri 40510 17388 40568 17446 ne
rect 40568 17388 40754 17446
tri 40754 17388 40812 17446 sw
rect 70813 17388 71000 17446
tri 40568 17368 40588 17388 ne
rect 40588 17368 40812 17388
tri 40812 17368 40832 17388 sw
tri 40588 17322 40634 17368 ne
rect 40634 17322 40710 17368
rect 40756 17342 40832 17368
tri 40832 17342 40858 17368 sw
rect 70813 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17322 40858 17342
tri 40858 17322 40878 17342 sw
tri 40634 17284 40672 17322 ne
rect 40672 17284 40878 17322
tri 40878 17284 40916 17322 sw
rect 70813 17284 71000 17342
tri 40672 17256 40700 17284 ne
rect 40700 17256 40916 17284
tri 40916 17256 40944 17284 sw
tri 40700 17238 40718 17256 ne
rect 40718 17238 40944 17256
tri 40944 17238 40962 17256 sw
rect 70813 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
tri 40718 17236 40720 17238 ne
rect 40720 17236 40962 17238
tri 40720 17190 40766 17236 ne
rect 40766 17190 40842 17236
rect 40888 17190 40962 17236
tri 40766 17180 40776 17190 ne
rect 40776 17180 40962 17190
tri 40962 17180 41020 17238 sw
rect 70813 17180 71000 17238
tri 40776 17134 40822 17180 ne
rect 40822 17134 41020 17180
tri 41020 17134 41066 17180 sw
rect 70813 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40822 17104 40852 17134 ne
rect 40852 17104 41066 17134
tri 41066 17104 41096 17134 sw
tri 40852 17058 40898 17104 ne
rect 40898 17058 40974 17104
rect 41020 17076 41096 17104
tri 41096 17076 41124 17104 sw
rect 70813 17076 71000 17134
rect 41020 17058 41124 17076
tri 41124 17058 41142 17076 sw
tri 40898 17030 40926 17058 ne
rect 40926 17030 41142 17058
tri 41142 17030 41170 17058 sw
rect 70813 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
tri 40926 17012 40944 17030 ne
rect 40944 17012 41170 17030
tri 41170 17012 41188 17030 sw
tri 40944 16972 40984 17012 ne
rect 40984 16972 41188 17012
tri 41188 16972 41228 17012 sw
rect 70813 16972 71000 17030
tri 40984 16926 41030 16972 ne
rect 41030 16926 41106 16972
rect 41152 16926 41228 16972
tri 41228 16926 41274 16972 sw
rect 70813 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41030 16868 41088 16926 ne
rect 41088 16868 41274 16926
tri 41274 16868 41332 16926 sw
rect 70813 16868 71000 16926
tri 41088 16840 41116 16868 ne
rect 41116 16840 41332 16868
tri 41332 16840 41360 16868 sw
tri 41116 16794 41162 16840 ne
rect 41162 16794 41238 16840
rect 41284 16822 41360 16840
tri 41360 16822 41378 16840 sw
rect 70813 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16794 41378 16822
tri 41378 16794 41406 16822 sw
tri 41162 16768 41188 16794 ne
rect 41188 16768 41406 16794
tri 41406 16768 41432 16794 sw
tri 41188 16764 41192 16768 ne
rect 41192 16764 41432 16768
tri 41432 16764 41436 16768 sw
rect 70813 16764 71000 16822
tri 41192 16718 41238 16764 ne
rect 41238 16718 41436 16764
tri 41436 16718 41482 16764 sw
rect 70813 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
tri 41238 16708 41248 16718 ne
rect 41248 16708 41482 16718
tri 41248 16662 41294 16708 ne
rect 41294 16662 41370 16708
rect 41416 16662 41482 16708
tri 41294 16660 41296 16662 ne
rect 41296 16660 41482 16662
tri 41482 16660 41540 16718 sw
rect 70813 16660 71000 16718
tri 41296 16614 41342 16660 ne
rect 41342 16614 41540 16660
tri 41540 16614 41586 16660 sw
rect 70813 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
tri 41342 16576 41380 16614 ne
rect 41380 16576 41586 16614
tri 41586 16576 41624 16614 sw
tri 41380 16530 41426 16576 ne
rect 41426 16530 41502 16576
rect 41548 16556 41624 16576
tri 41624 16556 41644 16576 sw
rect 70813 16556 71000 16614
rect 41548 16530 41644 16556
tri 41644 16530 41670 16556 sw
tri 41426 16524 41432 16530 ne
rect 41432 16524 41670 16530
tri 41670 16524 41676 16530 sw
tri 41432 16510 41446 16524 ne
rect 41446 16510 41676 16524
tri 41676 16510 41690 16524 sw
rect 70813 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41446 16452 41504 16510 ne
rect 41504 16452 41690 16510
tri 41690 16452 41748 16510 sw
rect 70813 16452 71000 16510
tri 41504 16444 41512 16452 ne
rect 41512 16444 41748 16452
tri 41748 16444 41756 16452 sw
tri 41512 16398 41558 16444 ne
rect 41558 16398 41634 16444
rect 41680 16406 41756 16444
tri 41756 16406 41794 16444 sw
rect 70813 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 41680 16398 41794 16406
tri 41794 16398 41802 16406 sw
tri 41558 16348 41608 16398 ne
rect 41608 16348 41802 16398
tri 41802 16348 41852 16398 sw
rect 70813 16348 71000 16406
tri 41608 16312 41644 16348 ne
rect 41644 16312 41852 16348
tri 41852 16312 41888 16348 sw
tri 41644 16280 41676 16312 ne
rect 41676 16280 41766 16312
tri 41676 16266 41690 16280 ne
rect 41690 16266 41766 16280
rect 41812 16302 41888 16312
tri 41888 16302 41898 16312 sw
rect 70813 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16280 41898 16302
tri 41898 16280 41920 16302 sw
rect 41812 16266 41920 16280
tri 41690 16244 41712 16266 ne
rect 41712 16244 41920 16266
tri 41920 16244 41956 16280 sw
rect 70813 16244 71000 16302
tri 41712 16198 41758 16244 ne
rect 41758 16198 41956 16244
tri 41956 16198 42002 16244 sw
rect 70813 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
tri 41758 16180 41776 16198 ne
rect 41776 16180 42002 16198
tri 42002 16180 42020 16198 sw
tri 41776 16134 41822 16180 ne
rect 41822 16134 41898 16180
rect 41944 16140 42020 16180
tri 42020 16140 42060 16180 sw
rect 70813 16140 71000 16198
rect 41944 16134 42060 16140
tri 42060 16134 42066 16140 sw
tri 41822 16094 41862 16134 ne
rect 41862 16094 42066 16134
tri 42066 16094 42106 16134 sw
rect 70813 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41862 16048 41908 16094 ne
rect 41908 16048 42106 16094
tri 42106 16048 42152 16094 sw
tri 41908 16036 41920 16048 ne
rect 41920 16036 42030 16048
tri 41920 16002 41954 16036 ne
rect 41954 16002 42030 16036
rect 42076 16036 42152 16048
tri 42152 16036 42164 16048 sw
rect 70813 16036 71000 16094
rect 42076 16002 42164 16036
tri 41954 15990 41966 16002 ne
rect 41966 15990 42164 16002
tri 42164 15990 42210 16036 sw
rect 70813 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
tri 41966 15932 42024 15990 ne
rect 42024 15932 42210 15990
tri 42210 15932 42268 15990 sw
rect 70813 15932 71000 15990
tri 42024 15916 42040 15932 ne
rect 42040 15916 42268 15932
tri 42268 15916 42284 15932 sw
tri 42040 15870 42086 15916 ne
rect 42086 15870 42162 15916
rect 42208 15886 42284 15916
tri 42284 15886 42314 15916 sw
rect 70813 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 42208 15870 42314 15886
tri 42314 15870 42330 15886 sw
tri 42086 15828 42128 15870 ne
rect 42128 15828 42330 15870
tri 42330 15828 42372 15870 sw
rect 70813 15828 71000 15886
tri 42128 15792 42164 15828 ne
rect 42164 15792 42372 15828
tri 42372 15792 42408 15828 sw
tri 42164 15784 42172 15792 ne
rect 42172 15784 42408 15792
tri 42172 15738 42218 15784 ne
rect 42218 15738 42294 15784
rect 42340 15782 42408 15784
tri 42408 15782 42418 15792 sw
rect 70813 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15738 42418 15782
tri 42218 15724 42232 15738 ne
rect 42232 15724 42418 15738
tri 42418 15724 42476 15782 sw
rect 70813 15724 71000 15782
tri 42232 15678 42278 15724 ne
rect 42278 15678 42476 15724
tri 42476 15678 42522 15724 sw
rect 70813 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
tri 42278 15652 42304 15678 ne
rect 42304 15652 42522 15678
tri 42522 15652 42548 15678 sw
tri 42304 15606 42350 15652 ne
rect 42350 15606 42426 15652
rect 42472 15620 42548 15652
tri 42548 15620 42580 15652 sw
rect 70813 15620 71000 15678
rect 42472 15606 42580 15620
tri 42580 15606 42594 15620 sw
tri 42350 15574 42382 15606 ne
rect 42382 15574 42594 15606
tri 42594 15574 42626 15606 sw
rect 70813 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
tri 42382 15548 42408 15574 ne
rect 42408 15548 42626 15574
tri 42626 15548 42652 15574 sw
tri 42408 15520 42436 15548 ne
rect 42436 15520 42652 15548
tri 42436 15474 42482 15520 ne
rect 42482 15474 42558 15520
rect 42604 15516 42652 15520
tri 42652 15516 42684 15548 sw
rect 70813 15516 71000 15574
rect 42604 15474 42684 15516
tri 42482 15470 42486 15474 ne
rect 42486 15470 42684 15474
tri 42684 15470 42730 15516 sw
rect 70813 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
tri 42486 15412 42544 15470 ne
rect 42544 15412 42730 15470
tri 42730 15412 42788 15470 sw
rect 70813 15412 71000 15470
tri 42544 15388 42568 15412 ne
rect 42568 15388 42788 15412
tri 42788 15388 42812 15412 sw
tri 42568 15342 42614 15388 ne
rect 42614 15342 42690 15388
rect 42736 15366 42812 15388
tri 42812 15366 42834 15388 sw
rect 70813 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15342 42834 15366
tri 42834 15342 42858 15366 sw
tri 42614 15308 42648 15342 ne
rect 42648 15308 42858 15342
tri 42858 15308 42892 15342 sw
rect 70813 15308 71000 15366
tri 42648 15304 42652 15308 ne
rect 42652 15304 42892 15308
tri 42892 15304 42896 15308 sw
tri 42652 15262 42694 15304 ne
rect 42694 15262 42896 15304
tri 42896 15262 42938 15304 sw
rect 70813 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
tri 42694 15256 42700 15262 ne
rect 42700 15256 42938 15262
tri 42700 15210 42746 15256 ne
rect 42746 15210 42822 15256
rect 42868 15210 42938 15256
tri 42746 15204 42752 15210 ne
rect 42752 15204 42938 15210
tri 42938 15204 42996 15262 sw
rect 70813 15204 71000 15262
tri 42752 15158 42798 15204 ne
rect 42798 15158 42996 15204
tri 42996 15158 43042 15204 sw
rect 70813 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42798 15124 42832 15158 ne
rect 42832 15124 43042 15158
tri 43042 15124 43076 15158 sw
tri 42832 15078 42878 15124 ne
rect 42878 15078 42954 15124
rect 43000 15100 43076 15124
tri 43076 15100 43100 15124 sw
rect 70813 15100 71000 15158
rect 43000 15078 43100 15100
tri 43100 15078 43122 15100 sw
tri 42878 15060 42896 15078 ne
rect 42896 15060 43122 15078
tri 43122 15060 43140 15078 sw
tri 42896 15054 42902 15060 ne
rect 42902 15054 43140 15060
tri 43140 15054 43146 15060 sw
rect 70813 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42902 14996 42960 15054 ne
rect 42960 14996 43146 15054
tri 43146 14996 43204 15054 sw
rect 70813 14996 71000 15054
tri 42960 14992 42964 14996 ne
rect 42964 14992 43204 14996
tri 42964 14946 43010 14992 ne
rect 43010 14946 43086 14992
rect 43132 14950 43204 14992
tri 43204 14950 43250 14996 sw
rect 70813 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 43132 14946 43250 14950
tri 43010 14892 43064 14946 ne
rect 43064 14892 43250 14946
tri 43250 14892 43308 14950 sw
rect 70813 14892 71000 14950
tri 43064 14860 43096 14892 ne
rect 43096 14860 43308 14892
tri 43308 14860 43340 14892 sw
tri 43096 14816 43140 14860 ne
rect 43140 14816 43218 14860
tri 43140 14814 43142 14816 ne
rect 43142 14814 43218 14816
rect 43264 14846 43340 14860
tri 43340 14846 43354 14860 sw
rect 70813 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 43264 14816 43354 14846
tri 43354 14816 43384 14846 sw
rect 43264 14814 43384 14816
tri 43142 14788 43168 14814 ne
rect 43168 14788 43384 14814
tri 43384 14788 43412 14816 sw
rect 70813 14788 71000 14846
tri 43168 14742 43214 14788 ne
rect 43214 14742 43412 14788
tri 43412 14742 43458 14788 sw
rect 70813 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
tri 43214 14728 43228 14742 ne
rect 43228 14728 43458 14742
tri 43458 14728 43472 14742 sw
tri 43228 14682 43274 14728 ne
rect 43274 14682 43350 14728
rect 43396 14684 43472 14728
tri 43472 14684 43516 14728 sw
rect 70813 14684 71000 14742
rect 43396 14682 43516 14684
tri 43516 14682 43518 14684 sw
tri 43274 14638 43318 14682 ne
rect 43318 14638 43518 14682
tri 43518 14638 43562 14682 sw
rect 70813 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43318 14596 43360 14638 ne
rect 43360 14596 43562 14638
tri 43562 14596 43604 14638 sw
tri 43360 14572 43384 14596 ne
rect 43384 14572 43482 14596
tri 43384 14550 43406 14572 ne
rect 43406 14550 43482 14572
rect 43528 14580 43604 14596
tri 43604 14580 43620 14596 sw
rect 70813 14580 71000 14638
rect 43528 14572 43620 14580
tri 43620 14572 43628 14580 sw
rect 43528 14550 43628 14572
tri 43406 14534 43422 14550 ne
rect 43422 14534 43628 14550
tri 43628 14534 43666 14572 sw
rect 70813 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
tri 43422 14476 43480 14534 ne
rect 43480 14476 43666 14534
tri 43666 14476 43724 14534 sw
rect 70813 14476 71000 14534
tri 43480 14464 43492 14476 ne
rect 43492 14464 43724 14476
tri 43724 14464 43736 14476 sw
tri 43492 14418 43538 14464 ne
rect 43538 14418 43614 14464
rect 43660 14430 43736 14464
tri 43736 14430 43770 14464 sw
rect 70813 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 43660 14418 43770 14430
tri 43770 14418 43782 14430 sw
tri 43538 14372 43584 14418 ne
rect 43584 14372 43782 14418
tri 43782 14372 43828 14418 sw
rect 70813 14372 71000 14430
tri 43584 14332 43624 14372 ne
rect 43624 14332 43828 14372
tri 43828 14332 43868 14372 sw
tri 43624 14328 43628 14332 ne
rect 43628 14328 43746 14332
tri 43628 14286 43670 14328 ne
rect 43670 14286 43746 14328
rect 43792 14328 43868 14332
tri 43868 14328 43872 14332 sw
rect 43792 14326 43872 14328
tri 43872 14326 43874 14328 sw
rect 70813 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43792 14286 43874 14326
tri 43670 14268 43688 14286 ne
rect 43688 14268 43874 14286
tri 43874 14268 43932 14326 sw
rect 70813 14268 71000 14326
tri 43688 14222 43734 14268 ne
rect 43734 14222 43932 14268
tri 43932 14222 43978 14268 sw
rect 70813 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43734 14200 43756 14222 ne
rect 43756 14200 43978 14222
tri 43978 14200 44000 14222 sw
tri 43756 14154 43802 14200 ne
rect 43802 14154 43878 14200
rect 43924 14164 44000 14200
tri 44000 14164 44036 14200 sw
rect 70813 14164 71000 14222
rect 43924 14154 44036 14164
tri 44036 14154 44046 14164 sw
tri 43802 14118 43838 14154 ne
rect 43838 14118 44046 14154
tri 44046 14118 44082 14154 sw
rect 70813 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
tri 43838 14084 43872 14118 ne
rect 43872 14084 44082 14118
tri 44082 14084 44116 14118 sw
tri 43872 14068 43888 14084 ne
rect 43888 14068 44116 14084
tri 43888 14022 43934 14068 ne
rect 43934 14022 44010 14068
rect 44056 14060 44116 14068
tri 44116 14060 44140 14084 sw
rect 70813 14060 71000 14118
rect 44056 14022 44140 14060
tri 43934 14014 43942 14022 ne
rect 43942 14014 44140 14022
tri 44140 14014 44186 14060 sw
rect 70813 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
tri 43942 13956 44000 14014 ne
rect 44000 13956 44186 14014
tri 44186 13956 44244 14014 sw
rect 70813 13956 71000 14014
tri 44000 13936 44020 13956 ne
rect 44020 13936 44244 13956
tri 44244 13936 44264 13956 sw
tri 44020 13890 44066 13936 ne
rect 44066 13890 44142 13936
rect 44188 13910 44264 13936
tri 44264 13910 44290 13936 sw
rect 70813 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 44188 13890 44290 13910
tri 44290 13890 44310 13910 sw
tri 44066 13852 44104 13890 ne
rect 44104 13852 44310 13890
tri 44310 13852 44348 13890 sw
rect 70813 13852 71000 13910
tri 44104 13840 44116 13852 ne
rect 44116 13840 44348 13852
tri 44348 13840 44360 13852 sw
tri 44116 13806 44150 13840 ne
rect 44150 13806 44360 13840
tri 44360 13806 44394 13840 sw
rect 70813 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
tri 44150 13804 44152 13806 ne
rect 44152 13804 44394 13806
tri 44152 13758 44198 13804 ne
rect 44198 13758 44274 13804
rect 44320 13758 44394 13804
tri 44198 13748 44208 13758 ne
rect 44208 13748 44394 13758
tri 44394 13748 44452 13806 sw
rect 70813 13748 71000 13806
tri 44208 13702 44254 13748 ne
rect 44254 13702 44452 13748
tri 44452 13702 44498 13748 sw
rect 70813 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
tri 44254 13672 44284 13702 ne
rect 44284 13672 44498 13702
tri 44498 13672 44528 13702 sw
tri 44284 13626 44330 13672 ne
rect 44330 13626 44406 13672
rect 44452 13644 44528 13672
tri 44528 13644 44556 13672 sw
rect 70813 13644 71000 13702
rect 44452 13626 44556 13644
tri 44556 13626 44574 13644 sw
tri 44330 13598 44358 13626 ne
rect 44358 13598 44574 13626
tri 44574 13598 44602 13626 sw
rect 70813 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
tri 44358 13596 44360 13598 ne
rect 44360 13596 44602 13598
tri 44602 13596 44604 13598 sw
tri 44360 13540 44416 13596 ne
rect 44416 13540 44604 13596
tri 44604 13540 44660 13596 sw
rect 70813 13540 71000 13598
tri 44416 13494 44462 13540 ne
rect 44462 13494 44538 13540
rect 44584 13494 44660 13540
tri 44660 13494 44706 13540 sw
rect 70813 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
tri 44462 13436 44520 13494 ne
rect 44520 13436 44706 13494
tri 44706 13436 44764 13494 sw
rect 70813 13436 71000 13494
tri 44520 13408 44548 13436 ne
rect 44548 13408 44764 13436
tri 44764 13408 44792 13436 sw
tri 44548 13362 44594 13408 ne
rect 44594 13362 44670 13408
rect 44716 13390 44792 13408
tri 44792 13390 44810 13408 sw
rect 70813 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13362 44810 13390
tri 44810 13362 44838 13390 sw
tri 44594 13352 44604 13362 ne
rect 44604 13352 44838 13362
tri 44838 13352 44848 13362 sw
tri 44604 13269 44687 13352 ne
rect 44687 13280 44848 13352
tri 44848 13280 44920 13352 sw
rect 70813 13280 71000 13390
rect 44687 13269 71000 13280
tri 44687 13256 44700 13269 ne
rect 44700 13256 45088 13269
tri 44700 13210 44746 13256 ne
rect 44746 13210 44850 13256
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
tri 44746 13165 44791 13210 ne
rect 44791 13165 71000 13210
tri 44791 13119 44837 13165 ne
rect 44837 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
tri 44837 13108 44848 13119 ne
rect 44848 13108 71000 13119
<< metal2 >>
rect 70584 68116 70702 68200
rect 70584 66916 70613 68116
rect 70669 66916 70702 68116
rect 70584 60120 70702 66916
rect 70584 58920 70613 60120
rect 70669 58920 70702 60120
rect 70584 56910 70702 58920
rect 70584 55710 70613 56910
rect 70669 55710 70702 56910
rect 70584 55302 70702 55710
rect 70584 54102 70613 55302
rect 70669 54102 70702 55302
rect 70584 53722 70702 54102
rect 70584 52522 70613 53722
rect 70669 52522 70702 53722
rect 70584 45739 70702 52522
rect 70584 42875 70613 45739
rect 70669 42875 70702 45739
rect 70584 42497 70702 42875
rect 70584 41297 70613 42497
rect 70669 41297 70702 42497
rect 70584 39332 70702 41297
rect 70584 36468 70613 39332
rect 70669 36468 70702 39332
rect 70584 36132 70702 36468
rect 70584 33268 70613 36132
rect 70669 33268 70702 36132
rect 70584 32920 70702 33268
rect 70584 30056 70613 32920
rect 70669 30056 70702 32920
rect 70584 29752 70702 30056
rect 70584 26888 70613 29752
rect 70669 26888 70702 29752
rect 70584 24906 70702 26888
rect 70584 23706 70613 24906
rect 70669 23706 70702 24906
rect 70584 23599 70702 23706
<< via2 >>
rect 70613 66916 70669 68116
rect 70613 58920 70669 60120
rect 70613 55710 70669 56910
rect 70613 54102 70669 55302
rect 70613 52522 70669 53722
rect 70613 42875 70669 45739
rect 70613 41297 70669 42497
rect 70613 36468 70669 39332
rect 70613 33268 70669 36132
rect 70613 30056 70669 32920
rect 70613 26888 70669 29752
rect 70613 23706 70669 24906
<< metal3 >>
rect 14000 47112 17000 71000
rect 17200 48448 20200 71000
rect 20400 49774 23400 71000
rect 23600 50451 25000 71000
rect 25200 51220 26600 71000
rect 26800 52454 29800 71000
rect 30000 53792 33000 71000
rect 33200 55124 36200 71000
rect 36400 56465 39400 71000
rect 39600 57138 41000 71000
rect 41200 57723 42600 71000
rect 42800 59150 45800 71000
rect 46000 60510 49000 71000
rect 49200 61175 50600 71000
rect 50800 61839 52200 71000
rect 52400 62507 53800 71000
rect 54000 63320 55400 71000
rect 55600 63836 57000 71000
rect 57200 64540 58600 71000
rect 58800 65166 60200 71000
rect 60400 65831 61800 71000
rect 62000 66494 63400 71000
rect 63600 67166 65000 71000
rect 65200 67829 66600 71000
rect 66800 68476 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68400 68693 68476 68769 ne
rect 68476 68693 71000 68769
tri 68200 68476 68417 68693 sw
tri 68476 68476 68693 68693 ne
rect 68693 68476 71000 68693
rect 66800 68200 68417 68476
tri 68417 68200 68693 68476 sw
tri 68693 68400 68769 68476 ne
rect 68769 68400 71000 68476
rect 66800 68116 71000 68200
rect 66800 68113 70613 68116
tri 66800 68029 66884 68113 ne
rect 66884 68029 70613 68113
tri 66600 67829 66800 68029 sw
tri 66884 67829 67084 68029 ne
rect 67084 67829 70613 68029
rect 65200 67545 66800 67829
tri 66800 67545 67084 67829 sw
tri 67084 67545 67368 67829 ne
rect 67368 67545 70613 67829
rect 65200 67449 67084 67545
tri 65200 67366 65283 67449 ne
rect 65283 67368 67084 67449
tri 67084 67368 67261 67545 sw
tri 67368 67368 67545 67545 ne
rect 67545 67368 70613 67545
rect 65283 67366 67261 67368
tri 65000 67166 65200 67366 sw
tri 65283 67166 65483 67366 ne
rect 65483 67166 67261 67366
rect 63600 66883 65200 67166
tri 65200 66883 65483 67166 sw
tri 65483 66883 65766 67166 ne
rect 65766 67084 67261 67166
tri 67261 67084 67545 67368 sw
tri 67545 67084 67829 67368 ne
rect 67829 67084 70613 67368
rect 65766 66883 67545 67084
rect 63600 66786 65483 66883
tri 63600 66694 63692 66786 ne
rect 63692 66694 65483 66786
tri 63400 66494 63600 66694 sw
tri 63692 66494 63892 66694 ne
rect 63892 66600 65483 66694
tri 65483 66600 65766 66883 sw
tri 65766 66600 66049 66883 ne
rect 66049 66800 67545 66883
tri 67545 66800 67829 67084 sw
tri 67829 66800 68113 67084 ne
rect 68113 66916 70613 67084
rect 70669 66916 71000 68116
rect 68113 66800 71000 66916
rect 66049 66600 67829 66800
tri 67829 66600 68029 66800 sw
rect 63892 66494 65766 66600
rect 62000 66202 63600 66494
tri 63600 66202 63892 66494 sw
tri 63892 66202 64184 66494 ne
rect 64184 66332 65766 66494
tri 65766 66332 66034 66600 sw
tri 66049 66332 66317 66600 ne
rect 66317 66332 71000 66600
rect 64184 66202 66034 66332
rect 62000 66114 63892 66202
tri 62000 66031 62083 66114 ne
rect 62083 66031 63892 66114
tri 61800 65831 62000 66031 sw
tri 62083 65831 62283 66031 ne
rect 62283 65964 63892 66031
tri 63892 65964 64130 66202 sw
tri 64184 65964 64422 66202 ne
rect 64422 66049 66034 66202
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64422 65964 66317 66049
rect 62283 65831 64130 65964
rect 60400 65663 62000 65831
tri 62000 65663 62168 65831 sw
tri 62283 65663 62451 65831 ne
rect 62451 65672 64130 65831
tri 64130 65672 64422 65964 sw
tri 64422 65672 64714 65964 ne
rect 64714 65766 66317 65964
tri 66317 65766 66600 66049 sw
tri 66600 65766 66883 66049 ne
rect 66883 65766 71000 66049
rect 64714 65672 66600 65766
rect 62451 65663 64422 65672
rect 60400 65451 62168 65663
tri 60400 65366 60485 65451 ne
rect 60485 65380 62168 65451
tri 62168 65380 62451 65663 sw
tri 62451 65380 62734 65663 ne
rect 62734 65380 64422 65663
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65483 66600 65672
tri 66600 65483 66883 65766 sw
tri 66883 65483 67166 65766 ne
rect 67166 65483 71000 65766
rect 65006 65380 66883 65483
rect 60485 65366 62451 65380
tri 60200 65166 60400 65366 sw
tri 60485 65166 60685 65366 ne
rect 60685 65166 62451 65366
rect 58800 64881 60400 65166
tri 60400 64881 60685 65166 sw
tri 60685 64881 60970 65166 ne
rect 60970 65097 62451 65166
tri 62451 65097 62734 65380 sw
tri 62734 65097 63017 65380 ne
rect 63017 65292 64714 65380
tri 64714 65292 64802 65380 sw
tri 65006 65292 65094 65380 ne
rect 65094 65292 66883 65380
rect 63017 65097 64802 65292
rect 60970 64997 62734 65097
tri 62734 64997 62834 65097 sw
tri 63017 64997 63117 65097 ne
rect 63117 65000 64802 65097
tri 64802 65000 65094 65292 sw
tri 65094 65000 65386 65292 ne
rect 65386 65200 66883 65292
tri 66883 65200 67166 65483 sw
tri 67166 65200 67449 65483 ne
rect 67449 65200 71000 65483
rect 65386 65000 67166 65200
tri 67166 65000 67366 65200 sw
rect 63117 64997 65094 65000
rect 60970 64881 62834 64997
rect 58800 64786 60685 64881
tri 58800 64699 58887 64786 ne
rect 58887 64730 60685 64786
tri 60685 64730 60836 64881 sw
tri 60970 64730 61121 64881 ne
rect 61121 64730 62834 64881
rect 58887 64699 60836 64730
tri 58600 64540 58759 64699 sw
tri 58887 64540 59046 64699 ne
rect 59046 64540 60836 64699
rect 57200 64499 58759 64540
tri 58759 64499 58800 64540 sw
tri 59046 64499 59087 64540 ne
rect 59087 64499 60836 64540
rect 57200 64447 58800 64499
tri 58800 64447 58852 64499 sw
tri 59087 64447 59139 64499 ne
rect 59139 64447 60836 64499
rect 57200 64160 58852 64447
tri 58852 64160 59139 64447 sw
tri 59139 64160 59426 64447 ne
rect 59426 64445 60836 64447
tri 60836 64445 61121 64730 sw
tri 61121 64445 61406 64730 ne
rect 61406 64714 62834 64730
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61406 64445 63117 64714
rect 59426 64160 61121 64445
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63117 64445
tri 63117 64431 63400 64714 sw
tri 63400 64431 63683 64714 ne
rect 63683 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63683 64431 65386 64708
rect 61691 64160 63400 64431
rect 57200 64119 59139 64160
tri 57200 64036 57283 64119 ne
rect 57283 64036 59139 64119
tri 57000 63836 57200 64036 sw
tri 57283 63836 57483 64036 ne
rect 57483 63873 59139 64036
tri 59139 63873 59426 64160 sw
tri 59426 63873 59713 64160 ne
rect 59713 64065 61406 64160
tri 61406 64065 61501 64160 sw
tri 61691 64065 61786 64160 ne
rect 61786 64148 63400 64160
tri 63400 64148 63683 64431 sw
tri 63683 64148 63966 64431 ne
rect 63966 64416 65386 64431
tri 65386 64416 65678 64708 sw
tri 65678 64416 65970 64708 ne
rect 65970 64416 71000 64708
rect 63966 64184 65678 64416
tri 65678 64184 65910 64416 sw
tri 65970 64184 66202 64416 ne
rect 66202 64184 71000 64416
rect 63966 64148 65910 64184
rect 61786 64065 63683 64148
rect 59713 63873 61501 64065
rect 57483 63836 59426 63873
rect 55600 63553 57200 63836
tri 57200 63553 57483 63836 sw
tri 57483 63553 57766 63836 ne
rect 57766 63673 59426 63836
tri 59426 63673 59626 63873 sw
tri 59713 63673 59913 63873 ne
rect 59913 63780 61501 63873
tri 61501 63780 61786 64065 sw
tri 61786 63780 62071 64065 ne
rect 62071 63966 63683 64065
tri 63683 63966 63865 64148 sw
tri 63966 63966 64148 64148 ne
rect 64148 63966 65910 64148
rect 62071 63780 63865 63966
rect 59913 63673 61786 63780
rect 57766 63553 59626 63673
rect 55600 63506 57483 63553
tri 57483 63506 57530 63553 sw
tri 57766 63506 57813 63553 ne
rect 57813 63506 59626 63553
rect 55600 63456 57530 63506
tri 55600 63373 55683 63456 ne
rect 55683 63373 57530 63456
tri 55400 63320 55453 63373 sw
tri 55683 63320 55736 63373 ne
rect 55736 63320 57530 63373
rect 54000 63173 55453 63320
tri 55453 63173 55600 63320 sw
tri 55736 63173 55883 63320 ne
rect 55883 63223 57530 63320
tri 57530 63223 57813 63506 sw
tri 57813 63223 58096 63506 ne
rect 58096 63386 59626 63506
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63683 63865 63780
tri 63865 63683 64148 63966 sw
tri 64148 63683 64431 63966 ne
rect 64431 63892 65910 63966
tri 65910 63892 66202 64184 sw
tri 66202 63892 66494 64184 ne
rect 66494 63892 71000 64184
rect 64431 63683 66202 63892
rect 62356 63495 64148 63683
rect 60200 63386 62071 63495
rect 58096 63223 59913 63386
rect 55883 63173 57813 63223
rect 54000 62940 55600 63173
tri 55600 62940 55833 63173 sw
tri 55883 62940 56116 63173 ne
rect 56116 62940 57813 63173
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59913 63223
tri 59913 63099 60200 63386 sw
tri 60200 63099 60487 63386 ne
rect 60487 63210 62071 63386
tri 62071 63210 62356 63495 sw
tri 62356 63210 62641 63495 ne
rect 62641 63400 64148 63495
tri 64148 63400 64431 63683 sw
tri 64431 63400 64714 63683 ne
rect 64714 63600 66202 63683
tri 66202 63600 66494 63892 sw
tri 66494 63600 66786 63892 ne
rect 66786 63600 71000 63892
rect 64714 63400 66494 63600
tri 66494 63400 66694 63600 sw
rect 62641 63210 64431 63400
rect 60487 63099 62356 63210
rect 58379 62940 60200 63099
rect 54000 62793 55833 62940
tri 54000 62707 54086 62793 ne
rect 54086 62707 55833 62793
tri 53800 62507 54000 62707 sw
tri 54086 62507 54286 62707 ne
rect 54286 62657 55833 62707
tri 55833 62657 56116 62940 sw
tri 56116 62657 56399 62940 ne
rect 56399 62843 58096 62940
tri 58096 62843 58193 62940 sw
tri 58379 62843 58476 62940 ne
rect 58476 62843 60200 62940
rect 56399 62657 58193 62843
rect 54286 62622 56116 62657
tri 56116 62622 56151 62657 sw
tri 56399 62622 56434 62657 ne
rect 56434 62622 58193 62657
rect 54286 62507 56151 62622
rect 52400 62221 54000 62507
tri 54000 62221 54286 62507 sw
tri 54286 62221 54572 62507 ne
rect 54572 62339 56151 62507
tri 56151 62339 56434 62622 sw
tri 56434 62339 56717 62622 ne
rect 56717 62560 58193 62622
tri 58193 62560 58476 62843 sw
tri 58476 62560 58759 62843 ne
rect 58759 62812 60200 62843
tri 60200 62812 60487 63099 sw
tri 60487 62812 60774 63099 ne
rect 60774 62925 62356 63099
tri 62356 62925 62641 63210 sw
tri 62641 62925 62926 63210 ne
rect 62926 63117 64431 63210
tri 64431 63117 64714 63400 sw
tri 64714 63117 64997 63400 ne
rect 64997 63117 71000 63400
rect 62926 62925 64714 63117
rect 60774 62812 62641 62925
rect 58759 62754 60487 62812
tri 60487 62754 60545 62812 sw
tri 60774 62754 60832 62812 ne
rect 60832 62754 62641 62812
rect 58759 62560 60545 62754
rect 56717 62339 58476 62560
rect 54572 62221 56434 62339
rect 52400 62127 54286 62221
tri 52400 62039 52488 62127 ne
rect 52488 62039 54286 62127
tri 52200 61839 52400 62039 sw
tri 52488 61839 52688 62039 ne
rect 52688 62006 54286 62039
tri 54286 62006 54501 62221 sw
tri 54572 62006 54787 62221 ne
rect 54787 62056 56434 62221
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62467 60545 62560
tri 60545 62467 60832 62754 sw
tri 60832 62467 61119 62754 ne
rect 61119 62750 62641 62754
tri 62641 62750 62816 62925 sw
tri 62926 62750 63101 62925 ne
rect 63101 62834 64714 62925
tri 64714 62834 64997 63117 sw
tri 64997 62834 65280 63117 ne
rect 65280 62834 71000 63117
rect 63101 62750 64997 62834
rect 61119 62467 62816 62750
rect 59042 62277 60832 62467
rect 57000 62056 58759 62277
rect 54787 62006 56717 62056
rect 52688 61839 54501 62006
rect 50800 61720 52400 61839
tri 52400 61720 52519 61839 sw
tri 52688 61720 52807 61839 ne
rect 52807 61720 54501 61839
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56717 62006
tri 56717 61773 57000 62056 sw
tri 57000 61773 57283 62056 ne
rect 57283 61994 58759 62056
tri 58759 61994 59042 62277 sw
tri 59042 61994 59325 62277 ne
rect 59325 62180 60832 62277
tri 60832 62180 61119 62467 sw
tri 61119 62180 61406 62467 ne
rect 61406 62465 62816 62467
tri 62816 62465 63101 62750 sw
tri 63101 62465 63386 62750 ne
rect 63386 62566 64997 62750
tri 64997 62566 65265 62834 sw
tri 65280 62566 65548 62834 ne
rect 65548 62566 71000 62834
rect 63386 62465 65265 62566
rect 61406 62180 63101 62465
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62283 65265 62465
tri 65265 62283 65548 62566 sw
tri 65548 62283 65831 62566 ne
rect 65831 62283 71000 62566
rect 63671 62180 65548 62283
rect 59325 61994 61119 62180
rect 57283 61773 59042 61994
rect 55073 61720 57000 61773
rect 50800 61459 52519 61720
tri 50800 61375 50884 61459 ne
rect 50884 61432 52519 61459
tri 52519 61432 52807 61720 sw
tri 52807 61432 53095 61720 ne
rect 53095 61626 54787 61720
tri 54787 61626 54881 61720 sw
tri 55073 61626 55167 61720 ne
rect 55167 61626 57000 61720
rect 53095 61432 54881 61626
rect 50884 61375 52807 61432
tri 50600 61175 50800 61375 sw
tri 50884 61175 51084 61375 ne
rect 51084 61303 52807 61375
tri 52807 61303 52936 61432 sw
tri 53095 61303 53224 61432 ne
rect 53224 61340 54881 61432
tri 54881 61340 55167 61626 sw
tri 55167 61340 55453 61626 ne
rect 55453 61490 57000 61626
tri 57000 61490 57283 61773 sw
tri 57283 61490 57566 61773 ne
rect 57566 61711 59042 61773
tri 59042 61711 59325 61994 sw
tri 59325 61711 59608 61994 ne
rect 59608 61893 61119 61994
tri 61119 61893 61406 62180 sw
tri 61406 61893 61693 62180 ne
rect 61693 62085 63386 62180
tri 63386 62085 63481 62180 sw
tri 63671 62085 63766 62180 ne
rect 63766 62085 65548 62180
rect 61693 61893 63481 62085
rect 59608 61711 61406 61893
rect 57566 61526 59325 61711
tri 59325 61526 59510 61711 sw
tri 59608 61526 59793 61711 ne
rect 59793 61606 61406 61711
tri 61406 61606 61693 61893 sw
tri 61693 61606 61980 61893 ne
rect 61980 61800 63481 61893
tri 63481 61800 63766 62085 sw
tri 63766 61800 64051 62085 ne
rect 64051 62000 65548 62085
tri 65548 62000 65831 62283 sw
tri 65831 62000 66114 62283 ne
rect 66114 62000 71000 62283
rect 64051 61800 65831 62000
tri 65831 61800 66031 62000 sw
rect 61980 61606 63766 61800
rect 59793 61526 61693 61606
rect 57566 61490 59510 61526
rect 55453 61340 57283 61490
rect 53224 61303 55167 61340
rect 51084 61175 52936 61303
rect 49200 60891 50800 61175
tri 50800 60891 51084 61175 sw
tri 51084 60891 51368 61175 ne
rect 51368 61015 52936 61175
tri 52936 61015 53224 61303 sw
tri 53224 61015 53512 61303 ne
rect 53512 61054 55167 61303
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61243 57283 61340
tri 57283 61243 57530 61490 sw
tri 57566 61243 57813 61490 ne
rect 57813 61243 59510 61490
tri 59510 61243 59793 61526 sw
tri 59793 61243 60076 61526 ne
rect 60076 61319 61693 61526
tri 61693 61319 61980 61606 sw
tri 61980 61319 62267 61606 ne
rect 62267 61515 63766 61606
tri 63766 61515 64051 61800 sw
tri 64051 61515 64336 61800 ne
rect 64336 61515 71000 61800
rect 62267 61319 64051 61515
rect 60076 61243 61980 61319
rect 55739 61054 57530 61243
rect 53512 61015 55453 61054
rect 51368 60891 53224 61015
rect 49200 60795 51084 60891
tri 49200 60710 49285 60795 ne
rect 49285 60784 51084 60795
tri 51084 60784 51191 60891 sw
tri 51368 60784 51475 60891 ne
rect 51475 60784 53224 60891
rect 49285 60710 51191 60784
tri 49000 60510 49200 60710 sw
tri 49285 60510 49485 60710 ne
rect 49485 60510 51191 60710
rect 46000 60500 49200 60510
tri 49200 60500 49210 60510 sw
tri 49485 60500 49495 60510 ne
rect 49495 60500 51191 60510
tri 51191 60500 51475 60784 sw
tri 51475 60500 51759 60784 ne
rect 51759 60727 53224 60784
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60768 55453 61015
tri 55453 60768 55739 61054 sw
tri 55739 60768 56025 61054 ne
rect 56025 60960 57530 61054
tri 57530 60960 57813 61243 sw
tri 57813 60960 58096 61243 ne
rect 58096 60960 59793 61243
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 61154 61980 61243
tri 61980 61154 62145 61319 sw
tri 62267 61154 62432 61319 ne
rect 62432 61230 64051 61319
tri 64051 61230 64336 61515 sw
tri 64336 61230 64621 61515 ne
rect 64621 61230 71000 61515
rect 62432 61154 64336 61230
rect 60359 60960 62145 61154
rect 56025 60768 57813 60960
rect 53800 60727 55739 60768
rect 51759 60500 53512 60727
rect 46000 60215 49210 60500
tri 49210 60215 49495 60500 sw
tri 49495 60215 49780 60500 ne
rect 49780 60404 51475 60500
tri 51475 60404 51571 60500 sw
tri 51759 60404 51855 60500 ne
rect 51855 60439 53512 60500
tri 53512 60439 53800 60727 sw
tri 53800 60439 54088 60727 ne
rect 54088 60482 55739 60727
tri 55739 60482 56025 60768 sw
tri 56025 60482 56311 60768 ne
rect 56311 60677 57813 60768
tri 57813 60677 58096 60960 sw
tri 58096 60677 58379 60960 ne
rect 58379 60863 60076 60960
tri 60076 60863 60173 60960 sw
tri 60359 60863 60456 60960 ne
rect 60456 60867 62145 60960
tri 62145 60867 62432 61154 sw
tri 62432 60867 62719 61154 ne
rect 62719 60970 64336 61154
tri 64336 60970 64596 61230 sw
tri 64621 60970 64881 61230 ne
rect 64881 60970 71000 61230
rect 62719 60867 64596 60970
rect 60456 60863 62432 60867
rect 58379 60677 60173 60863
rect 56311 60482 58096 60677
rect 54088 60439 56025 60482
rect 51855 60404 53800 60439
rect 49780 60215 51571 60404
rect 46000 59965 49495 60215
tri 49495 59965 49745 60215 sw
tri 49780 59965 50030 60215 ne
rect 50030 60120 51571 60215
tri 51571 60120 51855 60404 sw
tri 51855 60120 52139 60404 ne
rect 52139 60151 53800 60404
tri 53800 60151 54088 60439 sw
tri 54088 60151 54376 60439 ne
rect 54376 60312 56025 60439
tri 56025 60312 56195 60482 sw
tri 56311 60312 56481 60482 ne
rect 56481 60394 58096 60482
tri 58096 60394 58379 60677 sw
tri 58379 60394 58662 60677 ne
rect 58662 60580 60173 60677
tri 60173 60580 60456 60863 sw
tri 60456 60580 60739 60863 ne
rect 60739 60580 62432 60863
tri 62432 60580 62719 60867 sw
tri 62719 60580 63006 60867 ne
rect 63006 60685 64596 60867
tri 64596 60685 64881 60970 sw
tri 64881 60685 65166 60970 ne
rect 65166 60685 71000 60970
rect 63006 60580 64881 60685
rect 58662 60394 60456 60580
rect 56481 60312 58379 60394
rect 54376 60151 56195 60312
rect 52139 60120 54088 60151
rect 50030 60059 51855 60120
tri 51855 60059 51916 60120 sw
tri 52139 60059 52200 60120 ne
rect 52200 60059 54088 60120
rect 50030 59965 51916 60059
rect 46000 59680 49745 59965
tri 49745 59680 50030 59965 sw
tri 50030 59680 50315 59965 ne
rect 50315 59775 51916 59965
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 60028 54088 60059
tri 54088 60028 54211 60151 sw
tri 54376 60028 54499 60151 ne
rect 54499 60028 56195 60151
rect 52484 59775 54211 60028
rect 50315 59680 52200 59775
rect 46000 59461 50030 59680
tri 46000 59350 46111 59461 ne
rect 46111 59395 50030 59461
tri 50030 59395 50315 59680 sw
tri 50315 59395 50600 59680 ne
rect 50600 59491 52200 59680
tri 52200 59491 52484 59775 sw
tri 52484 59491 52768 59775 ne
rect 52768 59740 54211 59775
tri 54211 59740 54499 60028 sw
tri 54499 59740 54787 60028 ne
rect 54787 60026 56195 60028
tri 56195 60026 56481 60312 sw
tri 56481 60026 56767 60312 ne
rect 56767 60111 58379 60312
tri 58379 60111 58662 60394 sw
tri 58662 60111 58945 60394 ne
rect 58945 60297 60456 60394
tri 60456 60297 60739 60580 sw
tri 60739 60297 61022 60580 ne
rect 61022 60487 62719 60580
tri 62719 60487 62812 60580 sw
tri 63006 60487 63099 60580 ne
rect 63099 60487 64881 60580
rect 61022 60297 62812 60487
rect 58945 60111 60739 60297
rect 56767 60026 58662 60111
rect 54787 59740 56481 60026
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 59926 58662 60026
tri 58662 59926 58847 60111 sw
tri 58945 59926 59130 60111 ne
rect 59130 60014 60739 60111
tri 60739 60014 61022 60297 sw
tri 61022 60014 61305 60297 ne
rect 61305 60200 62812 60297
tri 62812 60200 63099 60487 sw
tri 63099 60200 63386 60487 ne
rect 63386 60400 64881 60487
tri 64881 60400 65166 60685 sw
tri 65166 60400 65451 60685 ne
rect 65451 60400 71000 60685
rect 63386 60200 65166 60400
tri 65166 60200 65366 60400 sw
rect 61305 60014 63099 60200
rect 59130 59926 61022 60014
rect 57053 59740 58847 59926
rect 52768 59491 54499 59740
rect 50600 59395 52484 59491
rect 46111 59350 50315 59395
tri 45800 59150 46000 59350 sw
tri 46111 59150 46311 59350 ne
rect 46311 59150 50315 59350
rect 42800 59058 46000 59150
tri 46000 59058 46092 59150 sw
tri 46311 59058 46403 59150 ne
rect 46403 59110 50315 59150
tri 50315 59110 50600 59395 sw
tri 50600 59110 50885 59395 ne
rect 50885 59207 52484 59395
tri 52484 59207 52768 59491 sw
tri 52768 59207 53052 59491 ne
rect 53052 59452 54499 59491
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59646 56767 59740
tri 56767 59646 56861 59740 sw
tri 57053 59646 57147 59740 ne
rect 57147 59646 58847 59740
rect 55075 59452 56861 59646
rect 53052 59207 54787 59452
rect 50885 59110 52768 59207
rect 46403 59058 50600 59110
rect 42800 58747 46092 59058
tri 46092 58747 46403 59058 sw
tri 46403 58747 46714 59058 ne
rect 46714 58825 50600 59058
tri 50600 58825 50885 59110 sw
tri 50885 58825 51170 59110 ne
rect 51170 59088 52768 59110
tri 52768 59088 52887 59207 sw
tri 53052 59088 53171 59207 ne
rect 53171 59164 54787 59207
tri 54787 59164 55075 59452 sw
tri 55075 59164 55363 59452 ne
rect 55363 59360 56861 59452
tri 56861 59360 57147 59646 sw
tri 57147 59360 57433 59646 ne
rect 57433 59643 58847 59646
tri 58847 59643 59130 59926 sw
tri 59130 59643 59413 59926 ne
rect 59413 59731 61022 59926
tri 61022 59731 61305 60014 sw
tri 61305 59731 61588 60014 ne
rect 61588 59913 63099 60014
tri 63099 59913 63386 60200 sw
tri 63386 59913 63673 60200 ne
rect 63673 60120 71000 60200
rect 63673 59913 70613 60120
rect 61588 59731 63386 59913
rect 59413 59643 61305 59731
rect 57433 59360 59130 59643
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59546 61305 59643
tri 61305 59546 61490 59731 sw
tri 61588 59546 61773 59731 ne
rect 61773 59626 63386 59731
tri 63386 59626 63673 59913 sw
tri 63673 59626 63960 59913 ne
rect 63960 59626 70613 59913
rect 61773 59546 63673 59626
rect 59696 59360 61490 59546
rect 55363 59164 57147 59360
rect 53171 59088 55075 59164
rect 51170 58825 52887 59088
rect 46714 58805 50885 58825
tri 50885 58805 50905 58825 sw
tri 51170 58805 51190 58825 ne
rect 51190 58805 52887 58825
rect 46714 58747 50905 58805
rect 42800 58436 46403 58747
tri 46403 58436 46714 58747 sw
tri 46714 58436 47025 58747 ne
rect 47025 58520 50905 58747
tri 50905 58520 51190 58805 sw
tri 51190 58520 51475 58805 ne
rect 51475 58804 52887 58805
tri 52887 58804 53171 59088 sw
tri 53171 58804 53455 59088 ne
rect 53455 58876 55075 59088
tri 55075 58876 55363 59164 sw
tri 55363 58876 55651 59164 ne
rect 55651 59074 57147 59164
tri 57147 59074 57433 59360 sw
tri 57433 59074 57719 59360 ne
rect 57719 59263 59413 59360
tri 59413 59263 59510 59360 sw
tri 59696 59263 59793 59360 ne
rect 59793 59263 61490 59360
tri 61490 59263 61773 59546 sw
tri 61773 59263 62056 59546 ne
rect 62056 59374 63673 59546
tri 63673 59374 63925 59626 sw
tri 63960 59374 64212 59626 ne
rect 64212 59374 70613 59626
rect 62056 59263 63925 59374
rect 57719 59074 59510 59263
rect 55651 58876 57433 59074
rect 53455 58804 55363 58876
rect 51475 58520 53171 58804
tri 53171 58520 53455 58804 sw
tri 53455 58520 53739 58804 ne
rect 53739 58716 55363 58804
tri 55363 58716 55523 58876 sw
tri 55651 58716 55811 58876 ne
rect 55811 58788 57433 58876
tri 57433 58788 57719 59074 sw
tri 57719 58788 58005 59074 ne
rect 58005 58980 59510 59074
tri 59510 58980 59793 59263 sw
tri 59793 58980 60076 59263 ne
rect 60076 58980 61773 59263
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 59087 63925 59263
tri 63925 59087 64212 59374 sw
tri 64212 59087 64499 59374 ne
rect 64499 59087 70613 59374
rect 62339 58980 64212 59087
rect 58005 58788 59793 58980
rect 55811 58716 57719 58788
rect 53739 58520 55523 58716
rect 47025 58436 51190 58520
rect 42800 58125 46714 58436
tri 46714 58125 47025 58436 sw
tri 47025 58125 47336 58436 ne
rect 47336 58235 51190 58436
tri 51190 58235 51475 58520 sw
tri 51475 58235 51760 58520 ne
rect 51760 58424 53455 58520
tri 53455 58424 53551 58520 sw
tri 53739 58424 53835 58520 ne
rect 53835 58428 55523 58520
tri 55523 58428 55811 58716 sw
tri 55811 58428 56099 58716 ne
rect 56099 58502 57719 58716
tri 57719 58502 58005 58788 sw
tri 58005 58502 58291 58788 ne
rect 58291 58697 59793 58788
tri 59793 58697 60076 58980 sw
tri 60076 58697 60359 58980 ne
rect 60359 58883 62056 58980
tri 62056 58883 62153 58980 sw
tri 62339 58883 62436 58980 ne
rect 62436 58883 64212 58980
rect 60359 58697 62153 58883
rect 58291 58502 60076 58697
rect 56099 58428 58005 58502
rect 53835 58424 55811 58428
rect 51760 58235 53551 58424
rect 47336 58125 51475 58235
rect 42800 58097 47025 58125
tri 42800 58010 42887 58097 ne
rect 42887 58010 47025 58097
tri 42600 57723 42887 58010 sw
tri 42887 57723 43174 58010 ne
rect 43174 57814 47025 58010
tri 47025 57814 47336 58125 sw
tri 47336 57814 47647 58125 ne
rect 47647 57950 51475 58125
tri 51475 57950 51760 58235 sw
tri 51760 57950 52045 58235 ne
rect 52045 58140 53551 58235
tri 53551 58140 53835 58424 sw
tri 53835 58140 54119 58424 ne
rect 54119 58140 55811 58424
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58332 58005 58428
tri 58005 58332 58175 58502 sw
tri 58291 58332 58461 58502 ne
rect 58461 58414 60076 58502
tri 60076 58414 60359 58697 sw
tri 60359 58414 60642 58697 ne
rect 60642 58600 62153 58697
tri 62153 58600 62436 58883 sw
tri 62436 58600 62719 58883 ne
rect 62719 58800 64212 58883
tri 64212 58800 64499 59087 sw
tri 64499 58800 64786 59087 ne
rect 64786 58920 70613 59087
rect 70669 58920 71000 60120
rect 64786 58800 71000 58920
rect 62719 58600 64499 58800
tri 64499 58600 64699 58800 sw
rect 60642 58414 62436 58600
rect 58461 58332 60359 58414
rect 56387 58140 58175 58332
rect 52045 57950 53835 58140
rect 47647 57814 51760 57950
rect 43174 57723 47336 57814
rect 41200 57436 42887 57723
tri 42887 57436 43174 57723 sw
tri 43174 57436 43461 57723 ne
rect 43461 57503 47336 57723
tri 47336 57503 47647 57814 sw
tri 47647 57503 47958 57814 ne
rect 47958 57665 51760 57814
tri 51760 57665 52045 57950 sw
tri 52045 57665 52330 57950 ne
rect 52330 57856 53835 57950
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 58048 56099 58140
tri 56099 58048 56191 58140 sw
tri 56387 58048 56479 58140 ne
rect 56479 58048 58175 58140
rect 54403 57856 56191 58048
rect 52330 57665 54119 57856
rect 47958 57503 52045 57665
rect 43461 57436 47647 57503
rect 41200 57430 43174 57436
tri 41200 57338 41292 57430 ne
rect 41292 57338 43174 57430
tri 41000 57138 41200 57338 sw
tri 41292 57138 41492 57338 ne
rect 41492 57321 43174 57338
tri 43174 57321 43289 57436 sw
tri 43461 57321 43576 57436 ne
rect 43576 57321 47647 57436
rect 41492 57138 43289 57321
rect 39600 57132 41200 57138
tri 41200 57132 41206 57138 sw
tri 41492 57132 41498 57138 ne
rect 41498 57132 43289 57138
rect 39600 56840 41206 57132
tri 41206 56840 41498 57132 sw
tri 41498 56840 41790 57132 ne
rect 41790 57034 43289 57132
tri 43289 57034 43576 57321 sw
tri 43576 57034 43863 57321 ne
rect 43863 57192 47647 57321
tri 47647 57192 47958 57503 sw
tri 47958 57192 48269 57503 ne
rect 48269 57395 52045 57503
tri 52045 57395 52315 57665 sw
tri 52330 57395 52600 57665 ne
rect 52600 57572 54119 57665
tri 54119 57572 54403 57856 sw
tri 54403 57572 54687 57856 ne
rect 54687 57760 56191 57856
tri 56191 57760 56479 58048 sw
tri 56479 57760 56767 58048 ne
rect 56767 58046 58175 58048
tri 58175 58046 58461 58332 sw
tri 58461 58046 58747 58332 ne
rect 58747 58131 60359 58332
tri 60359 58131 60642 58414 sw
tri 60642 58131 60925 58414 ne
rect 60925 58317 62436 58414
tri 62436 58317 62719 58600 sw
tri 62719 58317 63002 58600 ne
rect 63002 58317 71000 58600
rect 60925 58131 62719 58317
rect 58747 58046 60642 58131
rect 56767 57760 58461 58046
tri 58461 57760 58747 58046 sw
tri 58747 57760 59033 58046 ne
rect 59033 57946 60642 58046
tri 60642 57946 60827 58131 sw
tri 60925 57946 61110 58131 ne
rect 61110 58034 62719 58131
tri 62719 58034 63002 58317 sw
tri 63002 58034 63285 58317 ne
rect 63285 58034 71000 58317
rect 61110 57946 63002 58034
rect 59033 57760 60827 57946
rect 54687 57572 56479 57760
rect 52600 57395 54403 57572
rect 48269 57192 52315 57395
rect 43863 57114 47958 57192
tri 47958 57114 48036 57192 sw
tri 48269 57114 48347 57192 ne
rect 48347 57114 52315 57192
rect 43863 57034 48036 57114
rect 41790 56840 43576 57034
rect 39600 56758 41498 56840
tri 39600 56665 39693 56758 ne
rect 39693 56752 41498 56758
tri 41498 56752 41586 56840 sw
tri 41790 56752 41878 56840 ne
rect 41878 56752 43576 56840
rect 39693 56665 41586 56752
tri 39400 56465 39600 56665 sw
tri 39693 56465 39893 56665 ne
rect 39893 56465 41586 56665
rect 36400 56172 39600 56465
tri 39600 56172 39893 56465 sw
tri 39893 56172 40186 56465 ne
rect 40186 56460 41586 56465
tri 41586 56460 41878 56752 sw
tri 41878 56460 42170 56752 ne
rect 42170 56747 43576 56752
tri 43576 56747 43863 57034 sw
tri 43863 56747 44150 57034 ne
rect 44150 56803 48036 57034
tri 48036 56803 48347 57114 sw
tri 48347 56803 48658 57114 ne
rect 48658 57110 52315 57114
tri 52315 57110 52600 57395 sw
tri 52600 57110 52885 57395 ne
rect 52885 57288 54403 57395
tri 54403 57288 54687 57572 sw
tri 54687 57288 54971 57572 ne
rect 54971 57472 56479 57572
tri 56479 57472 56767 57760 sw
tri 56767 57472 57055 57760 ne
rect 57055 57666 58747 57760
tri 58747 57666 58841 57760 sw
tri 59033 57666 59127 57760 ne
rect 59127 57666 60827 57760
rect 57055 57472 58841 57666
rect 54971 57288 56767 57472
rect 52885 57110 54687 57288
rect 48658 56825 52600 57110
tri 52600 56825 52885 57110 sw
tri 52885 56825 53170 57110 ne
rect 53170 57108 54687 57110
tri 54687 57108 54867 57288 sw
tri 54971 57108 55151 57288 ne
rect 55151 57184 56767 57288
tri 56767 57184 57055 57472 sw
tri 57055 57184 57343 57472 ne
rect 57343 57380 58841 57472
tri 58841 57380 59127 57666 sw
tri 59127 57380 59413 57666 ne
rect 59413 57663 60827 57666
tri 60827 57663 61110 57946 sw
tri 61110 57663 61393 57946 ne
rect 61393 57766 63002 57946
tri 63002 57766 63270 58034 sw
tri 63285 57766 63553 58034 ne
rect 63553 57766 71000 58034
rect 61393 57663 63270 57766
rect 59413 57380 61110 57663
tri 61110 57380 61393 57663 sw
tri 61393 57380 61676 57663 ne
rect 61676 57483 63270 57663
tri 63270 57483 63553 57766 sw
tri 63553 57483 63836 57766 ne
rect 63836 57483 71000 57766
rect 61676 57380 63553 57483
rect 57343 57184 59127 57380
rect 55151 57108 57055 57184
rect 53170 56825 54867 57108
rect 48658 56803 52885 56825
rect 44150 56747 48347 56803
rect 42170 56460 43863 56747
tri 43863 56460 44150 56747 sw
tri 44150 56460 44437 56747 ne
rect 44437 56492 48347 56747
tri 48347 56492 48658 56803 sw
tri 48658 56492 48969 56803 ne
rect 48969 56540 52885 56803
tri 52885 56540 53170 56825 sw
tri 53170 56540 53455 56825 ne
rect 53455 56824 54867 56825
tri 54867 56824 55151 57108 sw
tri 55151 56824 55435 57108 ne
rect 55435 56896 57055 57108
tri 57055 56896 57343 57184 sw
tri 57343 56896 57631 57184 ne
rect 57631 57094 59127 57184
tri 59127 57094 59413 57380 sw
tri 59413 57094 59699 57380 ne
rect 59699 57283 61393 57380
tri 61393 57283 61490 57380 sw
tri 61676 57283 61773 57380 ne
rect 61773 57283 63553 57380
rect 59699 57094 61490 57283
rect 57631 56896 59413 57094
rect 55435 56824 57343 56896
rect 53455 56540 55151 56824
tri 55151 56540 55435 56824 sw
tri 55435 56540 55719 56824 ne
rect 55719 56736 57343 56824
tri 57343 56736 57503 56896 sw
tri 57631 56736 57791 56896 ne
rect 57791 56808 59413 56896
tri 59413 56808 59699 57094 sw
tri 59699 56808 59985 57094 ne
rect 59985 57000 61490 57094
tri 61490 57000 61773 57283 sw
tri 61773 57000 62056 57283 ne
rect 62056 57200 63553 57283
tri 63553 57200 63836 57483 sw
tri 63836 57200 64119 57483 ne
rect 64119 57200 71000 57483
rect 62056 57000 63836 57200
tri 63836 57000 64036 57200 sw
rect 59985 56808 61773 57000
rect 57791 56736 59699 56808
rect 55719 56540 57503 56736
rect 48969 56492 53170 56540
rect 44437 56460 48658 56492
rect 40186 56322 41878 56460
tri 41878 56322 42016 56460 sw
tri 42170 56322 42308 56460 ne
rect 42308 56322 44150 56460
rect 40186 56172 42016 56322
rect 36400 56145 39893 56172
tri 39893 56145 39920 56172 sw
tri 40186 56145 40213 56172 ne
rect 40213 56145 42016 56172
rect 36400 55852 39920 56145
tri 39920 55852 40213 56145 sw
tri 40213 55852 40506 56145 ne
rect 40506 56030 42016 56145
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56173 44150 56322
tri 44150 56173 44437 56460 sw
tri 44437 56173 44724 56460 ne
rect 44724 56181 48658 56460
tri 48658 56181 48969 56492 sw
tri 48969 56181 49280 56492 ne
rect 49280 56255 53170 56492
tri 53170 56255 53455 56540 sw
tri 53455 56255 53740 56540 ne
rect 53740 56444 55435 56540
tri 55435 56444 55531 56540 sw
tri 55719 56444 55815 56540 ne
rect 55815 56448 57503 56540
tri 57503 56448 57791 56736 sw
tri 57791 56448 58079 56736 ne
rect 58079 56522 59699 56736
tri 59699 56522 59985 56808 sw
tri 59985 56522 60271 56808 ne
rect 60271 56717 61773 56808
tri 61773 56717 62056 57000 sw
tri 62056 56717 62339 57000 ne
rect 62339 56910 71000 57000
rect 62339 56717 70613 56910
rect 60271 56522 62056 56717
rect 58079 56448 59985 56522
rect 55815 56444 57791 56448
rect 53740 56255 55531 56444
rect 49280 56181 53455 56255
rect 44724 56173 48969 56181
rect 42600 56030 44437 56173
rect 40506 55852 42308 56030
rect 36400 55559 40213 55852
tri 40213 55559 40506 55852 sw
tri 40506 55559 40799 55852 ne
rect 40799 55738 42308 55852
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55886 44437 56030
tri 44437 55886 44724 56173 sw
tri 44724 55886 45011 56173 ne
rect 45011 55886 48969 56173
rect 42892 55846 44724 55886
tri 44724 55846 44764 55886 sw
tri 45011 55846 45051 55886 ne
rect 45051 55870 48969 55886
tri 48969 55870 49280 56181 sw
tri 49280 55870 49591 56181 ne
rect 49591 55970 53455 56181
tri 53455 55970 53740 56255 sw
tri 53740 55970 54025 56255 ne
rect 54025 56160 55531 56255
tri 55531 56160 55815 56444 sw
tri 55815 56160 56099 56444 ne
rect 56099 56160 57791 56444
tri 57791 56160 58079 56448 sw
tri 58079 56160 58367 56448 ne
rect 58367 56352 59985 56448
tri 59985 56352 60155 56522 sw
tri 60271 56352 60441 56522 ne
rect 60441 56434 62056 56522
tri 62056 56434 62339 56717 sw
tri 62339 56434 62622 56717 ne
rect 62622 56434 70613 56717
rect 60441 56352 62339 56434
rect 58367 56160 60155 56352
rect 54025 55970 55815 56160
rect 49591 55870 53740 55970
rect 45051 55846 49280 55870
rect 42892 55738 44764 55846
rect 40799 55559 42600 55738
rect 36400 55421 40506 55559
tri 36400 55324 36497 55421 ne
rect 36497 55324 40506 55421
tri 36200 55124 36400 55324 sw
tri 36497 55124 36697 55324 ne
rect 36697 55266 40506 55324
tri 40506 55266 40799 55559 sw
tri 40799 55266 41092 55559 ne
rect 41092 55446 42600 55559
tri 42600 55446 42892 55738 sw
tri 42892 55446 43184 55738 ne
rect 43184 55559 44764 55738
tri 44764 55559 45051 55846 sw
tri 45051 55559 45338 55846 ne
rect 45338 55559 49280 55846
tri 49280 55559 49591 55870 sw
tri 49591 55559 49902 55870 ne
rect 49902 55685 53740 55870
tri 53740 55685 54025 55970 sw
tri 54025 55685 54310 55970 ne
rect 54310 55876 55815 55970
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 56068 58079 56160
tri 58079 56068 58171 56160 sw
tri 58367 56068 58459 56160 ne
rect 58459 56068 60155 56160
rect 56383 55876 58171 56068
rect 54310 55685 56099 55876
rect 49902 55559 54025 55685
rect 43184 55446 45051 55559
rect 41092 55266 42892 55446
rect 36697 55153 40799 55266
tri 40799 55153 40912 55266 sw
tri 41092 55153 41205 55266 ne
rect 41205 55154 42892 55266
tri 42892 55154 43184 55446 sw
tri 43184 55154 43476 55446 ne
rect 43476 55272 45051 55446
tri 45051 55272 45338 55559 sw
tri 45338 55272 45625 55559 ne
rect 45625 55272 49591 55559
rect 43476 55154 45338 55272
rect 41205 55153 43184 55154
rect 36697 55124 40912 55153
rect 33200 54827 36400 55124
tri 36400 54827 36697 55124 sw
tri 36697 54827 36994 55124 ne
rect 36994 54860 40912 55124
tri 40912 54860 41205 55153 sw
tri 41205 54860 41498 55153 ne
rect 41498 55064 43184 55153
tri 43184 55064 43274 55154 sw
tri 43476 55064 43566 55154 ne
rect 43566 55064 45338 55154
rect 41498 54860 43274 55064
rect 36994 54827 41205 54860
rect 33200 54674 36697 54827
tri 36697 54674 36850 54827 sw
tri 36994 54674 37147 54827 ne
rect 37147 54674 41205 54827
rect 33200 54377 36850 54674
tri 36850 54377 37147 54674 sw
tri 37147 54377 37444 54674 ne
rect 37444 54567 41205 54674
tri 41205 54567 41498 54860 sw
tri 41498 54567 41791 54860 ne
rect 41791 54772 43274 54860
tri 43274 54772 43566 55064 sw
tri 43566 54772 43858 55064 ne
rect 43858 55054 45338 55064
tri 45338 55054 45556 55272 sw
tri 45625 55054 45843 55272 ne
rect 45843 55248 49591 55272
tri 49591 55248 49902 55559 sw
tri 49902 55248 50213 55559 ne
rect 50213 55415 54025 55559
tri 54025 55415 54295 55685 sw
tri 54310 55415 54580 55685 ne
rect 54580 55592 56099 55685
tri 56099 55592 56383 55876 sw
tri 56383 55592 56667 55876 ne
rect 56667 55780 58171 55876
tri 58171 55780 58459 56068 sw
tri 58459 55780 58747 56068 ne
rect 58747 56066 60155 56068
tri 60155 56066 60441 56352 sw
tri 60441 56066 60727 56352 ne
rect 60727 56166 62339 56352
tri 62339 56166 62607 56434 sw
tri 62622 56166 62890 56434 ne
rect 62890 56166 70613 56434
rect 60727 56066 62607 56166
rect 58747 55780 60441 56066
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 55883 62607 56066
tri 62607 55883 62890 56166 sw
tri 62890 55883 63173 56166 ne
rect 63173 55883 70613 56166
rect 61013 55780 62890 55883
rect 56667 55592 58459 55780
rect 54580 55415 56383 55592
rect 50213 55248 54295 55415
rect 45843 55120 49902 55248
tri 49902 55120 50030 55248 sw
tri 50213 55120 50341 55248 ne
rect 50341 55130 54295 55248
tri 54295 55130 54580 55415 sw
tri 54580 55130 54865 55415 ne
rect 54865 55308 56383 55415
tri 56383 55308 56667 55592 sw
tri 56667 55308 56951 55592 ne
rect 56951 55492 58459 55592
tri 58459 55492 58747 55780 sw
tri 58747 55492 59035 55780 ne
rect 59035 55686 60727 55780
tri 60727 55686 60821 55780 sw
tri 61013 55686 61107 55780 ne
rect 61107 55686 62890 55780
rect 59035 55492 60821 55686
rect 56951 55308 58747 55492
rect 54865 55130 56667 55308
rect 50341 55120 54580 55130
rect 45843 55054 50030 55120
rect 43858 54772 45556 55054
rect 41791 54567 43566 54772
rect 37444 54377 41498 54567
rect 33200 54080 37147 54377
tri 37147 54080 37444 54377 sw
tri 37444 54080 37741 54377 ne
rect 37741 54274 41498 54377
tri 41498 54274 41791 54567 sw
tri 41791 54274 42084 54567 ne
rect 42084 54480 43566 54567
tri 43566 54480 43858 54772 sw
tri 43858 54480 44150 54772 ne
rect 44150 54767 45556 54772
tri 45556 54767 45843 55054 sw
tri 45843 54767 46130 55054 ne
rect 46130 54809 50030 55054
tri 50030 54809 50341 55120 sw
tri 50341 54809 50652 55120 ne
rect 50652 54845 54580 55120
tri 54580 54845 54865 55130 sw
tri 54865 54845 55150 55130 ne
rect 55150 55128 56667 55130
tri 56667 55128 56847 55308 sw
tri 56951 55128 57131 55308 ne
rect 57131 55204 58747 55308
tri 58747 55204 59035 55492 sw
tri 59035 55204 59323 55492 ne
rect 59323 55400 60821 55492
tri 60821 55400 61107 55686 sw
tri 61107 55400 61393 55686 ne
rect 61393 55600 62890 55686
tri 62890 55600 63173 55883 sw
tri 63173 55600 63456 55883 ne
rect 63456 55710 70613 55883
rect 70669 55710 71000 56910
rect 63456 55600 71000 55710
rect 61393 55400 63173 55600
tri 63173 55400 63373 55600 sw
rect 59323 55204 61107 55400
rect 57131 55128 59035 55204
rect 55150 54845 56847 55128
rect 50652 54809 54865 54845
rect 46130 54767 50341 54809
rect 44150 54480 45843 54767
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54498 50341 54767
tri 50341 54498 50652 54809 sw
tri 50652 54498 50963 54809 ne
rect 50963 54560 54865 54809
tri 54865 54560 55150 54845 sw
tri 55150 54560 55435 54845 ne
rect 55435 54844 56847 54845
tri 56847 54844 57131 55128 sw
tri 57131 54844 57415 55128 ne
rect 57415 54916 59035 55128
tri 59035 54916 59323 55204 sw
tri 59323 54916 59611 55204 ne
rect 59611 55114 61107 55204
tri 61107 55114 61393 55400 sw
tri 61393 55114 61679 55400 ne
rect 61679 55302 71000 55400
rect 61679 55114 70613 55302
rect 59611 54916 61393 55114
rect 57415 54844 59323 54916
rect 55435 54560 57131 54844
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54756 59323 54844
tri 59323 54756 59483 54916 sw
tri 59611 54756 59771 54916 ne
rect 59771 54828 61393 54916
tri 61393 54828 61679 55114 sw
tri 61679 54828 61965 55114 ne
rect 61965 54828 70613 55114
rect 59771 54756 61679 54828
rect 57699 54560 59483 54756
rect 50963 54498 55150 54560
rect 46417 54480 50652 54498
rect 42084 54274 43858 54480
rect 37741 54080 41791 54274
tri 33200 53992 33288 54080 ne
rect 33288 53992 37444 54080
tri 33000 53792 33200 53992 sw
tri 33288 53792 33488 53992 ne
rect 33488 53792 37444 53992
rect 30000 53504 33200 53792
tri 33200 53504 33488 53792 sw
tri 33488 53504 33776 53792 ne
rect 33776 53783 37444 53792
tri 37444 53783 37741 54080 sw
tri 37741 53783 38038 54080 ne
rect 38038 53981 41791 54080
tri 41791 53981 42084 54274 sw
tri 42084 53981 42377 54274 ne
rect 42377 54188 43858 54274
tri 43858 54188 44150 54480 sw
tri 44150 54188 44442 54480 ne
rect 44442 54193 46130 54480
tri 46130 54193 46417 54480 sw
tri 46417 54193 46704 54480 ne
rect 46704 54193 50652 54480
rect 44442 54188 46417 54193
rect 42377 53981 44150 54188
rect 38038 53783 42084 53981
rect 33776 53673 37741 53783
tri 37741 53673 37851 53783 sw
tri 38038 53673 38148 53783 ne
rect 38148 53759 42084 53783
tri 42084 53759 42306 53981 sw
tri 42377 53759 42599 53981 ne
rect 42599 53896 44150 53981
tri 44150 53896 44442 54188 sw
tri 44442 53896 44734 54188 ne
rect 44734 53906 46417 54188
tri 46417 53906 46704 54193 sw
tri 46704 53906 46991 54193 ne
rect 46991 54187 50652 54193
tri 50652 54187 50963 54498 sw
tri 50963 54187 51274 54498 ne
rect 51274 54275 55150 54498
tri 55150 54275 55435 54560 sw
tri 55435 54275 55720 54560 ne
rect 55720 54464 57415 54560
tri 57415 54464 57511 54560 sw
tri 57699 54464 57795 54560 ne
rect 57795 54468 59483 54560
tri 59483 54468 59771 54756 sw
tri 59771 54468 60059 54756 ne
rect 60059 54572 61679 54756
tri 61679 54572 61935 54828 sw
tri 61965 54572 62221 54828 ne
rect 62221 54572 70613 54828
rect 60059 54468 61935 54572
rect 57795 54464 59771 54468
rect 55720 54275 57511 54464
rect 51274 54187 55435 54275
rect 46991 53906 50963 54187
rect 44734 53896 46704 53906
rect 42599 53759 44442 53896
rect 38148 53673 42306 53759
rect 33776 53504 37851 53673
rect 30000 53216 33488 53504
tri 33488 53216 33776 53504 sw
tri 33776 53216 34064 53504 ne
rect 34064 53376 37851 53504
tri 37851 53376 38148 53673 sw
tri 38148 53376 38445 53673 ne
rect 38445 53466 42306 53673
tri 42306 53466 42599 53759 sw
tri 42599 53466 42892 53759 ne
rect 42892 53604 44442 53759
tri 44442 53604 44734 53896 sw
tri 44734 53604 45026 53896 ne
rect 45026 53619 46704 53896
tri 46704 53619 46991 53906 sw
tri 46991 53619 47278 53906 ne
rect 47278 53876 50963 53906
tri 50963 53876 51274 54187 sw
tri 51274 53876 51585 54187 ne
rect 51585 53990 55435 54187
tri 55435 53990 55720 54275 sw
tri 55720 53990 56005 54275 ne
rect 56005 54180 57511 54275
tri 57511 54180 57795 54464 sw
tri 57795 54180 58079 54464 ne
rect 58079 54180 59771 54464
tri 59771 54180 60059 54468 sw
tri 60059 54180 60347 54468 ne
rect 60347 54286 61935 54468
tri 61935 54286 62221 54572 sw
tri 62221 54286 62507 54572 ne
rect 62507 54286 70613 54572
rect 60347 54180 62221 54286
rect 56005 53990 57795 54180
rect 51585 53876 55720 53990
rect 47278 53619 51274 53876
rect 45026 53604 46991 53619
rect 42892 53466 44734 53604
rect 38445 53376 42599 53466
rect 34064 53216 38148 53376
rect 30000 52928 33776 53216
tri 33776 52928 34064 53216 sw
tri 34064 52928 34352 53216 ne
rect 34352 53079 38148 53216
tri 38148 53079 38445 53376 sw
tri 38445 53079 38742 53376 ne
rect 38742 53173 42599 53376
tri 42599 53173 42892 53466 sw
tri 42892 53173 43185 53466 ne
rect 43185 53464 44734 53466
tri 44734 53464 44874 53604 sw
tri 45026 53464 45166 53604 ne
rect 45166 53464 46991 53604
rect 43185 53173 44874 53464
rect 38742 53079 42892 53173
rect 34352 52928 38445 53079
rect 30000 52748 34064 52928
tri 30000 52654 30094 52748 ne
rect 30094 52654 34064 52748
tri 29800 52454 30000 52654 sw
tri 30094 52454 30294 52654 ne
rect 30294 52640 34064 52654
tri 34064 52640 34352 52928 sw
tri 34352 52640 34640 52928 ne
rect 34640 52782 38445 52928
tri 38445 52782 38742 53079 sw
tri 38742 52782 39039 53079 ne
rect 39039 52880 42892 53079
tri 42892 52880 43185 53173 sw
tri 43185 52880 43478 53173 ne
rect 43478 53172 44874 53173
tri 44874 53172 45166 53464 sw
tri 45166 53172 45458 53464 ne
rect 45458 53454 46991 53464
tri 46991 53454 47156 53619 sw
tri 47278 53454 47443 53619 ne
rect 47443 53565 51274 53619
tri 51274 53565 51585 53876 sw
tri 51585 53565 51896 53876 ne
rect 51896 53705 55720 53876
tri 55720 53705 56005 53990 sw
tri 56005 53705 56290 53990 ne
rect 56290 53896 57795 53990
tri 57795 53896 58079 54180 sw
tri 58079 53896 58363 54180 ne
rect 58363 54088 60059 54180
tri 60059 54088 60151 54180 sw
tri 60347 54088 60439 54180 ne
rect 60439 54088 62221 54180
rect 58363 53896 60151 54088
rect 56290 53705 58079 53896
rect 51896 53565 56005 53705
rect 47443 53454 51585 53565
rect 45458 53172 47156 53454
rect 43478 52880 45166 53172
tri 45166 52880 45458 53172 sw
tri 45458 52880 45750 53172 ne
rect 45750 53167 47156 53172
tri 47156 53167 47443 53454 sw
tri 47443 53167 47730 53454 ne
rect 47730 53254 51585 53454
tri 51585 53254 51896 53565 sw
tri 51896 53254 52207 53565 ne
rect 52207 53435 56005 53565
tri 56005 53435 56275 53705 sw
tri 56290 53435 56560 53705 ne
rect 56560 53612 58079 53705
tri 58079 53612 58363 53896 sw
tri 58363 53612 58647 53896 ne
rect 58647 53800 60151 53896
tri 60151 53800 60439 54088 sw
tri 60439 53800 60727 54088 ne
rect 60727 54000 62221 54088
tri 62221 54000 62507 54286 sw
tri 62507 54000 62793 54286 ne
rect 62793 54102 70613 54286
rect 70669 54102 71000 55302
rect 62793 54000 71000 54102
rect 60727 53800 62507 54000
tri 62507 53800 62707 54000 sw
rect 58647 53612 60439 53800
rect 56560 53435 58363 53612
rect 52207 53254 56275 53435
rect 47730 53167 51896 53254
rect 45750 52880 47443 53167
tri 47443 52880 47730 53167 sw
tri 47730 52880 48017 53167 ne
rect 48017 52943 51896 53167
tri 51896 52943 52207 53254 sw
tri 52207 52943 52518 53254 ne
rect 52518 53150 56275 53254
tri 56275 53150 56560 53435 sw
tri 56560 53150 56845 53435 ne
rect 56845 53328 58363 53435
tri 58363 53328 58647 53612 sw
tri 58647 53328 58931 53612 ne
rect 58931 53512 60439 53612
tri 60439 53512 60727 53800 sw
tri 60727 53512 61015 53800 ne
rect 61015 53722 71000 53800
rect 61015 53512 70613 53722
rect 58931 53328 60727 53512
rect 56845 53150 58647 53328
rect 52518 52943 56560 53150
rect 48017 52880 52207 52943
rect 39039 52782 43185 52880
rect 34640 52640 38742 52782
rect 30294 52454 34352 52640
rect 26800 52160 30000 52454
tri 30000 52160 30294 52454 sw
tri 30294 52160 30588 52454 ne
rect 30588 52372 34352 52454
tri 34352 52372 34620 52640 sw
tri 34640 52372 34908 52640 ne
rect 34908 52485 38742 52640
tri 38742 52485 39039 52782 sw
tri 39039 52485 39336 52782 ne
rect 39336 52587 43185 52782
tri 43185 52587 43478 52880 sw
tri 43478 52587 43771 52880 ne
rect 43771 52792 45458 52880
tri 45458 52792 45546 52880 sw
tri 45750 52792 45838 52880 ne
rect 45838 52792 47730 52880
rect 43771 52587 45546 52792
rect 39336 52485 43478 52587
rect 34908 52372 39039 52485
rect 30588 52160 34620 52372
rect 26800 51998 30294 52160
tri 30294 51998 30456 52160 sw
tri 30588 51998 30750 52160 ne
rect 30750 52084 34620 52160
tri 34620 52084 34908 52372 sw
tri 34908 52084 35196 52372 ne
rect 35196 52188 39039 52372
tri 39039 52188 39336 52485 sw
tri 39336 52188 39633 52485 ne
rect 39633 52294 43478 52485
tri 43478 52294 43771 52587 sw
tri 43771 52294 44064 52587 ne
rect 44064 52500 45546 52587
tri 45546 52500 45838 52792 sw
tri 45838 52500 46130 52792 ne
rect 46130 52787 47730 52792
tri 47730 52787 47823 52880 sw
tri 48017 52787 48110 52880 ne
rect 48110 52861 52207 52880
tri 52207 52861 52289 52943 sw
tri 52518 52861 52600 52943 ne
rect 52600 52865 56560 52943
tri 56560 52865 56845 53150 sw
tri 56845 52865 57130 53150 ne
rect 57130 53148 58647 53150
tri 58647 53148 58827 53328 sw
tri 58931 53148 59111 53328 ne
rect 59111 53224 60727 53328
tri 60727 53224 61015 53512 sw
tri 61015 53224 61303 53512 ne
rect 61303 53224 70613 53512
rect 59111 53148 61015 53224
rect 57130 52865 58827 53148
rect 52600 52861 56845 52865
rect 48110 52787 52289 52861
rect 46130 52500 47823 52787
tri 47823 52500 48110 52787 sw
tri 48110 52500 48397 52787 ne
rect 48397 52550 52289 52787
tri 52289 52550 52600 52861 sw
tri 52600 52550 52911 52861 ne
rect 52911 52580 56845 52861
tri 56845 52580 57130 52865 sw
tri 57130 52580 57415 52865 ne
rect 57415 52864 58827 52865
tri 58827 52864 59111 53148 sw
tri 59111 52864 59395 53148 ne
rect 59395 52976 61015 53148
tri 61015 52976 61263 53224 sw
tri 61303 52976 61551 53224 ne
rect 61551 52976 70613 53224
rect 59395 52864 61263 52976
rect 57415 52580 59111 52864
tri 59111 52580 59395 52864 sw
tri 59395 52580 59679 52864 ne
rect 59679 52688 61263 52864
tri 61263 52688 61551 52976 sw
tri 61551 52688 61839 52976 ne
rect 61839 52688 70613 52976
rect 59679 52580 61551 52688
rect 52911 52550 57130 52580
rect 48397 52500 52600 52550
rect 44064 52294 45838 52500
rect 39633 52188 43771 52294
rect 35196 52084 39336 52188
rect 30750 51998 34908 52084
rect 26800 51704 30456 51998
tri 30456 51704 30750 51998 sw
tri 30750 51704 31044 51998 ne
rect 31044 51796 34908 51998
tri 34908 51796 35196 52084 sw
tri 35196 51796 35484 52084 ne
rect 35484 51891 39336 52084
tri 39336 51891 39633 52188 sw
tri 39633 51891 39930 52188 ne
rect 39930 52001 43771 52188
tri 43771 52001 44064 52294 sw
tri 44064 52001 44357 52294 ne
rect 44357 52208 45838 52294
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52213 48110 52500
tri 48110 52213 48397 52500 sw
tri 48397 52213 48684 52500 ne
rect 48684 52239 52600 52500
tri 52600 52239 52911 52550 sw
tri 52911 52239 53222 52550 ne
rect 53222 52295 57130 52550
tri 57130 52295 57415 52580 sw
tri 57415 52295 57700 52580 ne
rect 57700 52484 59395 52580
tri 59395 52484 59491 52580 sw
tri 59679 52484 59775 52580 ne
rect 59775 52484 61551 52580
rect 57700 52295 59491 52484
rect 53222 52239 57415 52295
rect 48684 52213 52911 52239
rect 46422 52208 48397 52213
rect 44357 52001 46130 52208
rect 39930 51891 44064 52001
rect 35484 51796 39633 51891
rect 31044 51704 35196 51796
rect 26800 51410 30750 51704
tri 30750 51410 31044 51704 sw
tri 31044 51410 31338 51704 ne
rect 31338 51508 35196 51704
tri 35196 51508 35484 51796 sw
tri 35484 51508 35772 51796 ne
rect 35772 51661 39633 51796
tri 39633 51661 39863 51891 sw
tri 39930 51661 40160 51891 ne
rect 40160 51779 44064 51891
tri 44064 51779 44286 52001 sw
tri 44357 51779 44579 52001 ne
rect 44579 51916 46130 52001
tri 46130 51916 46422 52208 sw
tri 46422 51916 46714 52208 ne
rect 46714 51926 48397 52208
tri 48397 51926 48684 52213 sw
tri 48684 51926 48971 52213 ne
rect 48971 51928 52911 52213
tri 52911 51928 53222 52239 sw
tri 53222 51928 53533 52239 ne
rect 53533 52010 57415 52239
tri 57415 52010 57700 52295 sw
tri 57700 52010 57985 52295 ne
rect 57985 52200 59491 52295
tri 59491 52200 59775 52484 sw
tri 59775 52200 60059 52484 ne
rect 60059 52400 61551 52484
tri 61551 52400 61839 52688 sw
tri 61839 52400 62127 52688 ne
rect 62127 52522 70613 52688
rect 70669 52522 71000 53722
rect 62127 52400 71000 52522
rect 60059 52200 61839 52400
tri 61839 52200 62039 52400 sw
rect 57985 52010 59775 52200
rect 53533 51928 57700 52010
rect 48971 51926 53222 51928
rect 46714 51916 48684 51926
rect 44579 51779 46422 51916
rect 40160 51661 44286 51779
rect 35772 51508 39863 51661
rect 31338 51410 35484 51508
tri 26800 51320 26890 51410 ne
rect 26890 51320 31044 51410
tri 26600 51220 26700 51320 sw
tri 26890 51220 26990 51320 ne
rect 26990 51220 31044 51320
tri 31044 51220 31234 51410 sw
tri 31338 51220 31528 51410 ne
rect 31528 51220 35484 51410
tri 35484 51220 35772 51508 sw
tri 35772 51220 36060 51508 ne
rect 36060 51364 39863 51508
tri 39863 51364 40160 51661 sw
tri 40160 51364 40457 51661 ne
rect 40457 51486 44286 51661
tri 44286 51486 44579 51779 sw
tri 44579 51486 44872 51779 ne
rect 44872 51624 46422 51779
tri 46422 51624 46714 51916 sw
tri 46714 51624 47006 51916 ne
rect 47006 51880 48684 51916
tri 48684 51880 48730 51926 sw
tri 48971 51880 49017 51926 ne
rect 49017 51880 53222 51926
rect 47006 51624 48730 51880
rect 44872 51486 46714 51624
rect 40457 51364 44579 51486
rect 36060 51220 40160 51364
rect 25200 50930 26700 51220
tri 26700 50930 26990 51220 sw
tri 26990 50930 27280 51220 ne
rect 27280 50930 31234 51220
rect 25200 50740 26990 50930
tri 25200 50651 25289 50740 ne
rect 25289 50651 26990 50740
tri 25000 50451 25200 50651 sw
tri 25289 50451 25489 50651 ne
rect 25489 50650 26990 50651
tri 26990 50650 27270 50930 sw
tri 27280 50650 27560 50930 ne
rect 27560 50926 31234 50930
tri 31234 50926 31528 51220 sw
tri 31528 50926 31822 51220 ne
rect 31822 50932 35772 51220
tri 35772 50932 36060 51220 sw
tri 36060 50932 36348 51220 ne
rect 36348 51067 40160 51220
tri 40160 51067 40457 51364 sw
tri 40457 51067 40754 51364 ne
rect 40754 51193 44579 51364
tri 44579 51193 44872 51486 sw
tri 44872 51193 45165 51486 ne
rect 45165 51484 46714 51486
tri 46714 51484 46854 51624 sw
tri 47006 51484 47146 51624 ne
rect 47146 51593 48730 51624
tri 48730 51593 49017 51880 sw
tri 49017 51593 49304 51880 ne
rect 49304 51617 53222 51880
tri 53222 51617 53533 51928 sw
tri 53533 51617 53844 51928 ne
rect 53844 51725 57700 51928
tri 57700 51725 57985 52010 sw
tri 57985 51725 58270 52010 ne
rect 58270 51916 59775 52010
tri 59775 51916 60059 52200 sw
tri 60059 51916 60343 52200 ne
rect 60343 51916 71000 52200
rect 58270 51725 60059 51916
rect 53844 51617 57985 51725
rect 49304 51593 53533 51617
rect 47146 51484 49017 51593
rect 45165 51193 46854 51484
rect 40754 51067 44872 51193
rect 36348 50932 40457 51067
rect 31822 50926 36060 50932
rect 27560 50650 31528 50926
rect 25489 50451 27270 50650
rect 23600 50360 25200 50451
tri 25200 50360 25291 50451 sw
tri 25489 50360 25580 50451 ne
rect 25580 50360 27270 50451
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50632 31528 50650
tri 31528 50632 31822 50926 sw
tri 31822 50632 32116 50926 ne
rect 32116 50752 36060 50926
tri 36060 50752 36240 50932 sw
tri 36348 50752 36528 50932 ne
rect 36528 50770 40457 50932
tri 40457 50770 40754 51067 sw
tri 40754 50770 41051 51067 ne
rect 41051 50900 44872 51067
tri 44872 50900 45165 51193 sw
tri 45165 50900 45458 51193 ne
rect 45458 51192 46854 51193
tri 46854 51192 47146 51484 sw
tri 47146 51192 47438 51484 ne
rect 47438 51306 49017 51484
tri 49017 51306 49304 51593 sw
tri 49304 51306 49591 51593 ne
rect 49591 51306 53533 51593
tri 53533 51306 53844 51617 sw
tri 53844 51306 54155 51617 ne
rect 54155 51455 57985 51617
tri 57985 51455 58255 51725 sw
tri 58270 51455 58540 51725 ne
rect 58540 51632 60059 51725
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58540 51455 60343 51632
rect 54155 51306 58255 51455
rect 47438 51192 49304 51306
rect 45458 50900 47146 51192
tri 47146 50900 47438 51192 sw
tri 47438 50900 47730 51192 ne
rect 47730 51019 49304 51192
tri 49304 51019 49591 51306 sw
tri 49591 51019 49878 51306 ne
rect 49878 51019 53844 51306
rect 47730 50900 49591 51019
rect 41051 50770 45165 50900
rect 36528 50752 40754 50770
rect 32116 50632 36240 50752
rect 27850 50360 31822 50632
rect 23600 50071 25291 50360
tri 25291 50071 25580 50360 sw
tri 25580 50071 25869 50360 ne
rect 25869 50071 27560 50360
tri 23600 49974 23697 50071 ne
rect 23697 49974 25580 50071
tri 23400 49774 23600 49974 sw
tri 23697 49774 23897 49974 ne
rect 23897 49918 25580 49974
tri 25580 49918 25733 50071 sw
tri 25869 49918 26022 50071 ne
rect 26022 50070 27560 50071
tri 27560 50070 27850 50360 sw
tri 27850 50070 28140 50360 ne
rect 28140 50338 31822 50360
tri 31822 50338 32116 50632 sw
tri 32116 50338 32410 50632 ne
rect 32410 50464 36240 50632
tri 36240 50464 36528 50752 sw
tri 36528 50464 36816 50752 ne
rect 36816 50473 40754 50752
tri 40754 50473 41051 50770 sw
tri 41051 50473 41348 50770 ne
rect 41348 50607 45165 50770
tri 45165 50607 45458 50900 sw
tri 45458 50607 45751 50900 ne
rect 45751 50812 47438 50900
tri 47438 50812 47526 50900 sw
tri 47730 50812 47818 50900 ne
rect 47818 50812 49591 50900
rect 45751 50607 47526 50812
rect 41348 50473 45458 50607
rect 36816 50464 41051 50473
rect 32410 50338 36528 50464
rect 28140 50070 32116 50338
rect 26022 49918 27850 50070
rect 23897 49774 25733 49918
rect 20400 49477 23600 49774
tri 23600 49477 23897 49774 sw
tri 23897 49477 24194 49774 ne
rect 24194 49629 25733 49774
tri 25733 49629 26022 49918 sw
tri 26022 49629 26311 49918 ne
rect 26311 49780 27850 49918
tri 27850 49780 28140 50070 sw
tri 28140 49780 28430 50070 ne
rect 28430 50044 32116 50070
tri 32116 50044 32410 50338 sw
tri 32410 50044 32704 50338 ne
rect 32704 50176 36528 50338
tri 36528 50176 36816 50464 sw
tri 36816 50176 37104 50464 ne
rect 37104 50176 41051 50464
tri 41051 50176 41348 50473 sw
tri 41348 50176 41645 50473 ne
rect 41645 50314 45458 50473
tri 45458 50314 45751 50607 sw
tri 45751 50314 46044 50607 ne
rect 46044 50520 47526 50607
tri 47526 50520 47818 50812 sw
tri 47818 50520 48110 50812 ne
rect 48110 50807 49591 50812
tri 49591 50807 49803 51019 sw
tri 49878 50807 50090 51019 ne
rect 50090 50995 53844 51019
tri 53844 50995 54155 51306 sw
tri 54155 50995 54466 51306 ne
rect 54466 51170 58255 51306
tri 58255 51170 58540 51455 sw
tri 58540 51170 58825 51455 ne
rect 58825 51368 60343 51455
tri 60343 51368 60607 51632 sw
tri 60627 51368 60891 51632 ne
rect 60891 51368 71000 51632
rect 58825 51170 60607 51368
rect 54466 50995 58540 51170
rect 50090 50871 54155 50995
tri 54155 50871 54279 50995 sw
tri 54466 50871 54590 50995 ne
rect 54590 50885 58540 50995
tri 58540 50885 58825 51170 sw
tri 58825 50885 59110 51170 ne
rect 59110 51084 60607 51170
tri 60607 51084 60891 51368 sw
tri 60891 51084 61175 51368 ne
rect 61175 51084 71000 51368
rect 59110 50885 60891 51084
rect 54590 50871 58825 50885
rect 50090 50807 54279 50871
rect 48110 50520 49803 50807
tri 49803 50520 50090 50807 sw
tri 50090 50520 50377 50807 ne
rect 50377 50560 54279 50807
tri 54279 50560 54590 50871 sw
tri 54590 50560 54901 50871 ne
rect 54901 50600 58825 50871
tri 58825 50600 59110 50885 sw
tri 59110 50600 59395 50885 ne
rect 59395 50800 60891 50885
tri 60891 50800 61175 51084 sw
tri 61175 50800 61459 51084 ne
rect 61459 50800 71000 51084
rect 59395 50600 61175 50800
tri 61175 50600 61375 50800 sw
rect 54901 50560 59110 50600
rect 50377 50520 54590 50560
rect 46044 50314 47818 50520
rect 41645 50176 45751 50314
rect 32704 50044 36816 50176
rect 28430 49780 32410 50044
rect 26311 49629 28140 49780
rect 24194 49477 26022 49629
rect 20400 49354 23897 49477
tri 23897 49354 24020 49477 sw
tri 24194 49354 24317 49477 ne
rect 24317 49354 26022 49477
rect 20400 49057 24020 49354
tri 24020 49057 24317 49354 sw
tri 24317 49057 24614 49354 ne
rect 24614 49340 26022 49354
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49490 28140 49629
tri 28140 49490 28430 49780 sw
tri 28430 49490 28720 49780 ne
rect 28720 49750 32410 49780
tri 32410 49750 32704 50044 sw
tri 32704 49750 32998 50044 ne
rect 32998 49888 36816 50044
tri 36816 49888 37104 50176 sw
tri 37104 49888 37392 50176 ne
rect 37392 49888 41348 50176
rect 32998 49750 37104 49888
rect 28720 49490 32704 49750
tri 32704 49490 32964 49750 sw
tri 32998 49490 33258 49750 ne
rect 33258 49600 37104 49750
tri 37104 49600 37392 49888 sw
tri 37392 49600 37680 49888 ne
rect 37680 49879 41348 49888
tri 41348 49879 41645 50176 sw
tri 41645 49879 41942 50176 ne
rect 41942 50021 45751 50176
tri 45751 50021 46044 50314 sw
tri 46044 50021 46337 50314 ne
rect 46337 50228 47818 50314
tri 47818 50228 48110 50520 sw
tri 48110 50228 48402 50520 ne
rect 48402 50249 50090 50520
tri 50090 50249 50361 50520 sw
tri 50377 50249 50648 50520 ne
rect 50648 50249 54590 50520
tri 54590 50249 54901 50560 sw
tri 54901 50249 55212 50560 ne
rect 55212 50315 59110 50560
tri 59110 50315 59395 50600 sw
tri 59395 50315 59680 50600 ne
rect 59680 50315 71000 50600
rect 55212 50249 59395 50315
rect 48402 50228 50361 50249
rect 46337 50021 48110 50228
rect 41942 49879 46044 50021
rect 37680 49726 41645 49879
tri 41645 49726 41798 49879 sw
tri 41942 49726 42095 49879 ne
rect 42095 49799 46044 49879
tri 46044 49799 46266 50021 sw
tri 46337 49799 46559 50021 ne
rect 46559 49936 48110 50021
tri 48110 49936 48402 50228 sw
tri 48402 49936 48694 50228 ne
rect 48694 49962 50361 50228
tri 50361 49962 50648 50249 sw
tri 50648 49962 50935 50249 ne
rect 50935 49962 54901 50249
rect 48694 49936 50648 49962
rect 46559 49799 48402 49936
rect 42095 49726 46266 49799
rect 37680 49600 41798 49726
rect 33258 49490 37392 49600
rect 26600 49340 28430 49490
tri 28430 49340 28580 49490 sw
tri 28720 49340 28870 49490 ne
rect 28870 49340 32964 49490
rect 24614 49057 26311 49340
rect 20400 48760 24317 49057
tri 24317 48760 24614 49057 sw
tri 24614 48760 24911 49057 ne
rect 24911 49051 26311 49057
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49051 28580 49340
rect 24911 48762 26600 49051
tri 26600 48762 26889 49051 sw
tri 26889 48762 27178 49051 ne
rect 27178 49050 28580 49051
tri 28580 49050 28870 49340 sw
tri 28870 49050 29160 49340 ne
rect 29160 49196 32964 49340
tri 32964 49196 33258 49490 sw
tri 33258 49196 33552 49490 ne
rect 33552 49312 37392 49490
tri 37392 49312 37680 49600 sw
tri 37680 49312 37968 49600 ne
rect 37968 49429 41798 49600
tri 41798 49429 42095 49726 sw
tri 42095 49429 42392 49726 ne
rect 42392 49506 46266 49726
tri 46266 49506 46559 49799 sw
tri 46559 49506 46852 49799 ne
rect 46852 49644 48402 49799
tri 48402 49644 48694 49936 sw
tri 48694 49644 48986 49936 ne
rect 48986 49675 50648 49936
tri 50648 49675 50935 49962 sw
tri 50935 49675 51222 49962 ne
rect 51222 49938 54901 49962
tri 54901 49938 55212 50249 sw
tri 55212 49938 55523 50249 ne
rect 55523 50030 59395 50249
tri 59395 50030 59680 50315 sw
tri 59680 50030 59965 50315 ne
rect 59965 50030 71000 50315
rect 55523 49938 59680 50030
rect 51222 49675 55212 49938
rect 48986 49644 50935 49675
rect 46852 49506 48694 49644
rect 42392 49429 46559 49506
rect 37968 49312 42095 49429
rect 33552 49196 37680 49312
rect 29160 49050 33258 49196
rect 27178 48762 28870 49050
rect 24911 48760 26889 48762
rect 20400 48730 24614 48760
tri 20400 48648 20482 48730 ne
rect 20482 48671 24614 48730
tri 24614 48671 24703 48760 sw
tri 24911 48671 25000 48760 ne
rect 25000 48671 26889 48760
rect 20482 48648 24703 48671
tri 20200 48448 20400 48648 sw
tri 20482 48448 20682 48648 ne
rect 20682 48448 24703 48648
rect 17200 48166 20400 48448
tri 20400 48166 20682 48448 sw
tri 20682 48166 20964 48448 ne
rect 20964 48374 24703 48448
tri 24703 48374 25000 48671 sw
tri 25000 48374 25297 48671 ne
rect 25297 48669 26889 48671
tri 26889 48669 26982 48762 sw
tri 27178 48669 27271 48762 ne
rect 27271 48760 28870 48762
tri 28870 48760 29160 49050 sw
tri 29160 48760 29450 49050 ne
rect 29450 48902 33258 49050
tri 33258 48902 33552 49196 sw
tri 33552 48902 33846 49196 ne
rect 33846 49024 37680 49196
tri 37680 49024 37968 49312 sw
tri 37968 49024 38256 49312 ne
rect 38256 49132 42095 49312
tri 42095 49132 42392 49429 sw
tri 42392 49132 42689 49429 ne
rect 42689 49213 46559 49429
tri 46559 49213 46852 49506 sw
tri 46852 49213 47145 49506 ne
rect 47145 49504 48694 49506
tri 48694 49504 48834 49644 sw
tri 48986 49504 49126 49644 ne
rect 49126 49504 50935 49644
rect 47145 49213 48834 49504
rect 42689 49132 46852 49213
rect 38256 49024 42392 49132
rect 33846 48902 37968 49024
rect 29450 48760 33552 48902
rect 27271 48670 29160 48760
tri 29160 48670 29250 48760 sw
tri 29450 48670 29540 48760 ne
rect 29540 48670 33552 48760
rect 27271 48669 29250 48670
rect 25297 48380 26982 48669
tri 26982 48380 27271 48669 sw
tri 27271 48380 27560 48669 ne
rect 27560 48380 29250 48669
tri 29250 48380 29540 48670 sw
tri 29540 48380 29830 48670 ne
rect 29830 48608 33552 48670
tri 33552 48608 33846 48902 sw
tri 33846 48608 34140 48902 ne
rect 34140 48736 37968 48902
tri 37968 48736 38256 49024 sw
tri 38256 48736 38544 49024 ne
rect 38544 48835 42392 49024
tri 42392 48835 42689 49132 sw
tri 42689 48835 42986 49132 ne
rect 42986 48920 46852 49132
tri 46852 48920 47145 49213 sw
tri 47145 48920 47438 49213 ne
rect 47438 49212 48834 49213
tri 48834 49212 49126 49504 sw
tri 49126 49212 49418 49504 ne
rect 49418 49494 50935 49504
tri 50935 49494 51116 49675 sw
tri 51222 49494 51403 49675 ne
rect 51403 49627 55212 49675
tri 55212 49627 55523 49938 sw
tri 55523 49627 55834 49938 ne
rect 55834 49770 59680 49938
tri 59680 49770 59940 50030 sw
tri 59965 49770 60225 50030 ne
rect 60225 49770 71000 50030
rect 55834 49627 59940 49770
rect 51403 49494 55523 49627
rect 49418 49212 51116 49494
rect 47438 48920 49126 49212
tri 49126 48920 49418 49212 sw
tri 49418 48920 49710 49212 ne
rect 49710 49207 51116 49212
tri 51116 49207 51403 49494 sw
tri 51403 49207 51690 49494 ne
rect 51690 49316 55523 49494
tri 55523 49316 55834 49627 sw
tri 55834 49316 56145 49627 ne
rect 56145 49485 59940 49627
tri 59940 49485 60225 49770 sw
tri 60225 49485 60510 49770 ne
rect 60510 49485 71000 49770
rect 56145 49316 60225 49485
rect 51690 49207 55834 49316
rect 49710 48920 51403 49207
tri 51403 48920 51690 49207 sw
tri 51690 48920 51977 49207 ne
rect 51977 49005 55834 49207
tri 55834 49005 56145 49316 sw
tri 56145 49005 56456 49316 ne
rect 56456 49200 60225 49316
tri 60225 49200 60510 49485 sw
tri 60510 49200 60795 49485 ne
rect 60795 49200 71000 49485
rect 56456 49005 60510 49200
rect 51977 48920 56145 49005
rect 42986 48835 47145 48920
rect 38544 48736 42689 48835
rect 34140 48608 38256 48736
rect 29830 48380 33846 48608
rect 25297 48374 27271 48380
rect 20964 48166 25000 48374
rect 17200 47884 20682 48166
tri 20682 47884 20964 48166 sw
tri 20964 47884 21246 48166 ne
rect 21246 48077 25000 48166
tri 25000 48077 25297 48374 sw
tri 25297 48077 25594 48374 ne
rect 25594 48091 27271 48374
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48091 29540 48380
rect 25594 48077 27560 48091
rect 21246 47884 25297 48077
rect 17200 47602 20964 47884
tri 20964 47602 21246 47884 sw
tri 21246 47602 21528 47884 ne
rect 21528 47780 25297 47884
tri 25297 47780 25594 48077 sw
tri 25594 47780 25891 48077 ne
rect 25891 47802 27560 48077
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48090 29540 48091
tri 29540 48090 29830 48380 sw
tri 29830 48090 30120 48380 ne
rect 30120 48314 33846 48380
tri 33846 48314 34140 48608 sw
tri 34140 48314 34434 48608 ne
rect 34434 48448 38256 48608
tri 38256 48448 38544 48736 sw
tri 38544 48448 38832 48736 ne
rect 38832 48538 42689 48736
tri 42689 48538 42986 48835 sw
tri 42986 48538 43283 48835 ne
rect 43283 48627 47145 48835
tri 47145 48627 47438 48920 sw
tri 47438 48627 47731 48920 ne
rect 47731 48832 49418 48920
tri 49418 48832 49506 48920 sw
tri 49710 48832 49798 48920 ne
rect 49798 48832 51690 48920
rect 47731 48627 49506 48832
rect 43283 48538 47438 48627
rect 38832 48448 42986 48538
rect 34434 48416 38544 48448
tri 38544 48416 38576 48448 sw
tri 38832 48416 38864 48448 ne
rect 38864 48416 42986 48448
rect 34434 48314 38576 48416
rect 30120 48090 34140 48314
rect 28138 48020 29830 48090
tri 29830 48020 29900 48090 sw
tri 30120 48020 30190 48090 ne
rect 30190 48020 34140 48090
tri 34140 48020 34434 48314 sw
tri 34434 48020 34728 48314 ne
rect 34728 48128 38576 48314
tri 38576 48128 38864 48416 sw
tri 38864 48128 39152 48416 ne
rect 39152 48241 42986 48416
tri 42986 48241 43283 48538 sw
tri 43283 48241 43580 48538 ne
rect 43580 48334 47438 48538
tri 47438 48334 47731 48627 sw
tri 47731 48334 48024 48627 ne
rect 48024 48540 49506 48627
tri 49506 48540 49798 48832 sw
tri 49798 48540 50090 48832 ne
rect 50090 48827 51690 48832
tri 51690 48827 51783 48920 sw
tri 51977 48827 52070 48920 ne
rect 52070 48827 56145 48920
rect 50090 48540 51783 48827
tri 51783 48540 52070 48827 sw
tri 52070 48540 52357 48827 ne
rect 52357 48694 56145 48827
tri 56145 48694 56456 49005 sw
tri 56456 48694 56767 49005 ne
rect 56767 49000 60510 49005
tri 60510 49000 60710 49200 sw
rect 56767 48694 71000 49000
rect 52357 48608 56456 48694
tri 56456 48608 56542 48694 sw
tri 56767 48608 56853 48694 ne
rect 56853 48608 71000 48694
rect 52357 48540 56542 48608
rect 48024 48334 49798 48540
rect 43580 48241 47731 48334
rect 39152 48128 43283 48241
rect 34728 48020 38864 48128
rect 28138 47802 29900 48020
rect 25891 47780 27849 47802
rect 21528 47671 25594 47780
tri 25594 47671 25703 47780 sw
tri 25891 47671 26000 47780 ne
rect 26000 47671 27849 47780
rect 21528 47602 25703 47671
rect 17200 47404 21246 47602
tri 17200 47312 17292 47404 ne
rect 17292 47320 21246 47404
tri 21246 47320 21528 47602 sw
tri 21528 47320 21810 47602 ne
rect 21810 47374 25703 47602
tri 25703 47374 26000 47671 sw
tri 26000 47374 26297 47671 ne
rect 26297 47513 27849 47671
tri 27849 47513 28138 47802 sw
tri 28138 47513 28427 47802 ne
rect 28427 47730 29900 47802
tri 29900 47730 30190 48020 sw
tri 30190 47730 30480 48020 ne
rect 30480 47730 34434 48020
rect 28427 47513 30190 47730
rect 26297 47374 28138 47513
rect 21810 47320 26000 47374
rect 17292 47312 21528 47320
tri 17000 47112 17200 47312 sw
tri 17292 47112 17492 47312 ne
rect 17492 47274 21528 47312
tri 21528 47274 21574 47320 sw
tri 21810 47274 21856 47320 ne
rect 21856 47274 26000 47320
rect 17492 47112 21574 47274
rect 14000 46908 17200 47112
tri 17200 46908 17404 47112 sw
tri 17492 46908 17696 47112 ne
rect 17696 46992 21574 47112
tri 21574 46992 21856 47274 sw
tri 21856 46992 22138 47274 ne
rect 22138 47077 26000 47274
tri 26000 47077 26297 47374 sw
tri 26297 47077 26594 47374 ne
rect 26594 47358 28138 47374
tri 28138 47358 28293 47513 sw
tri 28427 47358 28582 47513 ne
rect 28582 47440 30190 47513
tri 30190 47440 30480 47730 sw
tri 30480 47440 30770 47730 ne
rect 30770 47726 34434 47730
tri 34434 47726 34728 48020 sw
tri 34728 47726 35022 48020 ne
rect 35022 47840 38864 48020
tri 38864 47840 39152 48128 sw
tri 39152 47840 39440 48128 ne
rect 39440 47944 43283 48128
tri 43283 47944 43580 48241 sw
tri 43580 47944 43877 48241 ne
rect 43877 48041 47731 48241
tri 47731 48041 48024 48334 sw
tri 48024 48041 48317 48334 ne
rect 48317 48248 49798 48334
tri 49798 48248 50090 48540 sw
tri 50090 48248 50382 48540 ne
rect 50382 48253 52070 48540
tri 52070 48253 52357 48540 sw
tri 52357 48253 52644 48540 ne
rect 52644 48297 56542 48540
tri 56542 48297 56853 48608 sw
tri 56853 48297 57164 48608 ne
rect 57164 48297 71000 48608
rect 52644 48253 56853 48297
rect 50382 48248 52357 48253
rect 48317 48041 50090 48248
rect 43877 47944 48024 48041
rect 39440 47840 43580 47944
rect 35022 47726 39152 47840
rect 30770 47564 34728 47726
tri 34728 47564 34890 47726 sw
tri 35022 47564 35184 47726 ne
rect 35184 47564 39152 47726
rect 30770 47440 34890 47564
rect 28582 47358 30480 47440
rect 26594 47077 28293 47358
rect 22138 46992 26297 47077
rect 17696 46908 21856 46992
rect 14000 46616 17404 46908
tri 17404 46616 17696 46908 sw
tri 17696 46616 17988 46908 ne
rect 17988 46710 21856 46908
tri 21856 46710 22138 46992 sw
tri 22138 46710 22420 46992 ne
rect 22420 46780 26297 46992
tri 26297 46780 26594 47077 sw
tri 26594 46780 26891 47077 ne
rect 26891 47069 28293 47077
tri 28293 47069 28582 47358 sw
tri 28582 47069 28871 47358 ne
rect 28871 47266 30480 47358
tri 30480 47266 30654 47440 sw
tri 30770 47266 30944 47440 ne
rect 30944 47270 34890 47440
tri 34890 47270 35184 47564 sw
tri 35184 47270 35478 47564 ne
rect 35478 47552 39152 47564
tri 39152 47552 39440 47840 sw
tri 39440 47552 39728 47840 ne
rect 39728 47647 43580 47840
tri 43580 47647 43877 47944 sw
tri 43877 47647 44174 47944 ne
rect 44174 47819 48024 47944
tri 48024 47819 48246 48041 sw
tri 48317 47819 48539 48041 ne
rect 48539 47956 50090 48041
tri 50090 47956 50382 48248 sw
tri 50382 47956 50674 48248 ne
rect 50674 47966 52357 48248
tri 52357 47966 52644 48253 sw
tri 52644 47966 52931 48253 ne
rect 52931 47986 56853 48253
tri 56853 47986 57164 48297 sw
tri 57164 47986 57475 48297 ne
rect 57475 47986 71000 48297
rect 52931 47966 57164 47986
rect 50674 47956 52644 47966
rect 48539 47819 50382 47956
rect 44174 47647 48246 47819
rect 39728 47552 43877 47647
rect 35478 47270 39440 47552
rect 30944 47266 35184 47270
rect 28871 47069 30654 47266
rect 26891 46780 28582 47069
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 46976 30654 47069
tri 30654 46976 30944 47266 sw
tri 30944 46976 31234 47266 ne
rect 31234 46976 35184 47266
tri 35184 46976 35478 47270 sw
tri 35478 46976 35772 47270 ne
rect 35772 47264 39440 47270
tri 39440 47264 39728 47552 sw
tri 39728 47264 40016 47552 ne
rect 40016 47417 43877 47552
tri 43877 47417 44107 47647 sw
tri 44174 47417 44404 47647 ne
rect 44404 47526 48246 47647
tri 48246 47526 48539 47819 sw
tri 48539 47526 48832 47819 ne
rect 48832 47664 50382 47819
tri 50382 47664 50674 47956 sw
tri 50674 47664 50966 47956 ne
rect 50966 47679 52644 47956
tri 52644 47679 52931 47966 sw
tri 52931 47679 53218 47966 ne
rect 53218 47679 57164 47966
rect 50966 47664 52931 47679
rect 48832 47526 50674 47664
rect 44404 47417 48539 47526
rect 40016 47264 44107 47417
rect 35772 46976 39728 47264
tri 39728 46976 40016 47264 sw
tri 40016 46976 40304 47264 ne
rect 40304 47120 44107 47264
tri 44107 47120 44404 47417 sw
tri 44404 47120 44701 47417 ne
rect 44701 47233 48539 47417
tri 48539 47233 48832 47526 sw
tri 48832 47233 49125 47526 ne
rect 49125 47524 50674 47526
tri 50674 47524 50814 47664 sw
tri 50966 47524 51106 47664 ne
rect 51106 47627 52931 47664
tri 52931 47627 52983 47679 sw
tri 53218 47627 53270 47679 ne
rect 53270 47675 57164 47679
tri 57164 47675 57475 47986 sw
tri 57475 47675 57786 47986 ne
rect 57786 47675 71000 47986
rect 53270 47627 57475 47675
rect 51106 47524 52983 47627
rect 49125 47233 50814 47524
rect 44701 47120 48832 47233
rect 40304 46976 44404 47120
rect 29160 46780 30944 46976
rect 22420 46710 26594 46780
rect 17988 46616 22138 46710
rect 14000 46324 17696 46616
tri 17696 46324 17988 46616 sw
tri 17988 46324 18280 46616 ne
rect 18280 46428 22138 46616
tri 22138 46428 22420 46710 sw
tri 22420 46428 22702 46710 ne
rect 22702 46483 26594 46710
tri 26594 46483 26891 46780 sw
tri 26891 46483 27188 46780 ne
rect 27188 46689 28871 46780
tri 28871 46689 28962 46780 sw
tri 29160 46689 29251 46780 ne
rect 29251 46690 30944 46780
tri 30944 46690 31230 46976 sw
tri 31234 46690 31520 46976 ne
rect 31520 46690 35478 46976
rect 29251 46689 31230 46690
rect 27188 46483 28962 46689
rect 22702 46428 26891 46483
rect 18280 46324 22420 46428
rect 14000 46068 17988 46324
tri 14000 43708 16360 46068 ne
rect 16360 46032 17988 46068
tri 17988 46032 18280 46324 sw
tri 18280 46032 18572 46324 ne
rect 18572 46146 22420 46324
tri 22420 46146 22702 46428 sw
tri 22702 46146 22984 46428 ne
rect 22984 46186 26891 46428
tri 26891 46186 27188 46483 sw
tri 27188 46186 27485 46483 ne
rect 27485 46400 28962 46483
tri 28962 46400 29251 46689 sw
tri 29251 46400 29540 46689 ne
rect 29540 46400 31230 46689
tri 31230 46400 31520 46690 sw
tri 31520 46400 31810 46690 ne
rect 31810 46682 35478 46690
tri 35478 46682 35772 46976 sw
tri 35772 46682 36066 46976 ne
rect 36066 46688 40016 46976
tri 40016 46688 40304 46976 sw
tri 40304 46688 40592 46976 ne
rect 40592 46823 44404 46976
tri 44404 46823 44701 47120 sw
tri 44701 46823 44998 47120 ne
rect 44998 46940 48832 47120
tri 48832 46940 49125 47233 sw
tri 49125 46940 49418 47233 ne
rect 49418 47232 50814 47233
tri 50814 47232 51106 47524 sw
tri 51106 47232 51398 47524 ne
rect 51398 47340 52983 47524
tri 52983 47340 53270 47627 sw
tri 53270 47340 53557 47627 ne
rect 53557 47364 57475 47627
tri 57475 47364 57786 47675 sw
tri 57786 47364 58097 47675 ne
rect 58097 47364 71000 47675
rect 53557 47340 57786 47364
rect 51398 47232 53270 47340
rect 49418 46940 51106 47232
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47053 53270 47232
tri 53270 47053 53557 47340 sw
tri 53557 47053 53844 47340 ne
rect 53844 47053 57786 47340
tri 57786 47053 58097 47364 sw
tri 58097 47053 58408 47364 ne
rect 58408 47053 71000 47364
rect 51690 46940 53557 47053
rect 44998 46823 49125 46940
rect 40592 46688 44701 46823
rect 36066 46682 40304 46688
rect 31810 46400 35772 46682
rect 27485 46186 29251 46400
rect 22984 46146 27188 46186
rect 18572 46032 22702 46146
rect 16360 45740 18280 46032
tri 18280 45740 18572 46032 sw
tri 18572 45740 18864 46032 ne
rect 18864 45864 22702 46032
tri 22702 45864 22984 46146 sw
tri 22984 45864 23266 46146 ne
rect 23266 45889 27188 46146
tri 27188 45889 27485 46186 sw
tri 27485 45889 27782 46186 ne
rect 27782 46111 29251 46186
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46111 31520 46400
rect 27782 45889 29540 46111
rect 23266 45864 27485 45889
rect 18864 45740 22984 45864
rect 16360 45448 18572 45740
tri 18572 45448 18864 45740 sw
tri 18864 45448 19156 45740 ne
rect 19156 45582 22984 45740
tri 22984 45582 23266 45864 sw
tri 23266 45582 23548 45864 ne
rect 23548 45691 27485 45864
tri 27485 45691 27683 45889 sw
tri 27782 45691 27980 45889 ne
rect 27980 45822 29540 45889
tri 29540 45822 29829 46111 sw
tri 29829 45822 30118 46111 ne
rect 30118 46110 31520 46111
tri 31520 46110 31810 46400 sw
tri 31810 46110 32100 46400 ne
rect 32100 46388 35772 46400
tri 35772 46388 36066 46682 sw
tri 36066 46388 36360 46682 ne
rect 36360 46508 40304 46682
tri 40304 46508 40484 46688 sw
tri 40592 46508 40772 46688 ne
rect 40772 46526 44701 46688
tri 44701 46526 44998 46823 sw
tri 44998 46526 45295 46823 ne
rect 45295 46647 49125 46823
tri 49125 46647 49418 46940 sw
tri 49418 46647 49711 46940 ne
rect 49711 46852 51398 46940
tri 51398 46852 51486 46940 sw
tri 51690 46852 51778 46940 ne
rect 51778 46852 53557 46940
rect 49711 46647 51486 46852
rect 45295 46526 49418 46647
rect 40772 46508 44998 46526
rect 36360 46388 40484 46508
rect 32100 46110 36066 46388
rect 30118 45822 31810 46110
rect 27980 45691 29829 45822
rect 23548 45582 27683 45691
rect 19156 45448 23266 45582
rect 16360 45168 18864 45448
tri 18864 45168 19144 45448 sw
tri 19156 45168 19436 45448 ne
rect 19436 45300 23266 45448
tri 23266 45300 23548 45582 sw
tri 23548 45300 23830 45582 ne
rect 23830 45394 27683 45582
tri 27683 45394 27980 45691 sw
tri 27980 45394 28277 45691 ne
rect 28277 45533 29829 45691
tri 29829 45533 30118 45822 sw
tri 30118 45533 30407 45822 ne
rect 30407 45820 31810 45822
tri 31810 45820 32100 46110 sw
tri 32100 45820 32390 46110 ne
rect 32390 46094 36066 46110
tri 36066 46094 36360 46388 sw
tri 36360 46094 36654 46388 ne
rect 36654 46220 40484 46388
tri 40484 46220 40772 46508 sw
tri 40772 46220 41060 46508 ne
rect 41060 46229 44998 46508
tri 44998 46229 45295 46526 sw
tri 45295 46229 45592 46526 ne
rect 45592 46354 49418 46526
tri 49418 46354 49711 46647 sw
tri 49711 46354 50004 46647 ne
rect 50004 46560 51486 46647
tri 51486 46560 51778 46852 sw
tri 51778 46560 52070 46852 ne
rect 52070 46847 53557 46852
tri 53557 46847 53763 47053 sw
tri 53844 46847 54050 47053 ne
rect 54050 46847 58097 47053
rect 52070 46560 53763 46847
tri 53763 46560 54050 46847 sw
tri 54050 46560 54337 46847 ne
rect 54337 46742 58097 46847
tri 58097 46742 58408 47053 sw
tri 58408 46742 58719 47053 ne
rect 58719 46742 71000 47053
rect 54337 46622 58408 46742
tri 58408 46622 58528 46742 sw
tri 58719 46622 58839 46742 ne
rect 58839 46622 71000 46742
rect 54337 46560 58528 46622
rect 50004 46354 51778 46560
rect 45592 46229 49711 46354
rect 41060 46220 45295 46229
rect 36654 46094 40772 46220
rect 32390 45820 36360 46094
rect 30407 45533 32100 45820
rect 28277 45394 30118 45533
rect 23830 45300 27980 45394
rect 19436 45168 23548 45300
rect 16360 44876 19144 45168
tri 19144 44876 19436 45168 sw
tri 19436 44876 19728 45168 ne
rect 19728 45018 23548 45168
tri 23548 45018 23830 45300 sw
tri 23830 45018 24112 45300 ne
rect 24112 45097 27980 45300
tri 27980 45097 28277 45394 sw
tri 28277 45097 28574 45394 ne
rect 28574 45378 30118 45394
tri 30118 45378 30273 45533 sw
tri 30407 45378 30562 45533 ne
rect 30562 45530 32100 45533
tri 32100 45530 32390 45820 sw
tri 32390 45530 32680 45820 ne
rect 32680 45800 36360 45820
tri 36360 45800 36654 46094 sw
tri 36654 45800 36948 46094 ne
rect 36948 45932 40772 46094
tri 40772 45932 41060 46220 sw
tri 41060 45932 41348 46220 ne
rect 41348 45932 45295 46220
tri 45295 45932 45592 46229 sw
tri 45592 45932 45889 46229 ne
rect 45889 46061 49711 46229
tri 49711 46061 50004 46354 sw
tri 50004 46061 50297 46354 ne
rect 50297 46268 51778 46354
tri 51778 46268 52070 46560 sw
tri 52070 46268 52362 46560 ne
rect 52362 46273 54050 46560
tri 54050 46273 54337 46560 sw
tri 54337 46273 54624 46560 ne
rect 54624 46311 58528 46560
tri 58528 46311 58839 46622 sw
tri 58839 46311 59150 46622 ne
rect 59150 46311 71000 46622
rect 54624 46273 58839 46311
rect 52362 46268 54337 46273
rect 50297 46061 52070 46268
rect 45889 45932 50004 46061
rect 36948 45800 41060 45932
rect 32680 45530 36654 45800
rect 30562 45380 32390 45530
tri 32390 45380 32540 45530 sw
tri 32680 45380 32830 45530 ne
rect 32830 45506 36654 45530
tri 36654 45506 36948 45800 sw
tri 36948 45506 37242 45800 ne
rect 37242 45644 41060 45800
tri 41060 45644 41348 45932 sw
tri 41348 45644 41636 45932 ne
rect 41636 45644 45592 45932
rect 37242 45506 41348 45644
rect 32830 45380 36948 45506
rect 30562 45378 32540 45380
rect 28574 45097 30273 45378
rect 24112 45018 28277 45097
rect 19728 44876 23830 45018
rect 16360 44584 19436 44876
tri 19436 44584 19728 44876 sw
tri 19728 44584 20020 44876 ne
rect 20020 44736 23830 44876
tri 23830 44736 24112 45018 sw
tri 24112 44736 24394 45018 ne
rect 24394 44800 28277 45018
tri 28277 44800 28574 45097 sw
tri 28574 44800 28871 45097 ne
rect 28871 45089 30273 45097
tri 30273 45089 30562 45378 sw
tri 30562 45089 30851 45378 ne
rect 30851 45090 32540 45378
tri 32540 45090 32830 45380 sw
tri 32830 45090 33120 45380 ne
rect 33120 45246 36948 45380
tri 36948 45246 37208 45506 sw
tri 37242 45246 37502 45506 ne
rect 37502 45356 41348 45506
tri 41348 45356 41636 45644 sw
tri 41636 45356 41924 45644 ne
rect 41924 45635 45592 45644
tri 45592 45635 45889 45932 sw
tri 45889 45635 46186 45932 ne
rect 46186 45839 50004 45932
tri 50004 45839 50226 46061 sw
tri 50297 45839 50519 46061 ne
rect 50519 45976 52070 46061
tri 52070 45976 52362 46268 sw
tri 52362 45976 52654 46268 ne
rect 52654 46000 54337 46268
tri 54337 46000 54610 46273 sw
tri 54624 46000 54897 46273 ne
rect 54897 46000 58839 46273
tri 58839 46000 59150 46311 sw
tri 59150 46000 59461 46311 ne
rect 59461 46000 71000 46311
rect 52654 45976 54610 46000
rect 50519 45839 52362 45976
rect 46186 45635 50226 45839
rect 41924 45482 45889 45635
tri 45889 45482 46042 45635 sw
tri 46186 45482 46339 45635 ne
rect 46339 45546 50226 45635
tri 50226 45546 50519 45839 sw
tri 50519 45546 50812 45839 ne
rect 50812 45684 52362 45839
tri 52362 45684 52654 45976 sw
tri 52654 45684 52946 45976 ne
rect 52946 45713 54610 45976
tri 54610 45713 54897 46000 sw
tri 54897 45713 55184 46000 ne
rect 55184 45799 59150 46000
tri 59150 45799 59351 46000 sw
rect 55184 45739 71000 45799
rect 55184 45713 70613 45739
rect 52946 45684 54897 45713
rect 50812 45546 52654 45684
rect 46339 45482 50519 45546
rect 41924 45356 46042 45482
rect 37502 45246 41636 45356
rect 33120 45090 37208 45246
rect 30851 45089 32830 45090
rect 28871 44800 30562 45089
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 44800 32830 45089
tri 32830 44800 33120 45090 sw
tri 33120 44800 33410 45090 ne
rect 33410 44952 37208 45090
tri 37208 44952 37502 45246 sw
tri 37502 44952 37796 45246 ne
rect 37796 45068 41636 45246
tri 41636 45068 41924 45356 sw
tri 41924 45068 42212 45356 ne
rect 42212 45185 46042 45356
tri 46042 45185 46339 45482 sw
tri 46339 45185 46636 45482 ne
rect 46636 45253 50519 45482
tri 50519 45253 50812 45546 sw
tri 50812 45253 51105 45546 ne
rect 51105 45544 52654 45546
tri 52654 45544 52794 45684 sw
tri 52946 45544 53086 45684 ne
rect 53086 45544 54897 45684
rect 51105 45253 52794 45544
rect 46636 45185 50812 45253
rect 42212 45068 46339 45185
rect 37796 44952 41924 45068
rect 33410 44800 37502 44952
rect 24394 44736 28574 44800
rect 20020 44584 24112 44736
rect 16360 44292 19728 44584
tri 19728 44292 20020 44584 sw
tri 20020 44292 20312 44584 ne
rect 20312 44454 24112 44584
tri 24112 44454 24394 44736 sw
tri 24394 44454 24676 44736 ne
rect 24676 44503 28574 44736
tri 28574 44503 28871 44800 sw
tri 28871 44503 29168 44800 ne
rect 29168 44709 30851 44800
tri 30851 44709 30942 44800 sw
tri 31140 44709 31231 44800 ne
rect 31231 44710 33120 44800
tri 33120 44710 33210 44800 sw
tri 33410 44710 33500 44800 ne
rect 33500 44710 37502 44800
rect 31231 44709 33210 44710
rect 29168 44503 30942 44709
rect 24676 44454 28871 44503
rect 20312 44292 24394 44454
rect 16360 44000 20020 44292
tri 20020 44000 20312 44292 sw
tri 20312 44000 20604 44292 ne
rect 20604 44172 24394 44292
tri 24394 44172 24676 44454 sw
tri 24676 44172 24958 44454 ne
rect 24958 44206 28871 44454
tri 28871 44206 29168 44503 sw
tri 29168 44206 29465 44503 ne
rect 29465 44420 30942 44503
tri 30942 44420 31231 44709 sw
tri 31231 44420 31520 44709 ne
rect 31520 44420 33210 44709
tri 33210 44420 33500 44710 sw
tri 33500 44420 33790 44710 ne
rect 33790 44658 37502 44710
tri 37502 44658 37796 44952 sw
tri 37796 44658 38090 44952 ne
rect 38090 44780 41924 44952
tri 41924 44780 42212 45068 sw
tri 42212 44780 42500 45068 ne
rect 42500 44888 46339 45068
tri 46339 44888 46636 45185 sw
tri 46636 44888 46933 45185 ne
rect 46933 44960 50812 45185
tri 50812 44960 51105 45253 sw
tri 51105 44960 51398 45253 ne
rect 51398 45252 52794 45253
tri 52794 45252 53086 45544 sw
tri 53086 45252 53378 45544 ne
rect 53378 45426 54897 45544
tri 54897 45426 55184 45713 sw
tri 55184 45426 55471 45713 ne
rect 55471 45426 70613 45713
rect 53378 45252 55184 45426
rect 51398 44960 53086 45252
tri 53086 44960 53378 45252 sw
tri 53378 44960 53670 45252 ne
rect 53670 45247 55184 45252
tri 55184 45247 55363 45426 sw
tri 55471 45247 55650 45426 ne
rect 55650 45247 70613 45426
rect 53670 44960 55363 45247
tri 55363 44960 55650 45247 sw
tri 55650 44960 55937 45247 ne
rect 55937 44960 70613 45247
rect 46933 44888 51105 44960
rect 42500 44780 46636 44888
rect 38090 44658 42212 44780
rect 33790 44420 37796 44658
rect 29465 44206 31231 44420
rect 24958 44172 29168 44206
rect 20604 44000 24676 44172
rect 16360 43708 20312 44000
tri 20312 43708 20604 44000 sw
tri 20604 43708 20896 44000 ne
rect 20896 43917 24676 44000
tri 24676 43917 24931 44172 sw
tri 24958 43917 25213 44172 ne
rect 25213 43917 29168 44172
rect 20896 43708 24931 43917
tri 16360 42664 17404 43708 ne
rect 17404 43416 20604 43708
tri 20604 43416 20896 43708 sw
tri 20896 43416 21188 43708 ne
rect 21188 43635 24931 43708
tri 24931 43635 25213 43917 sw
tri 25213 43635 25495 43917 ne
rect 25495 43909 29168 43917
tri 29168 43909 29465 44206 sw
tri 29465 43909 29762 44206 ne
rect 29762 44131 31231 44206
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44131 33500 44420
rect 29762 43909 31520 44131
rect 25495 43711 29465 43909
tri 29465 43711 29663 43909 sw
tri 29762 43711 29960 43909 ne
rect 29960 43842 31520 43909
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44130 33500 44131
tri 33500 44130 33790 44420 sw
tri 33790 44130 34080 44420 ne
rect 34080 44364 37796 44420
tri 37796 44364 38090 44658 sw
tri 38090 44364 38384 44658 ne
rect 38384 44492 42212 44658
tri 42212 44492 42500 44780 sw
tri 42500 44492 42788 44780 ne
rect 42788 44591 46636 44780
tri 46636 44591 46933 44888 sw
tri 46933 44591 47230 44888 ne
rect 47230 44667 51105 44888
tri 51105 44667 51398 44960 sw
tri 51398 44667 51691 44960 ne
rect 51691 44872 53378 44960
tri 53378 44872 53466 44960 sw
tri 53670 44872 53758 44960 ne
rect 53758 44872 55650 44960
rect 51691 44667 53466 44872
rect 47230 44591 51398 44667
rect 42788 44492 46933 44591
rect 38384 44364 42500 44492
rect 34080 44130 38090 44364
rect 32098 44066 33790 44130
tri 33790 44066 33854 44130 sw
tri 34080 44066 34144 44130 ne
rect 34144 44070 38090 44130
tri 38090 44070 38384 44364 sw
tri 38384 44070 38678 44364 ne
rect 38678 44204 42500 44364
tri 42500 44204 42788 44492 sw
tri 42788 44204 43076 44492 ne
rect 43076 44294 46933 44492
tri 46933 44294 47230 44591 sw
tri 47230 44294 47527 44591 ne
rect 47527 44374 51398 44591
tri 51398 44374 51691 44667 sw
tri 51691 44374 51984 44667 ne
rect 51984 44580 53466 44667
tri 53466 44580 53758 44872 sw
tri 53758 44580 54050 44872 ne
rect 54050 44867 55650 44872
tri 55650 44867 55743 44960 sw
tri 55937 44867 56030 44960 ne
rect 56030 44867 70613 44960
rect 54050 44580 55743 44867
tri 55743 44580 56030 44867 sw
tri 56030 44580 56317 44867 ne
rect 56317 44580 70613 44867
rect 51984 44374 53758 44580
rect 47527 44294 51691 44374
rect 43076 44204 47230 44294
rect 38678 44172 42788 44204
tri 42788 44172 42820 44204 sw
tri 43076 44172 43108 44204 ne
rect 43108 44172 47230 44204
rect 38678 44070 42820 44172
rect 34144 44066 38384 44070
rect 32098 43842 33854 44066
rect 29960 43711 31809 43842
rect 25495 43635 29663 43711
rect 21188 43416 25213 43635
rect 17404 43248 20896 43416
tri 20896 43248 21064 43416 sw
tri 21188 43248 21356 43416 ne
rect 21356 43353 25213 43416
tri 25213 43353 25495 43635 sw
tri 25495 43353 25777 43635 ne
rect 25777 43414 29663 43635
tri 29663 43414 29960 43711 sw
tri 29960 43414 30257 43711 ne
rect 30257 43553 31809 43711
tri 31809 43553 32098 43842 sw
tri 32098 43553 32387 43842 ne
rect 32387 43776 33854 43842
tri 33854 43776 34144 44066 sw
tri 34144 43776 34434 44066 ne
rect 34434 43776 38384 44066
tri 38384 43776 38678 44070 sw
tri 38678 43776 38972 44070 ne
rect 38972 43884 42820 44070
tri 42820 43884 43108 44172 sw
tri 43108 43884 43396 44172 ne
rect 43396 43997 47230 44172
tri 47230 43997 47527 44294 sw
tri 47527 43997 47824 44294 ne
rect 47824 44081 51691 44294
tri 51691 44081 51984 44374 sw
tri 51984 44081 52277 44374 ne
rect 52277 44288 53758 44374
tri 53758 44288 54050 44580 sw
tri 54050 44288 54342 44580 ne
rect 54342 44293 56030 44580
tri 56030 44293 56317 44580 sw
tri 56317 44293 56604 44580 ne
rect 56604 44293 70613 44580
rect 54342 44288 56317 44293
rect 52277 44081 54050 44288
rect 47824 43997 51984 44081
rect 43396 43884 47527 43997
rect 38972 43776 43108 43884
rect 32387 43553 34144 43776
rect 30257 43414 32098 43553
rect 25777 43353 29960 43414
rect 21356 43248 25495 43353
rect 17404 42956 21064 43248
tri 21064 42956 21356 43248 sw
tri 21356 42956 21648 43248 ne
rect 21648 43071 25495 43248
tri 25495 43071 25777 43353 sw
tri 25777 43071 26059 43353 ne
rect 26059 43117 29960 43353
tri 29960 43117 30257 43414 sw
tri 30257 43117 30554 43414 ne
rect 30554 43310 32098 43414
tri 32098 43310 32341 43553 sw
tri 32387 43310 32630 43553 ne
rect 32630 43486 34144 43553
tri 34144 43486 34434 43776 sw
tri 34434 43486 34724 43776 ne
rect 34724 43486 38678 43776
rect 32630 43310 34434 43486
rect 30554 43117 32341 43310
rect 26059 43071 30257 43117
rect 21648 42956 25777 43071
rect 17404 42664 21356 42956
tri 21356 42664 21648 42956 sw
tri 21648 42664 21940 42956 ne
rect 21940 42789 25777 42956
tri 25777 42789 26059 43071 sw
tri 26059 42789 26341 43071 ne
rect 26341 42820 30257 43071
tri 30257 42820 30554 43117 sw
tri 30554 42820 30851 43117 ne
rect 30851 43021 32341 43117
tri 32341 43021 32630 43310 sw
tri 32630 43021 32919 43310 ne
rect 32919 43196 34434 43310
tri 34434 43196 34724 43486 sw
tri 34724 43196 35014 43486 ne
rect 35014 43482 38678 43486
tri 38678 43482 38972 43776 sw
tri 38972 43482 39266 43776 ne
rect 39266 43596 43108 43776
tri 43108 43596 43396 43884 sw
tri 43396 43596 43684 43884 ne
rect 43684 43700 47527 43884
tri 47527 43700 47824 43997 sw
tri 47824 43700 48121 43997 ne
rect 48121 43859 51984 43997
tri 51984 43859 52206 44081 sw
tri 52277 43859 52499 44081 ne
rect 52499 43996 54050 44081
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44006 56317 44288
tri 56317 44006 56604 44293 sw
tri 56604 44006 56891 44293 ne
rect 56891 44006 70613 44293
rect 54634 43996 56604 44006
rect 52499 43859 54342 43996
rect 48121 43700 52206 43859
rect 43684 43596 47824 43700
rect 39266 43482 43396 43596
rect 35014 43320 38972 43482
tri 38972 43320 39134 43482 sw
tri 39266 43320 39428 43482 ne
rect 39428 43320 43396 43482
rect 35014 43196 39134 43320
rect 32919 43022 34724 43196
tri 34724 43022 34898 43196 sw
tri 35014 43022 35188 43196 ne
rect 35188 43026 39134 43196
tri 39134 43026 39428 43320 sw
tri 39428 43026 39722 43320 ne
rect 39722 43308 43396 43320
tri 43396 43308 43684 43596 sw
tri 43684 43308 43972 43596 ne
rect 43972 43403 47824 43596
tri 47824 43403 48121 43700 sw
tri 48121 43403 48418 43700 ne
rect 48418 43566 52206 43700
tri 52206 43566 52499 43859 sw
tri 52499 43566 52792 43859 ne
rect 52792 43704 54342 43859
tri 54342 43704 54634 43996 sw
tri 54634 43704 54926 43996 ne
rect 54926 43719 56604 43996
tri 56604 43719 56891 44006 sw
tri 56891 43719 57178 44006 ne
rect 57178 43719 70613 44006
rect 54926 43704 56891 43719
rect 52792 43566 54634 43704
rect 48418 43403 52499 43566
rect 43972 43308 48121 43403
rect 39722 43026 43684 43308
rect 35188 43022 39428 43026
rect 32919 43021 34898 43022
rect 30851 42820 32630 43021
rect 26341 42789 30554 42820
rect 21940 42664 26059 42789
tri 17404 38420 21648 42664 ne
tri 21648 42372 21940 42664 sw
tri 21940 42372 22232 42664 ne
rect 22232 42507 26059 42664
tri 26059 42507 26341 42789 sw
tri 26341 42507 26623 42789 ne
rect 26623 42523 30554 42789
tri 30554 42523 30851 42820 sw
tri 30851 42523 31148 42820 ne
rect 31148 42732 32630 42820
tri 32630 42732 32919 43021 sw
tri 32919 42732 33208 43021 ne
rect 33208 42732 34898 43021
tri 34898 42732 35188 43022 sw
tri 35188 42732 35478 43022 ne
rect 35478 42732 39428 43022
tri 39428 42732 39722 43026 sw
tri 39722 42732 40016 43026 ne
rect 40016 43020 43684 43026
tri 43684 43020 43972 43308 sw
tri 43972 43020 44260 43308 ne
rect 44260 43173 48121 43308
tri 48121 43173 48351 43403 sw
tri 48418 43173 48648 43403 ne
rect 48648 43273 52499 43403
tri 52499 43273 52792 43566 sw
tri 52792 43273 53085 43566 ne
rect 53085 43564 54634 43566
tri 54634 43564 54774 43704 sw
tri 54926 43564 55066 43704 ne
rect 55066 43564 56891 43704
rect 53085 43273 54774 43564
rect 48648 43173 52792 43273
rect 44260 43020 48351 43173
rect 40016 42732 43972 43020
tri 43972 42732 44260 43020 sw
tri 44260 42732 44548 43020 ne
rect 44548 42876 48351 43020
tri 48351 42876 48648 43173 sw
tri 48648 42876 48945 43173 ne
rect 48945 42980 52792 43173
tri 52792 42980 53085 43273 sw
tri 53085 42980 53378 43273 ne
rect 53378 43272 54774 43273
tri 54774 43272 55066 43564 sw
tri 55066 43272 55358 43564 ne
rect 55358 43554 56891 43564
tri 56891 43554 57056 43719 sw
tri 57178 43554 57343 43719 ne
rect 57343 43554 70613 43719
rect 55358 43272 57056 43554
rect 53378 42980 55066 43272
tri 55066 42980 55358 43272 sw
tri 55358 42980 55650 43272 ne
rect 55650 43267 57056 43272
tri 57056 43267 57343 43554 sw
tri 57343 43267 57630 43554 ne
rect 57630 43267 70613 43554
rect 55650 42980 57343 43267
tri 57343 42980 57630 43267 sw
tri 57630 42980 57917 43267 ne
rect 57917 42980 70613 43267
rect 48945 42876 53085 42980
rect 44548 42732 48648 42876
rect 31148 42729 32919 42732
tri 32919 42729 32922 42732 sw
tri 33208 42729 33211 42732 ne
rect 33211 42730 35188 42732
tri 35188 42730 35190 42732 sw
tri 35478 42730 35480 42732 ne
rect 35480 42730 39722 42732
rect 33211 42729 35190 42730
rect 31148 42523 32922 42729
rect 26623 42507 30851 42523
rect 22232 42372 26341 42507
rect 21648 42080 21940 42372
tri 21940 42080 22232 42372 sw
tri 22232 42080 22524 42372 ne
rect 22524 42225 26341 42372
tri 26341 42225 26623 42507 sw
tri 26623 42225 26905 42507 ne
rect 26905 42226 30851 42507
tri 30851 42226 31148 42523 sw
tri 31148 42226 31445 42523 ne
rect 31445 42440 32922 42523
tri 32922 42440 33211 42729 sw
tri 33211 42440 33500 42729 ne
rect 33500 42440 35190 42729
tri 35190 42440 35480 42730 sw
tri 35480 42440 35770 42730 ne
rect 35770 42440 39722 42730
rect 31445 42226 33211 42440
rect 26905 42225 31148 42226
rect 22524 42184 26623 42225
tri 26623 42184 26664 42225 sw
tri 26905 42184 26946 42225 ne
rect 26946 42184 31148 42225
rect 22524 42080 26664 42184
rect 21648 41788 22232 42080
tri 22232 41788 22524 42080 sw
tri 22524 41788 22816 42080 ne
rect 22816 41902 26664 42080
tri 26664 41902 26946 42184 sw
tri 26946 41902 27228 42184 ne
rect 27228 41929 31148 42184
tri 31148 41929 31445 42226 sw
tri 31445 41929 31742 42226 ne
rect 31742 42151 33211 42226
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42151 35480 42440
rect 31742 41929 33500 42151
rect 27228 41902 31445 41929
rect 22816 41788 26946 41902
rect 21648 41496 22524 41788
tri 22524 41496 22816 41788 sw
tri 22816 41496 23108 41788 ne
rect 23108 41620 26946 41788
tri 26946 41620 27228 41902 sw
tri 27228 41620 27510 41902 ne
rect 27510 41731 31445 41902
tri 31445 41731 31643 41929 sw
tri 31742 41731 31940 41929 ne
rect 31940 41862 33500 41929
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 42150 35480 42151
tri 35480 42150 35770 42440 sw
tri 35770 42150 36060 42440 ne
rect 36060 42438 39722 42440
tri 39722 42438 40016 42732 sw
tri 40016 42438 40310 42732 ne
rect 40310 42444 44260 42732
tri 44260 42444 44548 42732 sw
tri 44548 42444 44836 42732 ne
rect 44836 42579 48648 42732
tri 48648 42579 48945 42876 sw
tri 48945 42579 49242 42876 ne
rect 49242 42687 53085 42876
tri 53085 42687 53378 42980 sw
tri 53378 42687 53671 42980 ne
rect 53671 42892 55358 42980
tri 55358 42892 55446 42980 sw
tri 55650 42892 55738 42980 ne
rect 55738 42892 57630 42980
rect 53671 42687 55446 42892
rect 49242 42579 53378 42687
rect 44836 42444 48945 42579
rect 40310 42438 44548 42444
rect 36060 42150 40016 42438
rect 34078 41862 35770 42150
rect 31940 41731 33789 41862
rect 27510 41620 31643 41731
rect 23108 41496 27228 41620
rect 21648 41204 22816 41496
tri 22816 41204 23108 41496 sw
tri 23108 41204 23400 41496 ne
rect 23400 41338 27228 41496
tri 27228 41338 27510 41620 sw
tri 27510 41338 27792 41620 ne
rect 27792 41434 31643 41620
tri 31643 41434 31940 41731 sw
tri 31940 41434 32237 41731 ne
rect 32237 41573 33789 41731
tri 33789 41573 34078 41862 sw
tri 34078 41573 34367 41862 ne
rect 34367 41860 35770 41862
tri 35770 41860 36060 42150 sw
tri 36060 41860 36350 42150 ne
rect 36350 42144 40016 42150
tri 40016 42144 40310 42438 sw
tri 40310 42144 40604 42438 ne
rect 40604 42264 44548 42438
tri 44548 42264 44728 42444 sw
tri 44836 42264 45016 42444 ne
rect 45016 42282 48945 42444
tri 48945 42282 49242 42579 sw
tri 49242 42282 49539 42579 ne
rect 49539 42394 53378 42579
tri 53378 42394 53671 42687 sw
tri 53671 42394 53964 42687 ne
rect 53964 42600 55446 42687
tri 55446 42600 55738 42892 sw
tri 55738 42600 56030 42892 ne
rect 56030 42800 57630 42892
tri 57630 42800 57810 42980 sw
tri 57917 42800 58097 42980 ne
rect 58097 42875 70613 42980
rect 70669 42875 71000 45739
rect 58097 42800 71000 42875
rect 56030 42600 57810 42800
tri 57810 42600 58010 42800 sw
rect 53964 42394 55738 42600
rect 49539 42282 53671 42394
rect 45016 42264 49242 42282
rect 40604 42144 44728 42264
rect 36350 41860 40310 42144
rect 34367 41573 36060 41860
rect 32237 41434 34078 41573
rect 27792 41338 31940 41434
rect 23400 41204 27510 41338
rect 21648 40924 23108 41204
tri 23108 40924 23388 41204 sw
tri 23400 40924 23680 41204 ne
rect 23680 41056 27510 41204
tri 27510 41056 27792 41338 sw
tri 27792 41056 28074 41338 ne
rect 28074 41137 31940 41338
tri 31940 41137 32237 41434 sw
tri 32237 41137 32534 41434 ne
rect 32534 41418 34078 41434
tri 34078 41418 34233 41573 sw
tri 34367 41418 34522 41573 ne
rect 34522 41570 36060 41573
tri 36060 41570 36350 41860 sw
tri 36350 41570 36640 41860 ne
rect 36640 41850 40310 41860
tri 40310 41850 40604 42144 sw
tri 40604 41850 40898 42144 ne
rect 40898 41976 44728 42144
tri 44728 41976 45016 42264 sw
tri 45016 41976 45304 42264 ne
rect 45304 41985 49242 42264
tri 49242 41985 49539 42282 sw
tri 49539 41985 49836 42282 ne
rect 49836 42101 53671 42282
tri 53671 42101 53964 42394 sw
tri 53964 42101 54257 42394 ne
rect 54257 42308 55738 42394
tri 55738 42308 56030 42600 sw
tri 56030 42308 56322 42600 ne
rect 56322 42497 71000 42600
rect 56322 42308 70613 42497
rect 54257 42101 56030 42308
rect 49836 41985 53964 42101
rect 45304 41976 49539 41985
rect 40898 41850 45016 41976
rect 36640 41570 40604 41850
rect 34522 41420 36350 41570
tri 36350 41420 36500 41570 sw
tri 36640 41420 36790 41570 ne
rect 36790 41556 40604 41570
tri 40604 41556 40898 41850 sw
tri 40898 41556 41192 41850 ne
rect 41192 41688 45016 41850
tri 45016 41688 45304 41976 sw
tri 45304 41688 45592 41976 ne
rect 45592 41688 49539 41976
tri 49539 41688 49836 41985 sw
tri 49836 41688 50133 41985 ne
rect 50133 41879 53964 41985
tri 53964 41879 54186 42101 sw
tri 54257 41879 54479 42101 ne
rect 54479 42016 56030 42101
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 70613 42308
rect 54479 41879 56322 42016
rect 50133 41688 54186 41879
rect 41192 41556 45304 41688
rect 36790 41420 40898 41556
rect 34522 41418 36500 41420
rect 32534 41137 34233 41418
rect 28074 41056 32237 41137
rect 23680 40924 27792 41056
rect 21648 40632 23388 40924
tri 23388 40632 23680 40924 sw
tri 23680 40632 23972 40924 ne
rect 23972 40774 27792 40924
tri 27792 40774 28074 41056 sw
tri 28074 40774 28356 41056 ne
rect 28356 40840 32237 41056
tri 32237 40840 32534 41137 sw
tri 32534 40840 32831 41137 ne
rect 32831 41129 34233 41137
tri 34233 41129 34522 41418 sw
tri 34522 41129 34811 41418 ne
rect 34811 41130 36500 41418
tri 36500 41130 36790 41420 sw
tri 36790 41130 37080 41420 ne
rect 37080 41262 40898 41420
tri 40898 41262 41192 41556 sw
tri 41192 41262 41486 41556 ne
rect 41486 41400 45304 41556
tri 45304 41400 45592 41688 sw
tri 45592 41400 45880 41688 ne
rect 45880 41400 49836 41688
rect 41486 41262 45592 41400
rect 37080 41130 41192 41262
rect 34811 41129 36790 41130
rect 32831 40840 34522 41129
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 40840 36790 41129
tri 36790 40840 37080 41130 sw
tri 37080 40840 37370 41130 ne
rect 37370 41002 41192 41130
tri 41192 41002 41452 41262 sw
tri 41486 41002 41746 41262 ne
rect 41746 41112 45592 41262
tri 45592 41112 45880 41400 sw
tri 45880 41112 46168 41400 ne
rect 46168 41391 49836 41400
tri 49836 41391 50133 41688 sw
tri 50133 41391 50430 41688 ne
rect 50430 41586 54186 41688
tri 54186 41586 54479 41879 sw
tri 54479 41586 54772 41879 ne
rect 54772 41784 56322 41879
tri 56322 41784 56554 42016 sw
tri 56614 41784 56846 42016 ne
rect 56846 41784 70613 42016
rect 54772 41586 56554 41784
rect 50430 41391 54479 41586
rect 46168 41238 50133 41391
tri 50133 41238 50286 41391 sw
tri 50430 41238 50583 41391 ne
rect 50583 41293 54479 41391
tri 54479 41293 54772 41586 sw
tri 54772 41293 55065 41586 ne
rect 55065 41492 56554 41586
tri 56554 41492 56846 41784 sw
tri 56846 41492 57138 41784 ne
rect 57138 41492 70613 41784
rect 55065 41293 56846 41492
rect 50583 41238 54772 41293
rect 46168 41112 50286 41238
rect 41746 41002 45880 41112
rect 37370 40840 41452 41002
rect 28356 40774 32534 40840
rect 23972 40632 28074 40774
rect 21648 40340 23680 40632
tri 23680 40340 23972 40632 sw
tri 23972 40340 24264 40632 ne
rect 24264 40492 28074 40632
tri 28074 40492 28356 40774 sw
tri 28356 40492 28638 40774 ne
rect 28638 40543 32534 40774
tri 32534 40543 32831 40840 sw
tri 32831 40543 33128 40840 ne
rect 33128 40749 34811 40840
tri 34811 40749 34902 40840 sw
tri 35100 40749 35191 40840 ne
rect 35191 40750 37080 40840
tri 37080 40750 37170 40840 sw
tri 37370 40750 37460 40840 ne
rect 37460 40750 41452 40840
rect 35191 40749 37170 40750
rect 33128 40543 34902 40749
rect 28638 40492 32831 40543
rect 24264 40340 28356 40492
rect 21648 40048 23972 40340
tri 23972 40048 24264 40340 sw
tri 24264 40048 24556 40340 ne
rect 24556 40210 28356 40340
tri 28356 40210 28638 40492 sw
tri 28638 40210 28920 40492 ne
rect 28920 40246 32831 40492
tri 32831 40246 33128 40543 sw
tri 33128 40246 33425 40543 ne
rect 33425 40460 34902 40543
tri 34902 40460 35191 40749 sw
tri 35191 40460 35480 40749 ne
rect 35480 40460 37170 40749
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40708 41452 40750
tri 41452 40708 41746 41002 sw
tri 41746 40708 42040 41002 ne
rect 42040 40824 45880 41002
tri 45880 40824 46168 41112 sw
tri 46168 40824 46456 41112 ne
rect 46456 40941 50286 41112
tri 50286 40941 50583 41238 sw
tri 50583 40941 50880 41238 ne
rect 50880 41000 54772 41238
tri 54772 41000 55065 41293 sw
tri 55065 41000 55358 41293 ne
rect 55358 41200 56846 41293
tri 56846 41200 57138 41492 sw
tri 57138 41200 57430 41492 ne
rect 57430 41297 70613 41492
rect 70669 41297 71000 42497
rect 57430 41200 71000 41297
rect 55358 41000 57138 41200
tri 57138 41000 57338 41200 sw
rect 50880 40941 55065 41000
rect 46456 40824 50583 40941
rect 42040 40708 46168 40824
rect 37750 40460 41746 40708
rect 33425 40246 35191 40460
rect 28920 40210 33128 40246
rect 24556 40048 28638 40210
rect 21648 39756 24264 40048
tri 24264 39756 24556 40048 sw
tri 24556 39756 24848 40048 ne
rect 24848 39928 28638 40048
tri 28638 39928 28920 40210 sw
tri 28920 39928 29202 40210 ne
rect 29202 39949 33128 40210
tri 33128 39949 33425 40246 sw
tri 33425 39949 33722 40246 ne
rect 33722 40171 35191 40246
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40171 37460 40460
rect 33722 39949 35480 40171
rect 29202 39928 33425 39949
rect 24848 39830 28920 39928
tri 28920 39830 29018 39928 sw
tri 29202 39830 29300 39928 ne
rect 29300 39830 33425 39928
rect 24848 39756 29018 39830
rect 21648 39464 24556 39756
tri 24556 39464 24848 39756 sw
tri 24848 39464 25140 39756 ne
rect 25140 39548 29018 39756
tri 29018 39548 29300 39830 sw
tri 29300 39548 29582 39830 ne
rect 29582 39751 33425 39830
tri 33425 39751 33623 39949 sw
tri 33722 39751 33920 39949 ne
rect 33920 39882 35480 39949
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40170 37460 40171
tri 37460 40170 37750 40460 sw
tri 37750 40170 38040 40460 ne
rect 38040 40414 41746 40460
tri 41746 40414 42040 40708 sw
tri 42040 40414 42334 40708 ne
rect 42334 40536 46168 40708
tri 46168 40536 46456 40824 sw
tri 46456 40536 46744 40824 ne
rect 46744 40644 50583 40824
tri 50583 40644 50880 40941 sw
tri 50880 40644 51177 40941 ne
rect 51177 40707 55065 40941
tri 55065 40707 55358 41000 sw
tri 55358 40707 55651 41000 ne
rect 55651 40707 71000 41000
rect 51177 40644 55358 40707
rect 46744 40536 50880 40644
rect 42334 40414 46456 40536
rect 38040 40170 42040 40414
rect 36058 39882 37750 40170
rect 33920 39751 35769 39882
rect 29582 39548 33623 39751
rect 25140 39464 29300 39548
rect 21648 39172 24848 39464
tri 24848 39172 25140 39464 sw
tri 25140 39172 25432 39464 ne
rect 25432 39266 29300 39464
tri 29300 39266 29582 39548 sw
tri 29582 39266 29864 39548 ne
rect 29864 39454 33623 39548
tri 33623 39454 33920 39751 sw
tri 33920 39454 34217 39751 ne
rect 34217 39593 35769 39751
tri 35769 39593 36058 39882 sw
tri 36058 39593 36347 39882 ne
rect 36347 39880 37750 39882
tri 37750 39880 38040 40170 sw
tri 38040 39880 38330 40170 ne
rect 38330 40120 42040 40170
tri 42040 40120 42334 40414 sw
tri 42334 40120 42628 40414 ne
rect 42628 40248 46456 40414
tri 46456 40248 46744 40536 sw
tri 46744 40248 47032 40536 ne
rect 47032 40347 50880 40536
tri 50880 40347 51177 40644 sw
tri 51177 40347 51474 40644 ne
rect 51474 40414 55358 40644
tri 55358 40414 55651 40707 sw
tri 55651 40414 55944 40707 ne
rect 55944 40414 71000 40707
rect 51474 40347 55651 40414
rect 47032 40248 51177 40347
rect 42628 40120 46744 40248
rect 38330 39880 42334 40120
rect 36347 39822 38040 39880
tri 38040 39822 38098 39880 sw
tri 38330 39822 38388 39880 ne
rect 38388 39826 42334 39880
tri 42334 39826 42628 40120 sw
tri 42628 39826 42922 40120 ne
rect 42922 39960 46744 40120
tri 46744 39960 47032 40248 sw
tri 47032 39960 47320 40248 ne
rect 47320 40050 51177 40248
tri 51177 40050 51474 40347 sw
tri 51474 40050 51771 40347 ne
rect 51771 40186 55651 40347
tri 55651 40186 55879 40414 sw
tri 55944 40186 56172 40414 ne
rect 56172 40186 71000 40414
rect 51771 40050 55879 40186
rect 47320 39960 51474 40050
rect 42922 39928 47032 39960
tri 47032 39928 47064 39960 sw
tri 47320 39928 47352 39960 ne
rect 47352 39928 51474 39960
rect 42922 39826 47064 39928
rect 38388 39822 42628 39826
rect 36347 39593 38098 39822
rect 34217 39454 36058 39593
rect 29864 39266 33920 39454
rect 25432 39172 29582 39266
rect 21648 39004 25140 39172
tri 25140 39004 25308 39172 sw
tri 25432 39004 25600 39172 ne
rect 25600 39004 29582 39172
rect 21648 38712 25308 39004
tri 25308 38712 25600 39004 sw
tri 25600 38712 25892 39004 ne
rect 25892 38984 29582 39004
tri 29582 38984 29864 39266 sw
tri 29864 38984 30146 39266 ne
rect 30146 39157 33920 39266
tri 33920 39157 34217 39454 sw
tri 34217 39157 34514 39454 ne
rect 34514 39438 36058 39454
tri 36058 39438 36213 39593 sw
tri 36347 39438 36502 39593 ne
rect 36502 39532 38098 39593
tri 38098 39532 38388 39822 sw
tri 38388 39532 38678 39822 ne
rect 38678 39532 42628 39822
tri 42628 39532 42922 39826 sw
tri 42922 39532 43216 39826 ne
rect 43216 39640 47064 39826
tri 47064 39640 47352 39928 sw
tri 47352 39640 47640 39928 ne
rect 47640 39753 51474 39928
tri 51474 39753 51771 40050 sw
tri 51771 39753 52068 40050 ne
rect 52068 39893 55879 40050
tri 55879 39893 56172 40186 sw
tri 56172 39893 56465 40186 ne
rect 56465 39893 71000 40186
rect 52068 39753 56172 39893
rect 47640 39640 51771 39753
rect 43216 39532 47352 39640
rect 36502 39438 38388 39532
rect 34514 39157 36213 39438
rect 30146 38984 34217 39157
rect 25892 38712 29864 38984
rect 21648 38420 25600 38712
tri 25600 38420 25892 38712 sw
tri 25892 38420 26184 38712 ne
rect 26184 38702 29864 38712
tri 29864 38702 30146 38984 sw
tri 30146 38702 30428 38984 ne
rect 30428 38860 34217 38984
tri 34217 38860 34514 39157 sw
tri 34514 38860 34811 39157 ne
rect 34811 39149 36213 39157
tri 36213 39149 36502 39438 sw
tri 36502 39149 36791 39438 ne
rect 36791 39242 38388 39438
tri 38388 39242 38678 39532 sw
tri 38678 39242 38968 39532 ne
rect 38968 39242 42922 39532
rect 36791 39149 38678 39242
rect 34811 38860 36502 39149
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 39060 38678 39149
tri 38678 39060 38860 39242 sw
tri 38968 39060 39150 39242 ne
rect 39150 39238 42922 39242
tri 42922 39238 43216 39532 sw
tri 43216 39238 43510 39532 ne
rect 43510 39352 47352 39532
tri 47352 39352 47640 39640 sw
tri 47640 39352 47928 39640 ne
rect 47928 39456 51771 39640
tri 51771 39456 52068 39753 sw
tri 52068 39456 52365 39753 ne
rect 52365 39600 56172 39753
tri 56172 39600 56465 39893 sw
tri 56465 39600 56758 39893 ne
rect 56758 39600 71000 39893
rect 52365 39456 56465 39600
rect 47928 39352 52068 39456
rect 43510 39238 47640 39352
rect 39150 39076 43216 39238
tri 43216 39076 43378 39238 sw
tri 43510 39076 43672 39238 ne
rect 43672 39076 47640 39238
rect 39150 39060 43378 39076
rect 37080 38860 38860 39060
rect 30428 38702 34514 38860
rect 26184 38420 30146 38702
tri 30146 38420 30428 38702 sw
tri 30428 38420 30710 38702 ne
rect 30710 38563 34514 38702
tri 34514 38563 34811 38860 sw
tri 34811 38563 35108 38860 ne
rect 35108 38777 36791 38860
tri 36791 38777 36874 38860 sw
tri 37080 38777 37163 38860 ne
rect 37163 38777 38860 38860
rect 35108 38563 36874 38777
rect 30710 38420 34811 38563
tri 21648 34176 25892 38420 ne
tri 25892 38128 26184 38420 sw
tri 26184 38128 26476 38420 ne
rect 26476 38138 30428 38420
tri 30428 38138 30710 38420 sw
tri 30710 38138 30992 38420 ne
rect 30992 38266 34811 38420
tri 34811 38266 35108 38563 sw
tri 35108 38266 35405 38563 ne
rect 35405 38488 36874 38563
tri 36874 38488 37163 38777 sw
tri 37163 38488 37452 38777 ne
rect 37452 38770 38860 38777
tri 38860 38770 39150 39060 sw
tri 39150 38770 39440 39060 ne
rect 39440 38782 43378 39060
tri 43378 38782 43672 39076 sw
tri 43672 38782 43966 39076 ne
rect 43966 39064 47640 39076
tri 47640 39064 47928 39352 sw
tri 47928 39064 48216 39352 ne
rect 48216 39159 52068 39352
tri 52068 39159 52365 39456 sw
tri 52365 39159 52662 39456 ne
rect 52662 39400 56465 39456
tri 56465 39400 56665 39600 sw
rect 52662 39332 71000 39400
rect 52662 39159 70613 39332
rect 48216 39064 52365 39159
rect 43966 38782 47928 39064
rect 39440 38770 43672 38782
rect 37452 38488 39150 38770
rect 35405 38480 37163 38488
tri 37163 38480 37171 38488 sw
tri 37452 38480 37460 38488 ne
rect 37460 38480 39150 38488
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38488 43672 38770
tri 43672 38488 43966 38782 sw
tri 43966 38488 44260 38782 ne
rect 44260 38776 47928 38782
tri 47928 38776 48216 39064 sw
tri 48216 38776 48504 39064 ne
rect 48504 38929 52365 39064
tri 52365 38929 52595 39159 sw
tri 52662 38929 52892 39159 ne
rect 52892 38929 70613 39159
rect 48504 38776 52595 38929
rect 44260 38488 48216 38776
tri 48216 38488 48504 38776 sw
tri 48504 38488 48792 38776 ne
rect 48792 38632 52595 38776
tri 52595 38632 52892 38929 sw
tri 52892 38632 53189 38929 ne
rect 53189 38632 70613 38929
rect 48792 38488 52892 38632
rect 39730 38480 43966 38488
rect 35405 38266 37171 38480
rect 30992 38138 35108 38266
rect 26476 38128 30710 38138
rect 25892 37836 26184 38128
tri 26184 37836 26476 38128 sw
tri 26476 37836 26768 38128 ne
rect 26768 37940 30710 38128
tri 30710 37940 30908 38138 sw
tri 30992 37940 31190 38138 ne
rect 31190 37969 35108 38138
tri 35108 37969 35405 38266 sw
tri 35405 37969 35702 38266 ne
rect 35702 38191 37171 38266
tri 37171 38191 37460 38480 sw
tri 37460 38191 37749 38480 ne
rect 37749 38191 39440 38480
rect 35702 37969 37460 38191
rect 31190 37940 35405 37969
rect 26768 37836 30908 37940
rect 25892 37544 26476 37836
tri 26476 37544 26768 37836 sw
tri 26768 37544 27060 37836 ne
rect 27060 37658 30908 37836
tri 30908 37658 31190 37940 sw
tri 31190 37658 31472 37940 ne
rect 31472 37771 35405 37940
tri 35405 37771 35603 37969 sw
tri 35702 37771 35900 37969 ne
rect 35900 37902 37460 37969
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 38190 39440 38191
tri 39440 38190 39730 38480 sw
tri 39730 38190 40020 38480 ne
rect 40020 38194 43966 38480
tri 43966 38194 44260 38488 sw
tri 44260 38194 44554 38488 ne
rect 44554 38200 48504 38488
tri 48504 38200 48792 38488 sw
tri 48792 38200 49080 38488 ne
rect 49080 38335 52892 38488
tri 52892 38335 53189 38632 sw
tri 53189 38335 53486 38632 ne
rect 53486 38335 70613 38632
rect 49080 38200 53189 38335
rect 44554 38194 48792 38200
rect 40020 38190 44260 38194
rect 38038 37902 39730 38190
rect 35900 37771 37749 37902
rect 31472 37658 35603 37771
rect 27060 37544 31190 37658
rect 25892 37252 26768 37544
tri 26768 37252 27060 37544 sw
tri 27060 37252 27352 37544 ne
rect 27352 37376 31190 37544
tri 31190 37376 31472 37658 sw
tri 31472 37376 31754 37658 ne
rect 31754 37474 35603 37658
tri 35603 37474 35900 37771 sw
tri 35900 37474 36197 37771 ne
rect 36197 37613 37749 37771
tri 37749 37613 38038 37902 sw
tri 38038 37613 38327 37902 ne
rect 38327 37900 39730 37902
tri 39730 37900 40020 38190 sw
tri 40020 37900 40310 38190 ne
rect 40310 37900 44260 38190
tri 44260 37900 44554 38194 sw
tri 44554 37900 44848 38194 ne
rect 44848 38020 48792 38194
tri 48792 38020 48972 38200 sw
tri 49080 38020 49260 38200 ne
rect 49260 38038 53189 38200
tri 53189 38038 53486 38335 sw
tri 53486 38038 53783 38335 ne
rect 53783 38038 70613 38335
rect 49260 38020 53486 38038
rect 44848 37900 48972 38020
rect 38327 37613 40020 37900
rect 36197 37474 38038 37613
rect 31754 37376 35900 37474
rect 27352 37252 31472 37376
rect 25892 36960 27060 37252
tri 27060 36960 27352 37252 sw
tri 27352 36960 27644 37252 ne
rect 27644 37094 31472 37252
tri 31472 37094 31754 37376 sw
tri 31754 37094 32036 37376 ne
rect 32036 37177 35900 37376
tri 35900 37177 36197 37474 sw
tri 36197 37177 36494 37474 ne
rect 36494 37458 38038 37474
tri 38038 37458 38193 37613 sw
tri 38327 37458 38482 37613 ne
rect 38482 37610 40020 37613
tri 40020 37610 40310 37900 sw
tri 40310 37610 40600 37900 ne
rect 40600 37610 44554 37900
rect 38482 37460 40310 37610
tri 40310 37460 40460 37610 sw
tri 40600 37460 40750 37610 ne
rect 40750 37606 44554 37610
tri 44554 37606 44848 37900 sw
tri 44848 37606 45142 37900 ne
rect 45142 37732 48972 37900
tri 48972 37732 49260 38020 sw
tri 49260 37732 49548 38020 ne
rect 49548 37741 53486 38020
tri 53486 37741 53783 38038 sw
tri 53783 37741 54080 38038 ne
rect 54080 37741 70613 38038
rect 49548 37732 53783 37741
rect 45142 37606 49260 37732
rect 40750 37460 44848 37606
rect 38482 37458 40460 37460
rect 36494 37177 38193 37458
rect 32036 37094 36197 37177
rect 27644 36960 31754 37094
rect 25892 36680 27352 36960
tri 27352 36680 27632 36960 sw
tri 27644 36680 27924 36960 ne
rect 27924 36812 31754 36960
tri 31754 36812 32036 37094 sw
tri 32036 36812 32318 37094 ne
rect 32318 36880 36197 37094
tri 36197 36880 36494 37177 sw
tri 36494 36880 36791 37177 ne
rect 36791 37169 38193 37177
tri 38193 37169 38482 37458 sw
tri 38482 37169 38771 37458 ne
rect 38771 37170 40460 37458
tri 40460 37170 40750 37460 sw
tri 40750 37170 41040 37460 ne
rect 41040 37312 44848 37460
tri 44848 37312 45142 37606 sw
tri 45142 37312 45436 37606 ne
rect 45436 37444 49260 37606
tri 49260 37444 49548 37732 sw
tri 49548 37444 49836 37732 ne
rect 49836 37444 53783 37732
tri 53783 37444 54080 37741 sw
tri 54080 37444 54377 37741 ne
rect 54377 37444 70613 37741
rect 45436 37312 49548 37444
rect 41040 37170 45142 37312
rect 38771 37169 40750 37170
rect 36791 36880 38482 37169
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 36880 40750 37169
tri 40750 36880 41040 37170 sw
tri 41040 36880 41330 37170 ne
rect 41330 37018 45142 37170
tri 45142 37018 45436 37312 sw
tri 45436 37018 45730 37312 ne
rect 45730 37156 49548 37312
tri 49548 37156 49836 37444 sw
tri 49836 37156 50124 37444 ne
rect 50124 37156 54080 37444
rect 45730 37018 49836 37156
rect 41330 36880 45436 37018
rect 32318 36812 36494 36880
rect 27924 36680 32036 36812
rect 25892 36388 27632 36680
tri 27632 36388 27924 36680 sw
tri 27924 36388 28216 36680 ne
rect 28216 36530 32036 36680
tri 32036 36530 32318 36812 sw
tri 32318 36530 32600 36812 ne
rect 32600 36583 36494 36812
tri 36494 36583 36791 36880 sw
tri 36791 36583 37088 36880 ne
rect 37088 36789 38771 36880
tri 38771 36789 38862 36880 sw
tri 39060 36789 39151 36880 ne
rect 39151 36790 41040 36880
tri 41040 36790 41130 36880 sw
tri 41330 36790 41420 36880 ne
rect 41420 36790 45436 36880
rect 39151 36789 41130 36790
rect 37088 36583 38862 36789
rect 32600 36530 36791 36583
rect 28216 36388 32318 36530
rect 25892 36096 27924 36388
tri 27924 36096 28216 36388 sw
tri 28216 36096 28508 36388 ne
rect 28508 36248 32318 36388
tri 32318 36248 32600 36530 sw
tri 32600 36248 32882 36530 ne
rect 32882 36286 36791 36530
tri 36791 36286 37088 36583 sw
tri 37088 36286 37385 36583 ne
rect 37385 36500 38862 36583
tri 38862 36500 39151 36789 sw
tri 39151 36500 39440 36789 ne
rect 39440 36500 41130 36789
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36758 45436 36790
tri 45436 36758 45696 37018 sw
tri 45730 36758 45990 37018 ne
rect 45990 36868 49836 37018
tri 49836 36868 50124 37156 sw
tri 50124 36868 50412 37156 ne
rect 50412 37147 54080 37156
tri 54080 37147 54377 37444 sw
tri 54377 37147 54674 37444 ne
rect 54674 37147 70613 37444
rect 50412 36994 54377 37147
tri 54377 36994 54530 37147 sw
tri 54674 36994 54827 37147 ne
rect 54827 36994 70613 37147
rect 50412 36868 54530 36994
rect 45990 36758 50124 36868
rect 41710 36500 45696 36758
rect 37385 36286 39151 36500
rect 32882 36248 37088 36286
rect 28508 36096 32600 36248
rect 25892 35804 28216 36096
tri 28216 35804 28508 36096 sw
tri 28508 35804 28800 36096 ne
rect 28800 35966 32600 36096
tri 32600 35966 32882 36248 sw
tri 32882 35966 33164 36248 ne
rect 33164 35989 37088 36248
tri 37088 35989 37385 36286 sw
tri 37385 35989 37682 36286 ne
rect 37682 36211 39151 36286
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36211 41420 36500
rect 37682 35989 39440 36211
rect 33164 35966 37385 35989
rect 28800 35804 32882 35966
rect 25892 35512 28508 35804
tri 28508 35512 28800 35804 sw
tri 28800 35512 29092 35804 ne
rect 29092 35684 32882 35804
tri 32882 35684 33164 35966 sw
tri 33164 35684 33446 35966 ne
rect 33446 35791 37385 35966
tri 37385 35791 37583 35989 sw
tri 37682 35791 37880 35989 ne
rect 37880 35922 39440 35989
tri 39440 35922 39729 36211 sw
tri 39729 35922 40018 36211 ne
rect 40018 36210 41420 36211
tri 41420 36210 41710 36500 sw
tri 41710 36210 42000 36500 ne
rect 42000 36464 45696 36500
tri 45696 36464 45990 36758 sw
tri 45990 36464 46284 36758 ne
rect 46284 36580 50124 36758
tri 50124 36580 50412 36868 sw
tri 50412 36580 50700 36868 ne
rect 50700 36697 54530 36868
tri 54530 36697 54827 36994 sw
tri 54827 36697 55124 36994 ne
rect 55124 36697 70613 36994
rect 50700 36580 54827 36697
rect 46284 36464 50412 36580
rect 42000 36210 45990 36464
rect 40018 35922 41710 36210
rect 37880 35791 39729 35922
rect 33446 35684 37583 35791
rect 29092 35586 33164 35684
tri 33164 35586 33262 35684 sw
tri 33446 35586 33544 35684 ne
rect 33544 35586 37583 35684
rect 29092 35512 33262 35586
rect 25892 35220 28800 35512
tri 28800 35220 29092 35512 sw
tri 29092 35220 29384 35512 ne
rect 29384 35304 33262 35512
tri 33262 35304 33544 35586 sw
tri 33544 35304 33826 35586 ne
rect 33826 35494 37583 35586
tri 37583 35494 37880 35791 sw
tri 37880 35494 38177 35791 ne
rect 38177 35633 39729 35791
tri 39729 35633 40018 35922 sw
tri 40018 35633 40307 35922 ne
rect 40307 35920 41710 35922
tri 41710 35920 42000 36210 sw
tri 42000 35920 42290 36210 ne
rect 42290 36170 45990 36210
tri 45990 36170 46284 36464 sw
tri 46284 36170 46578 36464 ne
rect 46578 36292 50412 36464
tri 50412 36292 50700 36580 sw
tri 50700 36292 50988 36580 ne
rect 50988 36400 54827 36580
tri 54827 36400 55124 36697 sw
tri 55124 36400 55421 36697 ne
rect 55421 36468 70613 36697
rect 70669 36468 71000 39332
rect 55421 36400 71000 36468
rect 50988 36292 55124 36400
rect 46578 36170 50700 36292
rect 42290 35920 46284 36170
rect 40307 35868 42000 35920
tri 42000 35868 42052 35920 sw
tri 42290 35868 42342 35920 ne
rect 42342 35876 46284 35920
tri 46284 35876 46578 36170 sw
tri 46578 35876 46872 36170 ne
rect 46872 36004 50700 36170
tri 50700 36004 50988 36292 sw
tri 50988 36004 51276 36292 ne
rect 51276 36200 55124 36292
tri 55124 36200 55324 36400 sw
rect 51276 36132 71000 36200
rect 51276 36004 70613 36132
rect 46872 35876 50988 36004
rect 42342 35868 46578 35876
rect 40307 35633 42052 35868
rect 38177 35494 40018 35633
rect 33826 35304 37880 35494
rect 29384 35220 33544 35304
rect 25892 34928 29092 35220
tri 29092 34928 29384 35220 sw
tri 29384 34928 29676 35220 ne
rect 29676 35022 33544 35220
tri 33544 35022 33826 35304 sw
tri 33826 35022 34108 35304 ne
rect 34108 35197 37880 35304
tri 37880 35197 38177 35494 sw
tri 38177 35197 38474 35494 ne
rect 38474 35478 40018 35494
tri 40018 35478 40173 35633 sw
tri 40307 35478 40462 35633 ne
rect 40462 35578 42052 35633
tri 42052 35578 42342 35868 sw
tri 42342 35578 42632 35868 ne
rect 42632 35582 46578 35868
tri 46578 35582 46872 35876 sw
tri 46872 35582 47166 35876 ne
rect 47166 35716 50988 35876
tri 50988 35716 51276 36004 sw
tri 51276 35716 51564 36004 ne
rect 51564 35716 70613 36004
rect 47166 35684 51276 35716
tri 51276 35684 51308 35716 sw
tri 51564 35684 51596 35716 ne
rect 51596 35684 70613 35716
rect 47166 35582 51308 35684
rect 42632 35578 46872 35582
rect 40462 35478 42342 35578
rect 38474 35197 40173 35478
rect 34108 35022 38177 35197
rect 29676 34928 33826 35022
rect 25892 34760 29384 34928
tri 29384 34760 29552 34928 sw
tri 29676 34760 29844 34928 ne
rect 29844 34760 33826 34928
rect 25892 34468 29552 34760
tri 29552 34468 29844 34760 sw
tri 29844 34468 30136 34760 ne
rect 30136 34740 33826 34760
tri 33826 34740 34108 35022 sw
tri 34108 34740 34390 35022 ne
rect 34390 34900 38177 35022
tri 38177 34900 38474 35197 sw
tri 38474 34900 38771 35197 ne
rect 38771 35189 40173 35197
tri 40173 35189 40462 35478 sw
tri 40462 35189 40751 35478 ne
rect 40751 35288 42342 35478
tri 42342 35288 42632 35578 sw
tri 42632 35288 42922 35578 ne
rect 42922 35288 46872 35578
tri 46872 35288 47166 35582 sw
tri 47166 35288 47460 35582 ne
rect 47460 35396 51308 35582
tri 51308 35396 51596 35684 sw
tri 51596 35396 51884 35684 ne
rect 51884 35396 70613 35684
rect 47460 35288 51596 35396
rect 40751 35189 42632 35288
rect 38771 34900 40462 35189
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42632 35189
tri 42632 34998 42922 35288 sw
tri 42922 34998 43212 35288 ne
rect 43212 34998 47166 35288
rect 41040 34900 42922 34998
rect 34390 34740 38474 34900
rect 30136 34468 34108 34740
rect 25892 34176 29844 34468
tri 29844 34176 30136 34468 sw
tri 30136 34176 30428 34468 ne
rect 30428 34458 34108 34468
tri 34108 34458 34390 34740 sw
tri 34390 34458 34672 34740 ne
rect 34672 34603 38474 34740
tri 38474 34603 38771 34900 sw
tri 38771 34603 39068 34900 ne
rect 39068 34809 40751 34900
tri 40751 34809 40842 34900 sw
tri 41040 34809 41131 34900 ne
rect 41131 34810 42922 34900
tri 42922 34810 43110 34998 sw
tri 43212 34810 43400 34998 ne
rect 43400 34994 47166 34998
tri 47166 34994 47460 35288 sw
tri 47460 34994 47754 35288 ne
rect 47754 35108 51596 35288
tri 51596 35108 51884 35396 sw
tri 51884 35108 52172 35396 ne
rect 52172 35108 70613 35396
rect 47754 34994 51884 35108
rect 43400 34832 47460 34994
tri 47460 34832 47622 34994 sw
tri 47754 34832 47916 34994 ne
rect 47916 34832 51884 34994
rect 43400 34810 47622 34832
rect 41131 34809 43110 34810
rect 39068 34603 40842 34809
rect 34672 34458 38771 34603
rect 30428 34176 34390 34458
tri 34390 34176 34672 34458 sw
tri 34672 34176 34954 34458 ne
rect 34954 34306 38771 34458
tri 38771 34306 39068 34603 sw
tri 39068 34306 39365 34603 ne
rect 39365 34520 40842 34603
tri 40842 34520 41131 34809 sw
tri 41131 34520 41420 34809 ne
rect 41420 34520 43110 34809
tri 43110 34520 43400 34810 sw
tri 43400 34520 43690 34810 ne
rect 43690 34538 47622 34810
tri 47622 34538 47916 34832 sw
tri 47916 34538 48210 34832 ne
rect 48210 34820 51884 34832
tri 51884 34820 52172 35108 sw
tri 52172 34820 52460 35108 ne
rect 52460 34820 70613 35108
rect 48210 34538 52172 34820
rect 43690 34520 47916 34538
rect 39365 34306 41131 34520
rect 34954 34176 39068 34306
tri 25892 29932 30136 34176 ne
tri 30136 33884 30428 34176 sw
tri 30428 33884 30720 34176 ne
rect 30720 33894 34672 34176
tri 34672 33894 34954 34176 sw
tri 34954 33894 35236 34176 ne
rect 35236 34009 39068 34176
tri 39068 34009 39365 34306 sw
tri 39365 34009 39662 34306 ne
rect 39662 34231 41131 34306
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34244 43400 34520
tri 43400 34244 43676 34520 sw
tri 43690 34244 43966 34520 ne
rect 43966 34244 47916 34520
tri 47916 34244 48210 34538 sw
tri 48210 34244 48504 34538 ne
rect 48504 34532 52172 34538
tri 52172 34532 52460 34820 sw
tri 52460 34532 52748 34820 ne
rect 52748 34532 70613 34820
rect 48504 34244 52460 34532
tri 52460 34244 52748 34532 sw
tri 52748 34244 53036 34532 ne
rect 53036 34244 70613 34532
rect 41709 34231 43676 34244
rect 39662 34009 41420 34231
rect 35236 33894 39365 34009
rect 30720 33884 34954 33894
rect 30136 33592 30428 33884
tri 30428 33592 30720 33884 sw
tri 30720 33592 31012 33884 ne
rect 31012 33696 34954 33884
tri 34954 33696 35152 33894 sw
tri 35236 33696 35434 33894 ne
rect 35434 33811 39365 33894
tri 39365 33811 39563 34009 sw
tri 39662 33811 39860 34009 ne
rect 39860 33942 41420 34009
tri 41420 33942 41709 34231 sw
tri 41709 33942 41998 34231 ne
rect 41998 33954 43676 34231
tri 43676 33954 43966 34244 sw
tri 43966 33954 44256 34244 ne
rect 44256 33954 48210 34244
rect 41998 33942 43966 33954
rect 39860 33811 41709 33942
rect 35434 33696 39563 33811
rect 31012 33592 35152 33696
rect 30136 33300 30720 33592
tri 30720 33300 31012 33592 sw
tri 31012 33300 31304 33592 ne
rect 31304 33414 35152 33592
tri 35152 33414 35434 33696 sw
tri 35434 33414 35716 33696 ne
rect 35716 33514 39563 33696
tri 39563 33514 39860 33811 sw
tri 39860 33514 40157 33811 ne
rect 40157 33653 41709 33811
tri 41709 33653 41998 33942 sw
tri 41998 33653 42287 33942 ne
rect 42287 33664 43966 33942
tri 43966 33664 44256 33954 sw
tri 44256 33664 44546 33954 ne
rect 44546 33950 48210 33954
tri 48210 33950 48504 34244 sw
tri 48504 33950 48798 34244 ne
rect 48798 33956 52748 34244
tri 52748 33956 53036 34244 sw
tri 53036 33956 53324 34244 ne
rect 53324 33956 70613 34244
rect 48798 33950 53036 33956
rect 44546 33664 48504 33950
rect 42287 33653 44256 33664
rect 40157 33514 41998 33653
rect 35716 33414 39860 33514
rect 31304 33300 35434 33414
rect 30136 33008 31012 33300
tri 31012 33008 31304 33300 sw
tri 31304 33008 31596 33300 ne
rect 31596 33132 35434 33300
tri 35434 33132 35716 33414 sw
tri 35716 33132 35998 33414 ne
rect 35998 33217 39860 33414
tri 39860 33217 40157 33514 sw
tri 40157 33217 40454 33514 ne
rect 40454 33498 41998 33514
tri 41998 33498 42153 33653 sw
tri 42287 33498 42442 33653 ne
rect 42442 33500 44256 33653
tri 44256 33500 44420 33664 sw
tri 44546 33500 44710 33664 ne
rect 44710 33656 48504 33664
tri 48504 33656 48798 33950 sw
tri 48798 33656 49092 33950 ne
rect 49092 33776 53036 33950
tri 53036 33776 53216 33956 sw
tri 53324 33776 53504 33956 ne
rect 53504 33776 70613 33956
rect 49092 33656 53216 33776
rect 44710 33500 48798 33656
rect 42442 33498 44420 33500
rect 40454 33217 42153 33498
rect 35998 33132 40157 33217
rect 31596 33008 35716 33132
rect 30136 32716 31304 33008
tri 31304 32716 31596 33008 sw
tri 31596 32716 31888 33008 ne
rect 31888 32850 35716 33008
tri 35716 32850 35998 33132 sw
tri 35998 32850 36280 33132 ne
rect 36280 32920 40157 33132
tri 40157 32920 40454 33217 sw
tri 40454 32920 40751 33217 ne
rect 40751 33209 42153 33217
tri 42153 33209 42442 33498 sw
tri 42442 33209 42731 33498 ne
rect 42731 33210 44420 33498
tri 44420 33210 44710 33500 sw
tri 44710 33210 45000 33500 ne
rect 45000 33362 48798 33500
tri 48798 33362 49092 33656 sw
tri 49092 33362 49386 33656 ne
rect 49386 33488 53216 33656
tri 53216 33488 53504 33776 sw
tri 53504 33488 53792 33776 ne
rect 53792 33488 70613 33776
rect 49386 33362 53504 33488
rect 45000 33210 49092 33362
rect 42731 33209 44710 33210
rect 40751 32920 42442 33209
tri 42442 32920 42731 33209 sw
tri 42731 32920 43020 33209 ne
rect 43020 32920 44710 33209
tri 44710 32920 45000 33210 sw
tri 45000 32920 45290 33210 ne
rect 45290 33068 49092 33210
tri 49092 33068 49386 33362 sw
tri 49386 33068 49680 33362 ne
rect 49680 33200 53504 33362
tri 53504 33200 53792 33488 sw
tri 53792 33200 54080 33488 ne
rect 54080 33268 70613 33488
rect 70669 33268 71000 36132
rect 54080 33200 71000 33268
rect 49680 33068 53792 33200
rect 45290 32920 49386 33068
rect 36280 32850 40454 32920
rect 31888 32716 35998 32850
rect 30136 32436 31596 32716
tri 31596 32436 31876 32716 sw
tri 31888 32436 32168 32716 ne
rect 32168 32568 35998 32716
tri 35998 32568 36280 32850 sw
tri 36280 32568 36562 32850 ne
rect 36562 32623 40454 32850
tri 40454 32623 40751 32920 sw
tri 40751 32623 41048 32920 ne
rect 41048 32829 42731 32920
tri 42731 32829 42822 32920 sw
tri 43020 32829 43111 32920 ne
rect 43111 32830 45000 32920
tri 45000 32830 45090 32920 sw
tri 45290 32830 45380 32920 ne
rect 45380 32830 49386 32920
rect 43111 32829 45090 32830
rect 41048 32623 42822 32829
rect 36562 32568 40751 32623
rect 32168 32436 36280 32568
rect 30136 32144 31876 32436
tri 31876 32144 32168 32436 sw
tri 32168 32144 32460 32436 ne
rect 32460 32286 36280 32436
tri 36280 32286 36562 32568 sw
tri 36562 32286 36844 32568 ne
rect 36844 32326 40751 32568
tri 40751 32326 41048 32623 sw
tri 41048 32326 41345 32623 ne
rect 41345 32540 42822 32623
tri 42822 32540 43111 32829 sw
tri 43111 32540 43400 32829 ne
rect 43400 32540 45090 32829
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32774 49386 32830
tri 49386 32774 49680 33068 sw
tri 49680 32774 49974 33068 ne
rect 49974 33000 53792 33068
tri 53792 33000 53992 33200 sw
rect 49974 32920 71000 33000
rect 49974 32774 70613 32920
rect 45670 32540 49680 32774
rect 41345 32326 43111 32540
rect 36844 32286 41048 32326
rect 32460 32144 36562 32286
rect 30136 31852 32168 32144
tri 32168 31852 32460 32144 sw
tri 32460 31852 32752 32144 ne
rect 32752 32004 36562 32144
tri 36562 32004 36844 32286 sw
tri 36844 32004 37126 32286 ne
rect 37126 32029 41048 32286
tri 41048 32029 41345 32326 sw
tri 41345 32029 41642 32326 ne
rect 41642 32251 43111 32326
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32251 45380 32540
rect 41642 32029 43400 32251
rect 37126 32004 41345 32029
rect 32752 31852 36844 32004
rect 30136 31560 32460 31852
tri 32460 31560 32752 31852 sw
tri 32752 31560 33044 31852 ne
rect 33044 31722 36844 31852
tri 36844 31722 37126 32004 sw
tri 37126 31722 37408 32004 ne
rect 37408 31831 41345 32004
tri 41345 31831 41543 32029 sw
tri 41642 31831 41840 32029 ne
rect 41840 31962 43400 32029
tri 43400 31962 43689 32251 sw
tri 43689 31962 43978 32251 ne
rect 43978 32250 45380 32251
tri 45380 32250 45670 32540 sw
tri 45670 32250 45960 32540 ne
rect 45960 32514 49680 32540
tri 49680 32514 49940 32774 sw
tri 49974 32514 50234 32774 ne
rect 50234 32514 70613 32774
rect 45960 32250 49940 32514
rect 43978 31962 45670 32250
rect 41840 31831 43689 31962
rect 37408 31722 41543 31831
rect 33044 31560 37126 31722
rect 30136 31268 32752 31560
tri 32752 31268 33044 31560 sw
tri 33044 31268 33336 31560 ne
rect 33336 31440 37126 31560
tri 37126 31440 37408 31722 sw
tri 37408 31440 37690 31722 ne
rect 37690 31534 41543 31722
tri 41543 31534 41840 31831 sw
tri 41840 31534 42137 31831 ne
rect 42137 31673 43689 31831
tri 43689 31673 43978 31962 sw
tri 43978 31673 44267 31962 ne
rect 44267 31960 45670 31962
tri 45670 31960 45960 32250 sw
tri 45960 31960 46250 32250 ne
rect 46250 32220 49940 32250
tri 49940 32220 50234 32514 sw
tri 50234 32220 50528 32514 ne
rect 50528 32220 70613 32514
rect 46250 31960 50234 32220
rect 44267 31673 45960 31960
rect 42137 31534 43978 31673
rect 37690 31440 41840 31534
rect 33336 31342 37408 31440
tri 37408 31342 37506 31440 sw
tri 37690 31342 37788 31440 ne
rect 37788 31342 41840 31440
rect 33336 31268 37506 31342
rect 30136 30976 33044 31268
tri 33044 30976 33336 31268 sw
tri 33336 30976 33628 31268 ne
rect 33628 31060 37506 31268
tri 37506 31060 37788 31342 sw
tri 37788 31060 38070 31342 ne
rect 38070 31237 41840 31342
tri 41840 31237 42137 31534 sw
tri 42137 31237 42434 31534 ne
rect 42434 31518 43978 31534
tri 43978 31518 44133 31673 sw
tri 44267 31518 44422 31673 ne
rect 44422 31670 45960 31673
tri 45960 31670 46250 31960 sw
tri 46250 31670 46540 31960 ne
rect 46540 31926 50234 31960
tri 50234 31926 50528 32220 sw
tri 50528 31926 50822 32220 ne
rect 50822 31926 70613 32220
rect 46540 31670 50528 31926
rect 44422 31624 46250 31670
tri 46250 31624 46296 31670 sw
tri 46540 31624 46586 31670 ne
rect 46586 31632 50528 31670
tri 50528 31632 50822 31926 sw
tri 50822 31632 51116 31926 ne
rect 51116 31632 70613 31926
rect 46586 31624 50822 31632
rect 44422 31518 46296 31624
rect 42434 31237 44133 31518
rect 38070 31060 42137 31237
rect 33628 30976 37788 31060
rect 30136 30684 33336 30976
tri 33336 30684 33628 30976 sw
tri 33628 30684 33920 30976 ne
rect 33920 30778 37788 30976
tri 37788 30778 38070 31060 sw
tri 38070 30778 38352 31060 ne
rect 38352 30940 42137 31060
tri 42137 30940 42434 31237 sw
tri 42434 30940 42731 31237 ne
rect 42731 31229 44133 31237
tri 44133 31229 44422 31518 sw
tri 44422 31229 44711 31518 ne
rect 44711 31334 46296 31518
tri 46296 31334 46586 31624 sw
tri 46586 31334 46876 31624 ne
rect 46876 31338 50822 31624
tri 50822 31338 51116 31632 sw
tri 51116 31338 51410 31632 ne
rect 51410 31338 70613 31632
rect 46876 31334 51116 31338
rect 44711 31229 46586 31334
rect 42731 30940 44422 31229
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31044 46586 31229
tri 46586 31044 46876 31334 sw
tri 46876 31044 47166 31334 ne
rect 47166 31044 51116 31334
tri 51116 31044 51410 31338 sw
tri 51410 31044 51704 31338 ne
rect 51704 31044 70613 31338
rect 45000 30940 46876 31044
rect 38352 30778 42434 30940
rect 33920 30684 38070 30778
rect 30136 30516 33628 30684
tri 33628 30516 33796 30684 sw
tri 33920 30516 34088 30684 ne
rect 34088 30516 38070 30684
rect 30136 30224 33796 30516
tri 33796 30224 34088 30516 sw
tri 34088 30224 34380 30516 ne
rect 34380 30496 38070 30516
tri 38070 30496 38352 30778 sw
tri 38352 30496 38634 30778 ne
rect 38634 30643 42434 30778
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30849 44711 30940
tri 44711 30849 44802 30940 sw
tri 45000 30849 45091 30940 ne
rect 45091 30850 46876 30940
tri 46876 30850 47070 31044 sw
tri 47166 30850 47360 31044 ne
rect 47360 30850 51410 31044
rect 45091 30849 47070 30850
rect 43028 30643 44802 30849
rect 38634 30496 42731 30643
rect 34380 30224 38352 30496
rect 30136 29932 34088 30224
tri 34088 29932 34380 30224 sw
tri 34380 29932 34672 30224 ne
rect 34672 30214 38352 30224
tri 38352 30214 38634 30496 sw
tri 38634 30214 38916 30496 ne
rect 38916 30346 42731 30496
tri 42731 30346 43028 30643 sw
tri 43028 30346 43325 30643 ne
rect 43325 30560 44802 30643
tri 44802 30560 45091 30849 sw
tri 45091 30560 45380 30849 ne
rect 45380 30560 47070 30849
tri 47070 30560 47360 30850 sw
tri 47360 30560 47650 30850 ne
rect 47650 30750 51410 30850
tri 51410 30750 51704 31044 sw
tri 51704 30750 51998 31044 ne
rect 51998 30750 70613 31044
rect 47650 30588 51704 30750
tri 51704 30588 51866 30750 sw
tri 51998 30588 52160 30750 ne
rect 52160 30588 70613 30750
rect 47650 30560 51866 30588
rect 43325 30346 45091 30560
rect 38916 30214 43028 30346
rect 34672 29932 38634 30214
tri 38634 29932 38916 30214 sw
tri 38916 29932 39198 30214 ne
rect 39198 30049 43028 30214
tri 43028 30049 43325 30346 sw
tri 43325 30049 43622 30346 ne
rect 43622 30271 45091 30346
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30271 47360 30560
rect 43622 30049 45380 30271
rect 39198 29932 43325 30049
tri 30136 25688 34380 29932 ne
tri 34380 29640 34672 29932 sw
tri 34672 29640 34964 29932 ne
rect 34964 29650 38916 29932
tri 38916 29650 39198 29932 sw
tri 39198 29650 39480 29932 ne
rect 39480 29851 43325 29932
tri 43325 29851 43523 30049 sw
tri 43622 29851 43820 30049 ne
rect 43820 29982 45380 30049
tri 45380 29982 45669 30271 sw
tri 45669 29982 45958 30271 ne
rect 45958 30270 47360 30271
tri 47360 30270 47650 30560 sw
tri 47650 30270 47940 30560 ne
rect 47940 30294 51866 30560
tri 51866 30294 52160 30588 sw
tri 52160 30294 52454 30588 ne
rect 52454 30294 70613 30588
rect 47940 30270 52160 30294
rect 45958 30000 47650 30270
tri 47650 30000 47920 30270 sw
tri 47940 30000 48210 30270 ne
rect 48210 30000 52160 30270
tri 52160 30000 52454 30294 sw
tri 52454 30000 52748 30294 ne
rect 52748 30056 70613 30294
rect 70669 30056 71000 32920
rect 52748 30000 71000 30056
rect 45958 29982 47920 30000
rect 43820 29851 45669 29982
rect 39480 29650 43523 29851
rect 34964 29640 39198 29650
rect 34380 29348 34672 29640
tri 34672 29348 34964 29640 sw
tri 34964 29348 35256 29640 ne
rect 35256 29452 39198 29640
tri 39198 29452 39396 29650 sw
tri 39480 29452 39678 29650 ne
rect 39678 29554 43523 29650
tri 43523 29554 43820 29851 sw
tri 43820 29554 44117 29851 ne
rect 44117 29693 45669 29851
tri 45669 29693 45958 29982 sw
tri 45958 29693 46247 29982 ne
rect 46247 29710 47920 29982
tri 47920 29710 48210 30000 sw
tri 48210 29710 48500 30000 ne
rect 48500 29800 52454 30000
tri 52454 29800 52654 30000 sw
rect 48500 29752 71000 29800
rect 48500 29710 70613 29752
rect 46247 29693 48210 29710
rect 44117 29554 45958 29693
rect 39678 29452 43820 29554
rect 35256 29348 39396 29452
rect 34380 29056 34964 29348
tri 34964 29056 35256 29348 sw
tri 35256 29056 35548 29348 ne
rect 35548 29170 39396 29348
tri 39396 29170 39678 29452 sw
tri 39678 29170 39960 29452 ne
rect 39960 29257 43820 29452
tri 43820 29257 44117 29554 sw
tri 44117 29257 44414 29554 ne
rect 44414 29538 45958 29554
tri 45958 29538 46113 29693 sw
tri 46247 29538 46402 29693 ne
rect 46402 29538 48210 29693
rect 44414 29257 46113 29538
rect 39960 29170 44117 29257
rect 35548 29056 39678 29170
rect 34380 28764 35256 29056
tri 35256 28764 35548 29056 sw
tri 35548 28764 35840 29056 ne
rect 35840 28888 39678 29056
tri 39678 28888 39960 29170 sw
tri 39960 28888 40242 29170 ne
rect 40242 28960 44117 29170
tri 44117 28960 44414 29257 sw
tri 44414 28960 44711 29257 ne
rect 44711 29249 46113 29257
tri 46113 29249 46402 29538 sw
tri 46402 29249 46691 29538 ne
rect 46691 29420 48210 29538
tri 48210 29420 48500 29710 sw
tri 48500 29420 48790 29710 ne
rect 48790 29420 70613 29710
rect 46691 29250 48500 29420
tri 48500 29250 48670 29420 sw
tri 48790 29250 48960 29420 ne
rect 48960 29250 70613 29420
rect 46691 29249 48670 29250
rect 44711 28960 46402 29249
tri 46402 28960 46691 29249 sw
tri 46691 28960 46980 29249 ne
rect 46980 28960 48670 29249
tri 48670 28960 48960 29250 sw
tri 48960 28960 49250 29250 ne
rect 49250 28960 70613 29250
rect 40242 28888 44414 28960
rect 35840 28764 39960 28888
rect 34380 28472 35548 28764
tri 35548 28472 35840 28764 sw
tri 35840 28472 36132 28764 ne
rect 36132 28606 39960 28764
tri 39960 28606 40242 28888 sw
tri 40242 28606 40524 28888 ne
rect 40524 28663 44414 28888
tri 44414 28663 44711 28960 sw
tri 44711 28663 45008 28960 ne
rect 45008 28869 46691 28960
tri 46691 28869 46782 28960 sw
tri 46980 28869 47071 28960 ne
rect 47071 28870 48960 28960
tri 48960 28870 49050 28960 sw
tri 49250 28870 49340 28960 ne
rect 49340 28870 70613 28960
rect 47071 28869 49050 28870
rect 45008 28663 46782 28869
rect 40524 28606 44711 28663
rect 36132 28472 40242 28606
rect 34380 28192 35840 28472
tri 35840 28192 36120 28472 sw
tri 36132 28192 36412 28472 ne
rect 36412 28324 40242 28472
tri 40242 28324 40524 28606 sw
tri 40524 28324 40806 28606 ne
rect 40806 28366 44711 28606
tri 44711 28366 45008 28663 sw
tri 45008 28366 45305 28663 ne
rect 45305 28580 46782 28663
tri 46782 28580 47071 28869 sw
tri 47071 28580 47360 28869 ne
rect 47360 28580 49050 28869
tri 49050 28580 49340 28870 sw
tri 49340 28580 49630 28870 ne
rect 49630 28580 70613 28870
rect 45305 28366 47071 28580
rect 40806 28324 45008 28366
rect 36412 28192 40524 28324
rect 34380 27900 36120 28192
tri 36120 27900 36412 28192 sw
tri 36412 27900 36704 28192 ne
rect 36704 28042 40524 28192
tri 40524 28042 40806 28324 sw
tri 40806 28042 41088 28324 ne
rect 41088 28069 45008 28324
tri 45008 28069 45305 28366 sw
tri 45305 28069 45602 28366 ne
rect 45602 28291 47071 28366
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28291 49340 28580
rect 45602 28069 47360 28291
rect 41088 28042 45305 28069
rect 36704 27900 40806 28042
rect 34380 27608 36412 27900
tri 36412 27608 36704 27900 sw
tri 36704 27608 36996 27900 ne
rect 36996 27760 40806 27900
tri 40806 27760 41088 28042 sw
tri 41088 27760 41370 28042 ne
rect 41370 27871 45305 28042
tri 45305 27871 45503 28069 sw
tri 45602 27871 45800 28069 ne
rect 45800 28002 47360 28069
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28290 49340 28291
tri 49340 28290 49630 28580 sw
tri 49630 28290 49920 28580 ne
rect 49920 28290 70613 28580
rect 47938 28002 49630 28290
rect 45800 27871 47649 28002
rect 41370 27760 45503 27871
rect 36996 27608 41088 27760
rect 34380 27316 36704 27608
tri 36704 27316 36996 27608 sw
tri 36996 27316 37288 27608 ne
rect 37288 27478 41088 27608
tri 41088 27478 41370 27760 sw
tri 41370 27478 41652 27760 ne
rect 41652 27574 45503 27760
tri 45503 27574 45800 27871 sw
tri 45800 27574 46097 27871 ne
rect 46097 27713 47649 27871
tri 47649 27713 47938 28002 sw
tri 47938 27713 48227 28002 ne
rect 48227 28000 49630 28002
tri 49630 28000 49920 28290 sw
tri 49920 28000 50210 28290 ne
rect 50210 28000 70613 28290
rect 48227 27713 49920 28000
rect 46097 27574 47938 27713
rect 41652 27478 45800 27574
rect 37288 27316 41370 27478
rect 34380 27024 36996 27316
tri 36996 27024 37288 27316 sw
tri 37288 27024 37580 27316 ne
rect 37580 27196 41370 27316
tri 41370 27196 41652 27478 sw
tri 41652 27196 41934 27478 ne
rect 41934 27277 45800 27478
tri 45800 27277 46097 27574 sw
tri 46097 27277 46394 27574 ne
rect 46394 27558 47938 27574
tri 47938 27558 48093 27713 sw
tri 48227 27558 48382 27713 ne
rect 48382 27710 49920 27713
tri 49920 27710 50210 28000 sw
tri 50210 27710 50500 28000 ne
rect 50500 27710 70613 28000
rect 48382 27560 50210 27710
tri 50210 27560 50360 27710 sw
tri 50500 27560 50650 27710 ne
rect 50650 27560 70613 27710
rect 48382 27558 50360 27560
rect 46394 27277 48093 27558
rect 41934 27196 46097 27277
rect 37580 27098 41652 27196
tri 41652 27098 41750 27196 sw
tri 41934 27098 42032 27196 ne
rect 42032 27098 46097 27196
rect 37580 27024 41750 27098
rect 34380 26732 37288 27024
tri 37288 26732 37580 27024 sw
tri 37580 26732 37872 27024 ne
rect 37872 26816 41750 27024
tri 41750 26816 42032 27098 sw
tri 42032 26816 42314 27098 ne
rect 42314 26980 46097 27098
tri 46097 26980 46394 27277 sw
tri 46394 26980 46691 27277 ne
rect 46691 27269 48093 27277
tri 48093 27269 48382 27558 sw
tri 48382 27269 48671 27558 ne
rect 48671 27270 50360 27558
tri 50360 27270 50650 27560 sw
tri 50650 27270 50940 27560 ne
rect 50940 27270 70613 27560
rect 48671 27269 50650 27270
rect 46691 26980 48382 27269
tri 48382 26980 48671 27269 sw
tri 48671 26980 48960 27269 ne
rect 48960 26980 50650 27269
tri 50650 26980 50940 27270 sw
tri 50940 26980 51230 27270 ne
rect 51230 26980 70613 27270
rect 42314 26816 46394 26980
rect 37872 26732 42032 26816
rect 34380 26440 37580 26732
tri 37580 26440 37872 26732 sw
tri 37872 26440 38164 26732 ne
rect 38164 26534 42032 26732
tri 42032 26534 42314 26816 sw
tri 42314 26534 42596 26816 ne
rect 42596 26683 46394 26816
tri 46394 26683 46691 26980 sw
tri 46691 26683 46988 26980 ne
rect 46988 26889 48671 26980
tri 48671 26889 48762 26980 sw
tri 48960 26889 49051 26980 ne
rect 49051 26889 50940 26980
rect 46988 26683 48762 26889
rect 42596 26534 46691 26683
rect 38164 26440 42314 26534
rect 34380 26272 37872 26440
tri 37872 26272 38040 26440 sw
tri 38164 26272 38332 26440 ne
rect 38332 26272 42314 26440
rect 34380 25980 38040 26272
tri 38040 25980 38332 26272 sw
tri 38332 25980 38624 26272 ne
rect 38624 26252 42314 26272
tri 42314 26252 42596 26534 sw
tri 42596 26252 42878 26534 ne
rect 42878 26386 46691 26534
tri 46691 26386 46988 26683 sw
tri 46988 26386 47285 26683 ne
rect 47285 26600 48762 26683
tri 48762 26600 49051 26889 sw
tri 49051 26600 49340 26889 ne
rect 49340 26800 50940 26889
tri 50940 26800 51120 26980 sw
tri 51230 26800 51410 26980 ne
rect 51410 26888 70613 26980
rect 70669 26888 71000 29752
rect 51410 26800 71000 26888
rect 49340 26600 51120 26800
tri 51120 26600 51320 26800 sw
rect 47285 26386 49051 26600
rect 42878 26252 46988 26386
rect 38624 25980 42596 26252
rect 34380 25688 38332 25980
tri 38332 25688 38624 25980 sw
tri 38624 25688 38916 25980 ne
rect 38916 25970 42596 25980
tri 42596 25970 42878 26252 sw
tri 42878 25970 43160 26252 ne
rect 43160 26089 46988 26252
tri 46988 26089 47285 26386 sw
tri 47285 26089 47582 26386 ne
rect 47582 26311 49051 26386
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47582 26089 49340 26311
rect 43160 25970 47285 26089
rect 38916 25688 42878 25970
tri 42878 25688 43160 25970 sw
tri 43160 25688 43442 25970 ne
rect 43442 25891 47285 25970
tri 47285 25891 47483 26089 sw
tri 47582 25891 47780 26089 ne
rect 47780 26022 49340 26089
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47780 25891 49629 26022
rect 43442 25688 47483 25891
tri 34380 21444 38624 25688 ne
tri 38624 25396 38916 25688 sw
tri 38916 25396 39208 25688 ne
rect 39208 25406 43160 25688
tri 43160 25406 43442 25688 sw
tri 43442 25406 43724 25688 ne
rect 43724 25594 47483 25688
tri 47483 25594 47780 25891 sw
tri 47780 25594 48077 25891 ne
rect 48077 25778 49629 25891
tri 49629 25778 49873 26022 sw
tri 49918 25778 50162 26022 ne
rect 50162 25778 71000 26022
rect 48077 25594 49873 25778
rect 43724 25406 47780 25594
rect 39208 25396 43442 25406
rect 38624 25104 38916 25396
tri 38916 25104 39208 25396 sw
tri 39208 25104 39500 25396 ne
rect 39500 25208 43442 25396
tri 43442 25208 43640 25406 sw
tri 43724 25208 43922 25406 ne
rect 43922 25297 47780 25406
tri 47780 25297 48077 25594 sw
tri 48077 25297 48374 25594 ne
rect 48374 25489 49873 25594
tri 49873 25489 50162 25778 sw
tri 50162 25489 50451 25778 ne
rect 50451 25489 71000 25778
rect 48374 25297 50162 25489
rect 43922 25208 48077 25297
rect 39500 25104 43640 25208
rect 38624 24812 39208 25104
tri 39208 24812 39500 25104 sw
tri 39500 24812 39792 25104 ne
rect 39792 24926 43640 25104
tri 43640 24926 43922 25208 sw
tri 43922 24926 44204 25208 ne
rect 44204 25000 48077 25208
tri 48077 25000 48374 25297 sw
tri 48374 25000 48671 25297 ne
rect 48671 25200 50162 25297
tri 50162 25200 50451 25489 sw
tri 50451 25200 50740 25489 ne
rect 50740 25200 71000 25489
rect 48671 25000 50451 25200
tri 50451 25000 50651 25200 sw
rect 44204 24926 48374 25000
rect 39792 24812 43922 24926
rect 38624 24520 39500 24812
tri 39500 24520 39792 24812 sw
tri 39792 24520 40084 24812 ne
rect 40084 24644 43922 24812
tri 43922 24644 44204 24926 sw
tri 44204 24644 44486 24926 ne
rect 44486 24703 48374 24926
tri 48374 24703 48671 25000 sw
tri 48671 24703 48968 25000 ne
rect 48968 24906 71000 25000
rect 48968 24703 70613 24906
rect 44486 24644 48671 24703
rect 40084 24520 44204 24644
rect 38624 24228 39792 24520
tri 39792 24228 40084 24520 sw
tri 40084 24228 40376 24520 ne
rect 40376 24362 44204 24520
tri 44204 24362 44486 24644 sw
tri 44486 24362 44768 24644 ne
rect 44768 24406 48671 24644
tri 48671 24406 48968 24703 sw
tri 48968 24406 49265 24703 ne
rect 49265 24406 70613 24703
rect 44768 24362 48968 24406
rect 40376 24228 44486 24362
rect 38624 23948 40084 24228
tri 40084 23948 40364 24228 sw
tri 40376 23948 40656 24228 ne
rect 40656 24080 44486 24228
tri 44486 24080 44768 24362 sw
tri 44768 24080 45050 24362 ne
rect 45050 24194 48968 24362
tri 48968 24194 49180 24406 sw
tri 49265 24194 49477 24406 ne
rect 49477 24194 70613 24406
rect 45050 24080 49180 24194
rect 40656 23948 44768 24080
rect 38624 23656 40364 23948
tri 40364 23656 40656 23948 sw
tri 40656 23656 40948 23948 ne
rect 40948 23798 44768 23948
tri 44768 23798 45050 24080 sw
tri 45050 23798 45332 24080 ne
rect 45332 23897 49180 24080
tri 49180 23897 49477 24194 sw
tri 49477 23897 49774 24194 ne
rect 49774 23897 70613 24194
rect 45332 23798 49477 23897
rect 40948 23656 45050 23798
rect 38624 23364 40656 23656
tri 40656 23364 40948 23656 sw
tri 40948 23364 41240 23656 ne
rect 41240 23516 45050 23656
tri 45050 23516 45332 23798 sw
tri 45332 23516 45614 23798 ne
rect 45614 23600 49477 23798
tri 49477 23600 49774 23897 sw
tri 49774 23600 50071 23897 ne
rect 50071 23706 70613 23897
rect 70669 23706 71000 24906
rect 50071 23600 71000 23706
rect 45614 23516 49774 23600
rect 41240 23364 45332 23516
rect 38624 23072 40948 23364
tri 40948 23072 41240 23364 sw
tri 41240 23072 41532 23364 ne
rect 41532 23234 45332 23364
tri 45332 23234 45614 23516 sw
tri 45614 23234 45896 23516 ne
rect 45896 23400 49774 23516
tri 49774 23400 49974 23600 sw
rect 45896 23234 71000 23400
rect 41532 23072 45614 23234
rect 38624 22780 41240 23072
tri 41240 22780 41532 23072 sw
tri 41532 22780 41824 23072 ne
rect 41824 22952 45614 23072
tri 45614 22952 45896 23234 sw
tri 45896 22952 46178 23234 ne
rect 46178 22952 71000 23234
rect 41824 22854 45896 22952
tri 45896 22854 45994 22952 sw
tri 46178 22854 46276 22952 ne
rect 46276 22854 71000 22952
rect 41824 22780 45994 22854
rect 38624 22488 41532 22780
tri 41532 22488 41824 22780 sw
tri 41824 22488 42116 22780 ne
rect 42116 22572 45994 22780
tri 45994 22572 46276 22854 sw
tri 46276 22572 46558 22854 ne
rect 46558 22572 71000 22854
rect 42116 22488 46276 22572
rect 38624 22196 41824 22488
tri 41824 22196 42116 22488 sw
tri 42116 22196 42408 22488 ne
rect 42408 22290 46276 22488
tri 46276 22290 46558 22572 sw
tri 46558 22290 46840 22572 ne
rect 46840 22290 71000 22572
rect 42408 22196 46558 22290
rect 38624 22028 42116 22196
tri 42116 22028 42284 22196 sw
tri 42408 22028 42576 22196 ne
rect 42576 22028 46558 22196
rect 38624 21736 42284 22028
tri 42284 21736 42576 22028 sw
tri 42576 21736 42868 22028 ne
rect 42868 22008 46558 22028
tri 46558 22008 46840 22290 sw
tri 46840 22008 47122 22290 ne
rect 47122 22008 71000 22290
rect 42868 21736 46840 22008
rect 38624 21444 42576 21736
tri 42576 21444 42868 21736 sw
tri 42868 21444 43160 21736 ne
rect 43160 21726 46840 21736
tri 46840 21726 47122 22008 sw
tri 47122 21726 47404 22008 ne
rect 47404 21726 71000 22008
rect 43160 21444 47122 21726
tri 47122 21444 47404 21726 sw
tri 47404 21444 47686 21726 ne
rect 47686 21444 71000 21726
tri 38624 17200 42868 21444 ne
tri 42868 21152 43160 21444 sw
tri 43160 21152 43452 21444 ne
rect 43452 21162 47404 21444
tri 47404 21162 47686 21444 sw
tri 47686 21162 47968 21444 ne
rect 47968 21162 71000 21444
rect 43452 21152 47686 21162
rect 42868 20860 43160 21152
tri 43160 20860 43452 21152 sw
tri 43452 20860 43744 21152 ne
rect 43744 20964 47686 21152
tri 47686 20964 47884 21162 sw
tri 47968 20964 48166 21162 ne
rect 48166 20964 71000 21162
rect 43744 20860 47884 20964
rect 42868 20568 43452 20860
tri 43452 20568 43744 20860 sw
tri 43744 20568 44036 20860 ne
rect 44036 20682 47884 20860
tri 47884 20682 48166 20964 sw
tri 48166 20682 48448 20964 ne
rect 48448 20682 71000 20964
rect 44036 20568 48166 20682
rect 42868 20276 43744 20568
tri 43744 20276 44036 20568 sw
tri 44036 20276 44328 20568 ne
rect 44328 20400 48166 20568
tri 48166 20400 48448 20682 sw
tri 48448 20400 48730 20682 ne
rect 48730 20400 71000 20682
rect 44328 20276 48448 20400
rect 42868 19984 44036 20276
tri 44036 19984 44328 20276 sw
tri 44328 19984 44620 20276 ne
rect 44620 20200 48448 20276
tri 48448 20200 48648 20400 sw
rect 44620 19984 71000 20200
rect 42868 19704 44328 19984
tri 44328 19704 44608 19984 sw
tri 44620 19704 44900 19984 ne
rect 44900 19704 71000 19984
rect 42868 19412 44608 19704
tri 44608 19412 44900 19704 sw
tri 44900 19412 45192 19704 ne
rect 45192 19412 71000 19704
rect 42868 19120 44900 19412
tri 44900 19120 45192 19412 sw
tri 45192 19120 45484 19412 ne
rect 45484 19120 71000 19412
rect 42868 18828 45192 19120
tri 45192 18828 45484 19120 sw
tri 45484 18828 45776 19120 ne
rect 45776 18828 71000 19120
rect 42868 18536 45484 18828
tri 45484 18536 45776 18828 sw
tri 45776 18536 46068 18828 ne
rect 46068 18536 71000 18828
rect 42868 18244 45776 18536
tri 45776 18244 46068 18536 sw
tri 46068 18244 46360 18536 ne
rect 46360 18244 71000 18536
rect 42868 17952 46068 18244
tri 46068 17952 46360 18244 sw
tri 46360 17952 46652 18244 ne
rect 46652 17952 71000 18244
rect 42868 17784 46360 17952
tri 46360 17784 46528 17952 sw
tri 46652 17784 46820 17952 ne
rect 46820 17784 71000 17952
rect 42868 17492 46528 17784
tri 46528 17492 46820 17784 sw
tri 46820 17492 47112 17784 ne
rect 47112 17492 71000 17784
rect 42868 17200 46820 17492
tri 46820 17200 47112 17492 sw
tri 47112 17200 47404 17492 ne
rect 47404 17200 71000 17492
tri 42868 14000 46068 17200 ne
rect 46068 17000 47112 17200
tri 47112 17000 47312 17200 sw
rect 46068 14000 71000 17000
use M1_PSUB_CDNS_40661953145669  M1_PSUB_CDNS_40661953145669_0
timestamp 1759194789
transform -1 0 58007 0 -1 13194
box 0 0 1 1
use M1_PSUB_CDNS_40661953145670  M1_PSUB_CDNS_40661953145670_0
timestamp 1759194789
transform 0 -1 69871 1 0 70385
box 0 0 1 1
use M1_PSUB_CDNS_40661953145671  M1_PSUB_CDNS_40661953145671_0
timestamp 1759194789
transform 1 0 70235 0 1 69871
box 0 0 1 1
use M1_PSUB_CDNS_40661953145672  M1_PSUB_CDNS_40661953145672_0
timestamp 1759194789
transform 0 -1 70899 1 0 41649
box 0 0 1 1
use M1_PSUB_CDNS_40661953145672  M1_PSUB_CDNS_40661953145672_1
timestamp 1759194789
transform 1 0 41636 0 1 70900
box 0 0 1 1
use M1_PSUB_CDNS_40661953145673  M1_PSUB_CDNS_40661953145673_0
timestamp 1759194789
transform 0 -1 13194 1 0 58004
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_0
timestamp 1759194789
transform 1 0 42317 0 1 15761
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_1
timestamp 1759194789
transform 1 0 42185 0 1 15893
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_2
timestamp 1759194789
transform 1 0 42977 0 1 15101
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_3
timestamp 1759194789
transform 1 0 44873 0 1 13233
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_4
timestamp 1759194789
transform 1 0 44693 0 1 13385
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_5
timestamp 1759194789
transform 1 0 44561 0 1 13517
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_6
timestamp 1759194789
transform 1 0 44429 0 1 13649
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_7
timestamp 1759194789
transform 1 0 44297 0 1 13781
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_8
timestamp 1759194789
transform 1 0 44165 0 1 13913
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_9
timestamp 1759194789
transform 1 0 44033 0 1 14045
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_10
timestamp 1759194789
transform 1 0 43901 0 1 14177
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_11
timestamp 1759194789
transform 1 0 43769 0 1 14309
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_12
timestamp 1759194789
transform 1 0 43637 0 1 14441
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_13
timestamp 1759194789
transform 1 0 43505 0 1 14573
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_14
timestamp 1759194789
transform 1 0 43373 0 1 14705
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_15
timestamp 1759194789
transform 1 0 43241 0 1 14837
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_16
timestamp 1759194789
transform 1 0 43109 0 1 14969
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_17
timestamp 1759194789
transform 1 0 42845 0 1 15233
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_18
timestamp 1759194789
transform 1 0 42713 0 1 15365
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_19
timestamp 1759194789
transform 1 0 42581 0 1 15497
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_20
timestamp 1759194789
transform 1 0 42449 0 1 15629
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_21
timestamp 1759194789
transform 1 0 33605 0 1 24473
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_22
timestamp 1759194789
transform 1 0 39017 0 1 19061
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_23
timestamp 1759194789
transform 1 0 38885 0 1 19193
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_24
timestamp 1759194789
transform 1 0 38753 0 1 19325
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_25
timestamp 1759194789
transform 1 0 38621 0 1 19457
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_26
timestamp 1759194789
transform 1 0 38489 0 1 19589
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_27
timestamp 1759194789
transform 1 0 38357 0 1 19721
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_28
timestamp 1759194789
transform 1 0 33737 0 1 24341
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_29
timestamp 1759194789
transform 1 0 33869 0 1 24209
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_30
timestamp 1759194789
transform 1 0 34001 0 1 24077
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_31
timestamp 1759194789
transform 1 0 34133 0 1 23945
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_32
timestamp 1759194789
transform 1 0 34265 0 1 23813
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_33
timestamp 1759194789
transform 1 0 34397 0 1 23681
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_34
timestamp 1759194789
transform 1 0 34529 0 1 23549
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_35
timestamp 1759194789
transform 1 0 34661 0 1 23417
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_36
timestamp 1759194789
transform 1 0 34793 0 1 23285
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_37
timestamp 1759194789
transform 1 0 33209 0 1 24869
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_38
timestamp 1759194789
transform 1 0 39413 0 1 18665
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_39
timestamp 1759194789
transform 1 0 41261 0 1 16817
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_40
timestamp 1759194789
transform 1 0 36245 0 1 21833
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_41
timestamp 1759194789
transform 1 0 37301 0 1 20777
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_42
timestamp 1759194789
transform 1 0 37169 0 1 20909
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_43
timestamp 1759194789
transform 1 0 37037 0 1 21041
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_44
timestamp 1759194789
transform 1 0 36905 0 1 21173
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_45
timestamp 1759194789
transform 1 0 36773 0 1 21305
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_46
timestamp 1759194789
transform 1 0 36641 0 1 21437
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_47
timestamp 1759194789
transform 1 0 36509 0 1 21569
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_48
timestamp 1759194789
transform 1 0 36377 0 1 21701
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_49
timestamp 1759194789
transform 1 0 32945 0 1 25133
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_50
timestamp 1759194789
transform 1 0 32813 0 1 25265
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_51
timestamp 1759194789
transform 1 0 32681 0 1 25397
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_52
timestamp 1759194789
transform 1 0 32549 0 1 25529
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_53
timestamp 1759194789
transform 1 0 32417 0 1 25661
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_54
timestamp 1759194789
transform 1 0 32285 0 1 25793
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_55
timestamp 1759194789
transform 1 0 32153 0 1 25925
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_56
timestamp 1759194789
transform 1 0 32021 0 1 26057
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_57
timestamp 1759194789
transform 1 0 31889 0 1 26189
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_58
timestamp 1759194789
transform 1 0 31757 0 1 26321
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_59
timestamp 1759194789
transform 1 0 31625 0 1 26453
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_60
timestamp 1759194789
transform 1 0 31493 0 1 26585
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_61
timestamp 1759194789
transform 1 0 31361 0 1 26717
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_62
timestamp 1759194789
transform 1 0 31229 0 1 26849
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_63
timestamp 1759194789
transform 1 0 33077 0 1 25001
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_64
timestamp 1759194789
transform 1 0 30965 0 1 27113
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_65
timestamp 1759194789
transform 1 0 30833 0 1 27245
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_66
timestamp 1759194789
transform 1 0 30701 0 1 27377
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_67
timestamp 1759194789
transform 1 0 31097 0 1 26981
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_68
timestamp 1759194789
transform 1 0 36113 0 1 21965
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_69
timestamp 1759194789
transform 1 0 35981 0 1 22097
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_70
timestamp 1759194789
transform 1 0 35849 0 1 22229
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_71
timestamp 1759194789
transform 1 0 35717 0 1 22361
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_72
timestamp 1759194789
transform 1 0 35585 0 1 22493
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_73
timestamp 1759194789
transform 1 0 35453 0 1 22625
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_74
timestamp 1759194789
transform 1 0 35321 0 1 22757
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_75
timestamp 1759194789
transform 1 0 35189 0 1 22889
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_76
timestamp 1759194789
transform 1 0 34925 0 1 23153
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_77
timestamp 1759194789
transform 1 0 41921 0 1 16157
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_78
timestamp 1759194789
transform 1 0 41789 0 1 16289
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_79
timestamp 1759194789
transform 1 0 41657 0 1 16421
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_80
timestamp 1759194789
transform 1 0 41525 0 1 16553
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_81
timestamp 1759194789
transform 1 0 41393 0 1 16685
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_82
timestamp 1759194789
transform 1 0 39281 0 1 18797
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_83
timestamp 1759194789
transform 1 0 41129 0 1 16949
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_84
timestamp 1759194789
transform 1 0 40997 0 1 17081
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_85
timestamp 1759194789
transform 1 0 40865 0 1 17213
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_86
timestamp 1759194789
transform 1 0 40733 0 1 17345
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_87
timestamp 1759194789
transform 1 0 40601 0 1 17477
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_88
timestamp 1759194789
transform 1 0 40469 0 1 17609
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_89
timestamp 1759194789
transform 1 0 40337 0 1 17741
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_90
timestamp 1759194789
transform 1 0 40205 0 1 17873
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_91
timestamp 1759194789
transform 1 0 40073 0 1 18005
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_92
timestamp 1759194789
transform 1 0 39941 0 1 18137
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_93
timestamp 1759194789
transform 1 0 39809 0 1 18269
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_94
timestamp 1759194789
transform 1 0 39677 0 1 18401
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_95
timestamp 1759194789
transform 1 0 38225 0 1 19853
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_96
timestamp 1759194789
transform 1 0 38093 0 1 19985
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_97
timestamp 1759194789
transform 1 0 37961 0 1 20117
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_98
timestamp 1759194789
transform 1 0 37829 0 1 20249
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_99
timestamp 1759194789
transform 1 0 37697 0 1 20381
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_100
timestamp 1759194789
transform 1 0 37565 0 1 20513
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_101
timestamp 1759194789
transform 1 0 37433 0 1 20645
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_102
timestamp 1759194789
transform 1 0 39545 0 1 18533
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_103
timestamp 1759194789
transform 1 0 35057 0 1 23021
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_104
timestamp 1759194789
transform 1 0 39149 0 1 18929
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_105
timestamp 1759194789
transform 1 0 33341 0 1 24737
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_106
timestamp 1759194789
transform 1 0 33473 0 1 24605
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_107
timestamp 1759194789
transform 1 0 18689 0 1 39389
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_108
timestamp 1759194789
transform 1 0 23969 0 1 34109
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_109
timestamp 1759194789
transform 1 0 23045 0 1 35033
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_110
timestamp 1759194789
transform 1 0 23309 0 1 34769
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_111
timestamp 1759194789
transform 1 0 23441 0 1 34637
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_112
timestamp 1759194789
transform 1 0 23573 0 1 34505
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_113
timestamp 1759194789
transform 1 0 23705 0 1 34373
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_114
timestamp 1759194789
transform 1 0 23837 0 1 34241
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_115
timestamp 1759194789
transform 1 0 24101 0 1 33977
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_116
timestamp 1759194789
transform 1 0 24233 0 1 33845
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_117
timestamp 1759194789
transform 1 0 24365 0 1 33713
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_118
timestamp 1759194789
transform 1 0 24497 0 1 33581
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_119
timestamp 1759194789
transform 1 0 24629 0 1 33449
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_120
timestamp 1759194789
transform 1 0 24761 0 1 33317
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_121
timestamp 1759194789
transform 1 0 25025 0 1 33053
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_122
timestamp 1759194789
transform 1 0 23177 0 1 34901
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_123
timestamp 1759194789
transform 1 0 22913 0 1 35165
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_124
timestamp 1759194789
transform 1 0 22781 0 1 35297
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_125
timestamp 1759194789
transform 1 0 22649 0 1 35429
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_126
timestamp 1759194789
transform 1 0 22517 0 1 35561
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_127
timestamp 1759194789
transform 1 0 22385 0 1 35693
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_128
timestamp 1759194789
transform 1 0 22253 0 1 35825
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_129
timestamp 1759194789
transform 1 0 22121 0 1 35957
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_130
timestamp 1759194789
transform 1 0 21989 0 1 36089
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_131
timestamp 1759194789
transform 1 0 21857 0 1 36221
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_132
timestamp 1759194789
transform 1 0 21725 0 1 36353
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_133
timestamp 1759194789
transform 1 0 21593 0 1 36485
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_134
timestamp 1759194789
transform 1 0 21461 0 1 36617
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_135
timestamp 1759194789
transform 1 0 21329 0 1 36749
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_136
timestamp 1759194789
transform 1 0 21065 0 1 37013
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_137
timestamp 1759194789
transform 1 0 24893 0 1 33185
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_138
timestamp 1759194789
transform 1 0 18557 0 1 39521
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_139
timestamp 1759194789
transform 1 0 18425 0 1 39653
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_140
timestamp 1759194789
transform 1 0 18293 0 1 39785
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_141
timestamp 1759194789
transform 1 0 18161 0 1 39917
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_142
timestamp 1759194789
transform 1 0 16973 0 1 41105
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_143
timestamp 1759194789
transform 1 0 18029 0 1 40049
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_144
timestamp 1759194789
transform 1 0 17897 0 1 40181
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_145
timestamp 1759194789
transform 1 0 17765 0 1 40313
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_146
timestamp 1759194789
transform 1 0 17633 0 1 40445
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_147
timestamp 1759194789
transform 1 0 17501 0 1 40577
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_148
timestamp 1759194789
transform 1 0 17369 0 1 40709
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_149
timestamp 1759194789
transform 1 0 27401 0 1 30677
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_150
timestamp 1759194789
transform 1 0 27269 0 1 30809
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_151
timestamp 1759194789
transform 1 0 27137 0 1 30941
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_152
timestamp 1759194789
transform 1 0 21197 0 1 36881
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_153
timestamp 1759194789
transform 1 0 26873 0 1 31205
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_154
timestamp 1759194789
transform 1 0 26741 0 1 31337
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_155
timestamp 1759194789
transform 1 0 26609 0 1 31469
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_156
timestamp 1759194789
transform 1 0 26477 0 1 31601
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_157
timestamp 1759194789
transform 1 0 26345 0 1 31733
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_158
timestamp 1759194789
transform 1 0 26213 0 1 31865
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_159
timestamp 1759194789
transform 1 0 26081 0 1 31997
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_160
timestamp 1759194789
transform 1 0 25949 0 1 32129
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_161
timestamp 1759194789
transform 1 0 25817 0 1 32261
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_162
timestamp 1759194789
transform 1 0 25685 0 1 32393
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_163
timestamp 1759194789
transform 1 0 25553 0 1 32525
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_164
timestamp 1759194789
transform 1 0 25421 0 1 32657
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_165
timestamp 1759194789
transform 1 0 25289 0 1 32789
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_166
timestamp 1759194789
transform 1 0 25157 0 1 32921
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_167
timestamp 1759194789
transform 1 0 27005 0 1 31073
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_168
timestamp 1759194789
transform 1 0 17105 0 1 40973
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_169
timestamp 1759194789
transform 1 0 16841 0 1 41237
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_170
timestamp 1759194789
transform 1 0 16709 0 1 41369
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_171
timestamp 1759194789
transform 1 0 16577 0 1 41501
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_172
timestamp 1759194789
transform 1 0 16445 0 1 41633
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_173
timestamp 1759194789
transform 1 0 16313 0 1 41765
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_174
timestamp 1759194789
transform 1 0 16181 0 1 41897
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_175
timestamp 1759194789
transform 1 0 19085 0 1 38993
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_176
timestamp 1759194789
transform 1 0 20933 0 1 37145
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_177
timestamp 1759194789
transform 1 0 20801 0 1 37277
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_178
timestamp 1759194789
transform 1 0 20669 0 1 37409
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_179
timestamp 1759194789
transform 1 0 20537 0 1 37541
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_180
timestamp 1759194789
transform 1 0 20405 0 1 37673
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_181
timestamp 1759194789
transform 1 0 20273 0 1 37805
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_182
timestamp 1759194789
transform 1 0 20141 0 1 37937
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_183
timestamp 1759194789
transform 1 0 20009 0 1 38069
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_184
timestamp 1759194789
transform 1 0 19877 0 1 38201
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_185
timestamp 1759194789
transform 1 0 19745 0 1 38333
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_186
timestamp 1759194789
transform 1 0 19613 0 1 38465
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_187
timestamp 1759194789
transform 1 0 19481 0 1 38597
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_188
timestamp 1759194789
transform 1 0 19349 0 1 38729
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_189
timestamp 1759194789
transform 1 0 19217 0 1 38861
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_190
timestamp 1759194789
transform 1 0 17237 0 1 40841
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_191
timestamp 1759194789
transform 1 0 18953 0 1 39125
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_192
timestamp 1759194789
transform 1 0 18821 0 1 39257
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_193
timestamp 1759194789
transform 1 0 29117 0 1 28961
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_194
timestamp 1759194789
transform 1 0 28985 0 1 29093
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_195
timestamp 1759194789
transform 1 0 28721 0 1 29357
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_196
timestamp 1759194789
transform 1 0 28589 0 1 29489
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_197
timestamp 1759194789
transform 1 0 28457 0 1 29621
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_198
timestamp 1759194789
transform 1 0 28325 0 1 29753
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_199
timestamp 1759194789
transform 1 0 28193 0 1 29885
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_200
timestamp 1759194789
transform 1 0 28061 0 1 30017
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_201
timestamp 1759194789
transform 1 0 27929 0 1 30149
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_202
timestamp 1759194789
transform 1 0 27797 0 1 30281
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_203
timestamp 1759194789
transform 1 0 27665 0 1 30413
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_204
timestamp 1759194789
transform 1 0 29249 0 1 28829
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_205
timestamp 1759194789
transform 1 0 28853 0 1 29225
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_206
timestamp 1759194789
transform 1 0 29513 0 1 28565
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_207
timestamp 1759194789
transform 1 0 30437 0 1 27641
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_208
timestamp 1759194789
transform 1 0 30305 0 1 27773
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_209
timestamp 1759194789
transform 1 0 30173 0 1 27905
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_210
timestamp 1759194789
transform 1 0 30041 0 1 28037
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_211
timestamp 1759194789
transform 1 0 29909 0 1 28169
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_212
timestamp 1759194789
transform 1 0 29777 0 1 28301
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_213
timestamp 1759194789
transform 1 0 29645 0 1 28433
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_214
timestamp 1759194789
transform 1 0 29381 0 1 28697
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_215
timestamp 1759194789
transform 1 0 27533 0 1 30545
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_216
timestamp 1759194789
transform 1 0 30569 0 1 27509
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_217
timestamp 1759194789
transform 1 0 13937 0 1 44141
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_218
timestamp 1759194789
transform 1 0 13805 0 1 44273
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_219
timestamp 1759194789
transform 1 0 13673 0 1 44405
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_220
timestamp 1759194789
transform 1 0 13541 0 1 44537
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_221
timestamp 1759194789
transform 1 0 13409 0 1 44669
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_222
timestamp 1759194789
transform 1 0 13277 0 1 44801
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_223
timestamp 1759194789
transform 1 0 15125 0 1 42953
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_224
timestamp 1759194789
transform 1 0 15917 0 1 42161
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_225
timestamp 1759194789
transform 1 0 15785 0 1 42293
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_226
timestamp 1759194789
transform 1 0 15653 0 1 42425
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_227
timestamp 1759194789
transform 1 0 15521 0 1 42557
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_228
timestamp 1759194789
transform 1 0 15389 0 1 42689
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_229
timestamp 1759194789
transform 1 0 15257 0 1 42821
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_230
timestamp 1759194789
transform 1 0 14993 0 1 43085
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_231
timestamp 1759194789
transform 1 0 14861 0 1 43217
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_232
timestamp 1759194789
transform 1 0 14729 0 1 43349
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_233
timestamp 1759194789
transform 1 0 14597 0 1 43481
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_234
timestamp 1759194789
transform 1 0 14465 0 1 43613
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_235
timestamp 1759194789
transform 1 0 14333 0 1 43745
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_236
timestamp 1759194789
transform 1 0 14201 0 1 43877
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_237
timestamp 1759194789
transform 1 0 14069 0 1 44009
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_238
timestamp 1759194789
transform 1 0 16049 0 1 42029
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_239
timestamp 1759194789
transform 1 0 42053 0 1 16025
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_0
timestamp 1759194789
transform 1 0 70641 0 1 24306
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_1
timestamp 1759194789
transform 1 0 70641 0 1 67516
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_2
timestamp 1759194789
transform 1 0 70641 0 1 59520
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_3
timestamp 1759194789
transform 1 0 70641 0 1 54702
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_4
timestamp 1759194789
transform 1 0 70641 0 1 53122
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_5
timestamp 1759194789
transform 1 0 70641 0 1 56310
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_6
timestamp 1759194789
transform 1 0 70641 0 1 41897
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_0
timestamp 1759194789
transform 1 0 70641 0 1 28320
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_1
timestamp 1759194789
transform 1 0 70641 0 1 31488
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_2
timestamp 1759194789
transform 1 0 70641 0 1 34700
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_3
timestamp 1759194789
transform 1 0 70641 0 1 37900
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_4
timestamp 1759194789
transform 1 0 70641 0 1 44307
box 0 0 1 1
<< labels >>
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 1 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 2 nsew
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 4 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 4 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 4 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 4 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 4 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 2 nsew
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 1 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 4 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 4 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 4 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 4 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 4 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 4 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 4 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string GDS_END 17211668
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17193356
string path 1687.500 1775.000 1687.500 1710.075 1710.075 1687.500 1775.000 1687.500 
<< end >>
