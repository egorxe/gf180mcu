magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
use alatch_512x8m81  alatch_512x8m81_0
timestamp 1762296095
transform 1 0 70 0 1 -632
box -90 -1 1692 2968
use M1_NWELL14_512x8m81  M1_NWELL14_512x8m81_0
timestamp 1762296095
transform 1 0 334 0 1 5060
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_0
timestamp 1762296095
transform 1 0 1151 0 1 6529
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81  M1_POLY2$$46559276_512x8m81_1
timestamp 1762296095
transform 1 0 641 0 1 6529
box 0 0 1 1
use M1_PSUB$$47818796_512x8m81  M1_PSUB$$47818796_512x8m81_0
timestamp 1762296095
transform 1 0 395 0 1 7252
box 0 0 1 1
use M2_M1$$34864172_512x8m81  M2_M1$$34864172_512x8m81_0
timestamp 1762296095
transform 1 0 591 0 1 6529
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1762296095
transform 1 0 485 0 1 1489
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1762296095
transform 1 0 922 0 1 3852
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1762296095
transform 1 0 1436 0 1 3852
box 0 0 1 1
use M2_M1$$43377708_512x8m81  M2_M1$$43377708_512x8m81_0
timestamp 1762296095
transform 1 0 1219 0 1 5722
box 0 0 1 1
use M2_M1$$43377708_512x8m81  M2_M1$$43377708_512x8m81_1
timestamp 1762296095
transform 1 0 705 0 1 5722
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1762296095
transform 1 0 485 0 1 7424
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1762296095
transform 1 0 692 0 1 7424
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1762296095
transform 1 0 1212 0 1 7424
box 0 0 1 1
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_0
timestamp 1762296095
transform 1 0 1698 0 1 4096
box 0 0 1 1
use M3_M2$$43368492_512x8m81  M3_M2$$43368492_512x8m81_1
timestamp 1762296095
transform 1 0 1208 0 1 3620
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1762296095
transform 1 0 485 0 1 7424
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1762296095
transform 1 0 692 0 1 7424
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1762296095
transform 1 0 1212 0 1 7424
box 0 0 1 1
use M3_M2$$47334444_512x8m81  M3_M2$$47334444_512x8m81_0
timestamp 1762296095
transform 1 0 1219 0 1 5722
box 0 0 1 1
use M3_M2$$47334444_512x8m81  M3_M2$$47334444_512x8m81_1
timestamp 1762296095
transform 1 0 705 0 1 5722
box 0 0 1 1
use nmos_1p2$$47514668_512x8m81  nmos_1p2$$47514668_512x8m81_0
timestamp 1762296095
transform 1 0 1296 0 1 6670
box -31 0 -30 1
use nmos_1p2$$47514668_512x8m81  nmos_1p2$$47514668_512x8m81_1
timestamp 1762296095
transform 1 0 782 0 1 6670
box -31 0 -30 1
use pmos_1p2$$46887980_512x8m81  pmos_1p2$$46887980_512x8m81_0
timestamp 1762296095
transform 1 0 1296 0 1 3668
box -31 0 -30 1
use pmos_1p2$$46887980_512x8m81  pmos_1p2$$46887980_512x8m81_1
timestamp 1762296095
transform 1 0 782 0 1 3668
box -31 0 -30 1
<< properties >>
string GDS_END 827280
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 824622
<< end >>
