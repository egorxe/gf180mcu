magic
tech gf180mcuD
timestamp 1759194789
<< properties >>
string GDS_END 17594498
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17592126
<< end >>
