magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
<< metal1 >>
rect 2272 34614 2372 34659
rect 2272 33837 2296 34614
rect 2284 33834 2296 33837
rect 2348 33837 2372 34614
rect 7620 34632 7696 34644
rect 7620 34268 7632 34632
rect 7684 34268 7696 34632
rect 7620 34256 7696 34268
rect 13072 34614 13282 34659
rect 13072 33837 13096 34614
rect 2348 33834 2360 33837
rect 2284 33822 2360 33834
rect 13084 33834 13096 33837
rect 13148 33837 13282 34614
rect 18400 34632 18516 34659
rect 18400 34268 18432 34632
rect 18484 34268 18516 34632
rect 18400 33981 18516 34268
rect 23512 34614 23612 34659
rect 23512 33837 23536 34614
rect 13148 33834 13160 33837
rect 13084 33822 13160 33834
rect 23524 33834 23536 33837
rect 23588 33837 23612 34614
rect 61740 34614 61948 34659
rect 61740 33837 61872 34614
rect 23588 33834 23600 33837
rect 23524 33822 23600 33834
rect 61860 33834 61872 33837
rect 61924 33837 61948 34614
rect 67176 34632 67292 34659
rect 67176 34268 67208 34632
rect 67260 34268 67292 34632
rect 67176 33981 67292 34268
rect 72648 34614 72858 34659
rect 61924 33834 61936 33837
rect 61860 33822 61936 33834
rect 72648 33834 72672 34614
rect 72724 33834 72858 34614
rect 72648 33763 72858 33834
rect 77879 34632 78084 34659
rect 77879 34268 78008 34632
rect 78060 34268 78084 34632
rect 77879 33811 78084 34268
rect 83088 34614 83188 34659
rect 83088 34005 83112 34614
rect 82716 33834 83112 34005
rect 83164 33834 83188 34614
rect 82716 33722 83188 33834
<< via1 >>
rect 2296 33834 2348 34614
rect 7632 34268 7684 34632
rect 13096 33834 13148 34614
rect 18432 34268 18484 34632
rect 23536 33834 23588 34614
rect 61872 33834 61924 34614
rect 67208 34268 67260 34632
rect 72672 33834 72724 34614
rect 78008 34268 78060 34632
rect 83112 33834 83164 34614
<< metal2 >>
rect 7672 35034 7772 35222
rect 18472 35034 18572 35222
rect 67248 35034 67348 35222
rect 78048 35034 78148 35222
rect 7608 34934 7772 35034
rect 18408 34934 18572 35034
rect 67184 34934 67348 35034
rect 77984 34934 78148 35034
rect 7608 34632 7708 34934
rect 2284 34614 2360 34626
rect 2284 33834 2296 34614
rect 2348 33834 2360 34614
rect 7608 34268 7632 34632
rect 7684 34268 7708 34632
rect 18408 34632 18508 34934
rect 7608 34245 7708 34268
rect 13084 34614 13160 34626
rect 2284 33822 2360 33834
rect 13084 33834 13096 34614
rect 13148 33834 13160 34614
rect 18408 34268 18432 34632
rect 18484 34268 18508 34632
rect 18408 34245 18508 34268
rect 23524 34614 23600 34626
rect 13084 33822 13160 33834
rect 23524 33834 23536 34614
rect 23588 33834 23600 34614
rect 23524 33822 23600 33834
rect 1912 28330 2012 32592
rect 12712 32366 12812 32592
rect 12712 32266 13049 32366
rect 12955 31889 13049 32266
rect 23872 31965 23972 32592
rect 23755 31865 23972 31965
rect 1912 28274 1934 28330
rect 1990 28274 2012 28330
rect 1912 28214 2012 28274
rect 1912 28158 1934 28214
rect 1990 28158 2012 28214
rect 1912 28098 2012 28158
rect 1912 28042 1934 28098
rect 1990 28042 2012 28098
rect 1912 27982 2012 28042
rect 1912 27926 1934 27982
rect 1990 27926 2012 27982
rect 1912 27866 2012 27926
rect 1912 27810 1934 27866
rect 1990 27810 2012 27866
rect 1912 27750 2012 27810
rect 12571 28377 12647 28387
rect 12571 28321 12581 28377
rect 12637 28321 12647 28377
rect 12571 28265 12647 28321
rect 12571 28209 12581 28265
rect 12637 28209 12647 28265
rect 12571 28153 12647 28209
rect 12571 28097 12581 28153
rect 12637 28097 12647 28153
rect 12571 28041 12647 28097
rect 12571 27985 12581 28041
rect 12637 27985 12647 28041
rect 12571 27929 12647 27985
rect 12571 27873 12581 27929
rect 12637 27873 12647 27929
rect 12571 27817 12647 27873
rect 12571 27761 12581 27817
rect 12637 27761 12647 27817
rect 12571 27751 12647 27761
rect 12964 28377 13040 28387
rect 12964 28321 12974 28377
rect 13030 28321 13040 28377
rect 12964 28265 13040 28321
rect 12964 28209 12974 28265
rect 13030 28209 13040 28265
rect 12964 28153 13040 28209
rect 12964 28097 12974 28153
rect 13030 28097 13040 28153
rect 12964 28041 13040 28097
rect 12964 27985 12974 28041
rect 13030 27985 13040 28041
rect 12964 27929 13040 27985
rect 12964 27873 12974 27929
rect 13030 27873 13040 27929
rect 12964 27817 13040 27873
rect 12964 27761 12974 27817
rect 13030 27761 13040 27817
rect 12964 27751 13040 27761
rect 23371 28377 23447 28387
rect 23371 28321 23381 28377
rect 23437 28321 23447 28377
rect 23371 28265 23447 28321
rect 23371 28209 23381 28265
rect 23437 28209 23447 28265
rect 23371 28153 23447 28209
rect 23371 28097 23381 28153
rect 23437 28097 23447 28153
rect 23371 28041 23447 28097
rect 23371 27985 23381 28041
rect 23437 27985 23447 28041
rect 23371 27929 23447 27985
rect 23371 27873 23381 27929
rect 23437 27873 23447 27929
rect 23371 27817 23447 27873
rect 23371 27761 23381 27817
rect 23437 27761 23447 27817
rect 23371 27751 23447 27761
rect 23764 28377 23840 28387
rect 23764 28321 23774 28377
rect 23830 28321 23840 28377
rect 23764 28265 23840 28321
rect 23764 28209 23774 28265
rect 23830 28209 23840 28265
rect 23764 28153 23840 28209
rect 23764 28097 23774 28153
rect 23830 28097 23840 28153
rect 23764 28041 23840 28097
rect 23764 27985 23774 28041
rect 23830 27985 23840 28041
rect 23764 27929 23840 27985
rect 23764 27873 23774 27929
rect 23830 27873 23840 27929
rect 23764 27817 23840 27873
rect 23764 27761 23774 27817
rect 23830 27761 23840 27817
rect 23764 27751 23840 27761
rect 61487 28330 61587 34760
rect 67184 34632 67284 34934
rect 61860 34614 61936 34626
rect 61860 33834 61872 34614
rect 61924 33834 61936 34614
rect 67184 34268 67208 34632
rect 67260 34268 67284 34632
rect 67184 34245 67284 34268
rect 61860 33822 61936 33834
rect 72288 32366 72388 34758
rect 77984 34632 78084 34934
rect 72660 34614 72736 34626
rect 72660 33834 72672 34614
rect 72724 33834 72736 34614
rect 77984 34268 78008 34632
rect 78060 34268 78084 34632
rect 77984 34245 78084 34268
rect 83100 34614 83176 34626
rect 72660 33822 72736 33834
rect 83100 33834 83112 34614
rect 83164 33834 83176 34614
rect 83100 33822 83176 33834
rect 72288 32266 72625 32366
rect 72531 31889 72625 32266
rect 83448 31965 83548 32592
rect 83331 31865 83548 31965
rect 61487 28274 61509 28330
rect 61565 28274 61587 28330
rect 61487 28214 61587 28274
rect 61487 28158 61509 28214
rect 61565 28158 61587 28214
rect 61487 28098 61587 28158
rect 61487 28042 61509 28098
rect 61565 28042 61587 28098
rect 61487 27982 61587 28042
rect 61487 27926 61509 27982
rect 61565 27926 61587 27982
rect 61487 27866 61587 27926
rect 61487 27810 61509 27866
rect 61565 27810 61587 27866
rect 1912 27694 1934 27750
rect 1990 27694 2012 27750
rect 1912 27634 2012 27694
rect 1912 27578 1934 27634
rect 1990 27578 2012 27634
rect 1912 27518 2012 27578
rect 1912 27462 1934 27518
rect 1990 27462 2012 27518
rect 1912 27402 2012 27462
rect 1912 27346 1934 27402
rect 1990 27346 2012 27402
rect 1912 27286 2012 27346
rect 61487 27750 61587 27810
rect 72147 28377 72223 28387
rect 72147 28321 72157 28377
rect 72213 28321 72223 28377
rect 72147 28265 72223 28321
rect 72147 28209 72157 28265
rect 72213 28209 72223 28265
rect 72147 28153 72223 28209
rect 72147 28097 72157 28153
rect 72213 28097 72223 28153
rect 72147 28041 72223 28097
rect 72147 27985 72157 28041
rect 72213 27985 72223 28041
rect 72147 27929 72223 27985
rect 72147 27873 72157 27929
rect 72213 27873 72223 27929
rect 72147 27817 72223 27873
rect 72147 27761 72157 27817
rect 72213 27761 72223 27817
rect 72147 27751 72223 27761
rect 72540 28377 72616 28387
rect 72540 28321 72550 28377
rect 72606 28321 72616 28377
rect 72540 28265 72616 28321
rect 72540 28209 72550 28265
rect 72606 28209 72616 28265
rect 72540 28153 72616 28209
rect 72540 28097 72550 28153
rect 72606 28097 72616 28153
rect 72540 28041 72616 28097
rect 72540 27985 72550 28041
rect 72606 27985 72616 28041
rect 72540 27929 72616 27985
rect 72540 27873 72550 27929
rect 72606 27873 72616 27929
rect 72540 27817 72616 27873
rect 72540 27761 72550 27817
rect 72606 27761 72616 27817
rect 72540 27751 72616 27761
rect 82947 28377 83023 28387
rect 82947 28321 82957 28377
rect 83013 28321 83023 28377
rect 82947 28265 83023 28321
rect 82947 28209 82957 28265
rect 83013 28209 83023 28265
rect 82947 28153 83023 28209
rect 82947 28097 82957 28153
rect 83013 28097 83023 28153
rect 82947 28041 83023 28097
rect 82947 27985 82957 28041
rect 83013 27985 83023 28041
rect 82947 27929 83023 27985
rect 82947 27873 82957 27929
rect 83013 27873 83023 27929
rect 82947 27817 83023 27873
rect 82947 27761 82957 27817
rect 83013 27761 83023 27817
rect 82947 27751 83023 27761
rect 83340 28377 83416 28387
rect 83340 28321 83350 28377
rect 83406 28321 83416 28377
rect 83340 28265 83416 28321
rect 83340 28209 83350 28265
rect 83406 28209 83416 28265
rect 83340 28153 83416 28209
rect 83340 28097 83350 28153
rect 83406 28097 83416 28153
rect 83340 28041 83416 28097
rect 83340 27985 83350 28041
rect 83406 27985 83416 28041
rect 83340 27929 83416 27985
rect 83340 27873 83350 27929
rect 83406 27873 83416 27929
rect 83340 27817 83416 27873
rect 83340 27761 83350 27817
rect 83406 27761 83416 27817
rect 83340 27751 83416 27761
rect 61487 27694 61509 27750
rect 61565 27694 61587 27750
rect 61487 27634 61587 27694
rect 61487 27578 61509 27634
rect 61565 27578 61587 27634
rect 61487 27518 61587 27578
rect 61487 27462 61509 27518
rect 61565 27462 61587 27518
rect 61487 27402 61587 27462
rect 61487 27346 61509 27402
rect 61565 27346 61587 27402
rect 1912 27230 1934 27286
rect 1990 27230 2012 27286
rect 1912 27170 2012 27230
rect 1912 27114 1934 27170
rect 1990 27114 2012 27170
rect 1912 27054 2012 27114
rect 1912 26998 1934 27054
rect 1990 26998 2012 27054
rect 1912 26938 2012 26998
rect 1912 26882 1934 26938
rect 1990 26882 2012 26938
rect 1912 26822 2012 26882
rect 1912 26766 1934 26822
rect 1990 26766 2012 26822
rect 1912 26706 2012 26766
rect 1912 26650 1934 26706
rect 1990 26650 2012 26706
rect 1912 26590 2012 26650
rect 1912 26534 1934 26590
rect 1990 26534 2012 26590
rect 1912 26265 2012 26534
rect 12571 27302 12647 27312
rect 12571 27246 12581 27302
rect 12637 27246 12647 27302
rect 12571 27190 12647 27246
rect 12571 27134 12581 27190
rect 12637 27134 12647 27190
rect 12571 27078 12647 27134
rect 12571 27022 12581 27078
rect 12637 27022 12647 27078
rect 12571 26966 12647 27022
rect 12571 26910 12581 26966
rect 12637 26910 12647 26966
rect 12571 26854 12647 26910
rect 12571 26798 12581 26854
rect 12637 26798 12647 26854
rect 12571 26742 12647 26798
rect 12571 26686 12581 26742
rect 12637 26686 12647 26742
rect 12571 26630 12647 26686
rect 12571 26574 12581 26630
rect 12637 26574 12647 26630
rect 12571 26518 12647 26574
rect 12571 26462 12581 26518
rect 12637 26462 12647 26518
rect 12571 26452 12647 26462
rect 12964 27302 13040 27312
rect 12964 27246 12974 27302
rect 13030 27246 13040 27302
rect 12964 27190 13040 27246
rect 12964 27134 12974 27190
rect 13030 27134 13040 27190
rect 12964 27078 13040 27134
rect 12964 27022 12974 27078
rect 13030 27022 13040 27078
rect 12964 26966 13040 27022
rect 12964 26910 12974 26966
rect 13030 26910 13040 26966
rect 12964 26854 13040 26910
rect 12964 26798 12974 26854
rect 13030 26798 13040 26854
rect 12964 26742 13040 26798
rect 12964 26686 12974 26742
rect 13030 26686 13040 26742
rect 12964 26630 13040 26686
rect 12964 26574 12974 26630
rect 13030 26574 13040 26630
rect 12964 26518 13040 26574
rect 12964 26462 12974 26518
rect 13030 26462 13040 26518
rect 12964 26452 13040 26462
rect 23371 27302 23447 27312
rect 23371 27246 23381 27302
rect 23437 27246 23447 27302
rect 23371 27190 23447 27246
rect 23371 27134 23381 27190
rect 23437 27134 23447 27190
rect 23371 27078 23447 27134
rect 23371 27022 23381 27078
rect 23437 27022 23447 27078
rect 23371 26966 23447 27022
rect 23371 26910 23381 26966
rect 23437 26910 23447 26966
rect 23371 26854 23447 26910
rect 23371 26798 23381 26854
rect 23437 26798 23447 26854
rect 23371 26742 23447 26798
rect 23371 26686 23381 26742
rect 23437 26686 23447 26742
rect 23371 26630 23447 26686
rect 23371 26574 23381 26630
rect 23437 26574 23447 26630
rect 23371 26518 23447 26574
rect 23371 26462 23381 26518
rect 23437 26462 23447 26518
rect 23371 26452 23447 26462
rect 23764 27302 23840 27312
rect 23764 27246 23774 27302
rect 23830 27246 23840 27302
rect 23764 27190 23840 27246
rect 23764 27134 23774 27190
rect 23830 27134 23840 27190
rect 23764 27078 23840 27134
rect 23764 27022 23774 27078
rect 23830 27022 23840 27078
rect 23764 26966 23840 27022
rect 23764 26910 23774 26966
rect 23830 26910 23840 26966
rect 23764 26854 23840 26910
rect 23764 26798 23774 26854
rect 23830 26798 23840 26854
rect 23764 26742 23840 26798
rect 23764 26686 23774 26742
rect 23830 26686 23840 26742
rect 23764 26630 23840 26686
rect 23764 26574 23774 26630
rect 23830 26574 23840 26630
rect 23764 26518 23840 26574
rect 23764 26462 23774 26518
rect 23830 26462 23840 26518
rect 23764 26452 23840 26462
rect 61487 27286 61587 27346
rect 61487 27230 61509 27286
rect 61565 27230 61587 27286
rect 61487 27170 61587 27230
rect 61487 27114 61509 27170
rect 61565 27114 61587 27170
rect 61487 27054 61587 27114
rect 61487 26998 61509 27054
rect 61565 26998 61587 27054
rect 61487 26938 61587 26998
rect 61487 26882 61509 26938
rect 61565 26882 61587 26938
rect 61487 26822 61587 26882
rect 61487 26766 61509 26822
rect 61565 26766 61587 26822
rect 61487 26706 61587 26766
rect 61487 26650 61509 26706
rect 61565 26650 61587 26706
rect 61487 26590 61587 26650
rect 61487 26534 61509 26590
rect 61565 26534 61587 26590
rect 61487 26265 61587 26534
rect 72147 27302 72223 27312
rect 72147 27246 72157 27302
rect 72213 27246 72223 27302
rect 72147 27190 72223 27246
rect 72147 27134 72157 27190
rect 72213 27134 72223 27190
rect 72147 27078 72223 27134
rect 72147 27022 72157 27078
rect 72213 27022 72223 27078
rect 72147 26966 72223 27022
rect 72147 26910 72157 26966
rect 72213 26910 72223 26966
rect 72147 26854 72223 26910
rect 72147 26798 72157 26854
rect 72213 26798 72223 26854
rect 72147 26742 72223 26798
rect 72147 26686 72157 26742
rect 72213 26686 72223 26742
rect 72147 26630 72223 26686
rect 72147 26574 72157 26630
rect 72213 26574 72223 26630
rect 72147 26518 72223 26574
rect 72147 26462 72157 26518
rect 72213 26462 72223 26518
rect 72147 26452 72223 26462
rect 72540 27302 72616 27312
rect 72540 27246 72550 27302
rect 72606 27246 72616 27302
rect 72540 27190 72616 27246
rect 72540 27134 72550 27190
rect 72606 27134 72616 27190
rect 72540 27078 72616 27134
rect 72540 27022 72550 27078
rect 72606 27022 72616 27078
rect 72540 26966 72616 27022
rect 72540 26910 72550 26966
rect 72606 26910 72616 26966
rect 72540 26854 72616 26910
rect 72540 26798 72550 26854
rect 72606 26798 72616 26854
rect 72540 26742 72616 26798
rect 72540 26686 72550 26742
rect 72606 26686 72616 26742
rect 72540 26630 72616 26686
rect 72540 26574 72550 26630
rect 72606 26574 72616 26630
rect 72540 26518 72616 26574
rect 72540 26462 72550 26518
rect 72606 26462 72616 26518
rect 72540 26452 72616 26462
rect 82947 27302 83023 27312
rect 82947 27246 82957 27302
rect 83013 27246 83023 27302
rect 82947 27190 83023 27246
rect 82947 27134 82957 27190
rect 83013 27134 83023 27190
rect 82947 27078 83023 27134
rect 82947 27022 82957 27078
rect 83013 27022 83023 27078
rect 82947 26966 83023 27022
rect 82947 26910 82957 26966
rect 83013 26910 83023 26966
rect 82947 26854 83023 26910
rect 82947 26798 82957 26854
rect 83013 26798 83023 26854
rect 82947 26742 83023 26798
rect 82947 26686 82957 26742
rect 83013 26686 83023 26742
rect 82947 26630 83023 26686
rect 82947 26574 82957 26630
rect 83013 26574 83023 26630
rect 82947 26518 83023 26574
rect 82947 26462 82957 26518
rect 83013 26462 83023 26518
rect 82947 26452 83023 26462
rect 83340 27302 83416 27312
rect 83340 27246 83350 27302
rect 83406 27246 83416 27302
rect 83340 27190 83416 27246
rect 83340 27134 83350 27190
rect 83406 27134 83416 27190
rect 83340 27078 83416 27134
rect 83340 27022 83350 27078
rect 83406 27022 83416 27078
rect 83340 26966 83416 27022
rect 83340 26910 83350 26966
rect 83406 26910 83416 26966
rect 83340 26854 83416 26910
rect 83340 26798 83350 26854
rect 83406 26798 83416 26854
rect 83340 26742 83416 26798
rect 83340 26686 83350 26742
rect 83406 26686 83416 26742
rect 83340 26630 83416 26686
rect 83340 26574 83350 26630
rect 83406 26574 83416 26630
rect 83340 26518 83416 26574
rect 83340 26462 83350 26518
rect 83406 26462 83416 26518
rect 83340 26452 83416 26462
<< via2 >>
rect 1934 28274 1990 28330
rect 1934 28158 1990 28214
rect 1934 28042 1990 28098
rect 1934 27926 1990 27982
rect 1934 27810 1990 27866
rect 12581 28321 12637 28377
rect 12581 28209 12637 28265
rect 12581 28097 12637 28153
rect 12581 27985 12637 28041
rect 12581 27873 12637 27929
rect 12581 27761 12637 27817
rect 12974 28321 13030 28377
rect 12974 28209 13030 28265
rect 12974 28097 13030 28153
rect 12974 27985 13030 28041
rect 12974 27873 13030 27929
rect 12974 27761 13030 27817
rect 23381 28321 23437 28377
rect 23381 28209 23437 28265
rect 23381 28097 23437 28153
rect 23381 27985 23437 28041
rect 23381 27873 23437 27929
rect 23381 27761 23437 27817
rect 23774 28321 23830 28377
rect 23774 28209 23830 28265
rect 23774 28097 23830 28153
rect 23774 27985 23830 28041
rect 23774 27873 23830 27929
rect 23774 27761 23830 27817
rect 61509 28274 61565 28330
rect 61509 28158 61565 28214
rect 61509 28042 61565 28098
rect 61509 27926 61565 27982
rect 61509 27810 61565 27866
rect 1934 27694 1990 27750
rect 1934 27578 1990 27634
rect 1934 27462 1990 27518
rect 1934 27346 1990 27402
rect 72157 28321 72213 28377
rect 72157 28209 72213 28265
rect 72157 28097 72213 28153
rect 72157 27985 72213 28041
rect 72157 27873 72213 27929
rect 72157 27761 72213 27817
rect 72550 28321 72606 28377
rect 72550 28209 72606 28265
rect 72550 28097 72606 28153
rect 72550 27985 72606 28041
rect 72550 27873 72606 27929
rect 72550 27761 72606 27817
rect 82957 28321 83013 28377
rect 82957 28209 83013 28265
rect 82957 28097 83013 28153
rect 82957 27985 83013 28041
rect 82957 27873 83013 27929
rect 82957 27761 83013 27817
rect 83350 28321 83406 28377
rect 83350 28209 83406 28265
rect 83350 28097 83406 28153
rect 83350 27985 83406 28041
rect 83350 27873 83406 27929
rect 83350 27761 83406 27817
rect 61509 27694 61565 27750
rect 61509 27578 61565 27634
rect 61509 27462 61565 27518
rect 61509 27346 61565 27402
rect 1934 27230 1990 27286
rect 1934 27114 1990 27170
rect 1934 26998 1990 27054
rect 1934 26882 1990 26938
rect 1934 26766 1990 26822
rect 1934 26650 1990 26706
rect 1934 26534 1990 26590
rect 12581 27246 12637 27302
rect 12581 27134 12637 27190
rect 12581 27022 12637 27078
rect 12581 26910 12637 26966
rect 12581 26798 12637 26854
rect 12581 26686 12637 26742
rect 12581 26574 12637 26630
rect 12581 26462 12637 26518
rect 12974 27246 13030 27302
rect 12974 27134 13030 27190
rect 12974 27022 13030 27078
rect 12974 26910 13030 26966
rect 12974 26798 13030 26854
rect 12974 26686 13030 26742
rect 12974 26574 13030 26630
rect 12974 26462 13030 26518
rect 23381 27246 23437 27302
rect 23381 27134 23437 27190
rect 23381 27022 23437 27078
rect 23381 26910 23437 26966
rect 23381 26798 23437 26854
rect 23381 26686 23437 26742
rect 23381 26574 23437 26630
rect 23381 26462 23437 26518
rect 23774 27246 23830 27302
rect 23774 27134 23830 27190
rect 23774 27022 23830 27078
rect 23774 26910 23830 26966
rect 23774 26798 23830 26854
rect 23774 26686 23830 26742
rect 23774 26574 23830 26630
rect 23774 26462 23830 26518
rect 61509 27230 61565 27286
rect 61509 27114 61565 27170
rect 61509 26998 61565 27054
rect 61509 26882 61565 26938
rect 61509 26766 61565 26822
rect 61509 26650 61565 26706
rect 61509 26534 61565 26590
rect 72157 27246 72213 27302
rect 72157 27134 72213 27190
rect 72157 27022 72213 27078
rect 72157 26910 72213 26966
rect 72157 26798 72213 26854
rect 72157 26686 72213 26742
rect 72157 26574 72213 26630
rect 72157 26462 72213 26518
rect 72550 27246 72606 27302
rect 72550 27134 72606 27190
rect 72550 27022 72606 27078
rect 72550 26910 72606 26966
rect 72550 26798 72606 26854
rect 72550 26686 72606 26742
rect 72550 26574 72606 26630
rect 72550 26462 72606 26518
rect 82957 27246 83013 27302
rect 82957 27134 83013 27190
rect 82957 27022 83013 27078
rect 82957 26910 83013 26966
rect 82957 26798 83013 26854
rect 82957 26686 83013 26742
rect 82957 26574 83013 26630
rect 82957 26462 83013 26518
rect 83350 27246 83406 27302
rect 83350 27134 83406 27190
rect 83350 27022 83406 27078
rect 83350 26910 83406 26966
rect 83350 26798 83406 26854
rect 83350 26686 83406 26742
rect 83350 26574 83406 26630
rect 83350 26462 83406 26518
<< metal3 >>
rect 12571 28377 12647 28387
rect 1924 28330 2000 28340
rect 1924 28274 1934 28330
rect 1990 28274 2000 28330
rect 1924 28214 2000 28274
rect 1924 28158 1934 28214
rect 1990 28158 2000 28214
rect 1924 28098 2000 28158
rect 1924 28042 1934 28098
rect 1990 28042 2000 28098
rect 1924 27982 2000 28042
rect 1924 27926 1934 27982
rect 1990 27926 2000 27982
rect 1924 27866 2000 27926
rect 1924 27810 1934 27866
rect 1990 27810 2000 27866
rect 1924 27750 2000 27810
rect 12571 28321 12581 28377
rect 12637 28321 12647 28377
rect 12571 28265 12647 28321
rect 12571 28209 12581 28265
rect 12637 28209 12647 28265
rect 12571 28153 12647 28209
rect 12571 28097 12581 28153
rect 12637 28097 12647 28153
rect 12571 28041 12647 28097
rect 12571 27985 12581 28041
rect 12637 27985 12647 28041
rect 12571 27929 12647 27985
rect 12571 27873 12581 27929
rect 12637 27873 12647 27929
rect 12571 27817 12647 27873
rect 12571 27761 12581 27817
rect 12637 27761 12647 27817
rect 12571 27751 12647 27761
rect 12964 28377 13040 28387
rect 12964 28321 12974 28377
rect 13030 28321 13040 28377
rect 12964 28265 13040 28321
rect 12964 28209 12974 28265
rect 13030 28209 13040 28265
rect 12964 28153 13040 28209
rect 12964 28097 12974 28153
rect 13030 28097 13040 28153
rect 12964 28041 13040 28097
rect 12964 27985 12974 28041
rect 13030 27985 13040 28041
rect 12964 27929 13040 27985
rect 12964 27873 12974 27929
rect 13030 27873 13040 27929
rect 12964 27817 13040 27873
rect 12964 27761 12974 27817
rect 13030 27761 13040 27817
rect 12964 27751 13040 27761
rect 23371 28377 23447 28387
rect 23371 28321 23381 28377
rect 23437 28321 23447 28377
rect 23371 28265 23447 28321
rect 23371 28209 23381 28265
rect 23437 28209 23447 28265
rect 23371 28153 23447 28209
rect 23371 28097 23381 28153
rect 23437 28097 23447 28153
rect 23371 28041 23447 28097
rect 23371 27985 23381 28041
rect 23437 27985 23447 28041
rect 23371 27929 23447 27985
rect 23371 27873 23381 27929
rect 23437 27873 23447 27929
rect 23371 27817 23447 27873
rect 23371 27761 23381 27817
rect 23437 27761 23447 27817
rect 23371 27751 23447 27761
rect 23764 28377 23840 28387
rect 23764 28321 23774 28377
rect 23830 28321 23840 28377
rect 72147 28377 72223 28387
rect 23764 28265 23840 28321
rect 23764 28209 23774 28265
rect 23830 28209 23840 28265
rect 23764 28153 23840 28209
rect 23764 28097 23774 28153
rect 23830 28097 23840 28153
rect 23764 28041 23840 28097
rect 23764 27985 23774 28041
rect 23830 27985 23840 28041
rect 23764 27929 23840 27985
rect 23764 27873 23774 27929
rect 23830 27873 23840 27929
rect 23764 27817 23840 27873
rect 23764 27761 23774 27817
rect 23830 27761 23840 27817
rect 23764 27751 23840 27761
rect 61499 28330 61575 28340
rect 61499 28274 61509 28330
rect 61565 28274 61575 28330
rect 61499 28214 61575 28274
rect 61499 28158 61509 28214
rect 61565 28158 61575 28214
rect 61499 28098 61575 28158
rect 61499 28042 61509 28098
rect 61565 28042 61575 28098
rect 61499 27982 61575 28042
rect 61499 27926 61509 27982
rect 61565 27926 61575 27982
rect 61499 27866 61575 27926
rect 61499 27810 61509 27866
rect 61565 27810 61575 27866
rect 1924 27694 1934 27750
rect 1990 27694 2000 27750
rect 1924 27634 2000 27694
rect 1924 27578 1934 27634
rect 1990 27578 2000 27634
rect 1924 27518 2000 27578
rect 1924 27462 1934 27518
rect 1990 27462 2000 27518
rect 1924 27402 2000 27462
rect 1924 27346 1934 27402
rect 1990 27346 2000 27402
rect 1924 27286 2000 27346
rect 61499 27750 61575 27810
rect 72147 28321 72157 28377
rect 72213 28321 72223 28377
rect 72147 28265 72223 28321
rect 72147 28209 72157 28265
rect 72213 28209 72223 28265
rect 72147 28153 72223 28209
rect 72147 28097 72157 28153
rect 72213 28097 72223 28153
rect 72147 28041 72223 28097
rect 72147 27985 72157 28041
rect 72213 27985 72223 28041
rect 72147 27929 72223 27985
rect 72147 27873 72157 27929
rect 72213 27873 72223 27929
rect 72147 27817 72223 27873
rect 72147 27761 72157 27817
rect 72213 27761 72223 27817
rect 72147 27751 72223 27761
rect 72540 28377 72616 28387
rect 72540 28321 72550 28377
rect 72606 28321 72616 28377
rect 72540 28265 72616 28321
rect 72540 28209 72550 28265
rect 72606 28209 72616 28265
rect 72540 28153 72616 28209
rect 72540 28097 72550 28153
rect 72606 28097 72616 28153
rect 72540 28041 72616 28097
rect 72540 27985 72550 28041
rect 72606 27985 72616 28041
rect 72540 27929 72616 27985
rect 72540 27873 72550 27929
rect 72606 27873 72616 27929
rect 72540 27817 72616 27873
rect 72540 27761 72550 27817
rect 72606 27761 72616 27817
rect 72540 27751 72616 27761
rect 82947 28377 83023 28387
rect 82947 28321 82957 28377
rect 83013 28321 83023 28377
rect 82947 28265 83023 28321
rect 82947 28209 82957 28265
rect 83013 28209 83023 28265
rect 82947 28153 83023 28209
rect 82947 28097 82957 28153
rect 83013 28097 83023 28153
rect 82947 28041 83023 28097
rect 82947 27985 82957 28041
rect 83013 27985 83023 28041
rect 82947 27929 83023 27985
rect 82947 27873 82957 27929
rect 83013 27873 83023 27929
rect 82947 27817 83023 27873
rect 82947 27761 82957 27817
rect 83013 27761 83023 27817
rect 82947 27751 83023 27761
rect 83340 28377 83416 28387
rect 83340 28321 83350 28377
rect 83406 28321 83416 28377
rect 83340 28265 83416 28321
rect 83340 28209 83350 28265
rect 83406 28209 83416 28265
rect 83340 28153 83416 28209
rect 83340 28097 83350 28153
rect 83406 28097 83416 28153
rect 83340 28041 83416 28097
rect 83340 27985 83350 28041
rect 83406 27985 83416 28041
rect 83340 27929 83416 27985
rect 83340 27873 83350 27929
rect 83406 27873 83416 27929
rect 83340 27817 83416 27873
rect 83340 27761 83350 27817
rect 83406 27761 83416 27817
rect 83340 27751 83416 27761
rect 61499 27694 61509 27750
rect 61565 27694 61575 27750
rect 61499 27634 61575 27694
rect 61499 27578 61509 27634
rect 61565 27578 61575 27634
rect 61499 27518 61575 27578
rect 61499 27462 61509 27518
rect 61565 27462 61575 27518
rect 61499 27402 61575 27462
rect 61499 27346 61509 27402
rect 61565 27346 61575 27402
rect 1924 27230 1934 27286
rect 1990 27230 2000 27286
rect 1924 27170 2000 27230
rect 1924 27114 1934 27170
rect 1990 27114 2000 27170
rect 1924 27054 2000 27114
rect 1924 26998 1934 27054
rect 1990 26998 2000 27054
rect 1924 26938 2000 26998
rect 1924 26882 1934 26938
rect 1990 26882 2000 26938
rect 1924 26822 2000 26882
rect 1924 26766 1934 26822
rect 1990 26766 2000 26822
rect 1924 26706 2000 26766
rect 1924 26650 1934 26706
rect 1990 26650 2000 26706
rect 1924 26590 2000 26650
rect 1924 26534 1934 26590
rect 1990 26534 2000 26590
rect 1924 26524 2000 26534
rect 12571 27302 12647 27312
rect 12571 27246 12581 27302
rect 12637 27246 12647 27302
rect 12571 27190 12647 27246
rect 12571 27134 12581 27190
rect 12637 27134 12647 27190
rect 12571 27078 12647 27134
rect 12571 27022 12581 27078
rect 12637 27022 12647 27078
rect 12571 26966 12647 27022
rect 12571 26910 12581 26966
rect 12637 26910 12647 26966
rect 12571 26854 12647 26910
rect 12571 26798 12581 26854
rect 12637 26798 12647 26854
rect 12571 26742 12647 26798
rect 12571 26686 12581 26742
rect 12637 26686 12647 26742
rect 12571 26630 12647 26686
rect 12571 26574 12581 26630
rect 12637 26574 12647 26630
rect 12571 26518 12647 26574
rect 12571 26462 12581 26518
rect 12637 26462 12647 26518
rect 12571 26452 12647 26462
rect 12964 27302 13040 27312
rect 12964 27246 12974 27302
rect 13030 27246 13040 27302
rect 12964 27190 13040 27246
rect 12964 27134 12974 27190
rect 13030 27134 13040 27190
rect 12964 27078 13040 27134
rect 12964 27022 12974 27078
rect 13030 27022 13040 27078
rect 12964 26966 13040 27022
rect 12964 26910 12974 26966
rect 13030 26910 13040 26966
rect 12964 26854 13040 26910
rect 12964 26798 12974 26854
rect 13030 26798 13040 26854
rect 12964 26742 13040 26798
rect 12964 26686 12974 26742
rect 13030 26686 13040 26742
rect 12964 26630 13040 26686
rect 12964 26574 12974 26630
rect 13030 26574 13040 26630
rect 12964 26518 13040 26574
rect 12964 26462 12974 26518
rect 13030 26462 13040 26518
rect 12964 26452 13040 26462
rect 23371 27302 23447 27312
rect 23371 27246 23381 27302
rect 23437 27246 23447 27302
rect 23371 27190 23447 27246
rect 23371 27134 23381 27190
rect 23437 27134 23447 27190
rect 23371 27078 23447 27134
rect 23371 27022 23381 27078
rect 23437 27022 23447 27078
rect 23371 26966 23447 27022
rect 23371 26910 23381 26966
rect 23437 26910 23447 26966
rect 23371 26854 23447 26910
rect 23371 26798 23381 26854
rect 23437 26798 23447 26854
rect 23371 26742 23447 26798
rect 23371 26686 23381 26742
rect 23437 26686 23447 26742
rect 23371 26630 23447 26686
rect 23371 26574 23381 26630
rect 23437 26574 23447 26630
rect 23371 26518 23447 26574
rect 23371 26462 23381 26518
rect 23437 26462 23447 26518
rect 23371 26452 23447 26462
rect 23764 27302 23840 27312
rect 23764 27246 23774 27302
rect 23830 27246 23840 27302
rect 23764 27190 23840 27246
rect 23764 27134 23774 27190
rect 23830 27134 23840 27190
rect 23764 27078 23840 27134
rect 23764 27022 23774 27078
rect 23830 27022 23840 27078
rect 23764 26966 23840 27022
rect 23764 26910 23774 26966
rect 23830 26910 23840 26966
rect 23764 26854 23840 26910
rect 23764 26798 23774 26854
rect 23830 26798 23840 26854
rect 23764 26742 23840 26798
rect 23764 26686 23774 26742
rect 23830 26686 23840 26742
rect 23764 26630 23840 26686
rect 23764 26574 23774 26630
rect 23830 26574 23840 26630
rect 23764 26518 23840 26574
rect 61499 27286 61575 27346
rect 61499 27230 61509 27286
rect 61565 27230 61575 27286
rect 61499 27170 61575 27230
rect 61499 27114 61509 27170
rect 61565 27114 61575 27170
rect 61499 27054 61575 27114
rect 61499 26998 61509 27054
rect 61565 26998 61575 27054
rect 61499 26938 61575 26998
rect 61499 26882 61509 26938
rect 61565 26882 61575 26938
rect 61499 26822 61575 26882
rect 61499 26766 61509 26822
rect 61565 26766 61575 26822
rect 61499 26706 61575 26766
rect 61499 26650 61509 26706
rect 61565 26650 61575 26706
rect 61499 26590 61575 26650
rect 61499 26534 61509 26590
rect 61565 26534 61575 26590
rect 61499 26524 61575 26534
rect 72147 27302 72223 27312
rect 72147 27246 72157 27302
rect 72213 27246 72223 27302
rect 72147 27190 72223 27246
rect 72147 27134 72157 27190
rect 72213 27134 72223 27190
rect 72147 27078 72223 27134
rect 72147 27022 72157 27078
rect 72213 27022 72223 27078
rect 72147 26966 72223 27022
rect 72147 26910 72157 26966
rect 72213 26910 72223 26966
rect 72147 26854 72223 26910
rect 72147 26798 72157 26854
rect 72213 26798 72223 26854
rect 72147 26742 72223 26798
rect 72147 26686 72157 26742
rect 72213 26686 72223 26742
rect 72147 26630 72223 26686
rect 72147 26574 72157 26630
rect 72213 26574 72223 26630
rect 23764 26462 23774 26518
rect 23830 26462 23840 26518
rect 23764 26452 23840 26462
rect 72147 26518 72223 26574
rect 72147 26462 72157 26518
rect 72213 26462 72223 26518
rect 72147 26452 72223 26462
rect 72540 27302 72616 27312
rect 72540 27246 72550 27302
rect 72606 27246 72616 27302
rect 72540 27190 72616 27246
rect 72540 27134 72550 27190
rect 72606 27134 72616 27190
rect 72540 27078 72616 27134
rect 72540 27022 72550 27078
rect 72606 27022 72616 27078
rect 72540 26966 72616 27022
rect 72540 26910 72550 26966
rect 72606 26910 72616 26966
rect 72540 26854 72616 26910
rect 72540 26798 72550 26854
rect 72606 26798 72616 26854
rect 72540 26742 72616 26798
rect 72540 26686 72550 26742
rect 72606 26686 72616 26742
rect 72540 26630 72616 26686
rect 72540 26574 72550 26630
rect 72606 26574 72616 26630
rect 72540 26518 72616 26574
rect 72540 26462 72550 26518
rect 72606 26462 72616 26518
rect 72540 26452 72616 26462
rect 82947 27302 83023 27312
rect 82947 27246 82957 27302
rect 83013 27246 83023 27302
rect 82947 27190 83023 27246
rect 82947 27134 82957 27190
rect 83013 27134 83023 27190
rect 82947 27078 83023 27134
rect 82947 27022 82957 27078
rect 83013 27022 83023 27078
rect 82947 26966 83023 27022
rect 82947 26910 82957 26966
rect 83013 26910 83023 26966
rect 82947 26854 83023 26910
rect 82947 26798 82957 26854
rect 83013 26798 83023 26854
rect 82947 26742 83023 26798
rect 82947 26686 82957 26742
rect 83013 26686 83023 26742
rect 82947 26630 83023 26686
rect 82947 26574 82957 26630
rect 83013 26574 83023 26630
rect 82947 26518 83023 26574
rect 82947 26462 82957 26518
rect 83013 26462 83023 26518
rect 82947 26452 83023 26462
rect 83340 27302 83416 27312
rect 83340 27246 83350 27302
rect 83406 27246 83416 27302
rect 83340 27190 83416 27246
rect 83340 27134 83350 27190
rect 83406 27134 83416 27190
rect 83340 27078 83416 27134
rect 83340 27022 83350 27078
rect 83406 27022 83416 27078
rect 83340 26966 83416 27022
rect 83340 26910 83350 26966
rect 83406 26910 83416 26966
rect 83340 26854 83416 26910
rect 83340 26798 83350 26854
rect 83406 26798 83416 26854
rect 83340 26742 83416 26798
rect 83340 26686 83350 26742
rect 83406 26686 83416 26742
rect 83340 26630 83416 26686
rect 83340 26574 83350 26630
rect 83406 26574 83416 26630
rect 83340 26518 83416 26574
rect 83340 26462 83350 26518
rect 83406 26462 83416 26518
rect 83340 26452 83416 26462
rect 46982 15015 47947 16784
rect 27546 14936 47947 15015
rect 27546 14503 47683 14936
rect 41493 14491 47683 14503
rect 41493 13729 45977 14491
rect 41151 6592 51232 7392
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_0
timestamp 1762296095
transform 1 0 18458 0 1 34450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_1
timestamp 1762296095
transform 1 0 67234 0 1 34450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_2
timestamp 1762296095
transform 1 0 78034 0 1 34450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_3
timestamp 1762296095
transform 1 0 7658 0 1 34450
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_0
timestamp 1762296095
transform -1 0 72698 0 1 34224
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_1
timestamp 1762296095
transform -1 0 83138 0 1 34224
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_2
timestamp 1762296095
transform -1 0 61898 0 1 34224
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_3
timestamp 1762296095
transform 1 0 13122 0 1 34224
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_4
timestamp 1762296095
transform 1 0 2322 0 1 34224
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_5
timestamp 1762296095
transform 1 0 23562 0 1 34224
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_0
timestamp 1762296095
transform 1 0 12609 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_1
timestamp 1762296095
transform 1 0 23802 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_2
timestamp 1762296095
transform 1 0 23409 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_3
timestamp 1762296095
transform 1 0 72578 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_4
timestamp 1762296095
transform 1 0 72185 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_5
timestamp 1762296095
transform 1 0 83378 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_6
timestamp 1762296095
transform 1 0 82985 0 1 26882
box 0 0 1 1
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_7
timestamp 1762296095
transform 1 0 13002 0 1 26882
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_0
timestamp 1762296095
transform 1 0 12609 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_1
timestamp 1762296095
transform 1 0 23802 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_2
timestamp 1762296095
transform 1 0 23409 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_3
timestamp 1762296095
transform 1 0 72578 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_4
timestamp 1762296095
transform 1 0 72185 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_5
timestamp 1762296095
transform 1 0 83378 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_6
timestamp 1762296095
transform 1 0 82985 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_7
timestamp 1762296095
transform 1 0 13002 0 1 28069
box 0 0 1 1
use M3_M243105908781102_256x8m81  M3_M243105908781102_256x8m81_0
timestamp 1762296095
transform 1 0 61537 0 1 27432
box 0 0 1 1
use M3_M243105908781102_256x8m81  M3_M243105908781102_256x8m81_1
timestamp 1762296095
transform 1 0 1962 0 1 27432
box 0 0 1 1
<< properties >>
string GDS_END 2289122
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2286116
string path 205.755 34.960 256.160 34.960 
<< end >>
