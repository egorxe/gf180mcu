VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_fd_io__bi_t
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_fd_io__bi_t ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 264.460 69.780 350.000 ;
    END
  END A
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 328.545 3.740 350.000 ;
    END
  END CS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 166.000 75.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 334.000 1.000 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 294.000 1.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 262.000 1.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 270.000 1.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 278.000 1.000 285.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 206.000 1.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 214.000 1.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 134.000 1.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 150.000 1.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 166.000 1.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 182.000 1.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 1.000 125.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 342.000 75.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 342.000 1.000 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 326.000 1.000 333.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 302.000 1.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 286.000 1.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 230.000 1.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 198.000 1.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 126.000 1.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 70.000 1.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 86.000 1.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 1.000 117.000 ;
    END
  END DVSS
  PIN IE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.385 334.920 11.765 350.000 ;
    END
  END IE
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.799999 ;
    ANTENNADIFFAREA 7.776000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 266.340 70.510 350.000 ;
    END
  END OE
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 258.720001 ;
    PORT
      LAYER Metal5 ;
        RECT 25.000 20.000 50.000 45.000 ;
    END
  END PAD
  PIN PD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.500000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.330 330.100 10.710 350.000 ;
    END
  END PD
  PIN PDRV0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 2.592000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.110 264.665 7.490 350.000 ;
    END
  END PDRV0
  PIN PDRV1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.200000 ;
    ANTENNADIFFAREA 2.592000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.820 264.990 8.200 350.000 ;
    END
  END PDRV1
  PIN PU
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.350000 ;
    ANTENNADIFFAREA 2.980000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.965 330.420 6.345 350.000 ;
    END
  END PU
  PIN SL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.150000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.670 265.140 69.050 350.000 ;
    END
  END SL
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 310.000 75.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 310.000 1.000 317.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 1.000 261.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 246.000 75.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 74.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 7.800000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.860 319.900 71.240 350.000 ;
    END
  END Y
  OBS
      LAYER Nwell ;
        RECT 1.820 68.895 73.180 346.535 ;
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 328.245 3.060 348.375 ;
        RECT 4.040 330.120 5.665 348.375 ;
        RECT 6.645 330.120 6.810 348.375 ;
        RECT 4.040 328.245 6.810 330.120 ;
        RECT 0.000 264.365 6.810 328.245 ;
        RECT 8.500 329.800 10.030 348.375 ;
        RECT 11.010 334.620 11.085 348.375 ;
        RECT 12.065 334.620 68.370 348.375 ;
        RECT 11.010 329.800 68.370 334.620 ;
        RECT 8.500 264.840 68.370 329.800 ;
        RECT 71.540 319.600 75.000 348.375 ;
        RECT 70.810 266.040 75.000 319.600 ;
        RECT 8.500 264.690 69.100 264.840 ;
        RECT 7.790 264.365 69.100 264.690 ;
        RECT 0.000 264.160 69.100 264.365 ;
        RECT 70.080 264.160 75.000 266.040 ;
        RECT 0.000 0.000 75.000 264.160 ;
      LAYER Metal3 ;
        RECT 1.300 341.700 73.700 348.390 ;
        RECT 0.665 341.300 74.000 341.700 ;
        RECT 1.300 333.700 73.700 341.300 ;
        RECT 0.665 333.300 74.000 333.700 ;
        RECT 1.300 325.700 73.700 333.300 ;
        RECT 0.665 325.300 74.000 325.700 ;
        RECT 1.300 317.700 73.700 325.300 ;
        RECT 0.665 317.300 74.000 317.700 ;
        RECT 1.300 309.700 73.700 317.300 ;
        RECT 0.665 309.300 74.000 309.700 ;
        RECT 1.300 301.700 73.700 309.300 ;
        RECT 0.665 301.300 74.000 301.700 ;
        RECT 1.300 293.700 73.700 301.300 ;
        RECT 0.665 293.300 74.000 293.700 ;
        RECT 1.300 285.700 73.700 293.300 ;
        RECT 0.665 285.300 74.000 285.700 ;
        RECT 1.300 277.700 73.700 285.300 ;
        RECT 0.665 277.300 74.000 277.700 ;
        RECT 1.300 269.700 73.700 277.300 ;
        RECT 0.665 269.300 74.000 269.700 ;
        RECT 1.300 261.700 73.700 269.300 ;
        RECT 0.665 261.300 74.000 261.700 ;
        RECT 1.300 253.700 73.700 261.300 ;
        RECT 0.665 253.300 74.000 253.700 ;
        RECT 1.300 245.700 73.700 253.300 ;
        RECT 0.665 245.300 74.000 245.700 ;
        RECT 1.300 229.700 73.700 245.300 ;
        RECT 0.665 229.300 74.000 229.700 ;
        RECT 1.300 213.700 73.700 229.300 ;
        RECT 0.665 213.300 74.000 213.700 ;
        RECT 1.300 205.700 73.700 213.300 ;
        RECT 0.665 205.300 74.000 205.700 ;
        RECT 1.300 197.700 73.700 205.300 ;
        RECT 0.665 197.300 74.000 197.700 ;
        RECT 1.300 181.700 73.700 197.300 ;
        RECT 0.665 181.300 74.000 181.700 ;
        RECT 1.300 165.700 73.700 181.300 ;
        RECT 0.665 165.300 74.000 165.700 ;
        RECT 1.300 149.700 73.700 165.300 ;
        RECT 0.665 149.300 74.000 149.700 ;
        RECT 1.300 133.700 73.700 149.300 ;
        RECT 0.665 133.300 74.000 133.700 ;
        RECT 1.300 125.700 73.700 133.300 ;
        RECT 0.665 125.300 74.000 125.700 ;
        RECT 1.300 117.700 73.700 125.300 ;
        RECT 0.665 117.300 74.000 117.700 ;
        RECT 1.300 101.700 73.700 117.300 ;
        RECT 0.665 101.300 74.000 101.700 ;
        RECT 1.300 85.700 73.700 101.300 ;
        RECT 0.665 85.300 74.000 85.700 ;
        RECT 1.300 69.700 73.700 85.300 ;
        RECT 0.665 0.000 74.000 69.700 ;
      LAYER Metal4 ;
        RECT 1.300 341.700 73.700 348.390 ;
        RECT 1.000 341.300 74.000 341.700 ;
        RECT 1.300 333.700 73.700 341.300 ;
        RECT 1.000 333.300 74.000 333.700 ;
        RECT 1.300 325.700 73.700 333.300 ;
        RECT 1.000 325.300 74.000 325.700 ;
        RECT 1.300 317.700 73.700 325.300 ;
        RECT 1.000 317.300 74.000 317.700 ;
        RECT 1.300 309.700 73.700 317.300 ;
        RECT 1.000 309.300 74.000 309.700 ;
        RECT 1.300 301.700 73.700 309.300 ;
        RECT 1.000 301.300 74.000 301.700 ;
        RECT 1.300 293.700 73.700 301.300 ;
        RECT 1.000 293.300 74.000 293.700 ;
        RECT 1.300 285.700 73.700 293.300 ;
        RECT 1.000 285.300 74.000 285.700 ;
        RECT 1.300 277.700 73.700 285.300 ;
        RECT 1.000 277.300 74.000 277.700 ;
        RECT 1.300 269.700 73.700 277.300 ;
        RECT 1.000 269.300 74.000 269.700 ;
        RECT 1.300 261.700 73.700 269.300 ;
        RECT 1.000 261.300 74.000 261.700 ;
        RECT 1.300 253.700 73.700 261.300 ;
        RECT 1.000 253.300 74.000 253.700 ;
        RECT 1.300 245.700 73.700 253.300 ;
        RECT 1.000 245.300 74.000 245.700 ;
        RECT 1.300 229.700 73.700 245.300 ;
        RECT 1.000 229.300 74.000 229.700 ;
        RECT 1.300 213.700 73.700 229.300 ;
        RECT 1.000 213.300 74.000 213.700 ;
        RECT 1.300 205.700 73.700 213.300 ;
        RECT 1.000 205.300 74.000 205.700 ;
        RECT 1.300 197.700 73.700 205.300 ;
        RECT 1.000 197.300 74.000 197.700 ;
        RECT 1.300 181.700 73.700 197.300 ;
        RECT 1.000 181.300 74.000 181.700 ;
        RECT 1.300 165.700 73.700 181.300 ;
        RECT 1.000 165.300 74.000 165.700 ;
        RECT 1.300 149.700 73.700 165.300 ;
        RECT 1.000 149.300 74.000 149.700 ;
        RECT 1.300 133.700 73.700 149.300 ;
        RECT 1.000 133.300 74.000 133.700 ;
        RECT 1.300 125.700 73.700 133.300 ;
        RECT 1.000 125.300 74.000 125.700 ;
        RECT 1.300 117.700 73.700 125.300 ;
        RECT 1.000 117.300 74.000 117.700 ;
        RECT 1.300 101.700 73.700 117.300 ;
        RECT 1.000 101.300 74.000 101.700 ;
        RECT 1.300 85.700 73.700 101.300 ;
        RECT 1.000 85.300 74.000 85.700 ;
        RECT 1.300 69.700 73.700 85.300 ;
        RECT 1.000 0.000 74.000 69.700 ;
      LAYER Metal5 ;
        RECT 1.600 69.400 73.400 348.390 ;
        RECT 1.000 45.600 74.000 69.400 ;
        RECT 1.000 19.400 24.400 45.600 ;
        RECT 50.600 19.400 74.000 45.600 ;
        RECT 1.000 0.000 74.000 19.400 ;
  END
END gf180mcu_fd_io__bi_t
END LIBRARY

