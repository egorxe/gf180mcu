magic
tech gf180mcuD
magscale 1 10
timestamp 1759194789
<< metal3 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< metal4 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
<< metal5 >>
rect 14000 70800 17000 71000
rect 17200 70800 20200 71000
rect 20400 70800 23400 71000
rect 23600 70800 25000 71000
rect 25200 70800 26600 71000
rect 26800 70800 29800 71000
rect 30000 70800 33000 71000
rect 33200 70800 36200 71000
rect 36400 70800 39400 71000
rect 39600 70800 41000 71000
rect 41200 70800 42600 71000
rect 42800 70800 45800 71000
rect 46000 70800 49000 71000
rect 49200 70800 50600 71000
rect 50800 70800 52200 71000
rect 52400 70800 53800 71000
rect 54000 70800 55400 71000
rect 55600 70800 57000 71000
rect 57200 70800 58600 71000
rect 58800 70800 60200 71000
rect 60400 70800 61800 71000
rect 62000 70800 63400 71000
rect 63600 70800 65000 71000
rect 65200 70800 66600 71000
rect 66800 70800 68200 71000
rect 68400 70800 69678 71000
rect 70800 68400 71000 69678
rect 70800 66800 71000 68200
rect 70800 65200 71000 66600
rect 70800 63600 71000 65000
rect 70800 62000 71000 63400
rect 70800 60400 71000 61800
rect 70800 58800 71000 60200
rect 70800 57200 71000 58600
rect 70800 55600 71000 57000
rect 70800 54000 71000 55400
rect 70800 52400 71000 53800
rect 70800 50800 71000 52200
rect 70800 49200 71000 50600
rect 70800 46000 71000 49000
rect 70800 41200 71000 42600
rect 70800 39600 71000 41000
rect 70800 36400 71000 39400
rect 70800 33200 71000 36200
rect 70800 30000 71000 33000
rect 70800 26800 71000 29800
rect 70800 25200 71000 26600
rect 70800 23600 71000 25000
rect 70800 20400 71000 23400
rect 70800 17200 71000 20200
rect 70800 14000 71000 17000
use GF_NI_COR_BASE  GF_NI_COR_BASE_0
timestamp 1759194789
transform 1 0 12 0 1 0
box 12200 13361 70889 70890
use POWER_RAIL_COR  POWER_RAIL_COR_0
timestamp 1759194789
transform 1 0 0 0 1 0
box 13097 13097 71000 71000
<< labels >>
rlabel metal3 s 66800 70800 68200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 63600 70800 65000 71000 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 70800 66800 71000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 58800 70800 60200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 68400 70800 69678 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 58800 71000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 55600 70800 57000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 55600 71000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 54000 70800 55400 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 63600 71000 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 62000 70800 63400 71000 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 68400 71000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 54000 71000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 52400 70800 53800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 52400 71000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 42800 70800 45800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal3 s 41200 70800 42600 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 41200 71000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 36400 70800 39400 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 36400 71000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 33200 70800 36200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 33200 71000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 49200 70800 50600 71000 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 65200 70800 66600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 30000 70800 33000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 62000 71000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 65200 71000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 50800 70800 52200 71000 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 30000 71000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 60400 70800 61800 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 60400 71000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 57200 70800 58600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 26800 70800 29800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 57200 71000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 26800 71000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 46000 70800 49000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 46000 71000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 63600 70800 65000 71000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 62000 70800 63400 71000 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 23600 70800 25000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 39600 70800 41000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 39600 71000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 25200 70800 26600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 25200 71000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 20400 70800 23400 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 20400 71000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 17200 70800 20200 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 17200 71000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 14000 70800 17000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 68400 70800 69678 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 66800 70800 68200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 66800 71000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 68400 71000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 63600 71000 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 65200 70800 66600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 65200 71000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 60400 70800 61800 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 60400 71000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 57200 70800 58600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 49200 70800 50600 71000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 62000 71000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 58800 70800 60200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 58800 71000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 55600 70800 57000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 55600 71000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 54000 70800 55400 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 50800 70800 52200 71000 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 54000 71000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 52400 70800 53800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 57200 71000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 63600 70800 65000 71000 4 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 62000 70800 63400 71000 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 52400 71000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 42800 70800 45800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal4 s 46000 70800 49000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 41200 70800 42600 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 46000 71000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 62000 71000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal5 s 70800 63600 71000 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 39600 70800 41000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 41200 71000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 39600 71000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 49200 70800 50600 71000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 25200 70800 26600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 25200 71000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 20400 70800 23400 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 20400 71000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 17200 70800 20200 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 49200 71000 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 50800 70800 52200 71000 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 36400 70800 39400 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 36400 71000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 33200 70800 36200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 33200 71000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 30000 70800 33000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 50800 71000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 30000 71000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 26800 70800 29800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 17200 71000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 70800 49200 71000 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 70800 50800 71000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 70800 26800 71000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 23600 70800 25000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 66800 70800 68200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 14000 70800 17000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 66800 71000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 68400 70800 69678 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 70800 50800 71000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 70800 49200 71000 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 70800 68400 71000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal5 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal5 s 58800 70800 60200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 65200 70800 66600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 65200 71000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 60400 70800 61800 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 60400 71000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 57200 70800 58600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 57200 71000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 58800 71000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 55600 70800 57000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 55600 71000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54000 70800 55400 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 54000 71000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal5 s 52400 70800 53800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 52400 71000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 46000 70800 49000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal5 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal5 s 42800 70800 45800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal5 s 41200 70800 42600 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 46000 71000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 41200 71000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 39600 70800 41000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal5 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal5 s 70800 39600 71000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 25200 70800 26600 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 36400 70800 39400 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 36400 71000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 25200 71000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 33200 70800 36200 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 20400 70800 23400 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 20400 71000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 17200 70800 20200 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 33200 71000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 17200 71000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 14000 70800 17000 71000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 14000 71000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 30000 70800 33000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 70800 14000 71000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 30000 71000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 26800 70800 29800 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 70800 26800 71000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 23600 70800 25000 71000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 14000 71000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 70800 23600 71000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal4 s 70800 23600 71000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 70800 23600 71000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal5 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal5 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal5 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal5 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal5 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal5 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal5 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal5 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal5 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal5 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
rlabel metal5 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal5 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal5 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal5 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal5 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal5 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal5 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal4 s 69026 70220 69026 70220 4 DVSS
port 2 nsew
rlabel metal4 s 70548 51411 70548 51411 4 VDD
port 3 nsew
rlabel metal4 s 65891 70220 65891 70220 4 DVSS
port 2 nsew
rlabel metal4 s 62716 70220 62716 70220 4 VDD
port 3 nsew
rlabel metal4 s 59509 70220 59509 70220 4 DVDD
port 1 nsew
rlabel metal4 s 56327 70220 56327 70220 4 DVDD
port 1 nsew
rlabel metal4 s 53064 70220 53064 70220 4 DVDD
port 1 nsew
rlabel metal4 s 49849 70219 49849 70219 4 VSS
port 4 nsew
rlabel metal4 s 44292 70220 44292 70220 4 DVDD
port 1 nsew
rlabel metal4 s 40319 70220 40319 70220 4 DVSS
port 2 nsew
rlabel metal4 s 34449 70220 34449 70220 4 DVDD
port 1 nsew
rlabel metal4 s 28097 70220 28097 70220 4 DVDD
port 1 nsew
rlabel metal4 s 23985 70220 23985 70220 4 DVDD
port 1 nsew
rlabel metal4 s 18634 70150 18634 70150 4 DVSS
port 2 nsew
rlabel metal4 s 70444 67411 70444 67411 4 DVDD
port 1 nsew
rlabel metal4 s 70444 59576 70444 59576 4 DVDD
port 1 nsew
rlabel metal4 s 70444 54611 70444 54611 4 DVDD
port 1 nsew
rlabel metal4 s 70444 44321 70444 44321 4 DVDD
port 1 nsew
rlabel metal4 s 70444 37912 70444 37912 4 DVDD
port 1 nsew
rlabel metal4 s 70444 31562 70444 31562 4 DVDD
port 1 nsew
rlabel metal4 s 70444 24237 70444 24237 4 DVDD
port 1 nsew
rlabel metal4 s 70444 69002 70444 69002 4 DVSS
port 2 nsew
rlabel metal4 s 70444 61011 70444 61011 4 DVSS
port 2 nsew
rlabel metal4 s 70444 47548 70444 47548 4 DVSS
port 2 nsew
rlabel metal4 s 70444 26053 70444 26053 4 DVSS
port 2 nsew
rlabel metal4 s 70422 15703 70422 15703 4 DVSS
port 2 nsew
rlabel metal4 s 67482 70220 67482 70220 4 DVDD
port 1 nsew
rlabel metal4 s 70547 49976 70547 49976 4 VSS
port 4 nsew
rlabel metal4 s 64328 70220 64328 70220 4 VSS
port 4 nsew
rlabel metal4 s 61124 70220 61124 70220 4 DVSS
port 2 nsew
rlabel metal4 s 57931 70220 57931 70220 4 DVSS
port 2 nsew
rlabel metal4 s 54690 70220 54690 70220 4 DVDD
port 1 nsew
rlabel metal4 s 51498 70220 51498 70220 4 VDD
port 3 nsew
rlabel metal4 s 47523 70220 47523 70220 4 DVSS
port 2 nsew
rlabel metal4 s 41877 70220 41877 70220 4 DVDD
port 1 nsew
rlabel metal4 s 37671 70220 37671 70220 4 DVDD
port 1 nsew
rlabel metal4 s 31313 70220 31313 70220 4 DVDD
port 1 nsew
rlabel metal4 s 25800 70220 25800 70220 4 DVSS
port 2 nsew
rlabel metal4 s 21613 70220 21613 70220 4 DVSS
port 2 nsew
rlabel metal4 s 15448 70196 15448 70196 4 DVSS
port 2 nsew
rlabel metal4 s 70444 62776 70444 62776 4 VDD
port 3 nsew
rlabel metal4 s 70444 56376 70444 56376 4 DVDD
port 1 nsew
rlabel metal4 s 70444 53176 70444 53176 4 DVDD
port 1 nsew
rlabel metal4 s 70444 41930 70444 41930 4 DVDD
port 1 nsew
rlabel metal4 s 70444 34676 70444 34676 4 DVDD
port 1 nsew
rlabel metal4 s 70444 28347 70444 28347 4 DVDD
port 1 nsew
rlabel metal4 s 70444 64211 70444 64211 4 VSS
port 4 nsew
rlabel metal4 s 70444 65976 70444 65976 4 DVSS
port 2 nsew
rlabel metal4 s 70444 57811 70444 57811 4 DVSS
port 2 nsew
rlabel metal4 s 70444 40295 70444 40295 4 DVSS
port 2 nsew
rlabel metal4 s 70444 21860 70444 21860 4 DVSS
port 2 nsew
rlabel metal4 s 70375 18874 70375 18874 4 DVSS
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string GDS_END 17526940
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17516202
string LEFclass ENDCAP BOTTOMLEFT
string LEFsite GF_COR_Site
string LEFsymmetry X Y R90
<< end >>
