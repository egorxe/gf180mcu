magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
use M1_NWELL$$44998700_R90_256x8m81  M1_NWELL$$44998700_R90_256x8m81_0
timestamp 1762296095
transform 0 -1 2322 1 0 4888
box 0 0 1 1
use M1_NWELL$$44998700_R90_256x8m81  M1_NWELL$$44998700_R90_256x8m81_1
timestamp 1762296095
transform 0 -1 4475 1 0 4888
box 0 0 1 1
use M1_NWELL$$46278700_256x8m81  M1_NWELL$$46278700_256x8m81_0
timestamp 1762296095
transform 1 0 3667 0 1 601
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1762296095
transform -1 0 3887 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1762296095
transform -1 0 4179 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1762296095
transform 1 0 4515 0 1 3185
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1762296095
transform -1 0 2989 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1762296095
transform 1 0 2354 0 1 3185
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1762296095
transform 1 0 2686 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1762296095
transform -1 0 3435 0 1 2378
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1762296095
transform 1 0 3287 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_1
timestamp 1762296095
transform 1 0 3117 0 1 4268
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_2
timestamp 1762296095
transform 1 0 2741 0 1 4698
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_3
timestamp 1762296095
transform 1 0 2137 0 1 5193
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_4
timestamp 1762296095
transform 1 0 2718 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_5
timestamp 1762296095
transform 1 0 4677 0 1 5193
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_6
timestamp 1762296095
transform 1 0 3435 0 1 6717
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_7
timestamp 1762296095
transform 1 0 3762 0 1 4268
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_8
timestamp 1762296095
transform 1 0 3573 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_9
timestamp 1762296095
transform 1 0 4166 0 1 4484
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_10
timestamp 1762296095
transform 1 0 4079 0 1 4700
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_0
timestamp 1762296095
transform 1 0 3619 0 1 1551
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_1
timestamp 1762296095
transform 1 0 4360 0 1 1539
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_2
timestamp 1762296095
transform 1 0 2959 0 1 1551
box 0 0 1 1
use M1_PSUB$$46554156_R90_256x8m81  M1_PSUB$$46554156_R90_256x8m81_0
timestamp 1762296095
transform 0 -1 2547 1 0 1031
box 0 0 1 1
use M1_PSUB$$46555180_256x8m81  M1_PSUB$$46555180_256x8m81_0
timestamp 1762296095
transform 1 0 3439 0 1 7080
box 0 0 1 1
use M1_PSUB$$46556204_256x8m81  M1_PSUB$$46556204_256x8m81_0
timestamp 1762296095
transform 1 0 1915 0 1 4550
box 0 0 1 1
use M1_PSUB$$46557228_256x8m81  M1_PSUB$$46557228_256x8m81_0
timestamp 1762296095
transform 1 0 2231 0 1 2020
box 0 0 1 1
use M1_PSUB$$46558252_256x8m81  M1_PSUB$$46558252_256x8m81_0
timestamp 1762296095
transform 1 0 3674 0 1 152
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_0
timestamp 1762296095
transform 1 0 4337 0 1 3178
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_1
timestamp 1762296095
transform 1 0 2528 0 1 3178
box 0 0 1 1
use nmos_1p2$$45107244_256x8m81  nmos_1p2$$45107244_256x8m81_0
timestamp 1762296095
transform -1 0 4243 0 -1 2156
box -31 0 -30 1
use nmos_1p2$$46550060_256x8m81  nmos_1p2$$46550060_256x8m81_0
timestamp 1762296095
transform 1 0 2620 0 1 2510
box -31 0 -30 1
use nmos_1p2$$46551084_256x8m81  nmos_1p2$$46551084_256x8m81_0
timestamp 1762296095
transform -1 0 3123 0 -1 2156
box -31 0 -30 1
use nmos_1p2$$46552108_256x8m81  nmos_1p2$$46552108_256x8m81_0
timestamp 1762296095
transform 1 0 2587 0 1 3317
box -31 0 -30 1
use nmos_1p2$$46553132_256x8m81  nmos_1p2$$46553132_256x8m81_0
timestamp 1762296095
transform 1 0 4379 0 1 3317
box -31 0 -30 1
use nmos_1p2$$46553132_256x8m81  nmos_1p2$$46553132_256x8m81_1
timestamp 1762296095
transform 1 0 2363 0 1 3317
box -31 0 -30 1
use pmos_1p2$$46285868_256x8m81  pmos_1p2$$46285868_256x8m81_0
timestamp 1762296095
transform 1 0 3406 0 1 5266
box -31 0 -30 1
use pmos_1p2$$46286892_256x8m81  pmos_1p2$$46286892_256x8m81_0
timestamp 1762296095
transform 1 0 3182 0 1 6132
box -31 0 -30 1
use pmos_1p2$$46549036_256x8m81  pmos_1p2$$46549036_256x8m81_0
timestamp 1762296095
transform -1 0 4243 0 -1 1331
box -31 0 -30 1
use pmos_1p2$$46896172_256x8m81  pmos_1p2$$46896172_256x8m81_0
timestamp 1762296095
transform 1 0 3052 0 1 4802
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_0
timestamp 1762296095
transform 1 0 2495 0 1 6132
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_1
timestamp 1762296095
transform 1 0 2495 0 1 5266
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_2
timestamp 1762296095
transform 1 0 4080 0 1 6132
box -31 0 -30 1
use pmos_1p2$$46897196_256x8m81  pmos_1p2$$46897196_256x8m81_3
timestamp 1762296095
transform 1 0 4080 0 1 5266
box -31 0 -30 1
use pmos_1p2$$46898220_256x8m81  pmos_1p2$$46898220_256x8m81_0
timestamp 1762296095
transform 1 0 2828 0 1 4802
box -31 0 -30 1
use pmos_1p2$$46898220_256x8m81  pmos_1p2$$46898220_256x8m81_1
timestamp 1762296095
transform 1 0 3948 0 1 4802
box -31 0 -30 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_0
timestamp 1762296095
transform 1 0 3386 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_1
timestamp 1762296095
transform 1 0 4909 0 1 827
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_2
timestamp 1762296095
transform 1 0 3834 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_3
timestamp 1762296095
transform -1 0 3700 0 -1 2201
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_4
timestamp 1762296095
transform -1 0 4146 0 -1 2201
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_5
timestamp 1762296095
transform 1 0 4271 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_6
timestamp 1762296095
transform 1 0 2938 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_7
timestamp 1762296095
transform -1 0 3033 0 -1 2029
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_8
timestamp 1762296095
transform 1 0 2523 0 1 827
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_9
timestamp 1762296095
transform 1 0 2523 0 1 1630
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_10
timestamp 1762296095
transform 1 0 2501 0 1 2621
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_11
timestamp 1762296095
transform 1 0 3050 0 1 6225
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_12
timestamp 1762296095
transform 1 0 2701 0 1 4665
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_13
timestamp 1762296095
transform 1 0 3151 0 1 4722
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_14
timestamp 1762296095
transform 1 0 2287 0 1 4722
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_15
timestamp 1762296095
transform 1 0 3623 0 1 4722
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_16
timestamp 1762296095
transform 1 0 3722 0 1 6225
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_17
timestamp 1762296095
transform 1 0 4040 0 1 4665
box 0 0 1 1
use via1_2_x2_256x8m81  via1_2_x2_256x8m81_18
timestamp 1762296095
transform 1 0 4418 0 1 4722
box 0 0 1 1
use via1_2_x2_R90_256x8m81  via1_2_x2_R90_256x8m81_0
timestamp 1762296095
transform 0 -1 3259 1 0 7937
box 0 0 1 1
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_0
timestamp 1762296095
transform 0 1 4262 -1 0 544
box 0 0 1 1
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_1
timestamp 1762296095
transform 0 1 2723 -1 0 544
box 0 0 1 1
use via1_2_x2_R270_256x8m81  via1_2_x2_R270_256x8m81_2
timestamp 1762296095
transform 0 1 3182 -1 0 544
box 0 0 1 1
use via1_256x8m81  via1_256x8m81_0
timestamp 1762296095
transform 1 0 3388 0 -1 6790
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_0
timestamp 1762296095
transform 0 -1 4506 1 0 3149
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_1
timestamp 1762296095
transform 0 -1 2486 1 0 3149
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_2
timestamp 1762296095
transform 0 -1 2520 1 0 4226
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_3
timestamp 1762296095
transform 0 -1 4396 1 0 4437
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_4
timestamp 1762296095
transform 0 -1 4568 1 0 4226
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_5
timestamp 1762296095
transform 0 -1 3595 1 0 5792
box 0 0 1 1
use via1_R90_256x8m81  via1_R90_256x8m81_6
timestamp 1762296095
transform 0 1 3276 1 0 5964
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_0
timestamp 1762296095
transform 0 -1 2925 -1 0 6762
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_1
timestamp 1762296095
transform 0 1 3083 -1 0 4321
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_2
timestamp 1762296095
transform 0 1 3193 -1 0 4532
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_3
timestamp 1762296095
transform 0 -1 3500 -1 0 7361
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_4
timestamp 1762296095
transform 0 -1 4060 -1 0 6740
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_5
timestamp 1762296095
transform 0 1 3659 -1 0 4321
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_6
timestamp 1762296095
transform 0 1 3371 -1 0 4321
box 0 0 1 1
use via1_R270_256x8m81  via1_R270_256x8m81_7
timestamp 1762296095
transform 0 1 3549 -1 0 4532
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_0
timestamp 1762296095
transform -1 0 4153 0 1 1018
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_1
timestamp 1762296095
transform 1 0 4276 0 1 1712
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_2
timestamp 1762296095
transform 1 0 3601 0 1 1018
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_3
timestamp 1762296095
transform -1 0 3920 0 1 1712
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_4
timestamp 1762296095
transform -1 0 3478 0 1 1712
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_5
timestamp 1762296095
transform 1 0 2596 0 1 6146
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_6
timestamp 1762296095
transform 1 0 4181 0 1 6146
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_7
timestamp 1762296095
transform 1 0 3503 0 1 6146
box 0 0 1 1
use via1_x2_256x8m81  via1_x2_256x8m81_8
timestamp 1762296095
transform -1 0 3369 0 1 6146
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_0
timestamp 1762296095
transform 0 -1 4559 1 0 1494
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_1
timestamp 1762296095
transform 0 -1 3057 1 0 1505
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_2
timestamp 1762296095
transform 0 -1 2633 1 0 7937
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_3
timestamp 1762296095
transform 0 -1 3015 1 0 7728
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_4
timestamp 1762296095
transform 0 -1 3819 1 0 7728
box 0 0 1 1
use via1_x2_R90_256x8m81  via1_x2_R90_256x8m81_5
timestamp 1762296095
transform 0 -1 4497 1 0 7937
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_0
timestamp 1762296095
transform 0 1 2684 -1 0 4532
box 0 0 1 1
use via1_x2_R270_256x8m81  via1_x2_R270_256x8m81_1
timestamp 1762296095
transform 0 1 3883 -1 0 4532
box 0 0 1 1
use via2_x2_R90_256x8m81  via2_x2_R90_256x8m81_0
timestamp 1762296095
transform 0 -1 1992 1 0 7728
box 0 0 1 1
<< properties >>
string GDS_END 476260
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 462254
<< end >>
