magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
<< nwell >>
rect 29138 44674 56005 45190
rect 29138 43555 32850 44674
rect 29138 35918 33473 43555
rect 35260 43535 39818 44674
rect 42526 44185 43793 44475
rect 42526 44108 44118 44185
rect 42527 43535 44118 44108
rect 45169 43554 49764 44674
rect 35260 43505 39464 43535
rect 35124 43433 39464 43505
rect 35124 35949 37639 43433
rect 30658 35917 33473 35918
rect 31003 35899 33473 35917
rect 38864 35899 39464 43433
rect 44662 43504 49764 43554
rect 52285 43536 56005 44674
rect 44662 35950 50000 43504
rect 51652 43433 56005 43536
rect 44662 35900 48709 35950
rect 51652 35918 55985 43433
rect 54025 35917 54467 35918
<< pwell >>
rect 1774 44282 24710 44314
rect 1774 35138 24710 35170
<< mvnmos >>
rect 33001 43799 35023 43919
rect 40062 43799 40590 43919
rect 40963 43800 42281 43920
rect 44432 43799 44960 43919
rect 50001 43799 52023 43919
rect 33671 43155 34671 43275
rect 39727 43155 40167 43275
rect 43695 43144 44325 43264
rect 33671 42931 34671 43051
rect 50454 43155 51454 43275
rect 33671 42675 34671 42795
rect 37896 42844 38556 42964
rect 43695 42931 44325 43051
rect 37896 42620 38556 42740
rect 39598 42620 39730 42740
rect 43695 42707 44325 42827
rect 50454 42931 51454 43051
rect 50454 42675 51454 42795
rect 33671 42059 34671 42179
rect 33671 41803 34671 41923
rect 37896 42114 38556 42234
rect 37896 41890 38556 42010
rect 39598 42114 39730 42234
rect 43695 42027 44325 42147
rect 50454 42059 51454 42179
rect 43695 41803 44325 41923
rect 50454 41803 51454 41923
rect 33671 41579 34671 41699
rect 33671 41355 34671 41475
rect 39727 41579 40167 41699
rect 43695 41590 44325 41710
rect 39727 41355 40167 41475
rect 50454 41579 51454 41699
rect 43695 41344 44325 41464
rect 33671 41131 34671 41251
rect 50454 41355 51454 41475
rect 33671 40875 34671 40995
rect 37896 41044 38556 41164
rect 43695 41131 44325 41251
rect 37896 40820 38556 40940
rect 39598 40820 39730 40940
rect 43695 40907 44325 41027
rect 50454 41131 51454 41251
rect 50454 40875 51454 40995
rect 33671 40259 34671 40379
rect 33671 40003 34671 40123
rect 37896 40314 38556 40434
rect 37896 40090 38556 40210
rect 39598 40314 39730 40434
rect 43695 40227 44325 40347
rect 50454 40259 51454 40379
rect 43695 40003 44325 40123
rect 50454 40003 51454 40123
rect 33671 39779 34671 39899
rect 33671 39555 34671 39675
rect 39727 39779 40167 39899
rect 43695 39790 44325 39910
rect 39727 39555 40167 39675
rect 50454 39779 51454 39899
rect 43695 39544 44325 39664
rect 33671 39331 34671 39451
rect 50454 39555 51454 39675
rect 33671 39075 34671 39195
rect 37896 39244 38556 39364
rect 43695 39331 44325 39451
rect 37896 39020 38556 39140
rect 39598 39020 39730 39140
rect 43695 39107 44325 39227
rect 50454 39331 51454 39451
rect 50454 39075 51454 39195
rect 33671 38459 34671 38579
rect 33671 38203 34671 38323
rect 37896 38514 38556 38634
rect 37896 38290 38556 38410
rect 39598 38514 39730 38634
rect 43695 38427 44325 38547
rect 50454 38459 51454 38579
rect 43695 38203 44325 38323
rect 50454 38203 51454 38323
rect 33671 37979 34671 38099
rect 33671 37755 34671 37875
rect 39727 37979 40167 38099
rect 43695 37990 44325 38110
rect 39727 37755 40167 37875
rect 50454 37979 51454 38099
rect 43695 37744 44325 37864
rect 33671 37531 34671 37651
rect 50454 37755 51454 37875
rect 33671 37275 34671 37395
rect 37896 37444 38556 37564
rect 43695 37531 44325 37651
rect 37896 37220 38556 37340
rect 39598 37220 39730 37340
rect 43695 37307 44325 37427
rect 50454 37531 51454 37651
rect 50454 37275 51454 37395
rect 33671 36659 34671 36779
rect 33671 36403 34671 36523
rect 37896 36714 38556 36834
rect 37896 36490 38556 36610
rect 39598 36714 39730 36834
rect 43695 36627 44325 36747
rect 50454 36659 51454 36779
rect 43695 36403 44325 36523
rect 50454 36403 51454 36523
rect 33671 36179 34671 36299
rect 39727 36179 40167 36299
rect 43695 36190 44325 36310
rect 50454 36179 51454 36299
<< mvpmos >>
rect 29274 43383 30373 44171
rect 35396 44023 37922 44143
rect 35396 43799 37922 43919
rect 38363 43799 39681 43919
rect 42663 43799 43981 43919
rect 45333 43799 46651 43919
rect 47101 44023 49627 44143
rect 47101 43799 49627 43919
rect 29274 42483 30373 43271
rect 31336 43155 33336 43275
rect 31336 42931 33336 43051
rect 31336 42707 33336 42827
rect 44799 43155 45323 43275
rect 51789 43155 53789 43275
rect 54750 43383 55849 44171
rect 35260 42844 36360 42964
rect 35260 42620 36360 42740
rect 36841 42844 37501 42964
rect 44799 42931 45323 43051
rect 36841 42620 37501 42740
rect 39008 42620 39326 42740
rect 44799 42707 45323 42827
rect 48765 42844 49865 42964
rect 48765 42620 49865 42740
rect 51789 42931 53789 43051
rect 51789 42707 53789 42827
rect 29274 41583 30373 42371
rect 54750 42483 55849 43271
rect 31336 42027 33336 42147
rect 31336 41803 33336 41923
rect 29274 40683 30373 41471
rect 31336 41579 33336 41699
rect 35260 42114 36360 42234
rect 35260 41890 36360 42010
rect 36841 42114 37501 42234
rect 36841 41890 37501 42010
rect 39008 42114 39326 42234
rect 44799 42027 45323 42147
rect 48765 42114 49865 42234
rect 44799 41803 45323 41923
rect 48765 41890 49865 42010
rect 31336 41355 33336 41475
rect 31336 41131 33336 41251
rect 31336 40907 33336 41027
rect 44799 41579 45323 41699
rect 51789 42027 53789 42147
rect 51789 41803 53789 41923
rect 51789 41579 53789 41699
rect 44799 41355 45323 41475
rect 51789 41355 53789 41475
rect 54750 41583 55849 42371
rect 35260 41044 36360 41164
rect 35260 40820 36360 40940
rect 36841 41044 37501 41164
rect 44799 41131 45323 41251
rect 36841 40820 37501 40940
rect 39008 40820 39326 40940
rect 44799 40907 45323 41027
rect 48765 41044 49865 41164
rect 48765 40820 49865 40940
rect 51789 41131 53789 41251
rect 51789 40907 53789 41027
rect 29274 39783 30373 40571
rect 54750 40683 55849 41471
rect 31336 40227 33336 40347
rect 31336 40003 33336 40123
rect 29274 38883 30373 39671
rect 31336 39779 33336 39899
rect 35260 40314 36360 40434
rect 35260 40090 36360 40210
rect 36841 40314 37501 40434
rect 36841 40090 37501 40210
rect 39008 40314 39326 40434
rect 44799 40227 45323 40347
rect 48765 40314 49865 40434
rect 44799 40003 45323 40123
rect 48765 40090 49865 40210
rect 31336 39555 33336 39675
rect 31336 39331 33336 39451
rect 31336 39107 33336 39227
rect 44799 39779 45323 39899
rect 51789 40227 53789 40347
rect 51789 40003 53789 40123
rect 51789 39779 53789 39899
rect 44799 39555 45323 39675
rect 51789 39555 53789 39675
rect 54750 39783 55849 40571
rect 35260 39244 36360 39364
rect 35260 39020 36360 39140
rect 36841 39244 37501 39364
rect 44799 39331 45323 39451
rect 36841 39020 37501 39140
rect 39008 39020 39326 39140
rect 44799 39107 45323 39227
rect 48765 39244 49865 39364
rect 48765 39020 49865 39140
rect 51789 39331 53789 39451
rect 51789 39107 53789 39227
rect 29274 37983 30373 38771
rect 54750 38883 55849 39671
rect 31336 38427 33336 38547
rect 31336 38203 33336 38323
rect 29274 37083 30373 37871
rect 31336 37979 33336 38099
rect 35260 38514 36360 38634
rect 35260 38290 36360 38410
rect 36841 38514 37501 38634
rect 36841 38290 37501 38410
rect 39008 38514 39326 38634
rect 44799 38427 45323 38547
rect 48765 38514 49865 38634
rect 44799 38203 45323 38323
rect 48765 38290 49865 38410
rect 31336 37755 33336 37875
rect 31336 37531 33336 37651
rect 31336 37307 33336 37427
rect 44799 37979 45323 38099
rect 51789 38427 53789 38547
rect 51789 38203 53789 38323
rect 51789 37979 53789 38099
rect 44799 37755 45323 37875
rect 51789 37755 53789 37875
rect 54750 37983 55849 38771
rect 35260 37444 36360 37564
rect 35260 37220 36360 37340
rect 36841 37444 37501 37564
rect 44799 37531 45323 37651
rect 36841 37220 37501 37340
rect 39008 37220 39326 37340
rect 44799 37307 45323 37427
rect 48765 37444 49865 37564
rect 48765 37220 49865 37340
rect 51789 37531 53789 37651
rect 51789 37307 53789 37427
rect 29274 36183 30373 36971
rect 54750 37083 55849 37871
rect 31336 36627 33336 36747
rect 31336 36403 33336 36523
rect 31336 36179 33336 36299
rect 35260 36714 36360 36834
rect 35260 36490 36360 36610
rect 36841 36714 37501 36834
rect 36841 36490 37501 36610
rect 39008 36714 39326 36834
rect 44799 36627 45323 36747
rect 48765 36714 49865 36834
rect 44799 36403 45323 36523
rect 48765 36490 49865 36610
rect 44799 36179 45323 36299
rect 51789 36627 53789 36747
rect 51789 36403 53789 36523
rect 51789 36179 53789 36299
rect 54750 36183 55849 36971
<< mvndiff >>
rect 33001 43994 35023 44007
rect 33001 43948 33014 43994
rect 33774 43948 33831 43994
rect 33877 43948 33934 43994
rect 33980 43948 34037 43994
rect 34083 43948 34140 43994
rect 34186 43948 34243 43994
rect 34289 43948 34346 43994
rect 34392 43948 34449 43994
rect 34495 43948 34552 43994
rect 34598 43948 34655 43994
rect 34701 43948 34758 43994
rect 34804 43948 34861 43994
rect 34907 43948 34964 43994
rect 35010 43948 35023 43994
rect 33001 43919 35023 43948
rect 40062 43994 40590 44007
rect 40062 43948 40075 43994
rect 40121 43948 40189 43994
rect 40235 43948 40303 43994
rect 40349 43948 40417 43994
rect 40463 43948 40531 43994
rect 40577 43948 40590 43994
rect 40963 43995 42281 44008
rect 40062 43919 40590 43948
rect 40963 43949 40976 43995
rect 41022 43949 41079 43995
rect 41125 43949 41182 43995
rect 41228 43949 41286 43995
rect 41332 43949 41390 43995
rect 41436 43949 41494 43995
rect 41540 43949 41598 43995
rect 41644 43949 41702 43995
rect 41748 43949 41806 43995
rect 41852 43949 41910 43995
rect 41956 43949 42014 43995
rect 42060 43949 42118 43995
rect 42164 43949 42222 43995
rect 42268 43949 42281 43995
rect 40963 43920 42281 43949
rect 33001 43770 35023 43799
rect 33001 43724 33014 43770
rect 33774 43724 33831 43770
rect 33877 43724 33934 43770
rect 33980 43724 34037 43770
rect 34083 43724 34140 43770
rect 34186 43724 34243 43770
rect 34289 43724 34346 43770
rect 34392 43724 34449 43770
rect 34495 43724 34552 43770
rect 34598 43724 34655 43770
rect 34701 43724 34758 43770
rect 34804 43724 34861 43770
rect 34907 43724 34964 43770
rect 35010 43724 35023 43770
rect 33001 43711 35023 43724
rect 40062 43770 40590 43799
rect 40062 43724 40075 43770
rect 40121 43724 40189 43770
rect 40235 43724 40303 43770
rect 40349 43724 40417 43770
rect 40463 43724 40531 43770
rect 40577 43724 40590 43770
rect 40062 43711 40590 43724
rect 40963 43771 42281 43800
rect 44432 43994 44960 44007
rect 44432 43948 44445 43994
rect 44491 43948 44559 43994
rect 44605 43948 44673 43994
rect 44719 43948 44787 43994
rect 44833 43948 44901 43994
rect 44947 43948 44960 43994
rect 44432 43919 44960 43948
rect 50001 43994 52023 44007
rect 50001 43948 50014 43994
rect 50774 43948 50831 43994
rect 50877 43948 50934 43994
rect 50980 43948 51037 43994
rect 51083 43948 51140 43994
rect 51186 43948 51243 43994
rect 51289 43948 51346 43994
rect 51392 43948 51449 43994
rect 51495 43948 51552 43994
rect 51598 43948 51655 43994
rect 51701 43948 51758 43994
rect 51804 43948 51861 43994
rect 51907 43948 51964 43994
rect 52010 43948 52023 43994
rect 50001 43919 52023 43948
rect 40963 43725 40976 43771
rect 41022 43725 41079 43771
rect 41125 43725 41182 43771
rect 41228 43725 41286 43771
rect 41332 43725 41390 43771
rect 41436 43725 41494 43771
rect 41540 43725 41598 43771
rect 41644 43725 41702 43771
rect 41748 43725 41806 43771
rect 41852 43725 41910 43771
rect 41956 43725 42014 43771
rect 42060 43725 42118 43771
rect 42164 43725 42222 43771
rect 42268 43725 42281 43771
rect 40963 43712 42281 43725
rect 44432 43770 44960 43799
rect 44432 43724 44445 43770
rect 44491 43724 44559 43770
rect 44605 43724 44673 43770
rect 44719 43724 44787 43770
rect 44833 43724 44901 43770
rect 44947 43724 44960 43770
rect 44432 43711 44960 43724
rect 50001 43770 52023 43799
rect 50001 43724 50014 43770
rect 50774 43724 50831 43770
rect 50877 43724 50934 43770
rect 50980 43724 51037 43770
rect 51083 43724 51140 43770
rect 51186 43724 51243 43770
rect 51289 43724 51346 43770
rect 51392 43724 51449 43770
rect 51495 43724 51552 43770
rect 51598 43724 51655 43770
rect 51701 43724 51758 43770
rect 51804 43724 51861 43770
rect 51907 43724 51964 43770
rect 52010 43724 52023 43770
rect 50001 43711 52023 43724
rect 33671 43350 34671 43363
rect 33671 43304 33684 43350
rect 33730 43304 33787 43350
rect 33833 43304 33890 43350
rect 33936 43304 33993 43350
rect 34039 43304 34096 43350
rect 34142 43304 34199 43350
rect 34245 43304 34302 43350
rect 34348 43304 34405 43350
rect 34451 43304 34508 43350
rect 34554 43304 34612 43350
rect 34658 43304 34671 43350
rect 33671 43275 34671 43304
rect 39727 43350 40167 43363
rect 39727 43304 39740 43350
rect 39786 43304 39862 43350
rect 39908 43304 39985 43350
rect 40031 43304 40108 43350
rect 40154 43304 40167 43350
rect 39727 43275 40167 43304
rect 43695 43350 44325 43396
rect 43695 43304 43739 43350
rect 43785 43304 43906 43350
rect 43952 43304 44071 43350
rect 44117 43304 44236 43350
rect 44282 43304 44325 43350
rect 43695 43264 44325 43304
rect 33671 43126 34671 43155
rect 33671 43080 33684 43126
rect 33730 43080 33787 43126
rect 33833 43080 33890 43126
rect 33936 43080 33993 43126
rect 34039 43080 34096 43126
rect 34142 43080 34199 43126
rect 34245 43080 34302 43126
rect 34348 43080 34405 43126
rect 34451 43080 34508 43126
rect 34554 43080 34612 43126
rect 34658 43080 34671 43126
rect 33671 43051 34671 43080
rect 39727 43126 40167 43155
rect 39727 43080 39740 43126
rect 39786 43080 39862 43126
rect 39908 43080 39985 43126
rect 40031 43080 40108 43126
rect 40154 43080 40167 43126
rect 39727 43067 40167 43080
rect 50454 43350 51454 43363
rect 50454 43304 50467 43350
rect 50513 43304 50571 43350
rect 50617 43304 50674 43350
rect 50720 43304 50777 43350
rect 50823 43304 50880 43350
rect 50926 43304 50983 43350
rect 51029 43304 51086 43350
rect 51132 43304 51189 43350
rect 51235 43304 51292 43350
rect 51338 43304 51395 43350
rect 51441 43304 51454 43350
rect 50454 43275 51454 43304
rect 37896 43039 38556 43052
rect 43695 43051 44325 43144
rect 50454 43126 51454 43155
rect 50454 43080 50467 43126
rect 50513 43080 50571 43126
rect 50617 43080 50674 43126
rect 50720 43080 50777 43126
rect 50823 43080 50880 43126
rect 50926 43080 50983 43126
rect 51029 43080 51086 43126
rect 51132 43080 51189 43126
rect 51235 43080 51292 43126
rect 51338 43080 51395 43126
rect 51441 43080 51454 43126
rect 37896 42993 37909 43039
rect 37955 42993 38026 43039
rect 38072 42993 38143 43039
rect 38189 42993 38261 43039
rect 38307 42993 38379 43039
rect 38425 42993 38497 43039
rect 38543 42993 38556 43039
rect 37896 42964 38556 42993
rect 33671 42902 34671 42931
rect 33671 42856 33684 42902
rect 33730 42856 33787 42902
rect 33833 42856 33890 42902
rect 33936 42856 33993 42902
rect 34039 42856 34096 42902
rect 34142 42856 34199 42902
rect 34245 42856 34302 42902
rect 34348 42856 34405 42902
rect 34451 42856 34508 42902
rect 34554 42856 34612 42902
rect 34658 42856 34671 42902
rect 33671 42795 34671 42856
rect 33671 42643 34671 42675
rect 33671 42597 33816 42643
rect 33862 42597 34002 42643
rect 34048 42597 34189 42643
rect 34235 42597 34376 42643
rect 34422 42597 34562 42643
rect 34608 42597 34671 42643
rect 50454 43051 51454 43080
rect 37896 42815 38556 42844
rect 37896 42769 37909 42815
rect 37955 42769 38026 42815
rect 38072 42769 38143 42815
rect 38189 42769 38261 42815
rect 38307 42769 38379 42815
rect 38425 42769 38497 42815
rect 38543 42769 38556 42815
rect 37896 42740 38556 42769
rect 39598 42815 39730 42828
rect 43695 42827 44325 42931
rect 39598 42769 39641 42815
rect 39687 42769 39730 42815
rect 39598 42740 39730 42769
rect 50454 42902 51454 42931
rect 50454 42856 50467 42902
rect 50513 42856 50571 42902
rect 50617 42856 50674 42902
rect 50720 42856 50777 42902
rect 50823 42856 50880 42902
rect 50926 42856 50983 42902
rect 51029 42856 51086 42902
rect 51132 42856 51189 42902
rect 51235 42856 51292 42902
rect 51338 42856 51395 42902
rect 51441 42856 51454 42902
rect 50454 42795 51454 42856
rect 43695 42657 44325 42707
rect 33671 42551 34671 42597
rect 37896 42591 38556 42620
rect 37896 42545 37909 42591
rect 37955 42545 38026 42591
rect 38072 42545 38143 42591
rect 38189 42545 38261 42591
rect 38307 42545 38379 42591
rect 38425 42545 38497 42591
rect 38543 42545 38556 42591
rect 37896 42532 38556 42545
rect 39598 42591 39730 42620
rect 39598 42545 39641 42591
rect 39687 42545 39730 42591
rect 43695 42611 43739 42657
rect 43785 42611 43906 42657
rect 43952 42611 44071 42657
rect 44117 42611 44236 42657
rect 44282 42611 44325 42657
rect 50454 42643 51454 42675
rect 43695 42564 44325 42611
rect 39598 42532 39730 42545
rect 50454 42597 50516 42643
rect 50562 42597 50703 42643
rect 50749 42597 50890 42643
rect 50936 42597 51076 42643
rect 51122 42597 51263 42643
rect 51309 42597 51454 42643
rect 50454 42551 51454 42597
rect 33671 42257 34671 42303
rect 33671 42211 33816 42257
rect 33862 42211 34002 42257
rect 34048 42211 34189 42257
rect 34235 42211 34376 42257
rect 34422 42211 34562 42257
rect 34608 42211 34671 42257
rect 37896 42309 38556 42322
rect 37896 42263 37909 42309
rect 37955 42263 38026 42309
rect 38072 42263 38143 42309
rect 38189 42263 38261 42309
rect 38307 42263 38379 42309
rect 38425 42263 38497 42309
rect 38543 42263 38556 42309
rect 37896 42234 38556 42263
rect 39598 42309 39730 42322
rect 39598 42263 39641 42309
rect 39687 42263 39730 42309
rect 39598 42234 39730 42263
rect 43695 42243 44325 42290
rect 33671 42179 34671 42211
rect 33671 41998 34671 42059
rect 33671 41952 33684 41998
rect 33730 41952 33787 41998
rect 33833 41952 33890 41998
rect 33936 41952 33993 41998
rect 34039 41952 34096 41998
rect 34142 41952 34199 41998
rect 34245 41952 34302 41998
rect 34348 41952 34405 41998
rect 34451 41952 34508 41998
rect 34554 41952 34612 41998
rect 34658 41952 34671 41998
rect 33671 41923 34671 41952
rect 37896 42085 38556 42114
rect 37896 42039 37909 42085
rect 37955 42039 38026 42085
rect 38072 42039 38143 42085
rect 38189 42039 38261 42085
rect 38307 42039 38379 42085
rect 38425 42039 38497 42085
rect 38543 42039 38556 42085
rect 37896 42010 38556 42039
rect 43695 42197 43739 42243
rect 43785 42197 43906 42243
rect 43952 42197 44071 42243
rect 44117 42197 44236 42243
rect 44282 42197 44325 42243
rect 43695 42147 44325 42197
rect 50454 42257 51454 42303
rect 39598 42085 39730 42114
rect 39598 42039 39641 42085
rect 39687 42039 39730 42085
rect 39598 42026 39730 42039
rect 50454 42211 50516 42257
rect 50562 42211 50703 42257
rect 50749 42211 50890 42257
rect 50936 42211 51076 42257
rect 51122 42211 51263 42257
rect 51309 42211 51454 42257
rect 50454 42179 51454 42211
rect 43695 41923 44325 42027
rect 33671 41774 34671 41803
rect 37896 41861 38556 41890
rect 37896 41815 37909 41861
rect 37955 41815 38026 41861
rect 38072 41815 38143 41861
rect 38189 41815 38261 41861
rect 38307 41815 38379 41861
rect 38425 41815 38497 41861
rect 38543 41815 38556 41861
rect 37896 41802 38556 41815
rect 50454 41998 51454 42059
rect 50454 41952 50467 41998
rect 50513 41952 50571 41998
rect 50617 41952 50674 41998
rect 50720 41952 50777 41998
rect 50823 41952 50880 41998
rect 50926 41952 50983 41998
rect 51029 41952 51086 41998
rect 51132 41952 51189 41998
rect 51235 41952 51292 41998
rect 51338 41952 51395 41998
rect 51441 41952 51454 41998
rect 50454 41923 51454 41952
rect 33671 41728 33684 41774
rect 33730 41728 33787 41774
rect 33833 41728 33890 41774
rect 33936 41728 33993 41774
rect 34039 41728 34096 41774
rect 34142 41728 34199 41774
rect 34245 41728 34302 41774
rect 34348 41728 34405 41774
rect 34451 41728 34508 41774
rect 34554 41728 34612 41774
rect 34658 41728 34671 41774
rect 33671 41699 34671 41728
rect 39727 41774 40167 41787
rect 39727 41728 39740 41774
rect 39786 41728 39862 41774
rect 39908 41728 39985 41774
rect 40031 41728 40108 41774
rect 40154 41728 40167 41774
rect 39727 41699 40167 41728
rect 43695 41710 44325 41803
rect 50454 41774 51454 41803
rect 33671 41550 34671 41579
rect 33671 41504 33684 41550
rect 33730 41504 33787 41550
rect 33833 41504 33890 41550
rect 33936 41504 33993 41550
rect 34039 41504 34096 41550
rect 34142 41504 34199 41550
rect 34245 41504 34302 41550
rect 34348 41504 34405 41550
rect 34451 41504 34508 41550
rect 34554 41504 34612 41550
rect 34658 41504 34671 41550
rect 33671 41475 34671 41504
rect 39727 41550 40167 41579
rect 39727 41504 39740 41550
rect 39786 41504 39862 41550
rect 39908 41504 39985 41550
rect 40031 41504 40108 41550
rect 40154 41504 40167 41550
rect 39727 41475 40167 41504
rect 43695 41550 44325 41590
rect 50454 41728 50467 41774
rect 50513 41728 50571 41774
rect 50617 41728 50674 41774
rect 50720 41728 50777 41774
rect 50823 41728 50880 41774
rect 50926 41728 50983 41774
rect 51029 41728 51086 41774
rect 51132 41728 51189 41774
rect 51235 41728 51292 41774
rect 51338 41728 51395 41774
rect 51441 41728 51454 41774
rect 50454 41699 51454 41728
rect 43695 41504 43739 41550
rect 43785 41504 43906 41550
rect 43952 41504 44071 41550
rect 44117 41504 44236 41550
rect 44282 41504 44325 41550
rect 43695 41464 44325 41504
rect 33671 41326 34671 41355
rect 33671 41280 33684 41326
rect 33730 41280 33787 41326
rect 33833 41280 33890 41326
rect 33936 41280 33993 41326
rect 34039 41280 34096 41326
rect 34142 41280 34199 41326
rect 34245 41280 34302 41326
rect 34348 41280 34405 41326
rect 34451 41280 34508 41326
rect 34554 41280 34612 41326
rect 34658 41280 34671 41326
rect 33671 41251 34671 41280
rect 39727 41326 40167 41355
rect 39727 41280 39740 41326
rect 39786 41280 39862 41326
rect 39908 41280 39985 41326
rect 40031 41280 40108 41326
rect 40154 41280 40167 41326
rect 39727 41267 40167 41280
rect 50454 41550 51454 41579
rect 50454 41504 50467 41550
rect 50513 41504 50571 41550
rect 50617 41504 50674 41550
rect 50720 41504 50777 41550
rect 50823 41504 50880 41550
rect 50926 41504 50983 41550
rect 51029 41504 51086 41550
rect 51132 41504 51189 41550
rect 51235 41504 51292 41550
rect 51338 41504 51395 41550
rect 51441 41504 51454 41550
rect 50454 41475 51454 41504
rect 37896 41239 38556 41252
rect 43695 41251 44325 41344
rect 50454 41326 51454 41355
rect 50454 41280 50467 41326
rect 50513 41280 50571 41326
rect 50617 41280 50674 41326
rect 50720 41280 50777 41326
rect 50823 41280 50880 41326
rect 50926 41280 50983 41326
rect 51029 41280 51086 41326
rect 51132 41280 51189 41326
rect 51235 41280 51292 41326
rect 51338 41280 51395 41326
rect 51441 41280 51454 41326
rect 37896 41193 37909 41239
rect 37955 41193 38026 41239
rect 38072 41193 38143 41239
rect 38189 41193 38261 41239
rect 38307 41193 38379 41239
rect 38425 41193 38497 41239
rect 38543 41193 38556 41239
rect 37896 41164 38556 41193
rect 33671 41102 34671 41131
rect 33671 41056 33684 41102
rect 33730 41056 33787 41102
rect 33833 41056 33890 41102
rect 33936 41056 33993 41102
rect 34039 41056 34096 41102
rect 34142 41056 34199 41102
rect 34245 41056 34302 41102
rect 34348 41056 34405 41102
rect 34451 41056 34508 41102
rect 34554 41056 34612 41102
rect 34658 41056 34671 41102
rect 33671 40995 34671 41056
rect 33671 40843 34671 40875
rect 33671 40797 33816 40843
rect 33862 40797 34002 40843
rect 34048 40797 34189 40843
rect 34235 40797 34376 40843
rect 34422 40797 34562 40843
rect 34608 40797 34671 40843
rect 50454 41251 51454 41280
rect 37896 41015 38556 41044
rect 37896 40969 37909 41015
rect 37955 40969 38026 41015
rect 38072 40969 38143 41015
rect 38189 40969 38261 41015
rect 38307 40969 38379 41015
rect 38425 40969 38497 41015
rect 38543 40969 38556 41015
rect 37896 40940 38556 40969
rect 39598 41015 39730 41028
rect 43695 41027 44325 41131
rect 39598 40969 39641 41015
rect 39687 40969 39730 41015
rect 39598 40940 39730 40969
rect 50454 41102 51454 41131
rect 50454 41056 50467 41102
rect 50513 41056 50571 41102
rect 50617 41056 50674 41102
rect 50720 41056 50777 41102
rect 50823 41056 50880 41102
rect 50926 41056 50983 41102
rect 51029 41056 51086 41102
rect 51132 41056 51189 41102
rect 51235 41056 51292 41102
rect 51338 41056 51395 41102
rect 51441 41056 51454 41102
rect 50454 40995 51454 41056
rect 43695 40857 44325 40907
rect 33671 40751 34671 40797
rect 37896 40791 38556 40820
rect 37896 40745 37909 40791
rect 37955 40745 38026 40791
rect 38072 40745 38143 40791
rect 38189 40745 38261 40791
rect 38307 40745 38379 40791
rect 38425 40745 38497 40791
rect 38543 40745 38556 40791
rect 37896 40732 38556 40745
rect 39598 40791 39730 40820
rect 39598 40745 39641 40791
rect 39687 40745 39730 40791
rect 43695 40811 43739 40857
rect 43785 40811 43906 40857
rect 43952 40811 44071 40857
rect 44117 40811 44236 40857
rect 44282 40811 44325 40857
rect 50454 40843 51454 40875
rect 43695 40764 44325 40811
rect 39598 40732 39730 40745
rect 50454 40797 50516 40843
rect 50562 40797 50703 40843
rect 50749 40797 50890 40843
rect 50936 40797 51076 40843
rect 51122 40797 51263 40843
rect 51309 40797 51454 40843
rect 50454 40751 51454 40797
rect 33671 40457 34671 40503
rect 33671 40411 33816 40457
rect 33862 40411 34002 40457
rect 34048 40411 34189 40457
rect 34235 40411 34376 40457
rect 34422 40411 34562 40457
rect 34608 40411 34671 40457
rect 37896 40509 38556 40522
rect 37896 40463 37909 40509
rect 37955 40463 38026 40509
rect 38072 40463 38143 40509
rect 38189 40463 38261 40509
rect 38307 40463 38379 40509
rect 38425 40463 38497 40509
rect 38543 40463 38556 40509
rect 37896 40434 38556 40463
rect 39598 40509 39730 40522
rect 39598 40463 39641 40509
rect 39687 40463 39730 40509
rect 39598 40434 39730 40463
rect 43695 40443 44325 40490
rect 33671 40379 34671 40411
rect 33671 40198 34671 40259
rect 33671 40152 33684 40198
rect 33730 40152 33787 40198
rect 33833 40152 33890 40198
rect 33936 40152 33993 40198
rect 34039 40152 34096 40198
rect 34142 40152 34199 40198
rect 34245 40152 34302 40198
rect 34348 40152 34405 40198
rect 34451 40152 34508 40198
rect 34554 40152 34612 40198
rect 34658 40152 34671 40198
rect 33671 40123 34671 40152
rect 37896 40285 38556 40314
rect 37896 40239 37909 40285
rect 37955 40239 38026 40285
rect 38072 40239 38143 40285
rect 38189 40239 38261 40285
rect 38307 40239 38379 40285
rect 38425 40239 38497 40285
rect 38543 40239 38556 40285
rect 37896 40210 38556 40239
rect 43695 40397 43739 40443
rect 43785 40397 43906 40443
rect 43952 40397 44071 40443
rect 44117 40397 44236 40443
rect 44282 40397 44325 40443
rect 43695 40347 44325 40397
rect 50454 40457 51454 40503
rect 39598 40285 39730 40314
rect 39598 40239 39641 40285
rect 39687 40239 39730 40285
rect 39598 40226 39730 40239
rect 50454 40411 50516 40457
rect 50562 40411 50703 40457
rect 50749 40411 50890 40457
rect 50936 40411 51076 40457
rect 51122 40411 51263 40457
rect 51309 40411 51454 40457
rect 50454 40379 51454 40411
rect 43695 40123 44325 40227
rect 33671 39974 34671 40003
rect 37896 40061 38556 40090
rect 37896 40015 37909 40061
rect 37955 40015 38026 40061
rect 38072 40015 38143 40061
rect 38189 40015 38261 40061
rect 38307 40015 38379 40061
rect 38425 40015 38497 40061
rect 38543 40015 38556 40061
rect 37896 40002 38556 40015
rect 50454 40198 51454 40259
rect 50454 40152 50467 40198
rect 50513 40152 50571 40198
rect 50617 40152 50674 40198
rect 50720 40152 50777 40198
rect 50823 40152 50880 40198
rect 50926 40152 50983 40198
rect 51029 40152 51086 40198
rect 51132 40152 51189 40198
rect 51235 40152 51292 40198
rect 51338 40152 51395 40198
rect 51441 40152 51454 40198
rect 50454 40123 51454 40152
rect 33671 39928 33684 39974
rect 33730 39928 33787 39974
rect 33833 39928 33890 39974
rect 33936 39928 33993 39974
rect 34039 39928 34096 39974
rect 34142 39928 34199 39974
rect 34245 39928 34302 39974
rect 34348 39928 34405 39974
rect 34451 39928 34508 39974
rect 34554 39928 34612 39974
rect 34658 39928 34671 39974
rect 33671 39899 34671 39928
rect 39727 39974 40167 39987
rect 39727 39928 39740 39974
rect 39786 39928 39862 39974
rect 39908 39928 39985 39974
rect 40031 39928 40108 39974
rect 40154 39928 40167 39974
rect 39727 39899 40167 39928
rect 43695 39910 44325 40003
rect 50454 39974 51454 40003
rect 33671 39750 34671 39779
rect 33671 39704 33684 39750
rect 33730 39704 33787 39750
rect 33833 39704 33890 39750
rect 33936 39704 33993 39750
rect 34039 39704 34096 39750
rect 34142 39704 34199 39750
rect 34245 39704 34302 39750
rect 34348 39704 34405 39750
rect 34451 39704 34508 39750
rect 34554 39704 34612 39750
rect 34658 39704 34671 39750
rect 33671 39675 34671 39704
rect 39727 39750 40167 39779
rect 39727 39704 39740 39750
rect 39786 39704 39862 39750
rect 39908 39704 39985 39750
rect 40031 39704 40108 39750
rect 40154 39704 40167 39750
rect 39727 39675 40167 39704
rect 43695 39750 44325 39790
rect 50454 39928 50467 39974
rect 50513 39928 50571 39974
rect 50617 39928 50674 39974
rect 50720 39928 50777 39974
rect 50823 39928 50880 39974
rect 50926 39928 50983 39974
rect 51029 39928 51086 39974
rect 51132 39928 51189 39974
rect 51235 39928 51292 39974
rect 51338 39928 51395 39974
rect 51441 39928 51454 39974
rect 50454 39899 51454 39928
rect 43695 39704 43739 39750
rect 43785 39704 43906 39750
rect 43952 39704 44071 39750
rect 44117 39704 44236 39750
rect 44282 39704 44325 39750
rect 43695 39664 44325 39704
rect 33671 39526 34671 39555
rect 33671 39480 33684 39526
rect 33730 39480 33787 39526
rect 33833 39480 33890 39526
rect 33936 39480 33993 39526
rect 34039 39480 34096 39526
rect 34142 39480 34199 39526
rect 34245 39480 34302 39526
rect 34348 39480 34405 39526
rect 34451 39480 34508 39526
rect 34554 39480 34612 39526
rect 34658 39480 34671 39526
rect 33671 39451 34671 39480
rect 39727 39526 40167 39555
rect 39727 39480 39740 39526
rect 39786 39480 39862 39526
rect 39908 39480 39985 39526
rect 40031 39480 40108 39526
rect 40154 39480 40167 39526
rect 39727 39467 40167 39480
rect 50454 39750 51454 39779
rect 50454 39704 50467 39750
rect 50513 39704 50571 39750
rect 50617 39704 50674 39750
rect 50720 39704 50777 39750
rect 50823 39704 50880 39750
rect 50926 39704 50983 39750
rect 51029 39704 51086 39750
rect 51132 39704 51189 39750
rect 51235 39704 51292 39750
rect 51338 39704 51395 39750
rect 51441 39704 51454 39750
rect 50454 39675 51454 39704
rect 37896 39439 38556 39452
rect 43695 39451 44325 39544
rect 50454 39526 51454 39555
rect 50454 39480 50467 39526
rect 50513 39480 50571 39526
rect 50617 39480 50674 39526
rect 50720 39480 50777 39526
rect 50823 39480 50880 39526
rect 50926 39480 50983 39526
rect 51029 39480 51086 39526
rect 51132 39480 51189 39526
rect 51235 39480 51292 39526
rect 51338 39480 51395 39526
rect 51441 39480 51454 39526
rect 37896 39393 37909 39439
rect 37955 39393 38026 39439
rect 38072 39393 38143 39439
rect 38189 39393 38261 39439
rect 38307 39393 38379 39439
rect 38425 39393 38497 39439
rect 38543 39393 38556 39439
rect 37896 39364 38556 39393
rect 33671 39302 34671 39331
rect 33671 39256 33684 39302
rect 33730 39256 33787 39302
rect 33833 39256 33890 39302
rect 33936 39256 33993 39302
rect 34039 39256 34096 39302
rect 34142 39256 34199 39302
rect 34245 39256 34302 39302
rect 34348 39256 34405 39302
rect 34451 39256 34508 39302
rect 34554 39256 34612 39302
rect 34658 39256 34671 39302
rect 33671 39195 34671 39256
rect 33671 39043 34671 39075
rect 33671 38997 33816 39043
rect 33862 38997 34002 39043
rect 34048 38997 34189 39043
rect 34235 38997 34376 39043
rect 34422 38997 34562 39043
rect 34608 38997 34671 39043
rect 50454 39451 51454 39480
rect 37896 39215 38556 39244
rect 37896 39169 37909 39215
rect 37955 39169 38026 39215
rect 38072 39169 38143 39215
rect 38189 39169 38261 39215
rect 38307 39169 38379 39215
rect 38425 39169 38497 39215
rect 38543 39169 38556 39215
rect 37896 39140 38556 39169
rect 39598 39215 39730 39228
rect 43695 39227 44325 39331
rect 39598 39169 39641 39215
rect 39687 39169 39730 39215
rect 39598 39140 39730 39169
rect 50454 39302 51454 39331
rect 50454 39256 50467 39302
rect 50513 39256 50571 39302
rect 50617 39256 50674 39302
rect 50720 39256 50777 39302
rect 50823 39256 50880 39302
rect 50926 39256 50983 39302
rect 51029 39256 51086 39302
rect 51132 39256 51189 39302
rect 51235 39256 51292 39302
rect 51338 39256 51395 39302
rect 51441 39256 51454 39302
rect 50454 39195 51454 39256
rect 43695 39057 44325 39107
rect 33671 38951 34671 38997
rect 37896 38991 38556 39020
rect 37896 38945 37909 38991
rect 37955 38945 38026 38991
rect 38072 38945 38143 38991
rect 38189 38945 38261 38991
rect 38307 38945 38379 38991
rect 38425 38945 38497 38991
rect 38543 38945 38556 38991
rect 37896 38932 38556 38945
rect 39598 38991 39730 39020
rect 39598 38945 39641 38991
rect 39687 38945 39730 38991
rect 43695 39011 43739 39057
rect 43785 39011 43906 39057
rect 43952 39011 44071 39057
rect 44117 39011 44236 39057
rect 44282 39011 44325 39057
rect 50454 39043 51454 39075
rect 43695 38964 44325 39011
rect 39598 38932 39730 38945
rect 50454 38997 50516 39043
rect 50562 38997 50703 39043
rect 50749 38997 50890 39043
rect 50936 38997 51076 39043
rect 51122 38997 51263 39043
rect 51309 38997 51454 39043
rect 50454 38951 51454 38997
rect 33671 38657 34671 38703
rect 33671 38611 33816 38657
rect 33862 38611 34002 38657
rect 34048 38611 34189 38657
rect 34235 38611 34376 38657
rect 34422 38611 34562 38657
rect 34608 38611 34671 38657
rect 37896 38709 38556 38722
rect 37896 38663 37909 38709
rect 37955 38663 38026 38709
rect 38072 38663 38143 38709
rect 38189 38663 38261 38709
rect 38307 38663 38379 38709
rect 38425 38663 38497 38709
rect 38543 38663 38556 38709
rect 37896 38634 38556 38663
rect 39598 38709 39730 38722
rect 39598 38663 39641 38709
rect 39687 38663 39730 38709
rect 39598 38634 39730 38663
rect 43695 38643 44325 38690
rect 33671 38579 34671 38611
rect 33671 38398 34671 38459
rect 33671 38352 33684 38398
rect 33730 38352 33787 38398
rect 33833 38352 33890 38398
rect 33936 38352 33993 38398
rect 34039 38352 34096 38398
rect 34142 38352 34199 38398
rect 34245 38352 34302 38398
rect 34348 38352 34405 38398
rect 34451 38352 34508 38398
rect 34554 38352 34612 38398
rect 34658 38352 34671 38398
rect 33671 38323 34671 38352
rect 37896 38485 38556 38514
rect 37896 38439 37909 38485
rect 37955 38439 38026 38485
rect 38072 38439 38143 38485
rect 38189 38439 38261 38485
rect 38307 38439 38379 38485
rect 38425 38439 38497 38485
rect 38543 38439 38556 38485
rect 37896 38410 38556 38439
rect 43695 38597 43739 38643
rect 43785 38597 43906 38643
rect 43952 38597 44071 38643
rect 44117 38597 44236 38643
rect 44282 38597 44325 38643
rect 43695 38547 44325 38597
rect 50454 38657 51454 38703
rect 39598 38485 39730 38514
rect 39598 38439 39641 38485
rect 39687 38439 39730 38485
rect 39598 38426 39730 38439
rect 50454 38611 50516 38657
rect 50562 38611 50703 38657
rect 50749 38611 50890 38657
rect 50936 38611 51076 38657
rect 51122 38611 51263 38657
rect 51309 38611 51454 38657
rect 50454 38579 51454 38611
rect 43695 38323 44325 38427
rect 33671 38174 34671 38203
rect 37896 38261 38556 38290
rect 37896 38215 37909 38261
rect 37955 38215 38026 38261
rect 38072 38215 38143 38261
rect 38189 38215 38261 38261
rect 38307 38215 38379 38261
rect 38425 38215 38497 38261
rect 38543 38215 38556 38261
rect 37896 38202 38556 38215
rect 50454 38398 51454 38459
rect 50454 38352 50467 38398
rect 50513 38352 50571 38398
rect 50617 38352 50674 38398
rect 50720 38352 50777 38398
rect 50823 38352 50880 38398
rect 50926 38352 50983 38398
rect 51029 38352 51086 38398
rect 51132 38352 51189 38398
rect 51235 38352 51292 38398
rect 51338 38352 51395 38398
rect 51441 38352 51454 38398
rect 50454 38323 51454 38352
rect 33671 38128 33684 38174
rect 33730 38128 33787 38174
rect 33833 38128 33890 38174
rect 33936 38128 33993 38174
rect 34039 38128 34096 38174
rect 34142 38128 34199 38174
rect 34245 38128 34302 38174
rect 34348 38128 34405 38174
rect 34451 38128 34508 38174
rect 34554 38128 34612 38174
rect 34658 38128 34671 38174
rect 33671 38099 34671 38128
rect 39727 38174 40167 38187
rect 39727 38128 39740 38174
rect 39786 38128 39862 38174
rect 39908 38128 39985 38174
rect 40031 38128 40108 38174
rect 40154 38128 40167 38174
rect 39727 38099 40167 38128
rect 43695 38110 44325 38203
rect 50454 38174 51454 38203
rect 33671 37950 34671 37979
rect 33671 37904 33684 37950
rect 33730 37904 33787 37950
rect 33833 37904 33890 37950
rect 33936 37904 33993 37950
rect 34039 37904 34096 37950
rect 34142 37904 34199 37950
rect 34245 37904 34302 37950
rect 34348 37904 34405 37950
rect 34451 37904 34508 37950
rect 34554 37904 34612 37950
rect 34658 37904 34671 37950
rect 33671 37875 34671 37904
rect 39727 37950 40167 37979
rect 39727 37904 39740 37950
rect 39786 37904 39862 37950
rect 39908 37904 39985 37950
rect 40031 37904 40108 37950
rect 40154 37904 40167 37950
rect 39727 37875 40167 37904
rect 43695 37950 44325 37990
rect 50454 38128 50467 38174
rect 50513 38128 50571 38174
rect 50617 38128 50674 38174
rect 50720 38128 50777 38174
rect 50823 38128 50880 38174
rect 50926 38128 50983 38174
rect 51029 38128 51086 38174
rect 51132 38128 51189 38174
rect 51235 38128 51292 38174
rect 51338 38128 51395 38174
rect 51441 38128 51454 38174
rect 50454 38099 51454 38128
rect 43695 37904 43739 37950
rect 43785 37904 43906 37950
rect 43952 37904 44071 37950
rect 44117 37904 44236 37950
rect 44282 37904 44325 37950
rect 43695 37864 44325 37904
rect 33671 37726 34671 37755
rect 33671 37680 33684 37726
rect 33730 37680 33787 37726
rect 33833 37680 33890 37726
rect 33936 37680 33993 37726
rect 34039 37680 34096 37726
rect 34142 37680 34199 37726
rect 34245 37680 34302 37726
rect 34348 37680 34405 37726
rect 34451 37680 34508 37726
rect 34554 37680 34612 37726
rect 34658 37680 34671 37726
rect 33671 37651 34671 37680
rect 39727 37726 40167 37755
rect 39727 37680 39740 37726
rect 39786 37680 39862 37726
rect 39908 37680 39985 37726
rect 40031 37680 40108 37726
rect 40154 37680 40167 37726
rect 39727 37667 40167 37680
rect 50454 37950 51454 37979
rect 50454 37904 50467 37950
rect 50513 37904 50571 37950
rect 50617 37904 50674 37950
rect 50720 37904 50777 37950
rect 50823 37904 50880 37950
rect 50926 37904 50983 37950
rect 51029 37904 51086 37950
rect 51132 37904 51189 37950
rect 51235 37904 51292 37950
rect 51338 37904 51395 37950
rect 51441 37904 51454 37950
rect 50454 37875 51454 37904
rect 37896 37639 38556 37652
rect 43695 37651 44325 37744
rect 50454 37726 51454 37755
rect 50454 37680 50467 37726
rect 50513 37680 50571 37726
rect 50617 37680 50674 37726
rect 50720 37680 50777 37726
rect 50823 37680 50880 37726
rect 50926 37680 50983 37726
rect 51029 37680 51086 37726
rect 51132 37680 51189 37726
rect 51235 37680 51292 37726
rect 51338 37680 51395 37726
rect 51441 37680 51454 37726
rect 37896 37593 37909 37639
rect 37955 37593 38026 37639
rect 38072 37593 38143 37639
rect 38189 37593 38261 37639
rect 38307 37593 38379 37639
rect 38425 37593 38497 37639
rect 38543 37593 38556 37639
rect 37896 37564 38556 37593
rect 33671 37502 34671 37531
rect 33671 37456 33684 37502
rect 33730 37456 33787 37502
rect 33833 37456 33890 37502
rect 33936 37456 33993 37502
rect 34039 37456 34096 37502
rect 34142 37456 34199 37502
rect 34245 37456 34302 37502
rect 34348 37456 34405 37502
rect 34451 37456 34508 37502
rect 34554 37456 34612 37502
rect 34658 37456 34671 37502
rect 33671 37395 34671 37456
rect 33671 37243 34671 37275
rect 33671 37197 33816 37243
rect 33862 37197 34002 37243
rect 34048 37197 34189 37243
rect 34235 37197 34376 37243
rect 34422 37197 34562 37243
rect 34608 37197 34671 37243
rect 50454 37651 51454 37680
rect 37896 37415 38556 37444
rect 37896 37369 37909 37415
rect 37955 37369 38026 37415
rect 38072 37369 38143 37415
rect 38189 37369 38261 37415
rect 38307 37369 38379 37415
rect 38425 37369 38497 37415
rect 38543 37369 38556 37415
rect 37896 37340 38556 37369
rect 39598 37415 39730 37428
rect 43695 37427 44325 37531
rect 39598 37369 39641 37415
rect 39687 37369 39730 37415
rect 39598 37340 39730 37369
rect 50454 37502 51454 37531
rect 50454 37456 50467 37502
rect 50513 37456 50571 37502
rect 50617 37456 50674 37502
rect 50720 37456 50777 37502
rect 50823 37456 50880 37502
rect 50926 37456 50983 37502
rect 51029 37456 51086 37502
rect 51132 37456 51189 37502
rect 51235 37456 51292 37502
rect 51338 37456 51395 37502
rect 51441 37456 51454 37502
rect 50454 37395 51454 37456
rect 43695 37257 44325 37307
rect 33671 37151 34671 37197
rect 37896 37191 38556 37220
rect 37896 37145 37909 37191
rect 37955 37145 38026 37191
rect 38072 37145 38143 37191
rect 38189 37145 38261 37191
rect 38307 37145 38379 37191
rect 38425 37145 38497 37191
rect 38543 37145 38556 37191
rect 37896 37132 38556 37145
rect 39598 37191 39730 37220
rect 39598 37145 39641 37191
rect 39687 37145 39730 37191
rect 43695 37211 43739 37257
rect 43785 37211 43906 37257
rect 43952 37211 44071 37257
rect 44117 37211 44236 37257
rect 44282 37211 44325 37257
rect 50454 37243 51454 37275
rect 43695 37164 44325 37211
rect 39598 37132 39730 37145
rect 50454 37197 50516 37243
rect 50562 37197 50703 37243
rect 50749 37197 50890 37243
rect 50936 37197 51076 37243
rect 51122 37197 51263 37243
rect 51309 37197 51454 37243
rect 50454 37151 51454 37197
rect 33671 36857 34671 36903
rect 33671 36811 33816 36857
rect 33862 36811 34002 36857
rect 34048 36811 34189 36857
rect 34235 36811 34376 36857
rect 34422 36811 34562 36857
rect 34608 36811 34671 36857
rect 37896 36909 38556 36922
rect 37896 36863 37909 36909
rect 37955 36863 38026 36909
rect 38072 36863 38143 36909
rect 38189 36863 38261 36909
rect 38307 36863 38379 36909
rect 38425 36863 38497 36909
rect 38543 36863 38556 36909
rect 37896 36834 38556 36863
rect 39598 36909 39730 36922
rect 39598 36863 39641 36909
rect 39687 36863 39730 36909
rect 39598 36834 39730 36863
rect 43695 36843 44325 36890
rect 33671 36779 34671 36811
rect 33671 36598 34671 36659
rect 33671 36552 33684 36598
rect 33730 36552 33787 36598
rect 33833 36552 33890 36598
rect 33936 36552 33993 36598
rect 34039 36552 34096 36598
rect 34142 36552 34199 36598
rect 34245 36552 34302 36598
rect 34348 36552 34405 36598
rect 34451 36552 34508 36598
rect 34554 36552 34612 36598
rect 34658 36552 34671 36598
rect 33671 36523 34671 36552
rect 37896 36685 38556 36714
rect 37896 36639 37909 36685
rect 37955 36639 38026 36685
rect 38072 36639 38143 36685
rect 38189 36639 38261 36685
rect 38307 36639 38379 36685
rect 38425 36639 38497 36685
rect 38543 36639 38556 36685
rect 37896 36610 38556 36639
rect 43695 36797 43739 36843
rect 43785 36797 43906 36843
rect 43952 36797 44071 36843
rect 44117 36797 44236 36843
rect 44282 36797 44325 36843
rect 43695 36747 44325 36797
rect 50454 36857 51454 36903
rect 39598 36685 39730 36714
rect 39598 36639 39641 36685
rect 39687 36639 39730 36685
rect 39598 36626 39730 36639
rect 50454 36811 50516 36857
rect 50562 36811 50703 36857
rect 50749 36811 50890 36857
rect 50936 36811 51076 36857
rect 51122 36811 51263 36857
rect 51309 36811 51454 36857
rect 50454 36779 51454 36811
rect 43695 36523 44325 36627
rect 33671 36374 34671 36403
rect 37896 36461 38556 36490
rect 37896 36415 37909 36461
rect 37955 36415 38026 36461
rect 38072 36415 38143 36461
rect 38189 36415 38261 36461
rect 38307 36415 38379 36461
rect 38425 36415 38497 36461
rect 38543 36415 38556 36461
rect 37896 36402 38556 36415
rect 50454 36598 51454 36659
rect 50454 36552 50467 36598
rect 50513 36552 50571 36598
rect 50617 36552 50674 36598
rect 50720 36552 50777 36598
rect 50823 36552 50880 36598
rect 50926 36552 50983 36598
rect 51029 36552 51086 36598
rect 51132 36552 51189 36598
rect 51235 36552 51292 36598
rect 51338 36552 51395 36598
rect 51441 36552 51454 36598
rect 50454 36523 51454 36552
rect 33671 36328 33684 36374
rect 33730 36328 33787 36374
rect 33833 36328 33890 36374
rect 33936 36328 33993 36374
rect 34039 36328 34096 36374
rect 34142 36328 34199 36374
rect 34245 36328 34302 36374
rect 34348 36328 34405 36374
rect 34451 36328 34508 36374
rect 34554 36328 34612 36374
rect 34658 36328 34671 36374
rect 33671 36299 34671 36328
rect 39727 36374 40167 36387
rect 39727 36328 39740 36374
rect 39786 36328 39862 36374
rect 39908 36328 39985 36374
rect 40031 36328 40108 36374
rect 40154 36328 40167 36374
rect 39727 36299 40167 36328
rect 43695 36310 44325 36403
rect 50454 36374 51454 36403
rect 33671 36150 34671 36179
rect 33671 36104 33684 36150
rect 33730 36104 33787 36150
rect 33833 36104 33890 36150
rect 33936 36104 33993 36150
rect 34039 36104 34096 36150
rect 34142 36104 34199 36150
rect 34245 36104 34302 36150
rect 34348 36104 34405 36150
rect 34451 36104 34508 36150
rect 34554 36104 34612 36150
rect 34658 36104 34671 36150
rect 33671 36091 34671 36104
rect 39727 36150 40167 36179
rect 39727 36104 39740 36150
rect 39786 36104 39862 36150
rect 39908 36104 39985 36150
rect 40031 36104 40108 36150
rect 40154 36104 40167 36150
rect 39727 36091 40167 36104
rect 43695 36150 44325 36190
rect 50454 36328 50467 36374
rect 50513 36328 50571 36374
rect 50617 36328 50674 36374
rect 50720 36328 50777 36374
rect 50823 36328 50880 36374
rect 50926 36328 50983 36374
rect 51029 36328 51086 36374
rect 51132 36328 51189 36374
rect 51235 36328 51292 36374
rect 51338 36328 51395 36374
rect 51441 36328 51454 36374
rect 50454 36299 51454 36328
rect 43695 36104 43739 36150
rect 43785 36104 43906 36150
rect 43952 36104 44071 36150
rect 44117 36104 44236 36150
rect 44282 36104 44325 36150
rect 43695 36058 44325 36104
rect 50454 36150 51454 36179
rect 50454 36104 50467 36150
rect 50513 36104 50571 36150
rect 50617 36104 50674 36150
rect 50720 36104 50777 36150
rect 50823 36104 50880 36150
rect 50926 36104 50983 36150
rect 51029 36104 51086 36150
rect 51132 36104 51189 36150
rect 51235 36104 51292 36150
rect 51338 36104 51395 36150
rect 51441 36104 51454 36150
rect 50454 36091 51454 36104
<< mvpdiff >>
rect 29274 44250 30373 44296
rect 29274 44204 29317 44250
rect 29363 44204 29478 44250
rect 29524 44204 29638 44250
rect 29684 44204 29798 44250
rect 29844 44204 29959 44250
rect 30005 44204 30121 44250
rect 30167 44204 30284 44250
rect 30330 44204 30373 44250
rect 29274 44171 30373 44204
rect 35396 44218 37922 44231
rect 35396 44172 35409 44218
rect 37291 44172 37348 44218
rect 37394 44172 37451 44218
rect 37497 44172 37554 44218
rect 37600 44172 37657 44218
rect 37703 44172 37760 44218
rect 37806 44172 37863 44218
rect 37909 44172 37922 44218
rect 35396 44143 37922 44172
rect 35396 43994 37922 44023
rect 35396 43948 35409 43994
rect 37291 43948 37348 43994
rect 37394 43948 37451 43994
rect 37497 43948 37554 43994
rect 37600 43948 37657 43994
rect 37703 43948 37760 43994
rect 37806 43948 37863 43994
rect 37909 43948 37922 43994
rect 35396 43919 37922 43948
rect 38363 43994 39681 44007
rect 38363 43948 38376 43994
rect 38422 43948 38479 43994
rect 38525 43948 38582 43994
rect 38628 43948 38686 43994
rect 38732 43948 38790 43994
rect 38836 43948 38894 43994
rect 38940 43948 38998 43994
rect 39044 43948 39102 43994
rect 39148 43948 39206 43994
rect 39252 43948 39310 43994
rect 39356 43948 39414 43994
rect 39460 43948 39518 43994
rect 39564 43948 39622 43994
rect 39668 43948 39681 43994
rect 38363 43919 39681 43948
rect 42663 43994 43981 44007
rect 42663 43948 42676 43994
rect 42722 43948 42779 43994
rect 42825 43948 42882 43994
rect 42928 43948 42986 43994
rect 43032 43948 43090 43994
rect 43136 43948 43194 43994
rect 43240 43948 43298 43994
rect 43344 43948 43402 43994
rect 43448 43948 43506 43994
rect 43552 43948 43610 43994
rect 43656 43948 43714 43994
rect 43760 43948 43818 43994
rect 43864 43948 43922 43994
rect 43968 43948 43981 43994
rect 42663 43919 43981 43948
rect 47101 44218 49627 44231
rect 47101 44172 47114 44218
rect 48996 44172 49053 44218
rect 49099 44172 49156 44218
rect 49202 44172 49259 44218
rect 49305 44172 49362 44218
rect 49408 44172 49465 44218
rect 49511 44172 49568 44218
rect 49614 44172 49627 44218
rect 47101 44143 49627 44172
rect 35396 43770 37922 43799
rect 35396 43724 35409 43770
rect 37291 43724 37348 43770
rect 37394 43724 37451 43770
rect 37497 43724 37554 43770
rect 37600 43724 37657 43770
rect 37703 43724 37760 43770
rect 37806 43724 37863 43770
rect 37909 43724 37922 43770
rect 35396 43711 37922 43724
rect 38363 43770 39681 43799
rect 38363 43724 38376 43770
rect 38422 43724 38479 43770
rect 38525 43724 38582 43770
rect 38628 43724 38686 43770
rect 38732 43724 38790 43770
rect 38836 43724 38894 43770
rect 38940 43724 38998 43770
rect 39044 43724 39102 43770
rect 39148 43724 39206 43770
rect 39252 43724 39310 43770
rect 39356 43724 39414 43770
rect 39460 43724 39518 43770
rect 39564 43724 39622 43770
rect 39668 43724 39681 43770
rect 38363 43711 39681 43724
rect 45333 43994 46651 44007
rect 45333 43948 45346 43994
rect 45392 43948 45449 43994
rect 45495 43948 45552 43994
rect 45598 43948 45656 43994
rect 45702 43948 45760 43994
rect 45806 43948 45864 43994
rect 45910 43948 45968 43994
rect 46014 43948 46072 43994
rect 46118 43948 46176 43994
rect 46222 43948 46280 43994
rect 46326 43948 46384 43994
rect 46430 43948 46488 43994
rect 46534 43948 46592 43994
rect 46638 43948 46651 43994
rect 45333 43919 46651 43948
rect 47101 43994 49627 44023
rect 47101 43948 47114 43994
rect 48996 43948 49053 43994
rect 49099 43948 49156 43994
rect 49202 43948 49259 43994
rect 49305 43948 49362 43994
rect 49408 43948 49465 43994
rect 49511 43948 49568 43994
rect 49614 43948 49627 43994
rect 47101 43919 49627 43948
rect 54750 44250 55849 44296
rect 54750 44204 54793 44250
rect 54839 44204 54956 44250
rect 55002 44204 55118 44250
rect 55164 44204 55279 44250
rect 55325 44204 55439 44250
rect 55485 44204 55599 44250
rect 55645 44204 55760 44250
rect 55806 44204 55849 44250
rect 54750 44171 55849 44204
rect 42663 43770 43981 43799
rect 42663 43724 42676 43770
rect 42722 43724 42779 43770
rect 42825 43724 42882 43770
rect 42928 43724 42986 43770
rect 43032 43724 43090 43770
rect 43136 43724 43194 43770
rect 43240 43724 43298 43770
rect 43344 43724 43402 43770
rect 43448 43724 43506 43770
rect 43552 43724 43610 43770
rect 43656 43724 43714 43770
rect 43760 43724 43818 43770
rect 43864 43724 43922 43770
rect 43968 43724 43981 43770
rect 42663 43711 43981 43724
rect 45333 43770 46651 43799
rect 45333 43724 45346 43770
rect 45392 43724 45449 43770
rect 45495 43724 45552 43770
rect 45598 43724 45656 43770
rect 45702 43724 45760 43770
rect 45806 43724 45864 43770
rect 45910 43724 45968 43770
rect 46014 43724 46072 43770
rect 46118 43724 46176 43770
rect 46222 43724 46280 43770
rect 46326 43724 46384 43770
rect 46430 43724 46488 43770
rect 46534 43724 46592 43770
rect 46638 43724 46651 43770
rect 45333 43711 46651 43724
rect 47101 43770 49627 43799
rect 47101 43724 47114 43770
rect 48996 43724 49053 43770
rect 49099 43724 49156 43770
rect 49202 43724 49259 43770
rect 49305 43724 49362 43770
rect 49408 43724 49465 43770
rect 49511 43724 49568 43770
rect 49614 43724 49627 43770
rect 47101 43711 49627 43724
rect 29274 43350 30373 43383
rect 29274 43304 29317 43350
rect 29363 43304 29478 43350
rect 29524 43304 29638 43350
rect 29684 43304 29798 43350
rect 29844 43304 29959 43350
rect 30005 43304 30121 43350
rect 30167 43304 30284 43350
rect 30330 43304 30373 43350
rect 29274 43271 30373 43304
rect 31336 43350 33336 43363
rect 31336 43304 31349 43350
rect 33323 43304 33336 43350
rect 31336 43275 33336 43304
rect 31336 43126 33336 43155
rect 31336 43080 31349 43126
rect 33323 43080 33336 43126
rect 31336 43051 33336 43080
rect 31336 42902 33336 42931
rect 31336 42856 31349 42902
rect 33323 42856 33336 42902
rect 31336 42827 33336 42856
rect 44799 43350 45323 43363
rect 44799 43304 44812 43350
rect 44858 43304 44925 43350
rect 44971 43304 45038 43350
rect 45084 43304 45151 43350
rect 45197 43304 45264 43350
rect 45310 43304 45323 43350
rect 44799 43275 45323 43304
rect 51789 43350 53789 43363
rect 51789 43304 51802 43350
rect 53776 43304 53789 43350
rect 51789 43275 53789 43304
rect 35260 43039 36360 43052
rect 35260 42993 35273 43039
rect 35523 42993 35580 43039
rect 35626 42993 35683 43039
rect 35729 42993 35786 43039
rect 35832 42993 35889 43039
rect 35935 42993 35992 43039
rect 36038 42993 36095 43039
rect 36141 42993 36198 43039
rect 36244 42993 36301 43039
rect 36347 42993 36360 43039
rect 35260 42964 36360 42993
rect 36841 43039 37501 43052
rect 36841 42993 36854 43039
rect 36900 42993 36971 43039
rect 37017 42993 37088 43039
rect 37134 42993 37206 43039
rect 37252 42993 37324 43039
rect 37370 42993 37442 43039
rect 37488 42993 37501 43039
rect 36841 42964 37501 42993
rect 44799 43126 45323 43155
rect 44799 43080 44812 43126
rect 44858 43080 44925 43126
rect 44971 43080 45038 43126
rect 45084 43080 45151 43126
rect 45197 43080 45264 43126
rect 45310 43080 45323 43126
rect 54750 43350 55849 43383
rect 54750 43304 54793 43350
rect 54839 43304 54956 43350
rect 55002 43304 55118 43350
rect 55164 43304 55279 43350
rect 55325 43304 55439 43350
rect 55485 43304 55599 43350
rect 55645 43304 55760 43350
rect 55806 43304 55849 43350
rect 54750 43271 55849 43304
rect 44799 43051 45323 43080
rect 31336 42678 33336 42707
rect 31336 42632 31349 42678
rect 33323 42632 33336 42678
rect 35260 42815 36360 42844
rect 35260 42769 35273 42815
rect 35523 42769 35580 42815
rect 35626 42769 35683 42815
rect 35729 42769 35786 42815
rect 35832 42769 35889 42815
rect 35935 42769 35992 42815
rect 36038 42769 36095 42815
rect 36141 42769 36198 42815
rect 36244 42769 36301 42815
rect 36347 42769 36360 42815
rect 35260 42740 36360 42769
rect 31336 42619 33336 42632
rect 48765 43039 49865 43052
rect 48765 42993 48778 43039
rect 48824 42993 48881 43039
rect 48927 42993 48984 43039
rect 49030 42993 49087 43039
rect 49133 42993 49190 43039
rect 49236 42993 49293 43039
rect 49339 42993 49396 43039
rect 49442 42993 49499 43039
rect 49545 42993 49602 43039
rect 49852 42993 49865 43039
rect 48765 42964 49865 42993
rect 36841 42815 37501 42844
rect 36841 42769 36854 42815
rect 36900 42769 36971 42815
rect 37017 42769 37088 42815
rect 37134 42769 37206 42815
rect 37252 42769 37324 42815
rect 37370 42769 37442 42815
rect 37488 42769 37501 42815
rect 36841 42740 37501 42769
rect 39008 42815 39326 42828
rect 39008 42769 39021 42815
rect 39067 42769 39144 42815
rect 39190 42769 39267 42815
rect 39313 42769 39326 42815
rect 39008 42740 39326 42769
rect 44799 42902 45323 42931
rect 44799 42856 44812 42902
rect 44858 42856 44925 42902
rect 44971 42856 45038 42902
rect 45084 42856 45151 42902
rect 45197 42856 45264 42902
rect 45310 42856 45323 42902
rect 44799 42827 45323 42856
rect 48765 42815 49865 42844
rect 48765 42769 48778 42815
rect 48824 42769 48881 42815
rect 48927 42769 48984 42815
rect 49030 42769 49087 42815
rect 49133 42769 49190 42815
rect 49236 42769 49293 42815
rect 49339 42769 49396 42815
rect 49442 42769 49499 42815
rect 49545 42769 49602 42815
rect 49852 42769 49865 42815
rect 48765 42740 49865 42769
rect 35260 42591 36360 42620
rect 35260 42545 35273 42591
rect 35523 42545 35580 42591
rect 35626 42545 35683 42591
rect 35729 42545 35786 42591
rect 35832 42545 35889 42591
rect 35935 42545 35992 42591
rect 36038 42545 36095 42591
rect 36141 42545 36198 42591
rect 36244 42545 36301 42591
rect 36347 42545 36360 42591
rect 35260 42532 36360 42545
rect 36841 42591 37501 42620
rect 36841 42545 36854 42591
rect 36900 42545 36971 42591
rect 37017 42545 37088 42591
rect 37134 42545 37206 42591
rect 37252 42545 37324 42591
rect 37370 42545 37442 42591
rect 37488 42545 37501 42591
rect 36841 42532 37501 42545
rect 39008 42591 39326 42620
rect 39008 42545 39021 42591
rect 39067 42545 39144 42591
rect 39190 42545 39267 42591
rect 39313 42545 39326 42591
rect 39008 42532 39326 42545
rect 44799 42678 45323 42707
rect 44799 42632 44812 42678
rect 44858 42632 44925 42678
rect 44971 42632 45038 42678
rect 45084 42632 45151 42678
rect 45197 42632 45264 42678
rect 45310 42632 45323 42678
rect 44799 42619 45323 42632
rect 51789 43126 53789 43155
rect 51789 43080 51802 43126
rect 53776 43080 53789 43126
rect 51789 43051 53789 43080
rect 51789 42902 53789 42931
rect 51789 42856 51802 42902
rect 53776 42856 53789 42902
rect 51789 42827 53789 42856
rect 51789 42678 53789 42707
rect 48765 42591 49865 42620
rect 48765 42545 48778 42591
rect 48824 42545 48881 42591
rect 48927 42545 48984 42591
rect 49030 42545 49087 42591
rect 49133 42545 49190 42591
rect 49236 42545 49293 42591
rect 49339 42545 49396 42591
rect 49442 42545 49499 42591
rect 49545 42545 49602 42591
rect 49852 42545 49865 42591
rect 51789 42632 51802 42678
rect 53776 42632 53789 42678
rect 51789 42619 53789 42632
rect 48765 42532 49865 42545
rect 29274 42450 30373 42483
rect 29274 42404 29317 42450
rect 29363 42404 29478 42450
rect 29524 42404 29638 42450
rect 29684 42404 29798 42450
rect 29844 42404 29959 42450
rect 30005 42404 30121 42450
rect 30167 42404 30284 42450
rect 30330 42404 30373 42450
rect 29274 42371 30373 42404
rect 54750 42450 55849 42483
rect 54750 42404 54793 42450
rect 54839 42404 54956 42450
rect 55002 42404 55118 42450
rect 55164 42404 55279 42450
rect 55325 42404 55439 42450
rect 55485 42404 55599 42450
rect 55645 42404 55760 42450
rect 55806 42404 55849 42450
rect 54750 42371 55849 42404
rect 35260 42309 36360 42322
rect 31336 42222 33336 42235
rect 31336 42176 31349 42222
rect 33323 42176 33336 42222
rect 35260 42263 35273 42309
rect 35523 42263 35580 42309
rect 35626 42263 35683 42309
rect 35729 42263 35786 42309
rect 35832 42263 35889 42309
rect 35935 42263 35992 42309
rect 36038 42263 36095 42309
rect 36141 42263 36198 42309
rect 36244 42263 36301 42309
rect 36347 42263 36360 42309
rect 35260 42234 36360 42263
rect 36841 42309 37501 42322
rect 36841 42263 36854 42309
rect 36900 42263 36971 42309
rect 37017 42263 37088 42309
rect 37134 42263 37206 42309
rect 37252 42263 37324 42309
rect 37370 42263 37442 42309
rect 37488 42263 37501 42309
rect 36841 42234 37501 42263
rect 39008 42309 39326 42322
rect 39008 42263 39021 42309
rect 39067 42263 39144 42309
rect 39190 42263 39267 42309
rect 39313 42263 39326 42309
rect 39008 42234 39326 42263
rect 48765 42309 49865 42322
rect 31336 42147 33336 42176
rect 31336 41998 33336 42027
rect 31336 41952 31349 41998
rect 33323 41952 33336 41998
rect 31336 41923 33336 41952
rect 31336 41774 33336 41803
rect 31336 41728 31349 41774
rect 33323 41728 33336 41774
rect 31336 41699 33336 41728
rect 29274 41550 30373 41583
rect 29274 41504 29317 41550
rect 29363 41504 29478 41550
rect 29524 41504 29638 41550
rect 29684 41504 29798 41550
rect 29844 41504 29959 41550
rect 30005 41504 30121 41550
rect 30167 41504 30284 41550
rect 30330 41504 30373 41550
rect 29274 41471 30373 41504
rect 35260 42085 36360 42114
rect 35260 42039 35273 42085
rect 35523 42039 35580 42085
rect 35626 42039 35683 42085
rect 35729 42039 35786 42085
rect 35832 42039 35889 42085
rect 35935 42039 35992 42085
rect 36038 42039 36095 42085
rect 36141 42039 36198 42085
rect 36244 42039 36301 42085
rect 36347 42039 36360 42085
rect 35260 42010 36360 42039
rect 36841 42085 37501 42114
rect 36841 42039 36854 42085
rect 36900 42039 36971 42085
rect 37017 42039 37088 42085
rect 37134 42039 37206 42085
rect 37252 42039 37324 42085
rect 37370 42039 37442 42085
rect 37488 42039 37501 42085
rect 36841 42010 37501 42039
rect 48765 42263 48778 42309
rect 48824 42263 48881 42309
rect 48927 42263 48984 42309
rect 49030 42263 49087 42309
rect 49133 42263 49190 42309
rect 49236 42263 49293 42309
rect 49339 42263 49396 42309
rect 49442 42263 49499 42309
rect 49545 42263 49602 42309
rect 49852 42263 49865 42309
rect 44799 42222 45323 42235
rect 48765 42234 49865 42263
rect 44799 42176 44812 42222
rect 44858 42176 44925 42222
rect 44971 42176 45038 42222
rect 45084 42176 45151 42222
rect 45197 42176 45264 42222
rect 45310 42176 45323 42222
rect 44799 42147 45323 42176
rect 39008 42085 39326 42114
rect 39008 42039 39021 42085
rect 39067 42039 39144 42085
rect 39190 42039 39267 42085
rect 39313 42039 39326 42085
rect 39008 42026 39326 42039
rect 51789 42222 53789 42235
rect 44799 41998 45323 42027
rect 44799 41952 44812 41998
rect 44858 41952 44925 41998
rect 44971 41952 45038 41998
rect 45084 41952 45151 41998
rect 45197 41952 45264 41998
rect 45310 41952 45323 41998
rect 44799 41923 45323 41952
rect 48765 42085 49865 42114
rect 48765 42039 48778 42085
rect 48824 42039 48881 42085
rect 48927 42039 48984 42085
rect 49030 42039 49087 42085
rect 49133 42039 49190 42085
rect 49236 42039 49293 42085
rect 49339 42039 49396 42085
rect 49442 42039 49499 42085
rect 49545 42039 49602 42085
rect 49852 42039 49865 42085
rect 48765 42010 49865 42039
rect 51789 42176 51802 42222
rect 53776 42176 53789 42222
rect 51789 42147 53789 42176
rect 35260 41861 36360 41890
rect 35260 41815 35273 41861
rect 35523 41815 35580 41861
rect 35626 41815 35683 41861
rect 35729 41815 35786 41861
rect 35832 41815 35889 41861
rect 35935 41815 35992 41861
rect 36038 41815 36095 41861
rect 36141 41815 36198 41861
rect 36244 41815 36301 41861
rect 36347 41815 36360 41861
rect 35260 41802 36360 41815
rect 36841 41861 37501 41890
rect 36841 41815 36854 41861
rect 36900 41815 36971 41861
rect 37017 41815 37088 41861
rect 37134 41815 37206 41861
rect 37252 41815 37324 41861
rect 37370 41815 37442 41861
rect 37488 41815 37501 41861
rect 36841 41802 37501 41815
rect 48765 41861 49865 41890
rect 48765 41815 48778 41861
rect 48824 41815 48881 41861
rect 48927 41815 48984 41861
rect 49030 41815 49087 41861
rect 49133 41815 49190 41861
rect 49236 41815 49293 41861
rect 49339 41815 49396 41861
rect 49442 41815 49499 41861
rect 49545 41815 49602 41861
rect 49852 41815 49865 41861
rect 44799 41774 45323 41803
rect 48765 41802 49865 41815
rect 44799 41728 44812 41774
rect 44858 41728 44925 41774
rect 44971 41728 45038 41774
rect 45084 41728 45151 41774
rect 45197 41728 45264 41774
rect 45310 41728 45323 41774
rect 31336 41550 33336 41579
rect 31336 41504 31349 41550
rect 33323 41504 33336 41550
rect 31336 41475 33336 41504
rect 31336 41326 33336 41355
rect 31336 41280 31349 41326
rect 33323 41280 33336 41326
rect 31336 41251 33336 41280
rect 31336 41102 33336 41131
rect 31336 41056 31349 41102
rect 33323 41056 33336 41102
rect 31336 41027 33336 41056
rect 44799 41699 45323 41728
rect 51789 41998 53789 42027
rect 51789 41952 51802 41998
rect 53776 41952 53789 41998
rect 51789 41923 53789 41952
rect 51789 41774 53789 41803
rect 51789 41728 51802 41774
rect 53776 41728 53789 41774
rect 51789 41699 53789 41728
rect 44799 41550 45323 41579
rect 44799 41504 44812 41550
rect 44858 41504 44925 41550
rect 44971 41504 45038 41550
rect 45084 41504 45151 41550
rect 45197 41504 45264 41550
rect 45310 41504 45323 41550
rect 44799 41475 45323 41504
rect 51789 41550 53789 41579
rect 51789 41504 51802 41550
rect 53776 41504 53789 41550
rect 51789 41475 53789 41504
rect 35260 41239 36360 41252
rect 35260 41193 35273 41239
rect 35523 41193 35580 41239
rect 35626 41193 35683 41239
rect 35729 41193 35786 41239
rect 35832 41193 35889 41239
rect 35935 41193 35992 41239
rect 36038 41193 36095 41239
rect 36141 41193 36198 41239
rect 36244 41193 36301 41239
rect 36347 41193 36360 41239
rect 35260 41164 36360 41193
rect 36841 41239 37501 41252
rect 36841 41193 36854 41239
rect 36900 41193 36971 41239
rect 37017 41193 37088 41239
rect 37134 41193 37206 41239
rect 37252 41193 37324 41239
rect 37370 41193 37442 41239
rect 37488 41193 37501 41239
rect 36841 41164 37501 41193
rect 44799 41326 45323 41355
rect 44799 41280 44812 41326
rect 44858 41280 44925 41326
rect 44971 41280 45038 41326
rect 45084 41280 45151 41326
rect 45197 41280 45264 41326
rect 45310 41280 45323 41326
rect 54750 41550 55849 41583
rect 54750 41504 54793 41550
rect 54839 41504 54956 41550
rect 55002 41504 55118 41550
rect 55164 41504 55279 41550
rect 55325 41504 55439 41550
rect 55485 41504 55599 41550
rect 55645 41504 55760 41550
rect 55806 41504 55849 41550
rect 54750 41471 55849 41504
rect 44799 41251 45323 41280
rect 31336 40878 33336 40907
rect 31336 40832 31349 40878
rect 33323 40832 33336 40878
rect 35260 41015 36360 41044
rect 35260 40969 35273 41015
rect 35523 40969 35580 41015
rect 35626 40969 35683 41015
rect 35729 40969 35786 41015
rect 35832 40969 35889 41015
rect 35935 40969 35992 41015
rect 36038 40969 36095 41015
rect 36141 40969 36198 41015
rect 36244 40969 36301 41015
rect 36347 40969 36360 41015
rect 35260 40940 36360 40969
rect 31336 40819 33336 40832
rect 48765 41239 49865 41252
rect 48765 41193 48778 41239
rect 48824 41193 48881 41239
rect 48927 41193 48984 41239
rect 49030 41193 49087 41239
rect 49133 41193 49190 41239
rect 49236 41193 49293 41239
rect 49339 41193 49396 41239
rect 49442 41193 49499 41239
rect 49545 41193 49602 41239
rect 49852 41193 49865 41239
rect 48765 41164 49865 41193
rect 36841 41015 37501 41044
rect 36841 40969 36854 41015
rect 36900 40969 36971 41015
rect 37017 40969 37088 41015
rect 37134 40969 37206 41015
rect 37252 40969 37324 41015
rect 37370 40969 37442 41015
rect 37488 40969 37501 41015
rect 36841 40940 37501 40969
rect 39008 41015 39326 41028
rect 39008 40969 39021 41015
rect 39067 40969 39144 41015
rect 39190 40969 39267 41015
rect 39313 40969 39326 41015
rect 39008 40940 39326 40969
rect 44799 41102 45323 41131
rect 44799 41056 44812 41102
rect 44858 41056 44925 41102
rect 44971 41056 45038 41102
rect 45084 41056 45151 41102
rect 45197 41056 45264 41102
rect 45310 41056 45323 41102
rect 44799 41027 45323 41056
rect 48765 41015 49865 41044
rect 48765 40969 48778 41015
rect 48824 40969 48881 41015
rect 48927 40969 48984 41015
rect 49030 40969 49087 41015
rect 49133 40969 49190 41015
rect 49236 40969 49293 41015
rect 49339 40969 49396 41015
rect 49442 40969 49499 41015
rect 49545 40969 49602 41015
rect 49852 40969 49865 41015
rect 48765 40940 49865 40969
rect 35260 40791 36360 40820
rect 35260 40745 35273 40791
rect 35523 40745 35580 40791
rect 35626 40745 35683 40791
rect 35729 40745 35786 40791
rect 35832 40745 35889 40791
rect 35935 40745 35992 40791
rect 36038 40745 36095 40791
rect 36141 40745 36198 40791
rect 36244 40745 36301 40791
rect 36347 40745 36360 40791
rect 35260 40732 36360 40745
rect 36841 40791 37501 40820
rect 36841 40745 36854 40791
rect 36900 40745 36971 40791
rect 37017 40745 37088 40791
rect 37134 40745 37206 40791
rect 37252 40745 37324 40791
rect 37370 40745 37442 40791
rect 37488 40745 37501 40791
rect 36841 40732 37501 40745
rect 39008 40791 39326 40820
rect 39008 40745 39021 40791
rect 39067 40745 39144 40791
rect 39190 40745 39267 40791
rect 39313 40745 39326 40791
rect 39008 40732 39326 40745
rect 44799 40878 45323 40907
rect 44799 40832 44812 40878
rect 44858 40832 44925 40878
rect 44971 40832 45038 40878
rect 45084 40832 45151 40878
rect 45197 40832 45264 40878
rect 45310 40832 45323 40878
rect 44799 40819 45323 40832
rect 51789 41326 53789 41355
rect 51789 41280 51802 41326
rect 53776 41280 53789 41326
rect 51789 41251 53789 41280
rect 51789 41102 53789 41131
rect 51789 41056 51802 41102
rect 53776 41056 53789 41102
rect 51789 41027 53789 41056
rect 51789 40878 53789 40907
rect 48765 40791 49865 40820
rect 48765 40745 48778 40791
rect 48824 40745 48881 40791
rect 48927 40745 48984 40791
rect 49030 40745 49087 40791
rect 49133 40745 49190 40791
rect 49236 40745 49293 40791
rect 49339 40745 49396 40791
rect 49442 40745 49499 40791
rect 49545 40745 49602 40791
rect 49852 40745 49865 40791
rect 51789 40832 51802 40878
rect 53776 40832 53789 40878
rect 51789 40819 53789 40832
rect 48765 40732 49865 40745
rect 29274 40650 30373 40683
rect 29274 40604 29317 40650
rect 29363 40604 29478 40650
rect 29524 40604 29638 40650
rect 29684 40604 29798 40650
rect 29844 40604 29959 40650
rect 30005 40604 30121 40650
rect 30167 40604 30284 40650
rect 30330 40604 30373 40650
rect 29274 40571 30373 40604
rect 54750 40650 55849 40683
rect 54750 40604 54793 40650
rect 54839 40604 54956 40650
rect 55002 40604 55118 40650
rect 55164 40604 55279 40650
rect 55325 40604 55439 40650
rect 55485 40604 55599 40650
rect 55645 40604 55760 40650
rect 55806 40604 55849 40650
rect 54750 40571 55849 40604
rect 35260 40509 36360 40522
rect 31336 40422 33336 40435
rect 31336 40376 31349 40422
rect 33323 40376 33336 40422
rect 35260 40463 35273 40509
rect 35523 40463 35580 40509
rect 35626 40463 35683 40509
rect 35729 40463 35786 40509
rect 35832 40463 35889 40509
rect 35935 40463 35992 40509
rect 36038 40463 36095 40509
rect 36141 40463 36198 40509
rect 36244 40463 36301 40509
rect 36347 40463 36360 40509
rect 35260 40434 36360 40463
rect 36841 40509 37501 40522
rect 36841 40463 36854 40509
rect 36900 40463 36971 40509
rect 37017 40463 37088 40509
rect 37134 40463 37206 40509
rect 37252 40463 37324 40509
rect 37370 40463 37442 40509
rect 37488 40463 37501 40509
rect 36841 40434 37501 40463
rect 39008 40509 39326 40522
rect 39008 40463 39021 40509
rect 39067 40463 39144 40509
rect 39190 40463 39267 40509
rect 39313 40463 39326 40509
rect 39008 40434 39326 40463
rect 48765 40509 49865 40522
rect 31336 40347 33336 40376
rect 31336 40198 33336 40227
rect 31336 40152 31349 40198
rect 33323 40152 33336 40198
rect 31336 40123 33336 40152
rect 31336 39974 33336 40003
rect 31336 39928 31349 39974
rect 33323 39928 33336 39974
rect 31336 39899 33336 39928
rect 29274 39750 30373 39783
rect 29274 39704 29317 39750
rect 29363 39704 29478 39750
rect 29524 39704 29638 39750
rect 29684 39704 29798 39750
rect 29844 39704 29959 39750
rect 30005 39704 30121 39750
rect 30167 39704 30284 39750
rect 30330 39704 30373 39750
rect 29274 39671 30373 39704
rect 35260 40285 36360 40314
rect 35260 40239 35273 40285
rect 35523 40239 35580 40285
rect 35626 40239 35683 40285
rect 35729 40239 35786 40285
rect 35832 40239 35889 40285
rect 35935 40239 35992 40285
rect 36038 40239 36095 40285
rect 36141 40239 36198 40285
rect 36244 40239 36301 40285
rect 36347 40239 36360 40285
rect 35260 40210 36360 40239
rect 36841 40285 37501 40314
rect 36841 40239 36854 40285
rect 36900 40239 36971 40285
rect 37017 40239 37088 40285
rect 37134 40239 37206 40285
rect 37252 40239 37324 40285
rect 37370 40239 37442 40285
rect 37488 40239 37501 40285
rect 36841 40210 37501 40239
rect 48765 40463 48778 40509
rect 48824 40463 48881 40509
rect 48927 40463 48984 40509
rect 49030 40463 49087 40509
rect 49133 40463 49190 40509
rect 49236 40463 49293 40509
rect 49339 40463 49396 40509
rect 49442 40463 49499 40509
rect 49545 40463 49602 40509
rect 49852 40463 49865 40509
rect 44799 40422 45323 40435
rect 48765 40434 49865 40463
rect 44799 40376 44812 40422
rect 44858 40376 44925 40422
rect 44971 40376 45038 40422
rect 45084 40376 45151 40422
rect 45197 40376 45264 40422
rect 45310 40376 45323 40422
rect 44799 40347 45323 40376
rect 39008 40285 39326 40314
rect 39008 40239 39021 40285
rect 39067 40239 39144 40285
rect 39190 40239 39267 40285
rect 39313 40239 39326 40285
rect 39008 40226 39326 40239
rect 51789 40422 53789 40435
rect 44799 40198 45323 40227
rect 44799 40152 44812 40198
rect 44858 40152 44925 40198
rect 44971 40152 45038 40198
rect 45084 40152 45151 40198
rect 45197 40152 45264 40198
rect 45310 40152 45323 40198
rect 44799 40123 45323 40152
rect 48765 40285 49865 40314
rect 48765 40239 48778 40285
rect 48824 40239 48881 40285
rect 48927 40239 48984 40285
rect 49030 40239 49087 40285
rect 49133 40239 49190 40285
rect 49236 40239 49293 40285
rect 49339 40239 49396 40285
rect 49442 40239 49499 40285
rect 49545 40239 49602 40285
rect 49852 40239 49865 40285
rect 48765 40210 49865 40239
rect 51789 40376 51802 40422
rect 53776 40376 53789 40422
rect 51789 40347 53789 40376
rect 35260 40061 36360 40090
rect 35260 40015 35273 40061
rect 35523 40015 35580 40061
rect 35626 40015 35683 40061
rect 35729 40015 35786 40061
rect 35832 40015 35889 40061
rect 35935 40015 35992 40061
rect 36038 40015 36095 40061
rect 36141 40015 36198 40061
rect 36244 40015 36301 40061
rect 36347 40015 36360 40061
rect 35260 40002 36360 40015
rect 36841 40061 37501 40090
rect 36841 40015 36854 40061
rect 36900 40015 36971 40061
rect 37017 40015 37088 40061
rect 37134 40015 37206 40061
rect 37252 40015 37324 40061
rect 37370 40015 37442 40061
rect 37488 40015 37501 40061
rect 36841 40002 37501 40015
rect 48765 40061 49865 40090
rect 48765 40015 48778 40061
rect 48824 40015 48881 40061
rect 48927 40015 48984 40061
rect 49030 40015 49087 40061
rect 49133 40015 49190 40061
rect 49236 40015 49293 40061
rect 49339 40015 49396 40061
rect 49442 40015 49499 40061
rect 49545 40015 49602 40061
rect 49852 40015 49865 40061
rect 44799 39974 45323 40003
rect 48765 40002 49865 40015
rect 44799 39928 44812 39974
rect 44858 39928 44925 39974
rect 44971 39928 45038 39974
rect 45084 39928 45151 39974
rect 45197 39928 45264 39974
rect 45310 39928 45323 39974
rect 31336 39750 33336 39779
rect 31336 39704 31349 39750
rect 33323 39704 33336 39750
rect 31336 39675 33336 39704
rect 31336 39526 33336 39555
rect 31336 39480 31349 39526
rect 33323 39480 33336 39526
rect 31336 39451 33336 39480
rect 31336 39302 33336 39331
rect 31336 39256 31349 39302
rect 33323 39256 33336 39302
rect 31336 39227 33336 39256
rect 44799 39899 45323 39928
rect 51789 40198 53789 40227
rect 51789 40152 51802 40198
rect 53776 40152 53789 40198
rect 51789 40123 53789 40152
rect 51789 39974 53789 40003
rect 51789 39928 51802 39974
rect 53776 39928 53789 39974
rect 51789 39899 53789 39928
rect 44799 39750 45323 39779
rect 44799 39704 44812 39750
rect 44858 39704 44925 39750
rect 44971 39704 45038 39750
rect 45084 39704 45151 39750
rect 45197 39704 45264 39750
rect 45310 39704 45323 39750
rect 44799 39675 45323 39704
rect 51789 39750 53789 39779
rect 51789 39704 51802 39750
rect 53776 39704 53789 39750
rect 51789 39675 53789 39704
rect 35260 39439 36360 39452
rect 35260 39393 35273 39439
rect 35523 39393 35580 39439
rect 35626 39393 35683 39439
rect 35729 39393 35786 39439
rect 35832 39393 35889 39439
rect 35935 39393 35992 39439
rect 36038 39393 36095 39439
rect 36141 39393 36198 39439
rect 36244 39393 36301 39439
rect 36347 39393 36360 39439
rect 35260 39364 36360 39393
rect 36841 39439 37501 39452
rect 36841 39393 36854 39439
rect 36900 39393 36971 39439
rect 37017 39393 37088 39439
rect 37134 39393 37206 39439
rect 37252 39393 37324 39439
rect 37370 39393 37442 39439
rect 37488 39393 37501 39439
rect 36841 39364 37501 39393
rect 44799 39526 45323 39555
rect 44799 39480 44812 39526
rect 44858 39480 44925 39526
rect 44971 39480 45038 39526
rect 45084 39480 45151 39526
rect 45197 39480 45264 39526
rect 45310 39480 45323 39526
rect 54750 39750 55849 39783
rect 54750 39704 54793 39750
rect 54839 39704 54956 39750
rect 55002 39704 55118 39750
rect 55164 39704 55279 39750
rect 55325 39704 55439 39750
rect 55485 39704 55599 39750
rect 55645 39704 55760 39750
rect 55806 39704 55849 39750
rect 54750 39671 55849 39704
rect 44799 39451 45323 39480
rect 31336 39078 33336 39107
rect 31336 39032 31349 39078
rect 33323 39032 33336 39078
rect 35260 39215 36360 39244
rect 35260 39169 35273 39215
rect 35523 39169 35580 39215
rect 35626 39169 35683 39215
rect 35729 39169 35786 39215
rect 35832 39169 35889 39215
rect 35935 39169 35992 39215
rect 36038 39169 36095 39215
rect 36141 39169 36198 39215
rect 36244 39169 36301 39215
rect 36347 39169 36360 39215
rect 35260 39140 36360 39169
rect 31336 39019 33336 39032
rect 48765 39439 49865 39452
rect 48765 39393 48778 39439
rect 48824 39393 48881 39439
rect 48927 39393 48984 39439
rect 49030 39393 49087 39439
rect 49133 39393 49190 39439
rect 49236 39393 49293 39439
rect 49339 39393 49396 39439
rect 49442 39393 49499 39439
rect 49545 39393 49602 39439
rect 49852 39393 49865 39439
rect 48765 39364 49865 39393
rect 36841 39215 37501 39244
rect 36841 39169 36854 39215
rect 36900 39169 36971 39215
rect 37017 39169 37088 39215
rect 37134 39169 37206 39215
rect 37252 39169 37324 39215
rect 37370 39169 37442 39215
rect 37488 39169 37501 39215
rect 36841 39140 37501 39169
rect 39008 39215 39326 39228
rect 39008 39169 39021 39215
rect 39067 39169 39144 39215
rect 39190 39169 39267 39215
rect 39313 39169 39326 39215
rect 39008 39140 39326 39169
rect 44799 39302 45323 39331
rect 44799 39256 44812 39302
rect 44858 39256 44925 39302
rect 44971 39256 45038 39302
rect 45084 39256 45151 39302
rect 45197 39256 45264 39302
rect 45310 39256 45323 39302
rect 44799 39227 45323 39256
rect 48765 39215 49865 39244
rect 48765 39169 48778 39215
rect 48824 39169 48881 39215
rect 48927 39169 48984 39215
rect 49030 39169 49087 39215
rect 49133 39169 49190 39215
rect 49236 39169 49293 39215
rect 49339 39169 49396 39215
rect 49442 39169 49499 39215
rect 49545 39169 49602 39215
rect 49852 39169 49865 39215
rect 48765 39140 49865 39169
rect 35260 38991 36360 39020
rect 35260 38945 35273 38991
rect 35523 38945 35580 38991
rect 35626 38945 35683 38991
rect 35729 38945 35786 38991
rect 35832 38945 35889 38991
rect 35935 38945 35992 38991
rect 36038 38945 36095 38991
rect 36141 38945 36198 38991
rect 36244 38945 36301 38991
rect 36347 38945 36360 38991
rect 35260 38932 36360 38945
rect 36841 38991 37501 39020
rect 36841 38945 36854 38991
rect 36900 38945 36971 38991
rect 37017 38945 37088 38991
rect 37134 38945 37206 38991
rect 37252 38945 37324 38991
rect 37370 38945 37442 38991
rect 37488 38945 37501 38991
rect 36841 38932 37501 38945
rect 39008 38991 39326 39020
rect 39008 38945 39021 38991
rect 39067 38945 39144 38991
rect 39190 38945 39267 38991
rect 39313 38945 39326 38991
rect 39008 38932 39326 38945
rect 44799 39078 45323 39107
rect 44799 39032 44812 39078
rect 44858 39032 44925 39078
rect 44971 39032 45038 39078
rect 45084 39032 45151 39078
rect 45197 39032 45264 39078
rect 45310 39032 45323 39078
rect 44799 39019 45323 39032
rect 51789 39526 53789 39555
rect 51789 39480 51802 39526
rect 53776 39480 53789 39526
rect 51789 39451 53789 39480
rect 51789 39302 53789 39331
rect 51789 39256 51802 39302
rect 53776 39256 53789 39302
rect 51789 39227 53789 39256
rect 51789 39078 53789 39107
rect 48765 38991 49865 39020
rect 48765 38945 48778 38991
rect 48824 38945 48881 38991
rect 48927 38945 48984 38991
rect 49030 38945 49087 38991
rect 49133 38945 49190 38991
rect 49236 38945 49293 38991
rect 49339 38945 49396 38991
rect 49442 38945 49499 38991
rect 49545 38945 49602 38991
rect 49852 38945 49865 38991
rect 51789 39032 51802 39078
rect 53776 39032 53789 39078
rect 51789 39019 53789 39032
rect 48765 38932 49865 38945
rect 29274 38850 30373 38883
rect 29274 38804 29317 38850
rect 29363 38804 29478 38850
rect 29524 38804 29638 38850
rect 29684 38804 29798 38850
rect 29844 38804 29959 38850
rect 30005 38804 30121 38850
rect 30167 38804 30284 38850
rect 30330 38804 30373 38850
rect 29274 38771 30373 38804
rect 54750 38850 55849 38883
rect 54750 38804 54793 38850
rect 54839 38804 54956 38850
rect 55002 38804 55118 38850
rect 55164 38804 55279 38850
rect 55325 38804 55439 38850
rect 55485 38804 55599 38850
rect 55645 38804 55760 38850
rect 55806 38804 55849 38850
rect 54750 38771 55849 38804
rect 35260 38709 36360 38722
rect 31336 38622 33336 38635
rect 31336 38576 31349 38622
rect 33323 38576 33336 38622
rect 35260 38663 35273 38709
rect 35523 38663 35580 38709
rect 35626 38663 35683 38709
rect 35729 38663 35786 38709
rect 35832 38663 35889 38709
rect 35935 38663 35992 38709
rect 36038 38663 36095 38709
rect 36141 38663 36198 38709
rect 36244 38663 36301 38709
rect 36347 38663 36360 38709
rect 35260 38634 36360 38663
rect 36841 38709 37501 38722
rect 36841 38663 36854 38709
rect 36900 38663 36971 38709
rect 37017 38663 37088 38709
rect 37134 38663 37206 38709
rect 37252 38663 37324 38709
rect 37370 38663 37442 38709
rect 37488 38663 37501 38709
rect 36841 38634 37501 38663
rect 39008 38709 39326 38722
rect 39008 38663 39021 38709
rect 39067 38663 39144 38709
rect 39190 38663 39267 38709
rect 39313 38663 39326 38709
rect 39008 38634 39326 38663
rect 48765 38709 49865 38722
rect 31336 38547 33336 38576
rect 31336 38398 33336 38427
rect 31336 38352 31349 38398
rect 33323 38352 33336 38398
rect 31336 38323 33336 38352
rect 31336 38174 33336 38203
rect 31336 38128 31349 38174
rect 33323 38128 33336 38174
rect 31336 38099 33336 38128
rect 29274 37950 30373 37983
rect 29274 37904 29317 37950
rect 29363 37904 29478 37950
rect 29524 37904 29638 37950
rect 29684 37904 29798 37950
rect 29844 37904 29959 37950
rect 30005 37904 30121 37950
rect 30167 37904 30284 37950
rect 30330 37904 30373 37950
rect 29274 37871 30373 37904
rect 35260 38485 36360 38514
rect 35260 38439 35273 38485
rect 35523 38439 35580 38485
rect 35626 38439 35683 38485
rect 35729 38439 35786 38485
rect 35832 38439 35889 38485
rect 35935 38439 35992 38485
rect 36038 38439 36095 38485
rect 36141 38439 36198 38485
rect 36244 38439 36301 38485
rect 36347 38439 36360 38485
rect 35260 38410 36360 38439
rect 36841 38485 37501 38514
rect 36841 38439 36854 38485
rect 36900 38439 36971 38485
rect 37017 38439 37088 38485
rect 37134 38439 37206 38485
rect 37252 38439 37324 38485
rect 37370 38439 37442 38485
rect 37488 38439 37501 38485
rect 36841 38410 37501 38439
rect 48765 38663 48778 38709
rect 48824 38663 48881 38709
rect 48927 38663 48984 38709
rect 49030 38663 49087 38709
rect 49133 38663 49190 38709
rect 49236 38663 49293 38709
rect 49339 38663 49396 38709
rect 49442 38663 49499 38709
rect 49545 38663 49602 38709
rect 49852 38663 49865 38709
rect 44799 38622 45323 38635
rect 48765 38634 49865 38663
rect 44799 38576 44812 38622
rect 44858 38576 44925 38622
rect 44971 38576 45038 38622
rect 45084 38576 45151 38622
rect 45197 38576 45264 38622
rect 45310 38576 45323 38622
rect 44799 38547 45323 38576
rect 39008 38485 39326 38514
rect 39008 38439 39021 38485
rect 39067 38439 39144 38485
rect 39190 38439 39267 38485
rect 39313 38439 39326 38485
rect 39008 38426 39326 38439
rect 51789 38622 53789 38635
rect 44799 38398 45323 38427
rect 44799 38352 44812 38398
rect 44858 38352 44925 38398
rect 44971 38352 45038 38398
rect 45084 38352 45151 38398
rect 45197 38352 45264 38398
rect 45310 38352 45323 38398
rect 44799 38323 45323 38352
rect 48765 38485 49865 38514
rect 48765 38439 48778 38485
rect 48824 38439 48881 38485
rect 48927 38439 48984 38485
rect 49030 38439 49087 38485
rect 49133 38439 49190 38485
rect 49236 38439 49293 38485
rect 49339 38439 49396 38485
rect 49442 38439 49499 38485
rect 49545 38439 49602 38485
rect 49852 38439 49865 38485
rect 48765 38410 49865 38439
rect 51789 38576 51802 38622
rect 53776 38576 53789 38622
rect 51789 38547 53789 38576
rect 35260 38261 36360 38290
rect 35260 38215 35273 38261
rect 35523 38215 35580 38261
rect 35626 38215 35683 38261
rect 35729 38215 35786 38261
rect 35832 38215 35889 38261
rect 35935 38215 35992 38261
rect 36038 38215 36095 38261
rect 36141 38215 36198 38261
rect 36244 38215 36301 38261
rect 36347 38215 36360 38261
rect 35260 38202 36360 38215
rect 36841 38261 37501 38290
rect 36841 38215 36854 38261
rect 36900 38215 36971 38261
rect 37017 38215 37088 38261
rect 37134 38215 37206 38261
rect 37252 38215 37324 38261
rect 37370 38215 37442 38261
rect 37488 38215 37501 38261
rect 36841 38202 37501 38215
rect 48765 38261 49865 38290
rect 48765 38215 48778 38261
rect 48824 38215 48881 38261
rect 48927 38215 48984 38261
rect 49030 38215 49087 38261
rect 49133 38215 49190 38261
rect 49236 38215 49293 38261
rect 49339 38215 49396 38261
rect 49442 38215 49499 38261
rect 49545 38215 49602 38261
rect 49852 38215 49865 38261
rect 44799 38174 45323 38203
rect 48765 38202 49865 38215
rect 44799 38128 44812 38174
rect 44858 38128 44925 38174
rect 44971 38128 45038 38174
rect 45084 38128 45151 38174
rect 45197 38128 45264 38174
rect 45310 38128 45323 38174
rect 31336 37950 33336 37979
rect 31336 37904 31349 37950
rect 33323 37904 33336 37950
rect 31336 37875 33336 37904
rect 31336 37726 33336 37755
rect 31336 37680 31349 37726
rect 33323 37680 33336 37726
rect 31336 37651 33336 37680
rect 31336 37502 33336 37531
rect 31336 37456 31349 37502
rect 33323 37456 33336 37502
rect 31336 37427 33336 37456
rect 44799 38099 45323 38128
rect 51789 38398 53789 38427
rect 51789 38352 51802 38398
rect 53776 38352 53789 38398
rect 51789 38323 53789 38352
rect 51789 38174 53789 38203
rect 51789 38128 51802 38174
rect 53776 38128 53789 38174
rect 51789 38099 53789 38128
rect 44799 37950 45323 37979
rect 44799 37904 44812 37950
rect 44858 37904 44925 37950
rect 44971 37904 45038 37950
rect 45084 37904 45151 37950
rect 45197 37904 45264 37950
rect 45310 37904 45323 37950
rect 44799 37875 45323 37904
rect 51789 37950 53789 37979
rect 51789 37904 51802 37950
rect 53776 37904 53789 37950
rect 51789 37875 53789 37904
rect 35260 37639 36360 37652
rect 35260 37593 35273 37639
rect 35523 37593 35580 37639
rect 35626 37593 35683 37639
rect 35729 37593 35786 37639
rect 35832 37593 35889 37639
rect 35935 37593 35992 37639
rect 36038 37593 36095 37639
rect 36141 37593 36198 37639
rect 36244 37593 36301 37639
rect 36347 37593 36360 37639
rect 35260 37564 36360 37593
rect 36841 37639 37501 37652
rect 36841 37593 36854 37639
rect 36900 37593 36971 37639
rect 37017 37593 37088 37639
rect 37134 37593 37206 37639
rect 37252 37593 37324 37639
rect 37370 37593 37442 37639
rect 37488 37593 37501 37639
rect 36841 37564 37501 37593
rect 44799 37726 45323 37755
rect 44799 37680 44812 37726
rect 44858 37680 44925 37726
rect 44971 37680 45038 37726
rect 45084 37680 45151 37726
rect 45197 37680 45264 37726
rect 45310 37680 45323 37726
rect 54750 37950 55849 37983
rect 54750 37904 54793 37950
rect 54839 37904 54956 37950
rect 55002 37904 55118 37950
rect 55164 37904 55279 37950
rect 55325 37904 55439 37950
rect 55485 37904 55599 37950
rect 55645 37904 55760 37950
rect 55806 37904 55849 37950
rect 54750 37871 55849 37904
rect 44799 37651 45323 37680
rect 31336 37278 33336 37307
rect 31336 37232 31349 37278
rect 33323 37232 33336 37278
rect 35260 37415 36360 37444
rect 35260 37369 35273 37415
rect 35523 37369 35580 37415
rect 35626 37369 35683 37415
rect 35729 37369 35786 37415
rect 35832 37369 35889 37415
rect 35935 37369 35992 37415
rect 36038 37369 36095 37415
rect 36141 37369 36198 37415
rect 36244 37369 36301 37415
rect 36347 37369 36360 37415
rect 35260 37340 36360 37369
rect 31336 37219 33336 37232
rect 48765 37639 49865 37652
rect 48765 37593 48778 37639
rect 48824 37593 48881 37639
rect 48927 37593 48984 37639
rect 49030 37593 49087 37639
rect 49133 37593 49190 37639
rect 49236 37593 49293 37639
rect 49339 37593 49396 37639
rect 49442 37593 49499 37639
rect 49545 37593 49602 37639
rect 49852 37593 49865 37639
rect 48765 37564 49865 37593
rect 36841 37415 37501 37444
rect 36841 37369 36854 37415
rect 36900 37369 36971 37415
rect 37017 37369 37088 37415
rect 37134 37369 37206 37415
rect 37252 37369 37324 37415
rect 37370 37369 37442 37415
rect 37488 37369 37501 37415
rect 36841 37340 37501 37369
rect 39008 37415 39326 37428
rect 39008 37369 39021 37415
rect 39067 37369 39144 37415
rect 39190 37369 39267 37415
rect 39313 37369 39326 37415
rect 39008 37340 39326 37369
rect 44799 37502 45323 37531
rect 44799 37456 44812 37502
rect 44858 37456 44925 37502
rect 44971 37456 45038 37502
rect 45084 37456 45151 37502
rect 45197 37456 45264 37502
rect 45310 37456 45323 37502
rect 44799 37427 45323 37456
rect 48765 37415 49865 37444
rect 48765 37369 48778 37415
rect 48824 37369 48881 37415
rect 48927 37369 48984 37415
rect 49030 37369 49087 37415
rect 49133 37369 49190 37415
rect 49236 37369 49293 37415
rect 49339 37369 49396 37415
rect 49442 37369 49499 37415
rect 49545 37369 49602 37415
rect 49852 37369 49865 37415
rect 48765 37340 49865 37369
rect 35260 37191 36360 37220
rect 35260 37145 35273 37191
rect 35523 37145 35580 37191
rect 35626 37145 35683 37191
rect 35729 37145 35786 37191
rect 35832 37145 35889 37191
rect 35935 37145 35992 37191
rect 36038 37145 36095 37191
rect 36141 37145 36198 37191
rect 36244 37145 36301 37191
rect 36347 37145 36360 37191
rect 35260 37132 36360 37145
rect 36841 37191 37501 37220
rect 36841 37145 36854 37191
rect 36900 37145 36971 37191
rect 37017 37145 37088 37191
rect 37134 37145 37206 37191
rect 37252 37145 37324 37191
rect 37370 37145 37442 37191
rect 37488 37145 37501 37191
rect 36841 37132 37501 37145
rect 39008 37191 39326 37220
rect 39008 37145 39021 37191
rect 39067 37145 39144 37191
rect 39190 37145 39267 37191
rect 39313 37145 39326 37191
rect 39008 37132 39326 37145
rect 44799 37278 45323 37307
rect 44799 37232 44812 37278
rect 44858 37232 44925 37278
rect 44971 37232 45038 37278
rect 45084 37232 45151 37278
rect 45197 37232 45264 37278
rect 45310 37232 45323 37278
rect 44799 37219 45323 37232
rect 51789 37726 53789 37755
rect 51789 37680 51802 37726
rect 53776 37680 53789 37726
rect 51789 37651 53789 37680
rect 51789 37502 53789 37531
rect 51789 37456 51802 37502
rect 53776 37456 53789 37502
rect 51789 37427 53789 37456
rect 51789 37278 53789 37307
rect 48765 37191 49865 37220
rect 48765 37145 48778 37191
rect 48824 37145 48881 37191
rect 48927 37145 48984 37191
rect 49030 37145 49087 37191
rect 49133 37145 49190 37191
rect 49236 37145 49293 37191
rect 49339 37145 49396 37191
rect 49442 37145 49499 37191
rect 49545 37145 49602 37191
rect 49852 37145 49865 37191
rect 51789 37232 51802 37278
rect 53776 37232 53789 37278
rect 51789 37219 53789 37232
rect 48765 37132 49865 37145
rect 29274 37050 30373 37083
rect 29274 37004 29317 37050
rect 29363 37004 29478 37050
rect 29524 37004 29638 37050
rect 29684 37004 29798 37050
rect 29844 37004 29959 37050
rect 30005 37004 30121 37050
rect 30167 37004 30284 37050
rect 30330 37004 30373 37050
rect 29274 36971 30373 37004
rect 54750 37050 55849 37083
rect 54750 37004 54793 37050
rect 54839 37004 54956 37050
rect 55002 37004 55118 37050
rect 55164 37004 55279 37050
rect 55325 37004 55439 37050
rect 55485 37004 55599 37050
rect 55645 37004 55760 37050
rect 55806 37004 55849 37050
rect 54750 36971 55849 37004
rect 35260 36909 36360 36922
rect 31336 36822 33336 36835
rect 31336 36776 31349 36822
rect 33323 36776 33336 36822
rect 35260 36863 35273 36909
rect 35523 36863 35580 36909
rect 35626 36863 35683 36909
rect 35729 36863 35786 36909
rect 35832 36863 35889 36909
rect 35935 36863 35992 36909
rect 36038 36863 36095 36909
rect 36141 36863 36198 36909
rect 36244 36863 36301 36909
rect 36347 36863 36360 36909
rect 35260 36834 36360 36863
rect 36841 36909 37501 36922
rect 36841 36863 36854 36909
rect 36900 36863 36971 36909
rect 37017 36863 37088 36909
rect 37134 36863 37206 36909
rect 37252 36863 37324 36909
rect 37370 36863 37442 36909
rect 37488 36863 37501 36909
rect 36841 36834 37501 36863
rect 39008 36909 39326 36922
rect 39008 36863 39021 36909
rect 39067 36863 39144 36909
rect 39190 36863 39267 36909
rect 39313 36863 39326 36909
rect 39008 36834 39326 36863
rect 48765 36909 49865 36922
rect 31336 36747 33336 36776
rect 31336 36598 33336 36627
rect 31336 36552 31349 36598
rect 33323 36552 33336 36598
rect 31336 36523 33336 36552
rect 31336 36374 33336 36403
rect 31336 36328 31349 36374
rect 33323 36328 33336 36374
rect 31336 36299 33336 36328
rect 29274 36150 30373 36183
rect 29274 36104 29317 36150
rect 29363 36104 29478 36150
rect 29524 36104 29638 36150
rect 29684 36104 29798 36150
rect 29844 36104 29959 36150
rect 30005 36104 30121 36150
rect 30167 36104 30284 36150
rect 30330 36104 30373 36150
rect 29274 36058 30373 36104
rect 35260 36685 36360 36714
rect 35260 36639 35273 36685
rect 35523 36639 35580 36685
rect 35626 36639 35683 36685
rect 35729 36639 35786 36685
rect 35832 36639 35889 36685
rect 35935 36639 35992 36685
rect 36038 36639 36095 36685
rect 36141 36639 36198 36685
rect 36244 36639 36301 36685
rect 36347 36639 36360 36685
rect 35260 36610 36360 36639
rect 36841 36685 37501 36714
rect 36841 36639 36854 36685
rect 36900 36639 36971 36685
rect 37017 36639 37088 36685
rect 37134 36639 37206 36685
rect 37252 36639 37324 36685
rect 37370 36639 37442 36685
rect 37488 36639 37501 36685
rect 36841 36610 37501 36639
rect 48765 36863 48778 36909
rect 48824 36863 48881 36909
rect 48927 36863 48984 36909
rect 49030 36863 49087 36909
rect 49133 36863 49190 36909
rect 49236 36863 49293 36909
rect 49339 36863 49396 36909
rect 49442 36863 49499 36909
rect 49545 36863 49602 36909
rect 49852 36863 49865 36909
rect 44799 36822 45323 36835
rect 48765 36834 49865 36863
rect 44799 36776 44812 36822
rect 44858 36776 44925 36822
rect 44971 36776 45038 36822
rect 45084 36776 45151 36822
rect 45197 36776 45264 36822
rect 45310 36776 45323 36822
rect 44799 36747 45323 36776
rect 39008 36685 39326 36714
rect 39008 36639 39021 36685
rect 39067 36639 39144 36685
rect 39190 36639 39267 36685
rect 39313 36639 39326 36685
rect 39008 36626 39326 36639
rect 51789 36822 53789 36835
rect 44799 36598 45323 36627
rect 44799 36552 44812 36598
rect 44858 36552 44925 36598
rect 44971 36552 45038 36598
rect 45084 36552 45151 36598
rect 45197 36552 45264 36598
rect 45310 36552 45323 36598
rect 44799 36523 45323 36552
rect 48765 36685 49865 36714
rect 48765 36639 48778 36685
rect 48824 36639 48881 36685
rect 48927 36639 48984 36685
rect 49030 36639 49087 36685
rect 49133 36639 49190 36685
rect 49236 36639 49293 36685
rect 49339 36639 49396 36685
rect 49442 36639 49499 36685
rect 49545 36639 49602 36685
rect 49852 36639 49865 36685
rect 48765 36610 49865 36639
rect 51789 36776 51802 36822
rect 53776 36776 53789 36822
rect 51789 36747 53789 36776
rect 35260 36461 36360 36490
rect 35260 36415 35273 36461
rect 35523 36415 35580 36461
rect 35626 36415 35683 36461
rect 35729 36415 35786 36461
rect 35832 36415 35889 36461
rect 35935 36415 35992 36461
rect 36038 36415 36095 36461
rect 36141 36415 36198 36461
rect 36244 36415 36301 36461
rect 36347 36415 36360 36461
rect 35260 36402 36360 36415
rect 36841 36461 37501 36490
rect 36841 36415 36854 36461
rect 36900 36415 36971 36461
rect 37017 36415 37088 36461
rect 37134 36415 37206 36461
rect 37252 36415 37324 36461
rect 37370 36415 37442 36461
rect 37488 36415 37501 36461
rect 36841 36402 37501 36415
rect 48765 36461 49865 36490
rect 48765 36415 48778 36461
rect 48824 36415 48881 36461
rect 48927 36415 48984 36461
rect 49030 36415 49087 36461
rect 49133 36415 49190 36461
rect 49236 36415 49293 36461
rect 49339 36415 49396 36461
rect 49442 36415 49499 36461
rect 49545 36415 49602 36461
rect 49852 36415 49865 36461
rect 44799 36374 45323 36403
rect 48765 36402 49865 36415
rect 44799 36328 44812 36374
rect 44858 36328 44925 36374
rect 44971 36328 45038 36374
rect 45084 36328 45151 36374
rect 45197 36328 45264 36374
rect 45310 36328 45323 36374
rect 31336 36150 33336 36179
rect 31336 36104 31349 36150
rect 33323 36104 33336 36150
rect 31336 36091 33336 36104
rect 44799 36299 45323 36328
rect 51789 36598 53789 36627
rect 51789 36552 51802 36598
rect 53776 36552 53789 36598
rect 51789 36523 53789 36552
rect 51789 36374 53789 36403
rect 51789 36328 51802 36374
rect 53776 36328 53789 36374
rect 51789 36299 53789 36328
rect 44799 36150 45323 36179
rect 44799 36104 44812 36150
rect 44858 36104 44925 36150
rect 44971 36104 45038 36150
rect 45084 36104 45151 36150
rect 45197 36104 45264 36150
rect 45310 36104 45323 36150
rect 44799 36091 45323 36104
rect 51789 36150 53789 36179
rect 51789 36104 51802 36150
rect 53776 36104 53789 36150
rect 51789 36091 53789 36104
rect 54750 36150 55849 36183
rect 54750 36104 54793 36150
rect 54839 36104 54956 36150
rect 55002 36104 55118 36150
rect 55164 36104 55279 36150
rect 55325 36104 55439 36150
rect 55485 36104 55599 36150
rect 55645 36104 55760 36150
rect 55806 36104 55849 36150
rect 54750 36058 55849 36104
<< mvndiffc >>
rect 33014 43948 33774 43994
rect 33831 43948 33877 43994
rect 33934 43948 33980 43994
rect 34037 43948 34083 43994
rect 34140 43948 34186 43994
rect 34243 43948 34289 43994
rect 34346 43948 34392 43994
rect 34449 43948 34495 43994
rect 34552 43948 34598 43994
rect 34655 43948 34701 43994
rect 34758 43948 34804 43994
rect 34861 43948 34907 43994
rect 34964 43948 35010 43994
rect 40075 43948 40121 43994
rect 40189 43948 40235 43994
rect 40303 43948 40349 43994
rect 40417 43948 40463 43994
rect 40531 43948 40577 43994
rect 40976 43949 41022 43995
rect 41079 43949 41125 43995
rect 41182 43949 41228 43995
rect 41286 43949 41332 43995
rect 41390 43949 41436 43995
rect 41494 43949 41540 43995
rect 41598 43949 41644 43995
rect 41702 43949 41748 43995
rect 41806 43949 41852 43995
rect 41910 43949 41956 43995
rect 42014 43949 42060 43995
rect 42118 43949 42164 43995
rect 42222 43949 42268 43995
rect 33014 43724 33774 43770
rect 33831 43724 33877 43770
rect 33934 43724 33980 43770
rect 34037 43724 34083 43770
rect 34140 43724 34186 43770
rect 34243 43724 34289 43770
rect 34346 43724 34392 43770
rect 34449 43724 34495 43770
rect 34552 43724 34598 43770
rect 34655 43724 34701 43770
rect 34758 43724 34804 43770
rect 34861 43724 34907 43770
rect 34964 43724 35010 43770
rect 40075 43724 40121 43770
rect 40189 43724 40235 43770
rect 40303 43724 40349 43770
rect 40417 43724 40463 43770
rect 40531 43724 40577 43770
rect 44445 43948 44491 43994
rect 44559 43948 44605 43994
rect 44673 43948 44719 43994
rect 44787 43948 44833 43994
rect 44901 43948 44947 43994
rect 50014 43948 50774 43994
rect 50831 43948 50877 43994
rect 50934 43948 50980 43994
rect 51037 43948 51083 43994
rect 51140 43948 51186 43994
rect 51243 43948 51289 43994
rect 51346 43948 51392 43994
rect 51449 43948 51495 43994
rect 51552 43948 51598 43994
rect 51655 43948 51701 43994
rect 51758 43948 51804 43994
rect 51861 43948 51907 43994
rect 51964 43948 52010 43994
rect 40976 43725 41022 43771
rect 41079 43725 41125 43771
rect 41182 43725 41228 43771
rect 41286 43725 41332 43771
rect 41390 43725 41436 43771
rect 41494 43725 41540 43771
rect 41598 43725 41644 43771
rect 41702 43725 41748 43771
rect 41806 43725 41852 43771
rect 41910 43725 41956 43771
rect 42014 43725 42060 43771
rect 42118 43725 42164 43771
rect 42222 43725 42268 43771
rect 44445 43724 44491 43770
rect 44559 43724 44605 43770
rect 44673 43724 44719 43770
rect 44787 43724 44833 43770
rect 44901 43724 44947 43770
rect 50014 43724 50774 43770
rect 50831 43724 50877 43770
rect 50934 43724 50980 43770
rect 51037 43724 51083 43770
rect 51140 43724 51186 43770
rect 51243 43724 51289 43770
rect 51346 43724 51392 43770
rect 51449 43724 51495 43770
rect 51552 43724 51598 43770
rect 51655 43724 51701 43770
rect 51758 43724 51804 43770
rect 51861 43724 51907 43770
rect 51964 43724 52010 43770
rect 33684 43304 33730 43350
rect 33787 43304 33833 43350
rect 33890 43304 33936 43350
rect 33993 43304 34039 43350
rect 34096 43304 34142 43350
rect 34199 43304 34245 43350
rect 34302 43304 34348 43350
rect 34405 43304 34451 43350
rect 34508 43304 34554 43350
rect 34612 43304 34658 43350
rect 39740 43304 39786 43350
rect 39862 43304 39908 43350
rect 39985 43304 40031 43350
rect 40108 43304 40154 43350
rect 43739 43304 43785 43350
rect 43906 43304 43952 43350
rect 44071 43304 44117 43350
rect 44236 43304 44282 43350
rect 33684 43080 33730 43126
rect 33787 43080 33833 43126
rect 33890 43080 33936 43126
rect 33993 43080 34039 43126
rect 34096 43080 34142 43126
rect 34199 43080 34245 43126
rect 34302 43080 34348 43126
rect 34405 43080 34451 43126
rect 34508 43080 34554 43126
rect 34612 43080 34658 43126
rect 39740 43080 39786 43126
rect 39862 43080 39908 43126
rect 39985 43080 40031 43126
rect 40108 43080 40154 43126
rect 50467 43304 50513 43350
rect 50571 43304 50617 43350
rect 50674 43304 50720 43350
rect 50777 43304 50823 43350
rect 50880 43304 50926 43350
rect 50983 43304 51029 43350
rect 51086 43304 51132 43350
rect 51189 43304 51235 43350
rect 51292 43304 51338 43350
rect 51395 43304 51441 43350
rect 50467 43080 50513 43126
rect 50571 43080 50617 43126
rect 50674 43080 50720 43126
rect 50777 43080 50823 43126
rect 50880 43080 50926 43126
rect 50983 43080 51029 43126
rect 51086 43080 51132 43126
rect 51189 43080 51235 43126
rect 51292 43080 51338 43126
rect 51395 43080 51441 43126
rect 37909 42993 37955 43039
rect 38026 42993 38072 43039
rect 38143 42993 38189 43039
rect 38261 42993 38307 43039
rect 38379 42993 38425 43039
rect 38497 42993 38543 43039
rect 33684 42856 33730 42902
rect 33787 42856 33833 42902
rect 33890 42856 33936 42902
rect 33993 42856 34039 42902
rect 34096 42856 34142 42902
rect 34199 42856 34245 42902
rect 34302 42856 34348 42902
rect 34405 42856 34451 42902
rect 34508 42856 34554 42902
rect 34612 42856 34658 42902
rect 33816 42597 33862 42643
rect 34002 42597 34048 42643
rect 34189 42597 34235 42643
rect 34376 42597 34422 42643
rect 34562 42597 34608 42643
rect 37909 42769 37955 42815
rect 38026 42769 38072 42815
rect 38143 42769 38189 42815
rect 38261 42769 38307 42815
rect 38379 42769 38425 42815
rect 38497 42769 38543 42815
rect 39641 42769 39687 42815
rect 50467 42856 50513 42902
rect 50571 42856 50617 42902
rect 50674 42856 50720 42902
rect 50777 42856 50823 42902
rect 50880 42856 50926 42902
rect 50983 42856 51029 42902
rect 51086 42856 51132 42902
rect 51189 42856 51235 42902
rect 51292 42856 51338 42902
rect 51395 42856 51441 42902
rect 37909 42545 37955 42591
rect 38026 42545 38072 42591
rect 38143 42545 38189 42591
rect 38261 42545 38307 42591
rect 38379 42545 38425 42591
rect 38497 42545 38543 42591
rect 39641 42545 39687 42591
rect 43739 42611 43785 42657
rect 43906 42611 43952 42657
rect 44071 42611 44117 42657
rect 44236 42611 44282 42657
rect 50516 42597 50562 42643
rect 50703 42597 50749 42643
rect 50890 42597 50936 42643
rect 51076 42597 51122 42643
rect 51263 42597 51309 42643
rect 33816 42211 33862 42257
rect 34002 42211 34048 42257
rect 34189 42211 34235 42257
rect 34376 42211 34422 42257
rect 34562 42211 34608 42257
rect 37909 42263 37955 42309
rect 38026 42263 38072 42309
rect 38143 42263 38189 42309
rect 38261 42263 38307 42309
rect 38379 42263 38425 42309
rect 38497 42263 38543 42309
rect 39641 42263 39687 42309
rect 33684 41952 33730 41998
rect 33787 41952 33833 41998
rect 33890 41952 33936 41998
rect 33993 41952 34039 41998
rect 34096 41952 34142 41998
rect 34199 41952 34245 41998
rect 34302 41952 34348 41998
rect 34405 41952 34451 41998
rect 34508 41952 34554 41998
rect 34612 41952 34658 41998
rect 37909 42039 37955 42085
rect 38026 42039 38072 42085
rect 38143 42039 38189 42085
rect 38261 42039 38307 42085
rect 38379 42039 38425 42085
rect 38497 42039 38543 42085
rect 43739 42197 43785 42243
rect 43906 42197 43952 42243
rect 44071 42197 44117 42243
rect 44236 42197 44282 42243
rect 39641 42039 39687 42085
rect 50516 42211 50562 42257
rect 50703 42211 50749 42257
rect 50890 42211 50936 42257
rect 51076 42211 51122 42257
rect 51263 42211 51309 42257
rect 37909 41815 37955 41861
rect 38026 41815 38072 41861
rect 38143 41815 38189 41861
rect 38261 41815 38307 41861
rect 38379 41815 38425 41861
rect 38497 41815 38543 41861
rect 50467 41952 50513 41998
rect 50571 41952 50617 41998
rect 50674 41952 50720 41998
rect 50777 41952 50823 41998
rect 50880 41952 50926 41998
rect 50983 41952 51029 41998
rect 51086 41952 51132 41998
rect 51189 41952 51235 41998
rect 51292 41952 51338 41998
rect 51395 41952 51441 41998
rect 33684 41728 33730 41774
rect 33787 41728 33833 41774
rect 33890 41728 33936 41774
rect 33993 41728 34039 41774
rect 34096 41728 34142 41774
rect 34199 41728 34245 41774
rect 34302 41728 34348 41774
rect 34405 41728 34451 41774
rect 34508 41728 34554 41774
rect 34612 41728 34658 41774
rect 39740 41728 39786 41774
rect 39862 41728 39908 41774
rect 39985 41728 40031 41774
rect 40108 41728 40154 41774
rect 33684 41504 33730 41550
rect 33787 41504 33833 41550
rect 33890 41504 33936 41550
rect 33993 41504 34039 41550
rect 34096 41504 34142 41550
rect 34199 41504 34245 41550
rect 34302 41504 34348 41550
rect 34405 41504 34451 41550
rect 34508 41504 34554 41550
rect 34612 41504 34658 41550
rect 39740 41504 39786 41550
rect 39862 41504 39908 41550
rect 39985 41504 40031 41550
rect 40108 41504 40154 41550
rect 50467 41728 50513 41774
rect 50571 41728 50617 41774
rect 50674 41728 50720 41774
rect 50777 41728 50823 41774
rect 50880 41728 50926 41774
rect 50983 41728 51029 41774
rect 51086 41728 51132 41774
rect 51189 41728 51235 41774
rect 51292 41728 51338 41774
rect 51395 41728 51441 41774
rect 43739 41504 43785 41550
rect 43906 41504 43952 41550
rect 44071 41504 44117 41550
rect 44236 41504 44282 41550
rect 33684 41280 33730 41326
rect 33787 41280 33833 41326
rect 33890 41280 33936 41326
rect 33993 41280 34039 41326
rect 34096 41280 34142 41326
rect 34199 41280 34245 41326
rect 34302 41280 34348 41326
rect 34405 41280 34451 41326
rect 34508 41280 34554 41326
rect 34612 41280 34658 41326
rect 39740 41280 39786 41326
rect 39862 41280 39908 41326
rect 39985 41280 40031 41326
rect 40108 41280 40154 41326
rect 50467 41504 50513 41550
rect 50571 41504 50617 41550
rect 50674 41504 50720 41550
rect 50777 41504 50823 41550
rect 50880 41504 50926 41550
rect 50983 41504 51029 41550
rect 51086 41504 51132 41550
rect 51189 41504 51235 41550
rect 51292 41504 51338 41550
rect 51395 41504 51441 41550
rect 50467 41280 50513 41326
rect 50571 41280 50617 41326
rect 50674 41280 50720 41326
rect 50777 41280 50823 41326
rect 50880 41280 50926 41326
rect 50983 41280 51029 41326
rect 51086 41280 51132 41326
rect 51189 41280 51235 41326
rect 51292 41280 51338 41326
rect 51395 41280 51441 41326
rect 37909 41193 37955 41239
rect 38026 41193 38072 41239
rect 38143 41193 38189 41239
rect 38261 41193 38307 41239
rect 38379 41193 38425 41239
rect 38497 41193 38543 41239
rect 33684 41056 33730 41102
rect 33787 41056 33833 41102
rect 33890 41056 33936 41102
rect 33993 41056 34039 41102
rect 34096 41056 34142 41102
rect 34199 41056 34245 41102
rect 34302 41056 34348 41102
rect 34405 41056 34451 41102
rect 34508 41056 34554 41102
rect 34612 41056 34658 41102
rect 33816 40797 33862 40843
rect 34002 40797 34048 40843
rect 34189 40797 34235 40843
rect 34376 40797 34422 40843
rect 34562 40797 34608 40843
rect 37909 40969 37955 41015
rect 38026 40969 38072 41015
rect 38143 40969 38189 41015
rect 38261 40969 38307 41015
rect 38379 40969 38425 41015
rect 38497 40969 38543 41015
rect 39641 40969 39687 41015
rect 50467 41056 50513 41102
rect 50571 41056 50617 41102
rect 50674 41056 50720 41102
rect 50777 41056 50823 41102
rect 50880 41056 50926 41102
rect 50983 41056 51029 41102
rect 51086 41056 51132 41102
rect 51189 41056 51235 41102
rect 51292 41056 51338 41102
rect 51395 41056 51441 41102
rect 37909 40745 37955 40791
rect 38026 40745 38072 40791
rect 38143 40745 38189 40791
rect 38261 40745 38307 40791
rect 38379 40745 38425 40791
rect 38497 40745 38543 40791
rect 39641 40745 39687 40791
rect 43739 40811 43785 40857
rect 43906 40811 43952 40857
rect 44071 40811 44117 40857
rect 44236 40811 44282 40857
rect 50516 40797 50562 40843
rect 50703 40797 50749 40843
rect 50890 40797 50936 40843
rect 51076 40797 51122 40843
rect 51263 40797 51309 40843
rect 33816 40411 33862 40457
rect 34002 40411 34048 40457
rect 34189 40411 34235 40457
rect 34376 40411 34422 40457
rect 34562 40411 34608 40457
rect 37909 40463 37955 40509
rect 38026 40463 38072 40509
rect 38143 40463 38189 40509
rect 38261 40463 38307 40509
rect 38379 40463 38425 40509
rect 38497 40463 38543 40509
rect 39641 40463 39687 40509
rect 33684 40152 33730 40198
rect 33787 40152 33833 40198
rect 33890 40152 33936 40198
rect 33993 40152 34039 40198
rect 34096 40152 34142 40198
rect 34199 40152 34245 40198
rect 34302 40152 34348 40198
rect 34405 40152 34451 40198
rect 34508 40152 34554 40198
rect 34612 40152 34658 40198
rect 37909 40239 37955 40285
rect 38026 40239 38072 40285
rect 38143 40239 38189 40285
rect 38261 40239 38307 40285
rect 38379 40239 38425 40285
rect 38497 40239 38543 40285
rect 43739 40397 43785 40443
rect 43906 40397 43952 40443
rect 44071 40397 44117 40443
rect 44236 40397 44282 40443
rect 39641 40239 39687 40285
rect 50516 40411 50562 40457
rect 50703 40411 50749 40457
rect 50890 40411 50936 40457
rect 51076 40411 51122 40457
rect 51263 40411 51309 40457
rect 37909 40015 37955 40061
rect 38026 40015 38072 40061
rect 38143 40015 38189 40061
rect 38261 40015 38307 40061
rect 38379 40015 38425 40061
rect 38497 40015 38543 40061
rect 50467 40152 50513 40198
rect 50571 40152 50617 40198
rect 50674 40152 50720 40198
rect 50777 40152 50823 40198
rect 50880 40152 50926 40198
rect 50983 40152 51029 40198
rect 51086 40152 51132 40198
rect 51189 40152 51235 40198
rect 51292 40152 51338 40198
rect 51395 40152 51441 40198
rect 33684 39928 33730 39974
rect 33787 39928 33833 39974
rect 33890 39928 33936 39974
rect 33993 39928 34039 39974
rect 34096 39928 34142 39974
rect 34199 39928 34245 39974
rect 34302 39928 34348 39974
rect 34405 39928 34451 39974
rect 34508 39928 34554 39974
rect 34612 39928 34658 39974
rect 39740 39928 39786 39974
rect 39862 39928 39908 39974
rect 39985 39928 40031 39974
rect 40108 39928 40154 39974
rect 33684 39704 33730 39750
rect 33787 39704 33833 39750
rect 33890 39704 33936 39750
rect 33993 39704 34039 39750
rect 34096 39704 34142 39750
rect 34199 39704 34245 39750
rect 34302 39704 34348 39750
rect 34405 39704 34451 39750
rect 34508 39704 34554 39750
rect 34612 39704 34658 39750
rect 39740 39704 39786 39750
rect 39862 39704 39908 39750
rect 39985 39704 40031 39750
rect 40108 39704 40154 39750
rect 50467 39928 50513 39974
rect 50571 39928 50617 39974
rect 50674 39928 50720 39974
rect 50777 39928 50823 39974
rect 50880 39928 50926 39974
rect 50983 39928 51029 39974
rect 51086 39928 51132 39974
rect 51189 39928 51235 39974
rect 51292 39928 51338 39974
rect 51395 39928 51441 39974
rect 43739 39704 43785 39750
rect 43906 39704 43952 39750
rect 44071 39704 44117 39750
rect 44236 39704 44282 39750
rect 33684 39480 33730 39526
rect 33787 39480 33833 39526
rect 33890 39480 33936 39526
rect 33993 39480 34039 39526
rect 34096 39480 34142 39526
rect 34199 39480 34245 39526
rect 34302 39480 34348 39526
rect 34405 39480 34451 39526
rect 34508 39480 34554 39526
rect 34612 39480 34658 39526
rect 39740 39480 39786 39526
rect 39862 39480 39908 39526
rect 39985 39480 40031 39526
rect 40108 39480 40154 39526
rect 50467 39704 50513 39750
rect 50571 39704 50617 39750
rect 50674 39704 50720 39750
rect 50777 39704 50823 39750
rect 50880 39704 50926 39750
rect 50983 39704 51029 39750
rect 51086 39704 51132 39750
rect 51189 39704 51235 39750
rect 51292 39704 51338 39750
rect 51395 39704 51441 39750
rect 50467 39480 50513 39526
rect 50571 39480 50617 39526
rect 50674 39480 50720 39526
rect 50777 39480 50823 39526
rect 50880 39480 50926 39526
rect 50983 39480 51029 39526
rect 51086 39480 51132 39526
rect 51189 39480 51235 39526
rect 51292 39480 51338 39526
rect 51395 39480 51441 39526
rect 37909 39393 37955 39439
rect 38026 39393 38072 39439
rect 38143 39393 38189 39439
rect 38261 39393 38307 39439
rect 38379 39393 38425 39439
rect 38497 39393 38543 39439
rect 33684 39256 33730 39302
rect 33787 39256 33833 39302
rect 33890 39256 33936 39302
rect 33993 39256 34039 39302
rect 34096 39256 34142 39302
rect 34199 39256 34245 39302
rect 34302 39256 34348 39302
rect 34405 39256 34451 39302
rect 34508 39256 34554 39302
rect 34612 39256 34658 39302
rect 33816 38997 33862 39043
rect 34002 38997 34048 39043
rect 34189 38997 34235 39043
rect 34376 38997 34422 39043
rect 34562 38997 34608 39043
rect 37909 39169 37955 39215
rect 38026 39169 38072 39215
rect 38143 39169 38189 39215
rect 38261 39169 38307 39215
rect 38379 39169 38425 39215
rect 38497 39169 38543 39215
rect 39641 39169 39687 39215
rect 50467 39256 50513 39302
rect 50571 39256 50617 39302
rect 50674 39256 50720 39302
rect 50777 39256 50823 39302
rect 50880 39256 50926 39302
rect 50983 39256 51029 39302
rect 51086 39256 51132 39302
rect 51189 39256 51235 39302
rect 51292 39256 51338 39302
rect 51395 39256 51441 39302
rect 37909 38945 37955 38991
rect 38026 38945 38072 38991
rect 38143 38945 38189 38991
rect 38261 38945 38307 38991
rect 38379 38945 38425 38991
rect 38497 38945 38543 38991
rect 39641 38945 39687 38991
rect 43739 39011 43785 39057
rect 43906 39011 43952 39057
rect 44071 39011 44117 39057
rect 44236 39011 44282 39057
rect 50516 38997 50562 39043
rect 50703 38997 50749 39043
rect 50890 38997 50936 39043
rect 51076 38997 51122 39043
rect 51263 38997 51309 39043
rect 33816 38611 33862 38657
rect 34002 38611 34048 38657
rect 34189 38611 34235 38657
rect 34376 38611 34422 38657
rect 34562 38611 34608 38657
rect 37909 38663 37955 38709
rect 38026 38663 38072 38709
rect 38143 38663 38189 38709
rect 38261 38663 38307 38709
rect 38379 38663 38425 38709
rect 38497 38663 38543 38709
rect 39641 38663 39687 38709
rect 33684 38352 33730 38398
rect 33787 38352 33833 38398
rect 33890 38352 33936 38398
rect 33993 38352 34039 38398
rect 34096 38352 34142 38398
rect 34199 38352 34245 38398
rect 34302 38352 34348 38398
rect 34405 38352 34451 38398
rect 34508 38352 34554 38398
rect 34612 38352 34658 38398
rect 37909 38439 37955 38485
rect 38026 38439 38072 38485
rect 38143 38439 38189 38485
rect 38261 38439 38307 38485
rect 38379 38439 38425 38485
rect 38497 38439 38543 38485
rect 43739 38597 43785 38643
rect 43906 38597 43952 38643
rect 44071 38597 44117 38643
rect 44236 38597 44282 38643
rect 39641 38439 39687 38485
rect 50516 38611 50562 38657
rect 50703 38611 50749 38657
rect 50890 38611 50936 38657
rect 51076 38611 51122 38657
rect 51263 38611 51309 38657
rect 37909 38215 37955 38261
rect 38026 38215 38072 38261
rect 38143 38215 38189 38261
rect 38261 38215 38307 38261
rect 38379 38215 38425 38261
rect 38497 38215 38543 38261
rect 50467 38352 50513 38398
rect 50571 38352 50617 38398
rect 50674 38352 50720 38398
rect 50777 38352 50823 38398
rect 50880 38352 50926 38398
rect 50983 38352 51029 38398
rect 51086 38352 51132 38398
rect 51189 38352 51235 38398
rect 51292 38352 51338 38398
rect 51395 38352 51441 38398
rect 33684 38128 33730 38174
rect 33787 38128 33833 38174
rect 33890 38128 33936 38174
rect 33993 38128 34039 38174
rect 34096 38128 34142 38174
rect 34199 38128 34245 38174
rect 34302 38128 34348 38174
rect 34405 38128 34451 38174
rect 34508 38128 34554 38174
rect 34612 38128 34658 38174
rect 39740 38128 39786 38174
rect 39862 38128 39908 38174
rect 39985 38128 40031 38174
rect 40108 38128 40154 38174
rect 33684 37904 33730 37950
rect 33787 37904 33833 37950
rect 33890 37904 33936 37950
rect 33993 37904 34039 37950
rect 34096 37904 34142 37950
rect 34199 37904 34245 37950
rect 34302 37904 34348 37950
rect 34405 37904 34451 37950
rect 34508 37904 34554 37950
rect 34612 37904 34658 37950
rect 39740 37904 39786 37950
rect 39862 37904 39908 37950
rect 39985 37904 40031 37950
rect 40108 37904 40154 37950
rect 50467 38128 50513 38174
rect 50571 38128 50617 38174
rect 50674 38128 50720 38174
rect 50777 38128 50823 38174
rect 50880 38128 50926 38174
rect 50983 38128 51029 38174
rect 51086 38128 51132 38174
rect 51189 38128 51235 38174
rect 51292 38128 51338 38174
rect 51395 38128 51441 38174
rect 43739 37904 43785 37950
rect 43906 37904 43952 37950
rect 44071 37904 44117 37950
rect 44236 37904 44282 37950
rect 33684 37680 33730 37726
rect 33787 37680 33833 37726
rect 33890 37680 33936 37726
rect 33993 37680 34039 37726
rect 34096 37680 34142 37726
rect 34199 37680 34245 37726
rect 34302 37680 34348 37726
rect 34405 37680 34451 37726
rect 34508 37680 34554 37726
rect 34612 37680 34658 37726
rect 39740 37680 39786 37726
rect 39862 37680 39908 37726
rect 39985 37680 40031 37726
rect 40108 37680 40154 37726
rect 50467 37904 50513 37950
rect 50571 37904 50617 37950
rect 50674 37904 50720 37950
rect 50777 37904 50823 37950
rect 50880 37904 50926 37950
rect 50983 37904 51029 37950
rect 51086 37904 51132 37950
rect 51189 37904 51235 37950
rect 51292 37904 51338 37950
rect 51395 37904 51441 37950
rect 50467 37680 50513 37726
rect 50571 37680 50617 37726
rect 50674 37680 50720 37726
rect 50777 37680 50823 37726
rect 50880 37680 50926 37726
rect 50983 37680 51029 37726
rect 51086 37680 51132 37726
rect 51189 37680 51235 37726
rect 51292 37680 51338 37726
rect 51395 37680 51441 37726
rect 37909 37593 37955 37639
rect 38026 37593 38072 37639
rect 38143 37593 38189 37639
rect 38261 37593 38307 37639
rect 38379 37593 38425 37639
rect 38497 37593 38543 37639
rect 33684 37456 33730 37502
rect 33787 37456 33833 37502
rect 33890 37456 33936 37502
rect 33993 37456 34039 37502
rect 34096 37456 34142 37502
rect 34199 37456 34245 37502
rect 34302 37456 34348 37502
rect 34405 37456 34451 37502
rect 34508 37456 34554 37502
rect 34612 37456 34658 37502
rect 33816 37197 33862 37243
rect 34002 37197 34048 37243
rect 34189 37197 34235 37243
rect 34376 37197 34422 37243
rect 34562 37197 34608 37243
rect 37909 37369 37955 37415
rect 38026 37369 38072 37415
rect 38143 37369 38189 37415
rect 38261 37369 38307 37415
rect 38379 37369 38425 37415
rect 38497 37369 38543 37415
rect 39641 37369 39687 37415
rect 50467 37456 50513 37502
rect 50571 37456 50617 37502
rect 50674 37456 50720 37502
rect 50777 37456 50823 37502
rect 50880 37456 50926 37502
rect 50983 37456 51029 37502
rect 51086 37456 51132 37502
rect 51189 37456 51235 37502
rect 51292 37456 51338 37502
rect 51395 37456 51441 37502
rect 37909 37145 37955 37191
rect 38026 37145 38072 37191
rect 38143 37145 38189 37191
rect 38261 37145 38307 37191
rect 38379 37145 38425 37191
rect 38497 37145 38543 37191
rect 39641 37145 39687 37191
rect 43739 37211 43785 37257
rect 43906 37211 43952 37257
rect 44071 37211 44117 37257
rect 44236 37211 44282 37257
rect 50516 37197 50562 37243
rect 50703 37197 50749 37243
rect 50890 37197 50936 37243
rect 51076 37197 51122 37243
rect 51263 37197 51309 37243
rect 33816 36811 33862 36857
rect 34002 36811 34048 36857
rect 34189 36811 34235 36857
rect 34376 36811 34422 36857
rect 34562 36811 34608 36857
rect 37909 36863 37955 36909
rect 38026 36863 38072 36909
rect 38143 36863 38189 36909
rect 38261 36863 38307 36909
rect 38379 36863 38425 36909
rect 38497 36863 38543 36909
rect 39641 36863 39687 36909
rect 33684 36552 33730 36598
rect 33787 36552 33833 36598
rect 33890 36552 33936 36598
rect 33993 36552 34039 36598
rect 34096 36552 34142 36598
rect 34199 36552 34245 36598
rect 34302 36552 34348 36598
rect 34405 36552 34451 36598
rect 34508 36552 34554 36598
rect 34612 36552 34658 36598
rect 37909 36639 37955 36685
rect 38026 36639 38072 36685
rect 38143 36639 38189 36685
rect 38261 36639 38307 36685
rect 38379 36639 38425 36685
rect 38497 36639 38543 36685
rect 43739 36797 43785 36843
rect 43906 36797 43952 36843
rect 44071 36797 44117 36843
rect 44236 36797 44282 36843
rect 39641 36639 39687 36685
rect 50516 36811 50562 36857
rect 50703 36811 50749 36857
rect 50890 36811 50936 36857
rect 51076 36811 51122 36857
rect 51263 36811 51309 36857
rect 37909 36415 37955 36461
rect 38026 36415 38072 36461
rect 38143 36415 38189 36461
rect 38261 36415 38307 36461
rect 38379 36415 38425 36461
rect 38497 36415 38543 36461
rect 50467 36552 50513 36598
rect 50571 36552 50617 36598
rect 50674 36552 50720 36598
rect 50777 36552 50823 36598
rect 50880 36552 50926 36598
rect 50983 36552 51029 36598
rect 51086 36552 51132 36598
rect 51189 36552 51235 36598
rect 51292 36552 51338 36598
rect 51395 36552 51441 36598
rect 33684 36328 33730 36374
rect 33787 36328 33833 36374
rect 33890 36328 33936 36374
rect 33993 36328 34039 36374
rect 34096 36328 34142 36374
rect 34199 36328 34245 36374
rect 34302 36328 34348 36374
rect 34405 36328 34451 36374
rect 34508 36328 34554 36374
rect 34612 36328 34658 36374
rect 39740 36328 39786 36374
rect 39862 36328 39908 36374
rect 39985 36328 40031 36374
rect 40108 36328 40154 36374
rect 33684 36104 33730 36150
rect 33787 36104 33833 36150
rect 33890 36104 33936 36150
rect 33993 36104 34039 36150
rect 34096 36104 34142 36150
rect 34199 36104 34245 36150
rect 34302 36104 34348 36150
rect 34405 36104 34451 36150
rect 34508 36104 34554 36150
rect 34612 36104 34658 36150
rect 39740 36104 39786 36150
rect 39862 36104 39908 36150
rect 39985 36104 40031 36150
rect 40108 36104 40154 36150
rect 50467 36328 50513 36374
rect 50571 36328 50617 36374
rect 50674 36328 50720 36374
rect 50777 36328 50823 36374
rect 50880 36328 50926 36374
rect 50983 36328 51029 36374
rect 51086 36328 51132 36374
rect 51189 36328 51235 36374
rect 51292 36328 51338 36374
rect 51395 36328 51441 36374
rect 43739 36104 43785 36150
rect 43906 36104 43952 36150
rect 44071 36104 44117 36150
rect 44236 36104 44282 36150
rect 50467 36104 50513 36150
rect 50571 36104 50617 36150
rect 50674 36104 50720 36150
rect 50777 36104 50823 36150
rect 50880 36104 50926 36150
rect 50983 36104 51029 36150
rect 51086 36104 51132 36150
rect 51189 36104 51235 36150
rect 51292 36104 51338 36150
rect 51395 36104 51441 36150
<< mvpdiffc >>
rect 29317 44204 29363 44250
rect 29478 44204 29524 44250
rect 29638 44204 29684 44250
rect 29798 44204 29844 44250
rect 29959 44204 30005 44250
rect 30121 44204 30167 44250
rect 30284 44204 30330 44250
rect 35409 44172 37291 44218
rect 37348 44172 37394 44218
rect 37451 44172 37497 44218
rect 37554 44172 37600 44218
rect 37657 44172 37703 44218
rect 37760 44172 37806 44218
rect 37863 44172 37909 44218
rect 35409 43948 37291 43994
rect 37348 43948 37394 43994
rect 37451 43948 37497 43994
rect 37554 43948 37600 43994
rect 37657 43948 37703 43994
rect 37760 43948 37806 43994
rect 37863 43948 37909 43994
rect 38376 43948 38422 43994
rect 38479 43948 38525 43994
rect 38582 43948 38628 43994
rect 38686 43948 38732 43994
rect 38790 43948 38836 43994
rect 38894 43948 38940 43994
rect 38998 43948 39044 43994
rect 39102 43948 39148 43994
rect 39206 43948 39252 43994
rect 39310 43948 39356 43994
rect 39414 43948 39460 43994
rect 39518 43948 39564 43994
rect 39622 43948 39668 43994
rect 42676 43948 42722 43994
rect 42779 43948 42825 43994
rect 42882 43948 42928 43994
rect 42986 43948 43032 43994
rect 43090 43948 43136 43994
rect 43194 43948 43240 43994
rect 43298 43948 43344 43994
rect 43402 43948 43448 43994
rect 43506 43948 43552 43994
rect 43610 43948 43656 43994
rect 43714 43948 43760 43994
rect 43818 43948 43864 43994
rect 43922 43948 43968 43994
rect 47114 44172 48996 44218
rect 49053 44172 49099 44218
rect 49156 44172 49202 44218
rect 49259 44172 49305 44218
rect 49362 44172 49408 44218
rect 49465 44172 49511 44218
rect 49568 44172 49614 44218
rect 35409 43724 37291 43770
rect 37348 43724 37394 43770
rect 37451 43724 37497 43770
rect 37554 43724 37600 43770
rect 37657 43724 37703 43770
rect 37760 43724 37806 43770
rect 37863 43724 37909 43770
rect 38376 43724 38422 43770
rect 38479 43724 38525 43770
rect 38582 43724 38628 43770
rect 38686 43724 38732 43770
rect 38790 43724 38836 43770
rect 38894 43724 38940 43770
rect 38998 43724 39044 43770
rect 39102 43724 39148 43770
rect 39206 43724 39252 43770
rect 39310 43724 39356 43770
rect 39414 43724 39460 43770
rect 39518 43724 39564 43770
rect 39622 43724 39668 43770
rect 45346 43948 45392 43994
rect 45449 43948 45495 43994
rect 45552 43948 45598 43994
rect 45656 43948 45702 43994
rect 45760 43948 45806 43994
rect 45864 43948 45910 43994
rect 45968 43948 46014 43994
rect 46072 43948 46118 43994
rect 46176 43948 46222 43994
rect 46280 43948 46326 43994
rect 46384 43948 46430 43994
rect 46488 43948 46534 43994
rect 46592 43948 46638 43994
rect 47114 43948 48996 43994
rect 49053 43948 49099 43994
rect 49156 43948 49202 43994
rect 49259 43948 49305 43994
rect 49362 43948 49408 43994
rect 49465 43948 49511 43994
rect 49568 43948 49614 43994
rect 54793 44204 54839 44250
rect 54956 44204 55002 44250
rect 55118 44204 55164 44250
rect 55279 44204 55325 44250
rect 55439 44204 55485 44250
rect 55599 44204 55645 44250
rect 55760 44204 55806 44250
rect 42676 43724 42722 43770
rect 42779 43724 42825 43770
rect 42882 43724 42928 43770
rect 42986 43724 43032 43770
rect 43090 43724 43136 43770
rect 43194 43724 43240 43770
rect 43298 43724 43344 43770
rect 43402 43724 43448 43770
rect 43506 43724 43552 43770
rect 43610 43724 43656 43770
rect 43714 43724 43760 43770
rect 43818 43724 43864 43770
rect 43922 43724 43968 43770
rect 45346 43724 45392 43770
rect 45449 43724 45495 43770
rect 45552 43724 45598 43770
rect 45656 43724 45702 43770
rect 45760 43724 45806 43770
rect 45864 43724 45910 43770
rect 45968 43724 46014 43770
rect 46072 43724 46118 43770
rect 46176 43724 46222 43770
rect 46280 43724 46326 43770
rect 46384 43724 46430 43770
rect 46488 43724 46534 43770
rect 46592 43724 46638 43770
rect 47114 43724 48996 43770
rect 49053 43724 49099 43770
rect 49156 43724 49202 43770
rect 49259 43724 49305 43770
rect 49362 43724 49408 43770
rect 49465 43724 49511 43770
rect 49568 43724 49614 43770
rect 29317 43304 29363 43350
rect 29478 43304 29524 43350
rect 29638 43304 29684 43350
rect 29798 43304 29844 43350
rect 29959 43304 30005 43350
rect 30121 43304 30167 43350
rect 30284 43304 30330 43350
rect 31349 43304 33323 43350
rect 31349 43080 33323 43126
rect 31349 42856 33323 42902
rect 44812 43304 44858 43350
rect 44925 43304 44971 43350
rect 45038 43304 45084 43350
rect 45151 43304 45197 43350
rect 45264 43304 45310 43350
rect 51802 43304 53776 43350
rect 35273 42993 35523 43039
rect 35580 42993 35626 43039
rect 35683 42993 35729 43039
rect 35786 42993 35832 43039
rect 35889 42993 35935 43039
rect 35992 42993 36038 43039
rect 36095 42993 36141 43039
rect 36198 42993 36244 43039
rect 36301 42993 36347 43039
rect 36854 42993 36900 43039
rect 36971 42993 37017 43039
rect 37088 42993 37134 43039
rect 37206 42993 37252 43039
rect 37324 42993 37370 43039
rect 37442 42993 37488 43039
rect 44812 43080 44858 43126
rect 44925 43080 44971 43126
rect 45038 43080 45084 43126
rect 45151 43080 45197 43126
rect 45264 43080 45310 43126
rect 54793 43304 54839 43350
rect 54956 43304 55002 43350
rect 55118 43304 55164 43350
rect 55279 43304 55325 43350
rect 55439 43304 55485 43350
rect 55599 43304 55645 43350
rect 55760 43304 55806 43350
rect 31349 42632 33323 42678
rect 35273 42769 35523 42815
rect 35580 42769 35626 42815
rect 35683 42769 35729 42815
rect 35786 42769 35832 42815
rect 35889 42769 35935 42815
rect 35992 42769 36038 42815
rect 36095 42769 36141 42815
rect 36198 42769 36244 42815
rect 36301 42769 36347 42815
rect 48778 42993 48824 43039
rect 48881 42993 48927 43039
rect 48984 42993 49030 43039
rect 49087 42993 49133 43039
rect 49190 42993 49236 43039
rect 49293 42993 49339 43039
rect 49396 42993 49442 43039
rect 49499 42993 49545 43039
rect 49602 42993 49852 43039
rect 36854 42769 36900 42815
rect 36971 42769 37017 42815
rect 37088 42769 37134 42815
rect 37206 42769 37252 42815
rect 37324 42769 37370 42815
rect 37442 42769 37488 42815
rect 39021 42769 39067 42815
rect 39144 42769 39190 42815
rect 39267 42769 39313 42815
rect 44812 42856 44858 42902
rect 44925 42856 44971 42902
rect 45038 42856 45084 42902
rect 45151 42856 45197 42902
rect 45264 42856 45310 42902
rect 48778 42769 48824 42815
rect 48881 42769 48927 42815
rect 48984 42769 49030 42815
rect 49087 42769 49133 42815
rect 49190 42769 49236 42815
rect 49293 42769 49339 42815
rect 49396 42769 49442 42815
rect 49499 42769 49545 42815
rect 49602 42769 49852 42815
rect 35273 42545 35523 42591
rect 35580 42545 35626 42591
rect 35683 42545 35729 42591
rect 35786 42545 35832 42591
rect 35889 42545 35935 42591
rect 35992 42545 36038 42591
rect 36095 42545 36141 42591
rect 36198 42545 36244 42591
rect 36301 42545 36347 42591
rect 36854 42545 36900 42591
rect 36971 42545 37017 42591
rect 37088 42545 37134 42591
rect 37206 42545 37252 42591
rect 37324 42545 37370 42591
rect 37442 42545 37488 42591
rect 39021 42545 39067 42591
rect 39144 42545 39190 42591
rect 39267 42545 39313 42591
rect 44812 42632 44858 42678
rect 44925 42632 44971 42678
rect 45038 42632 45084 42678
rect 45151 42632 45197 42678
rect 45264 42632 45310 42678
rect 51802 43080 53776 43126
rect 51802 42856 53776 42902
rect 48778 42545 48824 42591
rect 48881 42545 48927 42591
rect 48984 42545 49030 42591
rect 49087 42545 49133 42591
rect 49190 42545 49236 42591
rect 49293 42545 49339 42591
rect 49396 42545 49442 42591
rect 49499 42545 49545 42591
rect 49602 42545 49852 42591
rect 51802 42632 53776 42678
rect 29317 42404 29363 42450
rect 29478 42404 29524 42450
rect 29638 42404 29684 42450
rect 29798 42404 29844 42450
rect 29959 42404 30005 42450
rect 30121 42404 30167 42450
rect 30284 42404 30330 42450
rect 54793 42404 54839 42450
rect 54956 42404 55002 42450
rect 55118 42404 55164 42450
rect 55279 42404 55325 42450
rect 55439 42404 55485 42450
rect 55599 42404 55645 42450
rect 55760 42404 55806 42450
rect 31349 42176 33323 42222
rect 35273 42263 35523 42309
rect 35580 42263 35626 42309
rect 35683 42263 35729 42309
rect 35786 42263 35832 42309
rect 35889 42263 35935 42309
rect 35992 42263 36038 42309
rect 36095 42263 36141 42309
rect 36198 42263 36244 42309
rect 36301 42263 36347 42309
rect 36854 42263 36900 42309
rect 36971 42263 37017 42309
rect 37088 42263 37134 42309
rect 37206 42263 37252 42309
rect 37324 42263 37370 42309
rect 37442 42263 37488 42309
rect 39021 42263 39067 42309
rect 39144 42263 39190 42309
rect 39267 42263 39313 42309
rect 31349 41952 33323 41998
rect 31349 41728 33323 41774
rect 29317 41504 29363 41550
rect 29478 41504 29524 41550
rect 29638 41504 29684 41550
rect 29798 41504 29844 41550
rect 29959 41504 30005 41550
rect 30121 41504 30167 41550
rect 30284 41504 30330 41550
rect 35273 42039 35523 42085
rect 35580 42039 35626 42085
rect 35683 42039 35729 42085
rect 35786 42039 35832 42085
rect 35889 42039 35935 42085
rect 35992 42039 36038 42085
rect 36095 42039 36141 42085
rect 36198 42039 36244 42085
rect 36301 42039 36347 42085
rect 36854 42039 36900 42085
rect 36971 42039 37017 42085
rect 37088 42039 37134 42085
rect 37206 42039 37252 42085
rect 37324 42039 37370 42085
rect 37442 42039 37488 42085
rect 48778 42263 48824 42309
rect 48881 42263 48927 42309
rect 48984 42263 49030 42309
rect 49087 42263 49133 42309
rect 49190 42263 49236 42309
rect 49293 42263 49339 42309
rect 49396 42263 49442 42309
rect 49499 42263 49545 42309
rect 49602 42263 49852 42309
rect 44812 42176 44858 42222
rect 44925 42176 44971 42222
rect 45038 42176 45084 42222
rect 45151 42176 45197 42222
rect 45264 42176 45310 42222
rect 39021 42039 39067 42085
rect 39144 42039 39190 42085
rect 39267 42039 39313 42085
rect 44812 41952 44858 41998
rect 44925 41952 44971 41998
rect 45038 41952 45084 41998
rect 45151 41952 45197 41998
rect 45264 41952 45310 41998
rect 48778 42039 48824 42085
rect 48881 42039 48927 42085
rect 48984 42039 49030 42085
rect 49087 42039 49133 42085
rect 49190 42039 49236 42085
rect 49293 42039 49339 42085
rect 49396 42039 49442 42085
rect 49499 42039 49545 42085
rect 49602 42039 49852 42085
rect 51802 42176 53776 42222
rect 35273 41815 35523 41861
rect 35580 41815 35626 41861
rect 35683 41815 35729 41861
rect 35786 41815 35832 41861
rect 35889 41815 35935 41861
rect 35992 41815 36038 41861
rect 36095 41815 36141 41861
rect 36198 41815 36244 41861
rect 36301 41815 36347 41861
rect 36854 41815 36900 41861
rect 36971 41815 37017 41861
rect 37088 41815 37134 41861
rect 37206 41815 37252 41861
rect 37324 41815 37370 41861
rect 37442 41815 37488 41861
rect 48778 41815 48824 41861
rect 48881 41815 48927 41861
rect 48984 41815 49030 41861
rect 49087 41815 49133 41861
rect 49190 41815 49236 41861
rect 49293 41815 49339 41861
rect 49396 41815 49442 41861
rect 49499 41815 49545 41861
rect 49602 41815 49852 41861
rect 44812 41728 44858 41774
rect 44925 41728 44971 41774
rect 45038 41728 45084 41774
rect 45151 41728 45197 41774
rect 45264 41728 45310 41774
rect 31349 41504 33323 41550
rect 31349 41280 33323 41326
rect 31349 41056 33323 41102
rect 51802 41952 53776 41998
rect 51802 41728 53776 41774
rect 44812 41504 44858 41550
rect 44925 41504 44971 41550
rect 45038 41504 45084 41550
rect 45151 41504 45197 41550
rect 45264 41504 45310 41550
rect 51802 41504 53776 41550
rect 35273 41193 35523 41239
rect 35580 41193 35626 41239
rect 35683 41193 35729 41239
rect 35786 41193 35832 41239
rect 35889 41193 35935 41239
rect 35992 41193 36038 41239
rect 36095 41193 36141 41239
rect 36198 41193 36244 41239
rect 36301 41193 36347 41239
rect 36854 41193 36900 41239
rect 36971 41193 37017 41239
rect 37088 41193 37134 41239
rect 37206 41193 37252 41239
rect 37324 41193 37370 41239
rect 37442 41193 37488 41239
rect 44812 41280 44858 41326
rect 44925 41280 44971 41326
rect 45038 41280 45084 41326
rect 45151 41280 45197 41326
rect 45264 41280 45310 41326
rect 54793 41504 54839 41550
rect 54956 41504 55002 41550
rect 55118 41504 55164 41550
rect 55279 41504 55325 41550
rect 55439 41504 55485 41550
rect 55599 41504 55645 41550
rect 55760 41504 55806 41550
rect 31349 40832 33323 40878
rect 35273 40969 35523 41015
rect 35580 40969 35626 41015
rect 35683 40969 35729 41015
rect 35786 40969 35832 41015
rect 35889 40969 35935 41015
rect 35992 40969 36038 41015
rect 36095 40969 36141 41015
rect 36198 40969 36244 41015
rect 36301 40969 36347 41015
rect 48778 41193 48824 41239
rect 48881 41193 48927 41239
rect 48984 41193 49030 41239
rect 49087 41193 49133 41239
rect 49190 41193 49236 41239
rect 49293 41193 49339 41239
rect 49396 41193 49442 41239
rect 49499 41193 49545 41239
rect 49602 41193 49852 41239
rect 36854 40969 36900 41015
rect 36971 40969 37017 41015
rect 37088 40969 37134 41015
rect 37206 40969 37252 41015
rect 37324 40969 37370 41015
rect 37442 40969 37488 41015
rect 39021 40969 39067 41015
rect 39144 40969 39190 41015
rect 39267 40969 39313 41015
rect 44812 41056 44858 41102
rect 44925 41056 44971 41102
rect 45038 41056 45084 41102
rect 45151 41056 45197 41102
rect 45264 41056 45310 41102
rect 48778 40969 48824 41015
rect 48881 40969 48927 41015
rect 48984 40969 49030 41015
rect 49087 40969 49133 41015
rect 49190 40969 49236 41015
rect 49293 40969 49339 41015
rect 49396 40969 49442 41015
rect 49499 40969 49545 41015
rect 49602 40969 49852 41015
rect 35273 40745 35523 40791
rect 35580 40745 35626 40791
rect 35683 40745 35729 40791
rect 35786 40745 35832 40791
rect 35889 40745 35935 40791
rect 35992 40745 36038 40791
rect 36095 40745 36141 40791
rect 36198 40745 36244 40791
rect 36301 40745 36347 40791
rect 36854 40745 36900 40791
rect 36971 40745 37017 40791
rect 37088 40745 37134 40791
rect 37206 40745 37252 40791
rect 37324 40745 37370 40791
rect 37442 40745 37488 40791
rect 39021 40745 39067 40791
rect 39144 40745 39190 40791
rect 39267 40745 39313 40791
rect 44812 40832 44858 40878
rect 44925 40832 44971 40878
rect 45038 40832 45084 40878
rect 45151 40832 45197 40878
rect 45264 40832 45310 40878
rect 51802 41280 53776 41326
rect 51802 41056 53776 41102
rect 48778 40745 48824 40791
rect 48881 40745 48927 40791
rect 48984 40745 49030 40791
rect 49087 40745 49133 40791
rect 49190 40745 49236 40791
rect 49293 40745 49339 40791
rect 49396 40745 49442 40791
rect 49499 40745 49545 40791
rect 49602 40745 49852 40791
rect 51802 40832 53776 40878
rect 29317 40604 29363 40650
rect 29478 40604 29524 40650
rect 29638 40604 29684 40650
rect 29798 40604 29844 40650
rect 29959 40604 30005 40650
rect 30121 40604 30167 40650
rect 30284 40604 30330 40650
rect 54793 40604 54839 40650
rect 54956 40604 55002 40650
rect 55118 40604 55164 40650
rect 55279 40604 55325 40650
rect 55439 40604 55485 40650
rect 55599 40604 55645 40650
rect 55760 40604 55806 40650
rect 31349 40376 33323 40422
rect 35273 40463 35523 40509
rect 35580 40463 35626 40509
rect 35683 40463 35729 40509
rect 35786 40463 35832 40509
rect 35889 40463 35935 40509
rect 35992 40463 36038 40509
rect 36095 40463 36141 40509
rect 36198 40463 36244 40509
rect 36301 40463 36347 40509
rect 36854 40463 36900 40509
rect 36971 40463 37017 40509
rect 37088 40463 37134 40509
rect 37206 40463 37252 40509
rect 37324 40463 37370 40509
rect 37442 40463 37488 40509
rect 39021 40463 39067 40509
rect 39144 40463 39190 40509
rect 39267 40463 39313 40509
rect 31349 40152 33323 40198
rect 31349 39928 33323 39974
rect 29317 39704 29363 39750
rect 29478 39704 29524 39750
rect 29638 39704 29684 39750
rect 29798 39704 29844 39750
rect 29959 39704 30005 39750
rect 30121 39704 30167 39750
rect 30284 39704 30330 39750
rect 35273 40239 35523 40285
rect 35580 40239 35626 40285
rect 35683 40239 35729 40285
rect 35786 40239 35832 40285
rect 35889 40239 35935 40285
rect 35992 40239 36038 40285
rect 36095 40239 36141 40285
rect 36198 40239 36244 40285
rect 36301 40239 36347 40285
rect 36854 40239 36900 40285
rect 36971 40239 37017 40285
rect 37088 40239 37134 40285
rect 37206 40239 37252 40285
rect 37324 40239 37370 40285
rect 37442 40239 37488 40285
rect 48778 40463 48824 40509
rect 48881 40463 48927 40509
rect 48984 40463 49030 40509
rect 49087 40463 49133 40509
rect 49190 40463 49236 40509
rect 49293 40463 49339 40509
rect 49396 40463 49442 40509
rect 49499 40463 49545 40509
rect 49602 40463 49852 40509
rect 44812 40376 44858 40422
rect 44925 40376 44971 40422
rect 45038 40376 45084 40422
rect 45151 40376 45197 40422
rect 45264 40376 45310 40422
rect 39021 40239 39067 40285
rect 39144 40239 39190 40285
rect 39267 40239 39313 40285
rect 44812 40152 44858 40198
rect 44925 40152 44971 40198
rect 45038 40152 45084 40198
rect 45151 40152 45197 40198
rect 45264 40152 45310 40198
rect 48778 40239 48824 40285
rect 48881 40239 48927 40285
rect 48984 40239 49030 40285
rect 49087 40239 49133 40285
rect 49190 40239 49236 40285
rect 49293 40239 49339 40285
rect 49396 40239 49442 40285
rect 49499 40239 49545 40285
rect 49602 40239 49852 40285
rect 51802 40376 53776 40422
rect 35273 40015 35523 40061
rect 35580 40015 35626 40061
rect 35683 40015 35729 40061
rect 35786 40015 35832 40061
rect 35889 40015 35935 40061
rect 35992 40015 36038 40061
rect 36095 40015 36141 40061
rect 36198 40015 36244 40061
rect 36301 40015 36347 40061
rect 36854 40015 36900 40061
rect 36971 40015 37017 40061
rect 37088 40015 37134 40061
rect 37206 40015 37252 40061
rect 37324 40015 37370 40061
rect 37442 40015 37488 40061
rect 48778 40015 48824 40061
rect 48881 40015 48927 40061
rect 48984 40015 49030 40061
rect 49087 40015 49133 40061
rect 49190 40015 49236 40061
rect 49293 40015 49339 40061
rect 49396 40015 49442 40061
rect 49499 40015 49545 40061
rect 49602 40015 49852 40061
rect 44812 39928 44858 39974
rect 44925 39928 44971 39974
rect 45038 39928 45084 39974
rect 45151 39928 45197 39974
rect 45264 39928 45310 39974
rect 31349 39704 33323 39750
rect 31349 39480 33323 39526
rect 31349 39256 33323 39302
rect 51802 40152 53776 40198
rect 51802 39928 53776 39974
rect 44812 39704 44858 39750
rect 44925 39704 44971 39750
rect 45038 39704 45084 39750
rect 45151 39704 45197 39750
rect 45264 39704 45310 39750
rect 51802 39704 53776 39750
rect 35273 39393 35523 39439
rect 35580 39393 35626 39439
rect 35683 39393 35729 39439
rect 35786 39393 35832 39439
rect 35889 39393 35935 39439
rect 35992 39393 36038 39439
rect 36095 39393 36141 39439
rect 36198 39393 36244 39439
rect 36301 39393 36347 39439
rect 36854 39393 36900 39439
rect 36971 39393 37017 39439
rect 37088 39393 37134 39439
rect 37206 39393 37252 39439
rect 37324 39393 37370 39439
rect 37442 39393 37488 39439
rect 44812 39480 44858 39526
rect 44925 39480 44971 39526
rect 45038 39480 45084 39526
rect 45151 39480 45197 39526
rect 45264 39480 45310 39526
rect 54793 39704 54839 39750
rect 54956 39704 55002 39750
rect 55118 39704 55164 39750
rect 55279 39704 55325 39750
rect 55439 39704 55485 39750
rect 55599 39704 55645 39750
rect 55760 39704 55806 39750
rect 31349 39032 33323 39078
rect 35273 39169 35523 39215
rect 35580 39169 35626 39215
rect 35683 39169 35729 39215
rect 35786 39169 35832 39215
rect 35889 39169 35935 39215
rect 35992 39169 36038 39215
rect 36095 39169 36141 39215
rect 36198 39169 36244 39215
rect 36301 39169 36347 39215
rect 48778 39393 48824 39439
rect 48881 39393 48927 39439
rect 48984 39393 49030 39439
rect 49087 39393 49133 39439
rect 49190 39393 49236 39439
rect 49293 39393 49339 39439
rect 49396 39393 49442 39439
rect 49499 39393 49545 39439
rect 49602 39393 49852 39439
rect 36854 39169 36900 39215
rect 36971 39169 37017 39215
rect 37088 39169 37134 39215
rect 37206 39169 37252 39215
rect 37324 39169 37370 39215
rect 37442 39169 37488 39215
rect 39021 39169 39067 39215
rect 39144 39169 39190 39215
rect 39267 39169 39313 39215
rect 44812 39256 44858 39302
rect 44925 39256 44971 39302
rect 45038 39256 45084 39302
rect 45151 39256 45197 39302
rect 45264 39256 45310 39302
rect 48778 39169 48824 39215
rect 48881 39169 48927 39215
rect 48984 39169 49030 39215
rect 49087 39169 49133 39215
rect 49190 39169 49236 39215
rect 49293 39169 49339 39215
rect 49396 39169 49442 39215
rect 49499 39169 49545 39215
rect 49602 39169 49852 39215
rect 35273 38945 35523 38991
rect 35580 38945 35626 38991
rect 35683 38945 35729 38991
rect 35786 38945 35832 38991
rect 35889 38945 35935 38991
rect 35992 38945 36038 38991
rect 36095 38945 36141 38991
rect 36198 38945 36244 38991
rect 36301 38945 36347 38991
rect 36854 38945 36900 38991
rect 36971 38945 37017 38991
rect 37088 38945 37134 38991
rect 37206 38945 37252 38991
rect 37324 38945 37370 38991
rect 37442 38945 37488 38991
rect 39021 38945 39067 38991
rect 39144 38945 39190 38991
rect 39267 38945 39313 38991
rect 44812 39032 44858 39078
rect 44925 39032 44971 39078
rect 45038 39032 45084 39078
rect 45151 39032 45197 39078
rect 45264 39032 45310 39078
rect 51802 39480 53776 39526
rect 51802 39256 53776 39302
rect 48778 38945 48824 38991
rect 48881 38945 48927 38991
rect 48984 38945 49030 38991
rect 49087 38945 49133 38991
rect 49190 38945 49236 38991
rect 49293 38945 49339 38991
rect 49396 38945 49442 38991
rect 49499 38945 49545 38991
rect 49602 38945 49852 38991
rect 51802 39032 53776 39078
rect 29317 38804 29363 38850
rect 29478 38804 29524 38850
rect 29638 38804 29684 38850
rect 29798 38804 29844 38850
rect 29959 38804 30005 38850
rect 30121 38804 30167 38850
rect 30284 38804 30330 38850
rect 54793 38804 54839 38850
rect 54956 38804 55002 38850
rect 55118 38804 55164 38850
rect 55279 38804 55325 38850
rect 55439 38804 55485 38850
rect 55599 38804 55645 38850
rect 55760 38804 55806 38850
rect 31349 38576 33323 38622
rect 35273 38663 35523 38709
rect 35580 38663 35626 38709
rect 35683 38663 35729 38709
rect 35786 38663 35832 38709
rect 35889 38663 35935 38709
rect 35992 38663 36038 38709
rect 36095 38663 36141 38709
rect 36198 38663 36244 38709
rect 36301 38663 36347 38709
rect 36854 38663 36900 38709
rect 36971 38663 37017 38709
rect 37088 38663 37134 38709
rect 37206 38663 37252 38709
rect 37324 38663 37370 38709
rect 37442 38663 37488 38709
rect 39021 38663 39067 38709
rect 39144 38663 39190 38709
rect 39267 38663 39313 38709
rect 31349 38352 33323 38398
rect 31349 38128 33323 38174
rect 29317 37904 29363 37950
rect 29478 37904 29524 37950
rect 29638 37904 29684 37950
rect 29798 37904 29844 37950
rect 29959 37904 30005 37950
rect 30121 37904 30167 37950
rect 30284 37904 30330 37950
rect 35273 38439 35523 38485
rect 35580 38439 35626 38485
rect 35683 38439 35729 38485
rect 35786 38439 35832 38485
rect 35889 38439 35935 38485
rect 35992 38439 36038 38485
rect 36095 38439 36141 38485
rect 36198 38439 36244 38485
rect 36301 38439 36347 38485
rect 36854 38439 36900 38485
rect 36971 38439 37017 38485
rect 37088 38439 37134 38485
rect 37206 38439 37252 38485
rect 37324 38439 37370 38485
rect 37442 38439 37488 38485
rect 48778 38663 48824 38709
rect 48881 38663 48927 38709
rect 48984 38663 49030 38709
rect 49087 38663 49133 38709
rect 49190 38663 49236 38709
rect 49293 38663 49339 38709
rect 49396 38663 49442 38709
rect 49499 38663 49545 38709
rect 49602 38663 49852 38709
rect 44812 38576 44858 38622
rect 44925 38576 44971 38622
rect 45038 38576 45084 38622
rect 45151 38576 45197 38622
rect 45264 38576 45310 38622
rect 39021 38439 39067 38485
rect 39144 38439 39190 38485
rect 39267 38439 39313 38485
rect 44812 38352 44858 38398
rect 44925 38352 44971 38398
rect 45038 38352 45084 38398
rect 45151 38352 45197 38398
rect 45264 38352 45310 38398
rect 48778 38439 48824 38485
rect 48881 38439 48927 38485
rect 48984 38439 49030 38485
rect 49087 38439 49133 38485
rect 49190 38439 49236 38485
rect 49293 38439 49339 38485
rect 49396 38439 49442 38485
rect 49499 38439 49545 38485
rect 49602 38439 49852 38485
rect 51802 38576 53776 38622
rect 35273 38215 35523 38261
rect 35580 38215 35626 38261
rect 35683 38215 35729 38261
rect 35786 38215 35832 38261
rect 35889 38215 35935 38261
rect 35992 38215 36038 38261
rect 36095 38215 36141 38261
rect 36198 38215 36244 38261
rect 36301 38215 36347 38261
rect 36854 38215 36900 38261
rect 36971 38215 37017 38261
rect 37088 38215 37134 38261
rect 37206 38215 37252 38261
rect 37324 38215 37370 38261
rect 37442 38215 37488 38261
rect 48778 38215 48824 38261
rect 48881 38215 48927 38261
rect 48984 38215 49030 38261
rect 49087 38215 49133 38261
rect 49190 38215 49236 38261
rect 49293 38215 49339 38261
rect 49396 38215 49442 38261
rect 49499 38215 49545 38261
rect 49602 38215 49852 38261
rect 44812 38128 44858 38174
rect 44925 38128 44971 38174
rect 45038 38128 45084 38174
rect 45151 38128 45197 38174
rect 45264 38128 45310 38174
rect 31349 37904 33323 37950
rect 31349 37680 33323 37726
rect 31349 37456 33323 37502
rect 51802 38352 53776 38398
rect 51802 38128 53776 38174
rect 44812 37904 44858 37950
rect 44925 37904 44971 37950
rect 45038 37904 45084 37950
rect 45151 37904 45197 37950
rect 45264 37904 45310 37950
rect 51802 37904 53776 37950
rect 35273 37593 35523 37639
rect 35580 37593 35626 37639
rect 35683 37593 35729 37639
rect 35786 37593 35832 37639
rect 35889 37593 35935 37639
rect 35992 37593 36038 37639
rect 36095 37593 36141 37639
rect 36198 37593 36244 37639
rect 36301 37593 36347 37639
rect 36854 37593 36900 37639
rect 36971 37593 37017 37639
rect 37088 37593 37134 37639
rect 37206 37593 37252 37639
rect 37324 37593 37370 37639
rect 37442 37593 37488 37639
rect 44812 37680 44858 37726
rect 44925 37680 44971 37726
rect 45038 37680 45084 37726
rect 45151 37680 45197 37726
rect 45264 37680 45310 37726
rect 54793 37904 54839 37950
rect 54956 37904 55002 37950
rect 55118 37904 55164 37950
rect 55279 37904 55325 37950
rect 55439 37904 55485 37950
rect 55599 37904 55645 37950
rect 55760 37904 55806 37950
rect 31349 37232 33323 37278
rect 35273 37369 35523 37415
rect 35580 37369 35626 37415
rect 35683 37369 35729 37415
rect 35786 37369 35832 37415
rect 35889 37369 35935 37415
rect 35992 37369 36038 37415
rect 36095 37369 36141 37415
rect 36198 37369 36244 37415
rect 36301 37369 36347 37415
rect 48778 37593 48824 37639
rect 48881 37593 48927 37639
rect 48984 37593 49030 37639
rect 49087 37593 49133 37639
rect 49190 37593 49236 37639
rect 49293 37593 49339 37639
rect 49396 37593 49442 37639
rect 49499 37593 49545 37639
rect 49602 37593 49852 37639
rect 36854 37369 36900 37415
rect 36971 37369 37017 37415
rect 37088 37369 37134 37415
rect 37206 37369 37252 37415
rect 37324 37369 37370 37415
rect 37442 37369 37488 37415
rect 39021 37369 39067 37415
rect 39144 37369 39190 37415
rect 39267 37369 39313 37415
rect 44812 37456 44858 37502
rect 44925 37456 44971 37502
rect 45038 37456 45084 37502
rect 45151 37456 45197 37502
rect 45264 37456 45310 37502
rect 48778 37369 48824 37415
rect 48881 37369 48927 37415
rect 48984 37369 49030 37415
rect 49087 37369 49133 37415
rect 49190 37369 49236 37415
rect 49293 37369 49339 37415
rect 49396 37369 49442 37415
rect 49499 37369 49545 37415
rect 49602 37369 49852 37415
rect 35273 37145 35523 37191
rect 35580 37145 35626 37191
rect 35683 37145 35729 37191
rect 35786 37145 35832 37191
rect 35889 37145 35935 37191
rect 35992 37145 36038 37191
rect 36095 37145 36141 37191
rect 36198 37145 36244 37191
rect 36301 37145 36347 37191
rect 36854 37145 36900 37191
rect 36971 37145 37017 37191
rect 37088 37145 37134 37191
rect 37206 37145 37252 37191
rect 37324 37145 37370 37191
rect 37442 37145 37488 37191
rect 39021 37145 39067 37191
rect 39144 37145 39190 37191
rect 39267 37145 39313 37191
rect 44812 37232 44858 37278
rect 44925 37232 44971 37278
rect 45038 37232 45084 37278
rect 45151 37232 45197 37278
rect 45264 37232 45310 37278
rect 51802 37680 53776 37726
rect 51802 37456 53776 37502
rect 48778 37145 48824 37191
rect 48881 37145 48927 37191
rect 48984 37145 49030 37191
rect 49087 37145 49133 37191
rect 49190 37145 49236 37191
rect 49293 37145 49339 37191
rect 49396 37145 49442 37191
rect 49499 37145 49545 37191
rect 49602 37145 49852 37191
rect 51802 37232 53776 37278
rect 29317 37004 29363 37050
rect 29478 37004 29524 37050
rect 29638 37004 29684 37050
rect 29798 37004 29844 37050
rect 29959 37004 30005 37050
rect 30121 37004 30167 37050
rect 30284 37004 30330 37050
rect 54793 37004 54839 37050
rect 54956 37004 55002 37050
rect 55118 37004 55164 37050
rect 55279 37004 55325 37050
rect 55439 37004 55485 37050
rect 55599 37004 55645 37050
rect 55760 37004 55806 37050
rect 31349 36776 33323 36822
rect 35273 36863 35523 36909
rect 35580 36863 35626 36909
rect 35683 36863 35729 36909
rect 35786 36863 35832 36909
rect 35889 36863 35935 36909
rect 35992 36863 36038 36909
rect 36095 36863 36141 36909
rect 36198 36863 36244 36909
rect 36301 36863 36347 36909
rect 36854 36863 36900 36909
rect 36971 36863 37017 36909
rect 37088 36863 37134 36909
rect 37206 36863 37252 36909
rect 37324 36863 37370 36909
rect 37442 36863 37488 36909
rect 39021 36863 39067 36909
rect 39144 36863 39190 36909
rect 39267 36863 39313 36909
rect 31349 36552 33323 36598
rect 31349 36328 33323 36374
rect 29317 36104 29363 36150
rect 29478 36104 29524 36150
rect 29638 36104 29684 36150
rect 29798 36104 29844 36150
rect 29959 36104 30005 36150
rect 30121 36104 30167 36150
rect 30284 36104 30330 36150
rect 35273 36639 35523 36685
rect 35580 36639 35626 36685
rect 35683 36639 35729 36685
rect 35786 36639 35832 36685
rect 35889 36639 35935 36685
rect 35992 36639 36038 36685
rect 36095 36639 36141 36685
rect 36198 36639 36244 36685
rect 36301 36639 36347 36685
rect 36854 36639 36900 36685
rect 36971 36639 37017 36685
rect 37088 36639 37134 36685
rect 37206 36639 37252 36685
rect 37324 36639 37370 36685
rect 37442 36639 37488 36685
rect 48778 36863 48824 36909
rect 48881 36863 48927 36909
rect 48984 36863 49030 36909
rect 49087 36863 49133 36909
rect 49190 36863 49236 36909
rect 49293 36863 49339 36909
rect 49396 36863 49442 36909
rect 49499 36863 49545 36909
rect 49602 36863 49852 36909
rect 44812 36776 44858 36822
rect 44925 36776 44971 36822
rect 45038 36776 45084 36822
rect 45151 36776 45197 36822
rect 45264 36776 45310 36822
rect 39021 36639 39067 36685
rect 39144 36639 39190 36685
rect 39267 36639 39313 36685
rect 44812 36552 44858 36598
rect 44925 36552 44971 36598
rect 45038 36552 45084 36598
rect 45151 36552 45197 36598
rect 45264 36552 45310 36598
rect 48778 36639 48824 36685
rect 48881 36639 48927 36685
rect 48984 36639 49030 36685
rect 49087 36639 49133 36685
rect 49190 36639 49236 36685
rect 49293 36639 49339 36685
rect 49396 36639 49442 36685
rect 49499 36639 49545 36685
rect 49602 36639 49852 36685
rect 51802 36776 53776 36822
rect 35273 36415 35523 36461
rect 35580 36415 35626 36461
rect 35683 36415 35729 36461
rect 35786 36415 35832 36461
rect 35889 36415 35935 36461
rect 35992 36415 36038 36461
rect 36095 36415 36141 36461
rect 36198 36415 36244 36461
rect 36301 36415 36347 36461
rect 36854 36415 36900 36461
rect 36971 36415 37017 36461
rect 37088 36415 37134 36461
rect 37206 36415 37252 36461
rect 37324 36415 37370 36461
rect 37442 36415 37488 36461
rect 48778 36415 48824 36461
rect 48881 36415 48927 36461
rect 48984 36415 49030 36461
rect 49087 36415 49133 36461
rect 49190 36415 49236 36461
rect 49293 36415 49339 36461
rect 49396 36415 49442 36461
rect 49499 36415 49545 36461
rect 49602 36415 49852 36461
rect 44812 36328 44858 36374
rect 44925 36328 44971 36374
rect 45038 36328 45084 36374
rect 45151 36328 45197 36374
rect 45264 36328 45310 36374
rect 31349 36104 33323 36150
rect 51802 36552 53776 36598
rect 51802 36328 53776 36374
rect 44812 36104 44858 36150
rect 44925 36104 44971 36150
rect 45038 36104 45084 36150
rect 45151 36104 45197 36150
rect 45264 36104 45310 36150
rect 51802 36104 53776 36150
rect 54793 36104 54839 36150
rect 54956 36104 55002 36150
rect 55118 36104 55164 36150
rect 55279 36104 55325 36150
rect 55439 36104 55485 36150
rect 55599 36104 55645 36150
rect 55760 36104 55806 36150
<< mvpsubdiff >>
rect 352 46083 86098 46102
rect 352 46037 371 46083
rect 417 46037 495 46083
rect 541 46037 619 46083
rect 665 46037 743 46083
rect 789 46037 867 46083
rect 913 46037 991 46083
rect 1037 46037 1115 46083
rect 1161 46037 1239 46083
rect 1285 46037 1363 46083
rect 1409 46037 1487 46083
rect 1533 46037 1611 46083
rect 1657 46037 1735 46083
rect 1781 46037 1859 46083
rect 1905 46037 1983 46083
rect 2029 46037 2107 46083
rect 2153 46037 2231 46083
rect 2277 46037 2355 46083
rect 2401 46037 2479 46083
rect 2525 46037 2603 46083
rect 2649 46037 2727 46083
rect 2773 46037 2851 46083
rect 2897 46037 2975 46083
rect 3021 46037 3099 46083
rect 3145 46037 3223 46083
rect 3269 46037 3347 46083
rect 3393 46037 3471 46083
rect 3517 46037 3595 46083
rect 3641 46037 3719 46083
rect 3765 46037 3843 46083
rect 3889 46037 3967 46083
rect 4013 46037 4091 46083
rect 4137 46037 4215 46083
rect 4261 46037 4339 46083
rect 4385 46037 4463 46083
rect 4509 46037 4587 46083
rect 4633 46037 4711 46083
rect 4757 46037 4835 46083
rect 4881 46037 4959 46083
rect 5005 46037 5083 46083
rect 5129 46037 5207 46083
rect 5253 46037 5331 46083
rect 5377 46037 5455 46083
rect 5501 46037 5579 46083
rect 5625 46037 5703 46083
rect 5749 46037 5827 46083
rect 5873 46037 5951 46083
rect 5997 46037 6075 46083
rect 6121 46037 6199 46083
rect 6245 46037 6323 46083
rect 6369 46037 6447 46083
rect 6493 46037 6571 46083
rect 6617 46037 6695 46083
rect 6741 46037 6819 46083
rect 6865 46037 6943 46083
rect 6989 46037 7067 46083
rect 7113 46037 7191 46083
rect 7237 46037 7315 46083
rect 7361 46037 7439 46083
rect 7485 46037 7563 46083
rect 7609 46037 7687 46083
rect 7733 46037 7811 46083
rect 7857 46037 7935 46083
rect 7981 46037 8059 46083
rect 8105 46037 8183 46083
rect 8229 46037 8307 46083
rect 8353 46037 8431 46083
rect 8477 46037 8555 46083
rect 8601 46037 8679 46083
rect 8725 46037 8803 46083
rect 8849 46037 8927 46083
rect 8973 46037 9051 46083
rect 9097 46037 9175 46083
rect 9221 46037 9299 46083
rect 9345 46037 9423 46083
rect 9469 46037 9547 46083
rect 9593 46037 9671 46083
rect 9717 46037 9795 46083
rect 9841 46037 9919 46083
rect 9965 46037 10043 46083
rect 10089 46037 10167 46083
rect 10213 46037 10291 46083
rect 10337 46037 10415 46083
rect 10461 46037 10539 46083
rect 10585 46037 10663 46083
rect 10709 46037 10787 46083
rect 10833 46037 10911 46083
rect 10957 46037 11035 46083
rect 11081 46037 11159 46083
rect 11205 46037 11283 46083
rect 11329 46037 11407 46083
rect 11453 46037 11531 46083
rect 11577 46037 11655 46083
rect 11701 46037 11779 46083
rect 11825 46037 11903 46083
rect 11949 46037 12027 46083
rect 12073 46037 12151 46083
rect 12197 46037 12275 46083
rect 12321 46037 12399 46083
rect 12445 46037 12523 46083
rect 12569 46037 12647 46083
rect 12693 46037 12771 46083
rect 12817 46037 12895 46083
rect 12941 46037 13019 46083
rect 13065 46037 13143 46083
rect 13189 46037 13267 46083
rect 13313 46037 13391 46083
rect 13437 46037 13515 46083
rect 13561 46037 13639 46083
rect 13685 46037 13763 46083
rect 13809 46037 13887 46083
rect 13933 46037 14011 46083
rect 14057 46037 14135 46083
rect 14181 46037 14259 46083
rect 14305 46037 14383 46083
rect 14429 46037 14507 46083
rect 14553 46037 14631 46083
rect 14677 46037 14755 46083
rect 14801 46037 14879 46083
rect 14925 46037 15003 46083
rect 15049 46037 15127 46083
rect 15173 46037 15251 46083
rect 15297 46037 15375 46083
rect 15421 46037 15499 46083
rect 15545 46037 15623 46083
rect 15669 46037 15747 46083
rect 15793 46037 15871 46083
rect 15917 46037 15995 46083
rect 16041 46037 16119 46083
rect 16165 46037 16243 46083
rect 16289 46037 16367 46083
rect 16413 46037 16491 46083
rect 16537 46037 16615 46083
rect 16661 46037 16739 46083
rect 16785 46037 16863 46083
rect 16909 46037 16987 46083
rect 17033 46037 17111 46083
rect 17157 46037 17235 46083
rect 17281 46037 17359 46083
rect 17405 46037 17483 46083
rect 17529 46037 17607 46083
rect 17653 46037 17731 46083
rect 17777 46037 17855 46083
rect 17901 46037 17979 46083
rect 18025 46037 18103 46083
rect 18149 46037 18227 46083
rect 18273 46037 18351 46083
rect 18397 46037 18475 46083
rect 18521 46037 18599 46083
rect 18645 46037 18723 46083
rect 18769 46037 18847 46083
rect 18893 46037 18971 46083
rect 19017 46037 19095 46083
rect 19141 46037 19219 46083
rect 19265 46037 19343 46083
rect 19389 46037 19467 46083
rect 19513 46037 19591 46083
rect 19637 46037 19715 46083
rect 19761 46037 19839 46083
rect 19885 46037 19963 46083
rect 20009 46037 20087 46083
rect 20133 46037 20211 46083
rect 20257 46037 20335 46083
rect 20381 46037 20459 46083
rect 20505 46037 20583 46083
rect 20629 46037 20707 46083
rect 20753 46037 20831 46083
rect 20877 46037 20955 46083
rect 21001 46037 21079 46083
rect 21125 46037 21203 46083
rect 21249 46037 21327 46083
rect 21373 46037 21451 46083
rect 21497 46037 21575 46083
rect 21621 46037 21699 46083
rect 21745 46037 21823 46083
rect 21869 46037 21947 46083
rect 21993 46037 22071 46083
rect 22117 46037 22195 46083
rect 22241 46037 22319 46083
rect 22365 46037 22443 46083
rect 22489 46037 22567 46083
rect 22613 46037 22691 46083
rect 22737 46037 22815 46083
rect 22861 46037 22939 46083
rect 22985 46037 23063 46083
rect 23109 46037 23187 46083
rect 23233 46037 23311 46083
rect 23357 46037 23435 46083
rect 23481 46037 23559 46083
rect 23605 46037 23683 46083
rect 23729 46037 23807 46083
rect 23853 46037 23931 46083
rect 23977 46037 24055 46083
rect 24101 46037 24179 46083
rect 24225 46037 24303 46083
rect 24349 46037 24427 46083
rect 24473 46037 24551 46083
rect 24597 46037 24675 46083
rect 24721 46037 24799 46083
rect 24845 46037 24923 46083
rect 24969 46037 25047 46083
rect 25093 46037 25171 46083
rect 25217 46037 25295 46083
rect 25341 46037 25419 46083
rect 25465 46037 25543 46083
rect 25589 46037 25667 46083
rect 25713 46037 25791 46083
rect 25837 46037 25915 46083
rect 25961 46037 26039 46083
rect 26085 46037 26163 46083
rect 26209 46037 26287 46083
rect 26333 46037 26411 46083
rect 26457 46037 26535 46083
rect 26581 46037 26659 46083
rect 26705 46037 26783 46083
rect 26829 46037 26907 46083
rect 26953 46037 27031 46083
rect 27077 46037 27155 46083
rect 27201 46037 27279 46083
rect 27325 46037 27403 46083
rect 27449 46037 27527 46083
rect 27573 46037 27651 46083
rect 27697 46037 27775 46083
rect 27821 46037 27899 46083
rect 27945 46037 28023 46083
rect 28069 46037 28147 46083
rect 28193 46037 28271 46083
rect 28317 46037 28395 46083
rect 28441 46037 28519 46083
rect 28565 46037 28643 46083
rect 28689 46037 28767 46083
rect 28813 46037 28891 46083
rect 28937 46037 29015 46083
rect 29061 46037 29139 46083
rect 29185 46037 29263 46083
rect 29309 46037 29387 46083
rect 29433 46037 29511 46083
rect 29557 46037 29635 46083
rect 29681 46037 29759 46083
rect 29805 46037 29883 46083
rect 29929 46037 30007 46083
rect 30053 46037 30131 46083
rect 30177 46037 30255 46083
rect 30301 46037 30379 46083
rect 30425 46037 30503 46083
rect 30549 46037 30627 46083
rect 30673 46037 30751 46083
rect 30797 46037 30875 46083
rect 30921 46037 30999 46083
rect 31045 46037 31123 46083
rect 31169 46037 31247 46083
rect 31293 46037 31371 46083
rect 31417 46037 31495 46083
rect 31541 46037 31619 46083
rect 31665 46037 31743 46083
rect 31789 46037 31867 46083
rect 31913 46037 31991 46083
rect 32037 46037 32115 46083
rect 32161 46037 32239 46083
rect 32285 46037 32363 46083
rect 32409 46037 32487 46083
rect 32533 46037 32611 46083
rect 32657 46037 32735 46083
rect 32781 46037 32859 46083
rect 32905 46037 32983 46083
rect 33029 46037 33107 46083
rect 33153 46037 33231 46083
rect 33277 46037 33355 46083
rect 33401 46037 33479 46083
rect 33525 46037 33603 46083
rect 33649 46037 33727 46083
rect 33773 46037 33851 46083
rect 33897 46037 33975 46083
rect 34021 46037 34099 46083
rect 34145 46037 34223 46083
rect 34269 46037 34347 46083
rect 34393 46037 34471 46083
rect 34517 46037 34595 46083
rect 34641 46037 34719 46083
rect 34765 46037 34843 46083
rect 34889 46037 34967 46083
rect 35013 46037 35091 46083
rect 35137 46037 35215 46083
rect 35261 46037 35339 46083
rect 35385 46037 35463 46083
rect 35509 46037 35587 46083
rect 35633 46037 35711 46083
rect 35757 46037 35835 46083
rect 35881 46037 35959 46083
rect 36005 46037 36083 46083
rect 36129 46037 36207 46083
rect 36253 46037 36331 46083
rect 36377 46037 36455 46083
rect 36501 46037 36579 46083
rect 36625 46037 36703 46083
rect 36749 46037 36827 46083
rect 36873 46037 36951 46083
rect 36997 46037 37075 46083
rect 37121 46037 37199 46083
rect 37245 46037 37323 46083
rect 37369 46037 37447 46083
rect 37493 46037 37571 46083
rect 37617 46037 37695 46083
rect 37741 46037 37819 46083
rect 37865 46037 37943 46083
rect 37989 46037 38067 46083
rect 38113 46037 38191 46083
rect 38237 46037 38315 46083
rect 38361 46037 38439 46083
rect 38485 46037 38563 46083
rect 38609 46037 38687 46083
rect 38733 46037 38811 46083
rect 38857 46037 38935 46083
rect 38981 46037 39059 46083
rect 39105 46037 39183 46083
rect 39229 46037 39307 46083
rect 39353 46037 39431 46083
rect 39477 46037 39555 46083
rect 39601 46037 39679 46083
rect 39725 46037 39803 46083
rect 39849 46037 39927 46083
rect 39973 46037 40051 46083
rect 40097 46037 40175 46083
rect 40221 46037 40299 46083
rect 40345 46037 40423 46083
rect 40469 46037 40547 46083
rect 40593 46037 40671 46083
rect 40717 46037 40795 46083
rect 40841 46037 40919 46083
rect 40965 46037 41043 46083
rect 41089 46037 41167 46083
rect 41213 46037 41291 46083
rect 41337 46037 41415 46083
rect 41461 46037 41539 46083
rect 41585 46037 41663 46083
rect 41709 46037 41787 46083
rect 41833 46037 41911 46083
rect 41957 46037 42035 46083
rect 42081 46037 42159 46083
rect 42205 46037 42283 46083
rect 42329 46037 42407 46083
rect 42453 46037 42531 46083
rect 42577 46037 42655 46083
rect 42701 46037 42779 46083
rect 42825 46037 42903 46083
rect 42949 46037 43027 46083
rect 43073 46037 43151 46083
rect 43197 46037 43275 46083
rect 43321 46037 43399 46083
rect 43445 46037 43523 46083
rect 43569 46037 43647 46083
rect 43693 46037 43771 46083
rect 43817 46037 43895 46083
rect 43941 46037 44019 46083
rect 44065 46037 44143 46083
rect 44189 46037 44267 46083
rect 44313 46037 44391 46083
rect 44437 46037 44515 46083
rect 44561 46037 44639 46083
rect 44685 46037 44763 46083
rect 44809 46037 44887 46083
rect 44933 46037 45011 46083
rect 45057 46037 45135 46083
rect 45181 46037 45259 46083
rect 45305 46037 45383 46083
rect 45429 46037 45507 46083
rect 45553 46037 45631 46083
rect 45677 46037 45755 46083
rect 45801 46037 45879 46083
rect 45925 46037 46003 46083
rect 46049 46037 46127 46083
rect 46173 46037 46251 46083
rect 46297 46037 46375 46083
rect 46421 46037 46499 46083
rect 46545 46037 46623 46083
rect 46669 46037 46747 46083
rect 46793 46037 46871 46083
rect 46917 46037 46995 46083
rect 47041 46037 47119 46083
rect 47165 46037 47243 46083
rect 47289 46037 47367 46083
rect 47413 46037 47491 46083
rect 47537 46037 47615 46083
rect 47661 46037 47739 46083
rect 47785 46037 47863 46083
rect 47909 46037 47987 46083
rect 48033 46037 48111 46083
rect 48157 46037 48235 46083
rect 48281 46037 48359 46083
rect 48405 46037 48483 46083
rect 48529 46037 48607 46083
rect 48653 46037 48731 46083
rect 48777 46037 48855 46083
rect 48901 46037 48979 46083
rect 49025 46037 49103 46083
rect 49149 46037 49227 46083
rect 49273 46037 49351 46083
rect 49397 46037 49475 46083
rect 49521 46037 49599 46083
rect 49645 46037 49723 46083
rect 49769 46037 49847 46083
rect 49893 46037 49971 46083
rect 50017 46037 50095 46083
rect 50141 46037 50219 46083
rect 50265 46037 50343 46083
rect 50389 46037 50467 46083
rect 50513 46037 50591 46083
rect 50637 46037 50715 46083
rect 50761 46037 50839 46083
rect 50885 46037 50963 46083
rect 51009 46037 51087 46083
rect 51133 46037 51211 46083
rect 51257 46037 51335 46083
rect 51381 46037 51459 46083
rect 51505 46037 51583 46083
rect 51629 46037 51707 46083
rect 51753 46037 51831 46083
rect 51877 46037 51955 46083
rect 52001 46037 52079 46083
rect 52125 46037 52203 46083
rect 52249 46037 52327 46083
rect 52373 46037 52451 46083
rect 52497 46037 52575 46083
rect 52621 46037 52699 46083
rect 52745 46037 52823 46083
rect 52869 46037 52947 46083
rect 52993 46037 53071 46083
rect 53117 46037 53195 46083
rect 53241 46037 53319 46083
rect 53365 46037 53443 46083
rect 53489 46037 53567 46083
rect 53613 46037 53691 46083
rect 53737 46037 53815 46083
rect 53861 46037 53939 46083
rect 53985 46037 54063 46083
rect 54109 46037 54187 46083
rect 54233 46037 54311 46083
rect 54357 46037 54435 46083
rect 54481 46037 54559 46083
rect 54605 46037 54683 46083
rect 54729 46037 54807 46083
rect 54853 46037 54931 46083
rect 54977 46037 55055 46083
rect 55101 46037 55179 46083
rect 55225 46037 55303 46083
rect 55349 46037 55427 46083
rect 55473 46037 55551 46083
rect 55597 46037 55675 46083
rect 55721 46037 55799 46083
rect 55845 46037 55923 46083
rect 55969 46037 56047 46083
rect 56093 46037 56171 46083
rect 56217 46037 56295 46083
rect 56341 46037 56419 46083
rect 56465 46037 56543 46083
rect 56589 46037 56667 46083
rect 56713 46037 56791 46083
rect 56837 46037 56915 46083
rect 56961 46037 57039 46083
rect 57085 46037 57163 46083
rect 57209 46037 57287 46083
rect 57333 46037 57411 46083
rect 57457 46037 57535 46083
rect 57581 46037 57659 46083
rect 57705 46037 57783 46083
rect 57829 46037 57907 46083
rect 57953 46037 58031 46083
rect 58077 46037 58155 46083
rect 58201 46037 58279 46083
rect 58325 46037 58403 46083
rect 58449 46037 58527 46083
rect 58573 46037 58651 46083
rect 58697 46037 58775 46083
rect 58821 46037 58899 46083
rect 58945 46037 59023 46083
rect 59069 46037 59147 46083
rect 59193 46037 59271 46083
rect 59317 46037 59395 46083
rect 59441 46037 59519 46083
rect 59565 46037 59643 46083
rect 59689 46037 59767 46083
rect 59813 46037 59891 46083
rect 59937 46037 60015 46083
rect 60061 46037 60139 46083
rect 60185 46037 60263 46083
rect 60309 46037 60387 46083
rect 60433 46037 60511 46083
rect 60557 46037 60635 46083
rect 60681 46037 60759 46083
rect 60805 46037 60883 46083
rect 60929 46037 61007 46083
rect 61053 46037 61131 46083
rect 61177 46037 61255 46083
rect 61301 46037 61379 46083
rect 61425 46037 61503 46083
rect 61549 46037 61627 46083
rect 61673 46037 61751 46083
rect 61797 46037 61875 46083
rect 61921 46037 61999 46083
rect 62045 46037 62123 46083
rect 62169 46037 62247 46083
rect 62293 46037 62371 46083
rect 62417 46037 62495 46083
rect 62541 46037 62619 46083
rect 62665 46037 62743 46083
rect 62789 46037 62867 46083
rect 62913 46037 62991 46083
rect 63037 46037 63115 46083
rect 63161 46037 63239 46083
rect 63285 46037 63363 46083
rect 63409 46037 63487 46083
rect 63533 46037 63611 46083
rect 63657 46037 63735 46083
rect 63781 46037 63859 46083
rect 63905 46037 63983 46083
rect 64029 46037 64107 46083
rect 64153 46037 64231 46083
rect 64277 46037 64355 46083
rect 64401 46037 64479 46083
rect 64525 46037 64603 46083
rect 64649 46037 64727 46083
rect 64773 46037 64851 46083
rect 64897 46037 64975 46083
rect 65021 46037 65099 46083
rect 65145 46037 65223 46083
rect 65269 46037 65347 46083
rect 65393 46037 65471 46083
rect 65517 46037 65595 46083
rect 65641 46037 65719 46083
rect 65765 46037 65843 46083
rect 65889 46037 65967 46083
rect 66013 46037 66091 46083
rect 66137 46037 66215 46083
rect 66261 46037 66339 46083
rect 66385 46037 66463 46083
rect 66509 46037 66587 46083
rect 66633 46037 66711 46083
rect 66757 46037 66835 46083
rect 66881 46037 66959 46083
rect 67005 46037 67083 46083
rect 67129 46037 67207 46083
rect 67253 46037 67331 46083
rect 67377 46037 67455 46083
rect 67501 46037 67579 46083
rect 67625 46037 67703 46083
rect 67749 46037 67827 46083
rect 67873 46037 67951 46083
rect 67997 46037 68075 46083
rect 68121 46037 68199 46083
rect 68245 46037 68323 46083
rect 68369 46037 68447 46083
rect 68493 46037 68571 46083
rect 68617 46037 68695 46083
rect 68741 46037 68819 46083
rect 68865 46037 68943 46083
rect 68989 46037 69067 46083
rect 69113 46037 69191 46083
rect 69237 46037 69315 46083
rect 69361 46037 69439 46083
rect 69485 46037 69563 46083
rect 69609 46037 69687 46083
rect 69733 46037 69811 46083
rect 69857 46037 69935 46083
rect 69981 46037 70059 46083
rect 70105 46037 70183 46083
rect 70229 46037 70307 46083
rect 70353 46037 70431 46083
rect 70477 46037 70555 46083
rect 70601 46037 70679 46083
rect 70725 46037 70803 46083
rect 70849 46037 70927 46083
rect 70973 46037 71051 46083
rect 71097 46037 71175 46083
rect 71221 46037 71299 46083
rect 71345 46037 71423 46083
rect 71469 46037 71547 46083
rect 71593 46037 71671 46083
rect 71717 46037 71795 46083
rect 71841 46037 71919 46083
rect 71965 46037 72043 46083
rect 72089 46037 72167 46083
rect 72213 46037 72291 46083
rect 72337 46037 72415 46083
rect 72461 46037 72539 46083
rect 72585 46037 72663 46083
rect 72709 46037 72787 46083
rect 72833 46037 72911 46083
rect 72957 46037 73035 46083
rect 73081 46037 73159 46083
rect 73205 46037 73283 46083
rect 73329 46037 73407 46083
rect 73453 46037 73531 46083
rect 73577 46037 73655 46083
rect 73701 46037 73779 46083
rect 73825 46037 73903 46083
rect 73949 46037 74027 46083
rect 74073 46037 74151 46083
rect 74197 46037 74275 46083
rect 74321 46037 74399 46083
rect 74445 46037 74523 46083
rect 74569 46037 74647 46083
rect 74693 46037 74771 46083
rect 74817 46037 74895 46083
rect 74941 46037 75019 46083
rect 75065 46037 75143 46083
rect 75189 46037 75267 46083
rect 75313 46037 75391 46083
rect 75437 46037 75515 46083
rect 75561 46037 75639 46083
rect 75685 46037 75763 46083
rect 75809 46037 75887 46083
rect 75933 46037 76011 46083
rect 76057 46037 76135 46083
rect 76181 46037 76259 46083
rect 76305 46037 76383 46083
rect 76429 46037 76507 46083
rect 76553 46037 76631 46083
rect 76677 46037 76755 46083
rect 76801 46037 76879 46083
rect 76925 46037 77003 46083
rect 77049 46037 77127 46083
rect 77173 46037 77251 46083
rect 77297 46037 77375 46083
rect 77421 46037 77499 46083
rect 77545 46037 77623 46083
rect 77669 46037 77747 46083
rect 77793 46037 77871 46083
rect 77917 46037 77995 46083
rect 78041 46037 78119 46083
rect 78165 46037 78243 46083
rect 78289 46037 78367 46083
rect 78413 46037 78491 46083
rect 78537 46037 78615 46083
rect 78661 46037 78739 46083
rect 78785 46037 78863 46083
rect 78909 46037 78987 46083
rect 79033 46037 79111 46083
rect 79157 46037 79235 46083
rect 79281 46037 79359 46083
rect 79405 46037 79483 46083
rect 79529 46037 79607 46083
rect 79653 46037 79731 46083
rect 79777 46037 79855 46083
rect 79901 46037 79979 46083
rect 80025 46037 80103 46083
rect 80149 46037 80227 46083
rect 80273 46037 80351 46083
rect 80397 46037 80475 46083
rect 80521 46037 80599 46083
rect 80645 46037 80723 46083
rect 80769 46037 80847 46083
rect 80893 46037 80971 46083
rect 81017 46037 81095 46083
rect 81141 46037 81219 46083
rect 81265 46037 81343 46083
rect 81389 46037 81467 46083
rect 81513 46037 81591 46083
rect 81637 46037 81715 46083
rect 81761 46037 81839 46083
rect 81885 46037 81963 46083
rect 82009 46037 82087 46083
rect 82133 46037 82211 46083
rect 82257 46037 82335 46083
rect 82381 46037 82459 46083
rect 82505 46037 82583 46083
rect 82629 46037 82707 46083
rect 82753 46037 82831 46083
rect 82877 46037 82955 46083
rect 83001 46037 83079 46083
rect 83125 46037 83203 46083
rect 83249 46037 83327 46083
rect 83373 46037 83451 46083
rect 83497 46037 83575 46083
rect 83621 46037 83699 46083
rect 83745 46037 83823 46083
rect 83869 46037 83947 46083
rect 83993 46037 84071 46083
rect 84117 46037 84195 46083
rect 84241 46037 84319 46083
rect 84365 46037 84443 46083
rect 84489 46037 84567 46083
rect 84613 46037 84691 46083
rect 84737 46037 84815 46083
rect 84861 46037 84939 46083
rect 84985 46037 85063 46083
rect 85109 46037 85187 46083
rect 85233 46037 85311 46083
rect 85357 46037 85435 46083
rect 85481 46037 85559 46083
rect 85605 46037 85683 46083
rect 85729 46037 85807 46083
rect 85853 46037 85931 46083
rect 85977 46037 86098 46083
rect 352 45959 86098 46037
rect 352 45913 371 45959
rect 417 45913 495 45959
rect 541 45913 619 45959
rect 665 45913 743 45959
rect 789 45913 867 45959
rect 913 45913 991 45959
rect 1037 45913 1115 45959
rect 1161 45913 1239 45959
rect 1285 45913 1363 45959
rect 1409 45913 1487 45959
rect 1533 45913 1611 45959
rect 1657 45913 1735 45959
rect 1781 45913 1859 45959
rect 1905 45913 1983 45959
rect 2029 45913 2107 45959
rect 2153 45913 2231 45959
rect 2277 45913 2355 45959
rect 2401 45913 2479 45959
rect 2525 45913 2603 45959
rect 2649 45913 2727 45959
rect 2773 45913 2851 45959
rect 2897 45913 2975 45959
rect 3021 45913 3099 45959
rect 3145 45913 3223 45959
rect 3269 45913 3347 45959
rect 3393 45913 3471 45959
rect 3517 45913 3595 45959
rect 3641 45913 3719 45959
rect 3765 45913 3843 45959
rect 3889 45913 3967 45959
rect 4013 45913 4091 45959
rect 4137 45913 4215 45959
rect 4261 45913 4339 45959
rect 4385 45913 4463 45959
rect 4509 45913 4587 45959
rect 4633 45913 4711 45959
rect 4757 45913 4835 45959
rect 4881 45913 4959 45959
rect 5005 45913 5083 45959
rect 5129 45913 5207 45959
rect 5253 45913 5331 45959
rect 5377 45913 5455 45959
rect 5501 45913 5579 45959
rect 5625 45913 5703 45959
rect 5749 45913 5827 45959
rect 5873 45913 5951 45959
rect 5997 45913 6075 45959
rect 6121 45913 6199 45959
rect 6245 45913 6323 45959
rect 6369 45913 6447 45959
rect 6493 45913 6571 45959
rect 6617 45913 6695 45959
rect 6741 45913 6819 45959
rect 6865 45913 6943 45959
rect 6989 45913 7067 45959
rect 7113 45913 7191 45959
rect 7237 45913 7315 45959
rect 7361 45913 7439 45959
rect 7485 45913 7563 45959
rect 7609 45913 7687 45959
rect 7733 45913 7811 45959
rect 7857 45913 7935 45959
rect 7981 45913 8059 45959
rect 8105 45913 8183 45959
rect 8229 45913 8307 45959
rect 8353 45913 8431 45959
rect 8477 45913 8555 45959
rect 8601 45913 8679 45959
rect 8725 45913 8803 45959
rect 8849 45913 8927 45959
rect 8973 45913 9051 45959
rect 9097 45913 9175 45959
rect 9221 45913 9299 45959
rect 9345 45913 9423 45959
rect 9469 45913 9547 45959
rect 9593 45913 9671 45959
rect 9717 45913 9795 45959
rect 9841 45913 9919 45959
rect 9965 45913 10043 45959
rect 10089 45913 10167 45959
rect 10213 45913 10291 45959
rect 10337 45913 10415 45959
rect 10461 45913 10539 45959
rect 10585 45913 10663 45959
rect 10709 45913 10787 45959
rect 10833 45913 10911 45959
rect 10957 45913 11035 45959
rect 11081 45913 11159 45959
rect 11205 45913 11283 45959
rect 11329 45913 11407 45959
rect 11453 45913 11531 45959
rect 11577 45913 11655 45959
rect 11701 45913 11779 45959
rect 11825 45913 11903 45959
rect 11949 45913 12027 45959
rect 12073 45913 12151 45959
rect 12197 45913 12275 45959
rect 12321 45913 12399 45959
rect 12445 45913 12523 45959
rect 12569 45913 12647 45959
rect 12693 45913 12771 45959
rect 12817 45913 12895 45959
rect 12941 45913 13019 45959
rect 13065 45913 13143 45959
rect 13189 45913 13267 45959
rect 13313 45913 13391 45959
rect 13437 45913 13515 45959
rect 13561 45913 13639 45959
rect 13685 45913 13763 45959
rect 13809 45913 13887 45959
rect 13933 45913 14011 45959
rect 14057 45913 14135 45959
rect 14181 45913 14259 45959
rect 14305 45913 14383 45959
rect 14429 45913 14507 45959
rect 14553 45913 14631 45959
rect 14677 45913 14755 45959
rect 14801 45913 14879 45959
rect 14925 45913 15003 45959
rect 15049 45913 15127 45959
rect 15173 45913 15251 45959
rect 15297 45913 15375 45959
rect 15421 45913 15499 45959
rect 15545 45913 15623 45959
rect 15669 45913 15747 45959
rect 15793 45913 15871 45959
rect 15917 45913 15995 45959
rect 16041 45913 16119 45959
rect 16165 45913 16243 45959
rect 16289 45913 16367 45959
rect 16413 45913 16491 45959
rect 16537 45913 16615 45959
rect 16661 45913 16739 45959
rect 16785 45913 16863 45959
rect 16909 45913 16987 45959
rect 17033 45913 17111 45959
rect 17157 45913 17235 45959
rect 17281 45913 17359 45959
rect 17405 45913 17483 45959
rect 17529 45913 17607 45959
rect 17653 45913 17731 45959
rect 17777 45913 17855 45959
rect 17901 45913 17979 45959
rect 18025 45913 18103 45959
rect 18149 45913 18227 45959
rect 18273 45913 18351 45959
rect 18397 45913 18475 45959
rect 18521 45913 18599 45959
rect 18645 45913 18723 45959
rect 18769 45913 18847 45959
rect 18893 45913 18971 45959
rect 19017 45913 19095 45959
rect 19141 45913 19219 45959
rect 19265 45913 19343 45959
rect 19389 45913 19467 45959
rect 19513 45913 19591 45959
rect 19637 45913 19715 45959
rect 19761 45913 19839 45959
rect 19885 45913 19963 45959
rect 20009 45913 20087 45959
rect 20133 45913 20211 45959
rect 20257 45913 20335 45959
rect 20381 45913 20459 45959
rect 20505 45913 20583 45959
rect 20629 45913 20707 45959
rect 20753 45913 20831 45959
rect 20877 45913 20955 45959
rect 21001 45913 21079 45959
rect 21125 45913 21203 45959
rect 21249 45913 21327 45959
rect 21373 45913 21451 45959
rect 21497 45913 21575 45959
rect 21621 45913 21699 45959
rect 21745 45913 21823 45959
rect 21869 45913 21947 45959
rect 21993 45913 22071 45959
rect 22117 45913 22195 45959
rect 22241 45913 22319 45959
rect 22365 45913 22443 45959
rect 22489 45913 22567 45959
rect 22613 45913 22691 45959
rect 22737 45913 22815 45959
rect 22861 45913 22939 45959
rect 22985 45913 23063 45959
rect 23109 45913 23187 45959
rect 23233 45913 23311 45959
rect 23357 45913 23435 45959
rect 23481 45913 23559 45959
rect 23605 45913 23683 45959
rect 23729 45913 23807 45959
rect 23853 45913 23931 45959
rect 23977 45913 24055 45959
rect 24101 45913 24179 45959
rect 24225 45913 24303 45959
rect 24349 45913 24427 45959
rect 24473 45913 24551 45959
rect 24597 45913 24675 45959
rect 24721 45913 24799 45959
rect 24845 45913 24923 45959
rect 24969 45913 25047 45959
rect 25093 45913 25171 45959
rect 25217 45913 25295 45959
rect 25341 45913 25419 45959
rect 25465 45913 25543 45959
rect 25589 45913 25667 45959
rect 25713 45913 25791 45959
rect 25837 45913 25915 45959
rect 25961 45913 26039 45959
rect 26085 45913 26163 45959
rect 26209 45913 26287 45959
rect 26333 45913 26411 45959
rect 26457 45913 26535 45959
rect 26581 45913 26659 45959
rect 26705 45913 26783 45959
rect 26829 45913 26907 45959
rect 26953 45913 27031 45959
rect 27077 45913 27155 45959
rect 27201 45913 27279 45959
rect 27325 45913 27403 45959
rect 27449 45913 27527 45959
rect 27573 45913 27651 45959
rect 27697 45913 27775 45959
rect 27821 45913 27899 45959
rect 27945 45913 28023 45959
rect 28069 45913 28147 45959
rect 28193 45913 28271 45959
rect 28317 45913 28395 45959
rect 28441 45913 28519 45959
rect 28565 45913 28643 45959
rect 28689 45913 28767 45959
rect 28813 45913 28891 45959
rect 28937 45913 29015 45959
rect 29061 45913 29139 45959
rect 29185 45913 29263 45959
rect 29309 45913 29387 45959
rect 29433 45913 29511 45959
rect 29557 45913 29635 45959
rect 29681 45913 29759 45959
rect 29805 45913 29883 45959
rect 29929 45913 30007 45959
rect 30053 45913 30131 45959
rect 30177 45913 30255 45959
rect 30301 45913 30379 45959
rect 30425 45913 30503 45959
rect 30549 45913 30627 45959
rect 30673 45913 30751 45959
rect 30797 45913 30875 45959
rect 30921 45913 30999 45959
rect 31045 45913 31123 45959
rect 31169 45913 31247 45959
rect 31293 45913 31371 45959
rect 31417 45913 31495 45959
rect 31541 45913 31619 45959
rect 31665 45913 31743 45959
rect 31789 45913 31867 45959
rect 31913 45913 31991 45959
rect 32037 45913 32115 45959
rect 32161 45913 32239 45959
rect 32285 45913 32363 45959
rect 32409 45913 32487 45959
rect 32533 45913 32611 45959
rect 32657 45913 32735 45959
rect 32781 45913 32859 45959
rect 32905 45913 32983 45959
rect 33029 45913 33107 45959
rect 33153 45913 33231 45959
rect 33277 45913 33355 45959
rect 33401 45913 33479 45959
rect 33525 45913 33603 45959
rect 33649 45913 33727 45959
rect 33773 45913 33851 45959
rect 33897 45913 33975 45959
rect 34021 45913 34099 45959
rect 34145 45913 34223 45959
rect 34269 45913 34347 45959
rect 34393 45913 34471 45959
rect 34517 45913 34595 45959
rect 34641 45913 34719 45959
rect 34765 45913 34843 45959
rect 34889 45913 34967 45959
rect 35013 45913 35091 45959
rect 35137 45913 35215 45959
rect 35261 45913 35339 45959
rect 35385 45913 35463 45959
rect 35509 45913 35587 45959
rect 35633 45913 35711 45959
rect 35757 45913 35835 45959
rect 35881 45913 35959 45959
rect 36005 45913 36083 45959
rect 36129 45913 36207 45959
rect 36253 45913 36331 45959
rect 36377 45913 36455 45959
rect 36501 45913 36579 45959
rect 36625 45913 36703 45959
rect 36749 45913 36827 45959
rect 36873 45913 36951 45959
rect 36997 45913 37075 45959
rect 37121 45913 37199 45959
rect 37245 45913 37323 45959
rect 37369 45913 37447 45959
rect 37493 45913 37571 45959
rect 37617 45913 37695 45959
rect 37741 45913 37819 45959
rect 37865 45913 37943 45959
rect 37989 45913 38067 45959
rect 38113 45913 38191 45959
rect 38237 45913 38315 45959
rect 38361 45913 38439 45959
rect 38485 45913 38563 45959
rect 38609 45913 38687 45959
rect 38733 45913 38811 45959
rect 38857 45913 38935 45959
rect 38981 45913 39059 45959
rect 39105 45913 39183 45959
rect 39229 45913 39307 45959
rect 39353 45913 39431 45959
rect 39477 45913 39555 45959
rect 39601 45913 39679 45959
rect 39725 45913 39803 45959
rect 39849 45913 39927 45959
rect 39973 45913 40051 45959
rect 40097 45913 40175 45959
rect 40221 45913 40299 45959
rect 40345 45913 40423 45959
rect 40469 45913 40547 45959
rect 40593 45913 40671 45959
rect 40717 45913 40795 45959
rect 40841 45913 40919 45959
rect 40965 45913 41043 45959
rect 41089 45913 41167 45959
rect 41213 45913 41291 45959
rect 41337 45913 41415 45959
rect 41461 45913 41539 45959
rect 41585 45913 41663 45959
rect 41709 45913 41787 45959
rect 41833 45913 41911 45959
rect 41957 45913 42035 45959
rect 42081 45913 42159 45959
rect 42205 45913 42283 45959
rect 42329 45913 42407 45959
rect 42453 45913 42531 45959
rect 42577 45913 42655 45959
rect 42701 45913 42779 45959
rect 42825 45913 42903 45959
rect 42949 45913 43027 45959
rect 43073 45913 43151 45959
rect 43197 45913 43275 45959
rect 43321 45913 43399 45959
rect 43445 45913 43523 45959
rect 43569 45913 43647 45959
rect 43693 45913 43771 45959
rect 43817 45913 43895 45959
rect 43941 45913 44019 45959
rect 44065 45913 44143 45959
rect 44189 45913 44267 45959
rect 44313 45913 44391 45959
rect 44437 45913 44515 45959
rect 44561 45913 44639 45959
rect 44685 45913 44763 45959
rect 44809 45913 44887 45959
rect 44933 45913 45011 45959
rect 45057 45913 45135 45959
rect 45181 45913 45259 45959
rect 45305 45913 45383 45959
rect 45429 45913 45507 45959
rect 45553 45913 45631 45959
rect 45677 45913 45755 45959
rect 45801 45913 45879 45959
rect 45925 45913 46003 45959
rect 46049 45913 46127 45959
rect 46173 45913 46251 45959
rect 46297 45913 46375 45959
rect 46421 45913 46499 45959
rect 46545 45913 46623 45959
rect 46669 45913 46747 45959
rect 46793 45913 46871 45959
rect 46917 45913 46995 45959
rect 47041 45913 47119 45959
rect 47165 45913 47243 45959
rect 47289 45913 47367 45959
rect 47413 45913 47491 45959
rect 47537 45913 47615 45959
rect 47661 45913 47739 45959
rect 47785 45913 47863 45959
rect 47909 45913 47987 45959
rect 48033 45913 48111 45959
rect 48157 45913 48235 45959
rect 48281 45913 48359 45959
rect 48405 45913 48483 45959
rect 48529 45913 48607 45959
rect 48653 45913 48731 45959
rect 48777 45913 48855 45959
rect 48901 45913 48979 45959
rect 49025 45913 49103 45959
rect 49149 45913 49227 45959
rect 49273 45913 49351 45959
rect 49397 45913 49475 45959
rect 49521 45913 49599 45959
rect 49645 45913 49723 45959
rect 49769 45913 49847 45959
rect 49893 45913 49971 45959
rect 50017 45913 50095 45959
rect 50141 45913 50219 45959
rect 50265 45913 50343 45959
rect 50389 45913 50467 45959
rect 50513 45913 50591 45959
rect 50637 45913 50715 45959
rect 50761 45913 50839 45959
rect 50885 45913 50963 45959
rect 51009 45913 51087 45959
rect 51133 45913 51211 45959
rect 51257 45913 51335 45959
rect 51381 45913 51459 45959
rect 51505 45913 51583 45959
rect 51629 45913 51707 45959
rect 51753 45913 51831 45959
rect 51877 45913 51955 45959
rect 52001 45913 52079 45959
rect 52125 45913 52203 45959
rect 52249 45913 52327 45959
rect 52373 45913 52451 45959
rect 52497 45913 52575 45959
rect 52621 45913 52699 45959
rect 52745 45913 52823 45959
rect 52869 45913 52947 45959
rect 52993 45913 53071 45959
rect 53117 45913 53195 45959
rect 53241 45913 53319 45959
rect 53365 45913 53443 45959
rect 53489 45913 53567 45959
rect 53613 45913 53691 45959
rect 53737 45913 53815 45959
rect 53861 45913 53939 45959
rect 53985 45913 54063 45959
rect 54109 45913 54187 45959
rect 54233 45913 54311 45959
rect 54357 45913 54435 45959
rect 54481 45913 54559 45959
rect 54605 45913 54683 45959
rect 54729 45913 54807 45959
rect 54853 45913 54931 45959
rect 54977 45913 55055 45959
rect 55101 45913 55179 45959
rect 55225 45913 55303 45959
rect 55349 45913 55427 45959
rect 55473 45913 55551 45959
rect 55597 45913 55675 45959
rect 55721 45913 55799 45959
rect 55845 45913 55923 45959
rect 55969 45913 56047 45959
rect 56093 45913 56171 45959
rect 56217 45913 56295 45959
rect 56341 45913 56419 45959
rect 56465 45913 56543 45959
rect 56589 45913 56667 45959
rect 56713 45913 56791 45959
rect 56837 45913 56915 45959
rect 56961 45913 57039 45959
rect 57085 45913 57163 45959
rect 57209 45913 57287 45959
rect 57333 45913 57411 45959
rect 57457 45913 57535 45959
rect 57581 45913 57659 45959
rect 57705 45913 57783 45959
rect 57829 45913 57907 45959
rect 57953 45913 58031 45959
rect 58077 45913 58155 45959
rect 58201 45913 58279 45959
rect 58325 45913 58403 45959
rect 58449 45913 58527 45959
rect 58573 45913 58651 45959
rect 58697 45913 58775 45959
rect 58821 45913 58899 45959
rect 58945 45913 59023 45959
rect 59069 45913 59147 45959
rect 59193 45913 59271 45959
rect 59317 45913 59395 45959
rect 59441 45913 59519 45959
rect 59565 45913 59643 45959
rect 59689 45913 59767 45959
rect 59813 45913 59891 45959
rect 59937 45913 60015 45959
rect 60061 45913 60139 45959
rect 60185 45913 60263 45959
rect 60309 45913 60387 45959
rect 60433 45913 60511 45959
rect 60557 45913 60635 45959
rect 60681 45913 60759 45959
rect 60805 45913 60883 45959
rect 60929 45913 61007 45959
rect 61053 45913 61131 45959
rect 61177 45913 61255 45959
rect 61301 45913 61379 45959
rect 61425 45913 61503 45959
rect 61549 45913 61627 45959
rect 61673 45913 61751 45959
rect 61797 45913 61875 45959
rect 61921 45913 61999 45959
rect 62045 45913 62123 45959
rect 62169 45913 62247 45959
rect 62293 45913 62371 45959
rect 62417 45913 62495 45959
rect 62541 45913 62619 45959
rect 62665 45913 62743 45959
rect 62789 45913 62867 45959
rect 62913 45913 62991 45959
rect 63037 45913 63115 45959
rect 63161 45913 63239 45959
rect 63285 45913 63363 45959
rect 63409 45913 63487 45959
rect 63533 45913 63611 45959
rect 63657 45913 63735 45959
rect 63781 45913 63859 45959
rect 63905 45913 63983 45959
rect 64029 45913 64107 45959
rect 64153 45913 64231 45959
rect 64277 45913 64355 45959
rect 64401 45913 64479 45959
rect 64525 45913 64603 45959
rect 64649 45913 64727 45959
rect 64773 45913 64851 45959
rect 64897 45913 64975 45959
rect 65021 45913 65099 45959
rect 65145 45913 65223 45959
rect 65269 45913 65347 45959
rect 65393 45913 65471 45959
rect 65517 45913 65595 45959
rect 65641 45913 65719 45959
rect 65765 45913 65843 45959
rect 65889 45913 65967 45959
rect 66013 45913 66091 45959
rect 66137 45913 66215 45959
rect 66261 45913 66339 45959
rect 66385 45913 66463 45959
rect 66509 45913 66587 45959
rect 66633 45913 66711 45959
rect 66757 45913 66835 45959
rect 66881 45913 66959 45959
rect 67005 45913 67083 45959
rect 67129 45913 67207 45959
rect 67253 45913 67331 45959
rect 67377 45913 67455 45959
rect 67501 45913 67579 45959
rect 67625 45913 67703 45959
rect 67749 45913 67827 45959
rect 67873 45913 67951 45959
rect 67997 45913 68075 45959
rect 68121 45913 68199 45959
rect 68245 45913 68323 45959
rect 68369 45913 68447 45959
rect 68493 45913 68571 45959
rect 68617 45913 68695 45959
rect 68741 45913 68819 45959
rect 68865 45913 68943 45959
rect 68989 45913 69067 45959
rect 69113 45913 69191 45959
rect 69237 45913 69315 45959
rect 69361 45913 69439 45959
rect 69485 45913 69563 45959
rect 69609 45913 69687 45959
rect 69733 45913 69811 45959
rect 69857 45913 69935 45959
rect 69981 45913 70059 45959
rect 70105 45913 70183 45959
rect 70229 45913 70307 45959
rect 70353 45913 70431 45959
rect 70477 45913 70555 45959
rect 70601 45913 70679 45959
rect 70725 45913 70803 45959
rect 70849 45913 70927 45959
rect 70973 45913 71051 45959
rect 71097 45913 71175 45959
rect 71221 45913 71299 45959
rect 71345 45913 71423 45959
rect 71469 45913 71547 45959
rect 71593 45913 71671 45959
rect 71717 45913 71795 45959
rect 71841 45913 71919 45959
rect 71965 45913 72043 45959
rect 72089 45913 72167 45959
rect 72213 45913 72291 45959
rect 72337 45913 72415 45959
rect 72461 45913 72539 45959
rect 72585 45913 72663 45959
rect 72709 45913 72787 45959
rect 72833 45913 72911 45959
rect 72957 45913 73035 45959
rect 73081 45913 73159 45959
rect 73205 45913 73283 45959
rect 73329 45913 73407 45959
rect 73453 45913 73531 45959
rect 73577 45913 73655 45959
rect 73701 45913 73779 45959
rect 73825 45913 73903 45959
rect 73949 45913 74027 45959
rect 74073 45913 74151 45959
rect 74197 45913 74275 45959
rect 74321 45913 74399 45959
rect 74445 45913 74523 45959
rect 74569 45913 74647 45959
rect 74693 45913 74771 45959
rect 74817 45913 74895 45959
rect 74941 45913 75019 45959
rect 75065 45913 75143 45959
rect 75189 45913 75267 45959
rect 75313 45913 75391 45959
rect 75437 45913 75515 45959
rect 75561 45913 75639 45959
rect 75685 45913 75763 45959
rect 75809 45913 75887 45959
rect 75933 45913 76011 45959
rect 76057 45913 76135 45959
rect 76181 45913 76259 45959
rect 76305 45913 76383 45959
rect 76429 45913 76507 45959
rect 76553 45913 76631 45959
rect 76677 45913 76755 45959
rect 76801 45913 76879 45959
rect 76925 45913 77003 45959
rect 77049 45913 77127 45959
rect 77173 45913 77251 45959
rect 77297 45913 77375 45959
rect 77421 45913 77499 45959
rect 77545 45913 77623 45959
rect 77669 45913 77747 45959
rect 77793 45913 77871 45959
rect 77917 45913 77995 45959
rect 78041 45913 78119 45959
rect 78165 45913 78243 45959
rect 78289 45913 78367 45959
rect 78413 45913 78491 45959
rect 78537 45913 78615 45959
rect 78661 45913 78739 45959
rect 78785 45913 78863 45959
rect 78909 45913 78987 45959
rect 79033 45913 79111 45959
rect 79157 45913 79235 45959
rect 79281 45913 79359 45959
rect 79405 45913 79483 45959
rect 79529 45913 79607 45959
rect 79653 45913 79731 45959
rect 79777 45913 79855 45959
rect 79901 45913 79979 45959
rect 80025 45913 80103 45959
rect 80149 45913 80227 45959
rect 80273 45913 80351 45959
rect 80397 45913 80475 45959
rect 80521 45913 80599 45959
rect 80645 45913 80723 45959
rect 80769 45913 80847 45959
rect 80893 45913 80971 45959
rect 81017 45913 81095 45959
rect 81141 45913 81219 45959
rect 81265 45913 81343 45959
rect 81389 45913 81467 45959
rect 81513 45913 81591 45959
rect 81637 45913 81715 45959
rect 81761 45913 81839 45959
rect 81885 45913 81963 45959
rect 82009 45913 82087 45959
rect 82133 45913 82211 45959
rect 82257 45913 82335 45959
rect 82381 45913 82459 45959
rect 82505 45913 82583 45959
rect 82629 45913 82707 45959
rect 82753 45913 82831 45959
rect 82877 45913 82955 45959
rect 83001 45913 83079 45959
rect 83125 45913 83203 45959
rect 83249 45913 83327 45959
rect 83373 45913 83451 45959
rect 83497 45913 83575 45959
rect 83621 45913 83699 45959
rect 83745 45913 83823 45959
rect 83869 45913 83947 45959
rect 83993 45913 84071 45959
rect 84117 45913 84195 45959
rect 84241 45913 84319 45959
rect 84365 45913 84443 45959
rect 84489 45913 84567 45959
rect 84613 45913 84691 45959
rect 84737 45913 84815 45959
rect 84861 45913 84939 45959
rect 84985 45913 85063 45959
rect 85109 45913 85187 45959
rect 85233 45913 85311 45959
rect 85357 45913 85435 45959
rect 85481 45913 85559 45959
rect 85605 45913 85683 45959
rect 85729 45913 85807 45959
rect 85853 45913 85931 45959
rect 85977 45913 86098 45959
rect 352 45835 86098 45913
rect 352 45789 371 45835
rect 417 45789 495 45835
rect 541 45789 619 45835
rect 665 45789 743 45835
rect 789 45789 867 45835
rect 913 45789 991 45835
rect 1037 45789 1115 45835
rect 1161 45789 1239 45835
rect 1285 45789 1363 45835
rect 1409 45789 1487 45835
rect 1533 45789 1611 45835
rect 1657 45789 1735 45835
rect 1781 45789 1859 45835
rect 1905 45789 1983 45835
rect 2029 45789 2107 45835
rect 2153 45789 2231 45835
rect 2277 45789 2355 45835
rect 2401 45789 2479 45835
rect 2525 45789 2603 45835
rect 2649 45789 2727 45835
rect 2773 45789 2851 45835
rect 2897 45789 2975 45835
rect 3021 45789 3099 45835
rect 3145 45789 3223 45835
rect 3269 45789 3347 45835
rect 3393 45789 3471 45835
rect 3517 45789 3595 45835
rect 3641 45789 3719 45835
rect 3765 45789 3843 45835
rect 3889 45789 3967 45835
rect 4013 45789 4091 45835
rect 4137 45789 4215 45835
rect 4261 45789 4339 45835
rect 4385 45789 4463 45835
rect 4509 45789 4587 45835
rect 4633 45789 4711 45835
rect 4757 45789 4835 45835
rect 4881 45789 4959 45835
rect 5005 45789 5083 45835
rect 5129 45789 5207 45835
rect 5253 45789 5331 45835
rect 5377 45789 5455 45835
rect 5501 45789 5579 45835
rect 5625 45789 5703 45835
rect 5749 45789 5827 45835
rect 5873 45789 5951 45835
rect 5997 45789 6075 45835
rect 6121 45789 6199 45835
rect 6245 45789 6323 45835
rect 6369 45789 6447 45835
rect 6493 45789 6571 45835
rect 6617 45789 6695 45835
rect 6741 45789 6819 45835
rect 6865 45789 6943 45835
rect 6989 45789 7067 45835
rect 7113 45789 7191 45835
rect 7237 45789 7315 45835
rect 7361 45789 7439 45835
rect 7485 45789 7563 45835
rect 7609 45789 7687 45835
rect 7733 45789 7811 45835
rect 7857 45789 7935 45835
rect 7981 45789 8059 45835
rect 8105 45789 8183 45835
rect 8229 45789 8307 45835
rect 8353 45789 8431 45835
rect 8477 45789 8555 45835
rect 8601 45789 8679 45835
rect 8725 45789 8803 45835
rect 8849 45789 8927 45835
rect 8973 45789 9051 45835
rect 9097 45789 9175 45835
rect 9221 45789 9299 45835
rect 9345 45789 9423 45835
rect 9469 45789 9547 45835
rect 9593 45789 9671 45835
rect 9717 45789 9795 45835
rect 9841 45789 9919 45835
rect 9965 45789 10043 45835
rect 10089 45789 10167 45835
rect 10213 45789 10291 45835
rect 10337 45789 10415 45835
rect 10461 45789 10539 45835
rect 10585 45789 10663 45835
rect 10709 45789 10787 45835
rect 10833 45789 10911 45835
rect 10957 45789 11035 45835
rect 11081 45789 11159 45835
rect 11205 45789 11283 45835
rect 11329 45789 11407 45835
rect 11453 45789 11531 45835
rect 11577 45789 11655 45835
rect 11701 45789 11779 45835
rect 11825 45789 11903 45835
rect 11949 45789 12027 45835
rect 12073 45789 12151 45835
rect 12197 45789 12275 45835
rect 12321 45789 12399 45835
rect 12445 45789 12523 45835
rect 12569 45789 12647 45835
rect 12693 45789 12771 45835
rect 12817 45789 12895 45835
rect 12941 45789 13019 45835
rect 13065 45789 13143 45835
rect 13189 45789 13267 45835
rect 13313 45789 13391 45835
rect 13437 45789 13515 45835
rect 13561 45789 13639 45835
rect 13685 45789 13763 45835
rect 13809 45789 13887 45835
rect 13933 45789 14011 45835
rect 14057 45789 14135 45835
rect 14181 45789 14259 45835
rect 14305 45789 14383 45835
rect 14429 45789 14507 45835
rect 14553 45789 14631 45835
rect 14677 45789 14755 45835
rect 14801 45789 14879 45835
rect 14925 45789 15003 45835
rect 15049 45789 15127 45835
rect 15173 45789 15251 45835
rect 15297 45789 15375 45835
rect 15421 45789 15499 45835
rect 15545 45789 15623 45835
rect 15669 45789 15747 45835
rect 15793 45789 15871 45835
rect 15917 45789 15995 45835
rect 16041 45789 16119 45835
rect 16165 45789 16243 45835
rect 16289 45789 16367 45835
rect 16413 45789 16491 45835
rect 16537 45789 16615 45835
rect 16661 45789 16739 45835
rect 16785 45789 16863 45835
rect 16909 45789 16987 45835
rect 17033 45789 17111 45835
rect 17157 45789 17235 45835
rect 17281 45789 17359 45835
rect 17405 45789 17483 45835
rect 17529 45789 17607 45835
rect 17653 45789 17731 45835
rect 17777 45789 17855 45835
rect 17901 45789 17979 45835
rect 18025 45789 18103 45835
rect 18149 45789 18227 45835
rect 18273 45789 18351 45835
rect 18397 45789 18475 45835
rect 18521 45789 18599 45835
rect 18645 45789 18723 45835
rect 18769 45789 18847 45835
rect 18893 45789 18971 45835
rect 19017 45789 19095 45835
rect 19141 45789 19219 45835
rect 19265 45789 19343 45835
rect 19389 45789 19467 45835
rect 19513 45789 19591 45835
rect 19637 45789 19715 45835
rect 19761 45789 19839 45835
rect 19885 45789 19963 45835
rect 20009 45789 20087 45835
rect 20133 45789 20211 45835
rect 20257 45789 20335 45835
rect 20381 45789 20459 45835
rect 20505 45789 20583 45835
rect 20629 45789 20707 45835
rect 20753 45789 20831 45835
rect 20877 45789 20955 45835
rect 21001 45789 21079 45835
rect 21125 45789 21203 45835
rect 21249 45789 21327 45835
rect 21373 45789 21451 45835
rect 21497 45789 21575 45835
rect 21621 45789 21699 45835
rect 21745 45789 21823 45835
rect 21869 45789 21947 45835
rect 21993 45789 22071 45835
rect 22117 45789 22195 45835
rect 22241 45789 22319 45835
rect 22365 45789 22443 45835
rect 22489 45789 22567 45835
rect 22613 45789 22691 45835
rect 22737 45789 22815 45835
rect 22861 45789 22939 45835
rect 22985 45789 23063 45835
rect 23109 45789 23187 45835
rect 23233 45789 23311 45835
rect 23357 45789 23435 45835
rect 23481 45789 23559 45835
rect 23605 45789 23683 45835
rect 23729 45789 23807 45835
rect 23853 45789 23931 45835
rect 23977 45789 24055 45835
rect 24101 45789 24179 45835
rect 24225 45789 24303 45835
rect 24349 45789 24427 45835
rect 24473 45789 24551 45835
rect 24597 45789 24675 45835
rect 24721 45789 24799 45835
rect 24845 45789 24923 45835
rect 24969 45789 25047 45835
rect 25093 45789 25171 45835
rect 25217 45789 25295 45835
rect 25341 45789 25419 45835
rect 25465 45789 25543 45835
rect 25589 45789 25667 45835
rect 25713 45789 25791 45835
rect 25837 45789 25915 45835
rect 25961 45789 26039 45835
rect 26085 45789 26163 45835
rect 26209 45789 26287 45835
rect 26333 45789 26411 45835
rect 26457 45789 26535 45835
rect 26581 45789 26659 45835
rect 26705 45789 26783 45835
rect 26829 45789 26907 45835
rect 26953 45789 27031 45835
rect 27077 45789 27155 45835
rect 27201 45789 27279 45835
rect 27325 45789 27403 45835
rect 27449 45789 27527 45835
rect 27573 45789 27651 45835
rect 27697 45789 27775 45835
rect 27821 45789 27899 45835
rect 27945 45789 28023 45835
rect 28069 45789 28147 45835
rect 28193 45789 28271 45835
rect 28317 45789 28395 45835
rect 28441 45789 28519 45835
rect 28565 45789 28643 45835
rect 28689 45789 28767 45835
rect 28813 45789 28891 45835
rect 28937 45789 29015 45835
rect 29061 45789 29139 45835
rect 29185 45789 29263 45835
rect 29309 45789 29387 45835
rect 29433 45789 29511 45835
rect 29557 45789 29635 45835
rect 29681 45789 29759 45835
rect 29805 45789 29883 45835
rect 29929 45789 30007 45835
rect 30053 45789 30131 45835
rect 30177 45789 30255 45835
rect 30301 45789 30379 45835
rect 30425 45789 30503 45835
rect 30549 45789 30627 45835
rect 30673 45789 30751 45835
rect 30797 45789 30875 45835
rect 30921 45789 30999 45835
rect 31045 45789 31123 45835
rect 31169 45789 31247 45835
rect 31293 45789 31371 45835
rect 31417 45789 31495 45835
rect 31541 45789 31619 45835
rect 31665 45789 31743 45835
rect 31789 45789 31867 45835
rect 31913 45789 31991 45835
rect 32037 45789 32115 45835
rect 32161 45789 32239 45835
rect 32285 45789 32363 45835
rect 32409 45789 32487 45835
rect 32533 45789 32611 45835
rect 32657 45789 32735 45835
rect 32781 45789 32859 45835
rect 32905 45789 32983 45835
rect 33029 45789 33107 45835
rect 33153 45789 33231 45835
rect 33277 45789 33355 45835
rect 33401 45789 33479 45835
rect 33525 45789 33603 45835
rect 33649 45789 33727 45835
rect 33773 45789 33851 45835
rect 33897 45789 33975 45835
rect 34021 45789 34099 45835
rect 34145 45789 34223 45835
rect 34269 45789 34347 45835
rect 34393 45789 34471 45835
rect 34517 45789 34595 45835
rect 34641 45789 34719 45835
rect 34765 45789 34843 45835
rect 34889 45789 34967 45835
rect 35013 45789 35091 45835
rect 35137 45789 35215 45835
rect 35261 45789 35339 45835
rect 35385 45789 35463 45835
rect 35509 45789 35587 45835
rect 35633 45789 35711 45835
rect 35757 45789 35835 45835
rect 35881 45789 35959 45835
rect 36005 45789 36083 45835
rect 36129 45789 36207 45835
rect 36253 45789 36331 45835
rect 36377 45789 36455 45835
rect 36501 45789 36579 45835
rect 36625 45789 36703 45835
rect 36749 45789 36827 45835
rect 36873 45789 36951 45835
rect 36997 45789 37075 45835
rect 37121 45789 37199 45835
rect 37245 45789 37323 45835
rect 37369 45789 37447 45835
rect 37493 45789 37571 45835
rect 37617 45789 37695 45835
rect 37741 45789 37819 45835
rect 37865 45789 37943 45835
rect 37989 45789 38067 45835
rect 38113 45789 38191 45835
rect 38237 45789 38315 45835
rect 38361 45789 38439 45835
rect 38485 45789 38563 45835
rect 38609 45789 38687 45835
rect 38733 45789 38811 45835
rect 38857 45789 38935 45835
rect 38981 45789 39059 45835
rect 39105 45789 39183 45835
rect 39229 45789 39307 45835
rect 39353 45789 39431 45835
rect 39477 45789 39555 45835
rect 39601 45789 39679 45835
rect 39725 45789 39803 45835
rect 39849 45789 39927 45835
rect 39973 45789 40051 45835
rect 40097 45789 40175 45835
rect 40221 45789 40299 45835
rect 40345 45789 40423 45835
rect 40469 45789 40547 45835
rect 40593 45789 40671 45835
rect 40717 45789 40795 45835
rect 40841 45789 40919 45835
rect 40965 45789 41043 45835
rect 41089 45789 41167 45835
rect 41213 45789 41291 45835
rect 41337 45789 41415 45835
rect 41461 45789 41539 45835
rect 41585 45789 41663 45835
rect 41709 45789 41787 45835
rect 41833 45789 41911 45835
rect 41957 45789 42035 45835
rect 42081 45789 42159 45835
rect 42205 45789 42283 45835
rect 42329 45789 42407 45835
rect 42453 45789 42531 45835
rect 42577 45789 42655 45835
rect 42701 45789 42779 45835
rect 42825 45789 42903 45835
rect 42949 45789 43027 45835
rect 43073 45789 43151 45835
rect 43197 45789 43275 45835
rect 43321 45789 43399 45835
rect 43445 45789 43523 45835
rect 43569 45789 43647 45835
rect 43693 45789 43771 45835
rect 43817 45789 43895 45835
rect 43941 45789 44019 45835
rect 44065 45789 44143 45835
rect 44189 45789 44267 45835
rect 44313 45789 44391 45835
rect 44437 45789 44515 45835
rect 44561 45789 44639 45835
rect 44685 45789 44763 45835
rect 44809 45789 44887 45835
rect 44933 45789 45011 45835
rect 45057 45789 45135 45835
rect 45181 45789 45259 45835
rect 45305 45789 45383 45835
rect 45429 45789 45507 45835
rect 45553 45789 45631 45835
rect 45677 45789 45755 45835
rect 45801 45789 45879 45835
rect 45925 45789 46003 45835
rect 46049 45789 46127 45835
rect 46173 45789 46251 45835
rect 46297 45789 46375 45835
rect 46421 45789 46499 45835
rect 46545 45789 46623 45835
rect 46669 45789 46747 45835
rect 46793 45789 46871 45835
rect 46917 45789 46995 45835
rect 47041 45789 47119 45835
rect 47165 45789 47243 45835
rect 47289 45789 47367 45835
rect 47413 45789 47491 45835
rect 47537 45789 47615 45835
rect 47661 45789 47739 45835
rect 47785 45789 47863 45835
rect 47909 45789 47987 45835
rect 48033 45789 48111 45835
rect 48157 45789 48235 45835
rect 48281 45789 48359 45835
rect 48405 45789 48483 45835
rect 48529 45789 48607 45835
rect 48653 45789 48731 45835
rect 48777 45789 48855 45835
rect 48901 45789 48979 45835
rect 49025 45789 49103 45835
rect 49149 45789 49227 45835
rect 49273 45789 49351 45835
rect 49397 45789 49475 45835
rect 49521 45789 49599 45835
rect 49645 45789 49723 45835
rect 49769 45789 49847 45835
rect 49893 45789 49971 45835
rect 50017 45789 50095 45835
rect 50141 45789 50219 45835
rect 50265 45789 50343 45835
rect 50389 45789 50467 45835
rect 50513 45789 50591 45835
rect 50637 45789 50715 45835
rect 50761 45789 50839 45835
rect 50885 45789 50963 45835
rect 51009 45789 51087 45835
rect 51133 45789 51211 45835
rect 51257 45789 51335 45835
rect 51381 45789 51459 45835
rect 51505 45789 51583 45835
rect 51629 45789 51707 45835
rect 51753 45789 51831 45835
rect 51877 45789 51955 45835
rect 52001 45789 52079 45835
rect 52125 45789 52203 45835
rect 52249 45789 52327 45835
rect 52373 45789 52451 45835
rect 52497 45789 52575 45835
rect 52621 45789 52699 45835
rect 52745 45789 52823 45835
rect 52869 45789 52947 45835
rect 52993 45789 53071 45835
rect 53117 45789 53195 45835
rect 53241 45789 53319 45835
rect 53365 45789 53443 45835
rect 53489 45789 53567 45835
rect 53613 45789 53691 45835
rect 53737 45789 53815 45835
rect 53861 45789 53939 45835
rect 53985 45789 54063 45835
rect 54109 45789 54187 45835
rect 54233 45789 54311 45835
rect 54357 45789 54435 45835
rect 54481 45789 54559 45835
rect 54605 45789 54683 45835
rect 54729 45789 54807 45835
rect 54853 45789 54931 45835
rect 54977 45789 55055 45835
rect 55101 45789 55179 45835
rect 55225 45789 55303 45835
rect 55349 45789 55427 45835
rect 55473 45789 55551 45835
rect 55597 45789 55675 45835
rect 55721 45789 55799 45835
rect 55845 45789 55923 45835
rect 55969 45789 56047 45835
rect 56093 45789 56171 45835
rect 56217 45789 56295 45835
rect 56341 45789 56419 45835
rect 56465 45789 56543 45835
rect 56589 45789 56667 45835
rect 56713 45789 56791 45835
rect 56837 45789 56915 45835
rect 56961 45789 57039 45835
rect 57085 45789 57163 45835
rect 57209 45789 57287 45835
rect 57333 45789 57411 45835
rect 57457 45789 57535 45835
rect 57581 45789 57659 45835
rect 57705 45789 57783 45835
rect 57829 45789 57907 45835
rect 57953 45789 58031 45835
rect 58077 45789 58155 45835
rect 58201 45789 58279 45835
rect 58325 45789 58403 45835
rect 58449 45789 58527 45835
rect 58573 45789 58651 45835
rect 58697 45789 58775 45835
rect 58821 45789 58899 45835
rect 58945 45789 59023 45835
rect 59069 45789 59147 45835
rect 59193 45789 59271 45835
rect 59317 45789 59395 45835
rect 59441 45789 59519 45835
rect 59565 45789 59643 45835
rect 59689 45789 59767 45835
rect 59813 45789 59891 45835
rect 59937 45789 60015 45835
rect 60061 45789 60139 45835
rect 60185 45789 60263 45835
rect 60309 45789 60387 45835
rect 60433 45789 60511 45835
rect 60557 45789 60635 45835
rect 60681 45789 60759 45835
rect 60805 45789 60883 45835
rect 60929 45789 61007 45835
rect 61053 45789 61131 45835
rect 61177 45789 61255 45835
rect 61301 45789 61379 45835
rect 61425 45789 61503 45835
rect 61549 45789 61627 45835
rect 61673 45789 61751 45835
rect 61797 45789 61875 45835
rect 61921 45789 61999 45835
rect 62045 45789 62123 45835
rect 62169 45789 62247 45835
rect 62293 45789 62371 45835
rect 62417 45789 62495 45835
rect 62541 45789 62619 45835
rect 62665 45789 62743 45835
rect 62789 45789 62867 45835
rect 62913 45789 62991 45835
rect 63037 45789 63115 45835
rect 63161 45789 63239 45835
rect 63285 45789 63363 45835
rect 63409 45789 63487 45835
rect 63533 45789 63611 45835
rect 63657 45789 63735 45835
rect 63781 45789 63859 45835
rect 63905 45789 63983 45835
rect 64029 45789 64107 45835
rect 64153 45789 64231 45835
rect 64277 45789 64355 45835
rect 64401 45789 64479 45835
rect 64525 45789 64603 45835
rect 64649 45789 64727 45835
rect 64773 45789 64851 45835
rect 64897 45789 64975 45835
rect 65021 45789 65099 45835
rect 65145 45789 65223 45835
rect 65269 45789 65347 45835
rect 65393 45789 65471 45835
rect 65517 45789 65595 45835
rect 65641 45789 65719 45835
rect 65765 45789 65843 45835
rect 65889 45789 65967 45835
rect 66013 45789 66091 45835
rect 66137 45789 66215 45835
rect 66261 45789 66339 45835
rect 66385 45789 66463 45835
rect 66509 45789 66587 45835
rect 66633 45789 66711 45835
rect 66757 45789 66835 45835
rect 66881 45789 66959 45835
rect 67005 45789 67083 45835
rect 67129 45789 67207 45835
rect 67253 45789 67331 45835
rect 67377 45789 67455 45835
rect 67501 45789 67579 45835
rect 67625 45789 67703 45835
rect 67749 45789 67827 45835
rect 67873 45789 67951 45835
rect 67997 45789 68075 45835
rect 68121 45789 68199 45835
rect 68245 45789 68323 45835
rect 68369 45789 68447 45835
rect 68493 45789 68571 45835
rect 68617 45789 68695 45835
rect 68741 45789 68819 45835
rect 68865 45789 68943 45835
rect 68989 45789 69067 45835
rect 69113 45789 69191 45835
rect 69237 45789 69315 45835
rect 69361 45789 69439 45835
rect 69485 45789 69563 45835
rect 69609 45789 69687 45835
rect 69733 45789 69811 45835
rect 69857 45789 69935 45835
rect 69981 45789 70059 45835
rect 70105 45789 70183 45835
rect 70229 45789 70307 45835
rect 70353 45789 70431 45835
rect 70477 45789 70555 45835
rect 70601 45789 70679 45835
rect 70725 45789 70803 45835
rect 70849 45789 70927 45835
rect 70973 45789 71051 45835
rect 71097 45789 71175 45835
rect 71221 45789 71299 45835
rect 71345 45789 71423 45835
rect 71469 45789 71547 45835
rect 71593 45789 71671 45835
rect 71717 45789 71795 45835
rect 71841 45789 71919 45835
rect 71965 45789 72043 45835
rect 72089 45789 72167 45835
rect 72213 45789 72291 45835
rect 72337 45789 72415 45835
rect 72461 45789 72539 45835
rect 72585 45789 72663 45835
rect 72709 45789 72787 45835
rect 72833 45789 72911 45835
rect 72957 45789 73035 45835
rect 73081 45789 73159 45835
rect 73205 45789 73283 45835
rect 73329 45789 73407 45835
rect 73453 45789 73531 45835
rect 73577 45789 73655 45835
rect 73701 45789 73779 45835
rect 73825 45789 73903 45835
rect 73949 45789 74027 45835
rect 74073 45789 74151 45835
rect 74197 45789 74275 45835
rect 74321 45789 74399 45835
rect 74445 45789 74523 45835
rect 74569 45789 74647 45835
rect 74693 45789 74771 45835
rect 74817 45789 74895 45835
rect 74941 45789 75019 45835
rect 75065 45789 75143 45835
rect 75189 45789 75267 45835
rect 75313 45789 75391 45835
rect 75437 45789 75515 45835
rect 75561 45789 75639 45835
rect 75685 45789 75763 45835
rect 75809 45789 75887 45835
rect 75933 45789 76011 45835
rect 76057 45789 76135 45835
rect 76181 45789 76259 45835
rect 76305 45789 76383 45835
rect 76429 45789 76507 45835
rect 76553 45789 76631 45835
rect 76677 45789 76755 45835
rect 76801 45789 76879 45835
rect 76925 45789 77003 45835
rect 77049 45789 77127 45835
rect 77173 45789 77251 45835
rect 77297 45789 77375 45835
rect 77421 45789 77499 45835
rect 77545 45789 77623 45835
rect 77669 45789 77747 45835
rect 77793 45789 77871 45835
rect 77917 45789 77995 45835
rect 78041 45789 78119 45835
rect 78165 45789 78243 45835
rect 78289 45789 78367 45835
rect 78413 45789 78491 45835
rect 78537 45789 78615 45835
rect 78661 45789 78739 45835
rect 78785 45789 78863 45835
rect 78909 45789 78987 45835
rect 79033 45789 79111 45835
rect 79157 45789 79235 45835
rect 79281 45789 79359 45835
rect 79405 45789 79483 45835
rect 79529 45789 79607 45835
rect 79653 45789 79731 45835
rect 79777 45789 79855 45835
rect 79901 45789 79979 45835
rect 80025 45789 80103 45835
rect 80149 45789 80227 45835
rect 80273 45789 80351 45835
rect 80397 45789 80475 45835
rect 80521 45789 80599 45835
rect 80645 45789 80723 45835
rect 80769 45789 80847 45835
rect 80893 45789 80971 45835
rect 81017 45789 81095 45835
rect 81141 45789 81219 45835
rect 81265 45789 81343 45835
rect 81389 45789 81467 45835
rect 81513 45789 81591 45835
rect 81637 45789 81715 45835
rect 81761 45789 81839 45835
rect 81885 45789 81963 45835
rect 82009 45789 82087 45835
rect 82133 45789 82211 45835
rect 82257 45789 82335 45835
rect 82381 45789 82459 45835
rect 82505 45789 82583 45835
rect 82629 45789 82707 45835
rect 82753 45789 82831 45835
rect 82877 45789 82955 45835
rect 83001 45789 83079 45835
rect 83125 45789 83203 45835
rect 83249 45789 83327 45835
rect 83373 45789 83451 45835
rect 83497 45789 83575 45835
rect 83621 45789 83699 45835
rect 83745 45789 83823 45835
rect 83869 45789 83947 45835
rect 83993 45789 84071 45835
rect 84117 45789 84195 45835
rect 84241 45789 84319 45835
rect 84365 45789 84443 45835
rect 84489 45789 84567 45835
rect 84613 45789 84691 45835
rect 84737 45789 84815 45835
rect 84861 45789 84939 45835
rect 84985 45789 85063 45835
rect 85109 45789 85187 45835
rect 85233 45789 85311 45835
rect 85357 45789 85435 45835
rect 85481 45789 85559 45835
rect 85605 45789 85683 45835
rect 85729 45789 85807 45835
rect 85853 45789 85931 45835
rect 85977 45789 86098 45835
rect 352 45711 86098 45789
rect 352 45665 371 45711
rect 417 45665 495 45711
rect 541 45665 619 45711
rect 665 45665 743 45711
rect 789 45665 867 45711
rect 913 45665 991 45711
rect 1037 45665 1115 45711
rect 1161 45665 1239 45711
rect 1285 45665 1363 45711
rect 1409 45665 1487 45711
rect 1533 45665 1611 45711
rect 1657 45665 1735 45711
rect 1781 45665 1859 45711
rect 1905 45665 1983 45711
rect 2029 45665 2107 45711
rect 2153 45665 2231 45711
rect 2277 45665 2355 45711
rect 2401 45665 2479 45711
rect 2525 45665 2603 45711
rect 2649 45665 2727 45711
rect 2773 45665 2851 45711
rect 2897 45665 2975 45711
rect 3021 45665 3099 45711
rect 3145 45665 3223 45711
rect 3269 45665 3347 45711
rect 3393 45665 3471 45711
rect 3517 45665 3595 45711
rect 3641 45665 3719 45711
rect 3765 45665 3843 45711
rect 3889 45665 3967 45711
rect 4013 45665 4091 45711
rect 4137 45665 4215 45711
rect 4261 45665 4339 45711
rect 4385 45665 4463 45711
rect 4509 45665 4587 45711
rect 4633 45665 4711 45711
rect 4757 45665 4835 45711
rect 4881 45665 4959 45711
rect 5005 45665 5083 45711
rect 5129 45665 5207 45711
rect 5253 45665 5331 45711
rect 5377 45665 5455 45711
rect 5501 45665 5579 45711
rect 5625 45665 5703 45711
rect 5749 45665 5827 45711
rect 5873 45665 5951 45711
rect 5997 45665 6075 45711
rect 6121 45665 6199 45711
rect 6245 45665 6323 45711
rect 6369 45665 6447 45711
rect 6493 45665 6571 45711
rect 6617 45665 6695 45711
rect 6741 45665 6819 45711
rect 6865 45665 6943 45711
rect 6989 45665 7067 45711
rect 7113 45665 7191 45711
rect 7237 45665 7315 45711
rect 7361 45665 7439 45711
rect 7485 45665 7563 45711
rect 7609 45665 7687 45711
rect 7733 45665 7811 45711
rect 7857 45665 7935 45711
rect 7981 45665 8059 45711
rect 8105 45665 8183 45711
rect 8229 45665 8307 45711
rect 8353 45665 8431 45711
rect 8477 45665 8555 45711
rect 8601 45665 8679 45711
rect 8725 45665 8803 45711
rect 8849 45665 8927 45711
rect 8973 45665 9051 45711
rect 9097 45665 9175 45711
rect 9221 45665 9299 45711
rect 9345 45665 9423 45711
rect 9469 45665 9547 45711
rect 9593 45665 9671 45711
rect 9717 45665 9795 45711
rect 9841 45665 9919 45711
rect 9965 45665 10043 45711
rect 10089 45665 10167 45711
rect 10213 45665 10291 45711
rect 10337 45665 10415 45711
rect 10461 45665 10539 45711
rect 10585 45665 10663 45711
rect 10709 45665 10787 45711
rect 10833 45665 10911 45711
rect 10957 45665 11035 45711
rect 11081 45665 11159 45711
rect 11205 45665 11283 45711
rect 11329 45665 11407 45711
rect 11453 45665 11531 45711
rect 11577 45665 11655 45711
rect 11701 45665 11779 45711
rect 11825 45665 11903 45711
rect 11949 45665 12027 45711
rect 12073 45665 12151 45711
rect 12197 45665 12275 45711
rect 12321 45665 12399 45711
rect 12445 45665 12523 45711
rect 12569 45665 12647 45711
rect 12693 45665 12771 45711
rect 12817 45665 12895 45711
rect 12941 45665 13019 45711
rect 13065 45665 13143 45711
rect 13189 45665 13267 45711
rect 13313 45665 13391 45711
rect 13437 45665 13515 45711
rect 13561 45665 13639 45711
rect 13685 45665 13763 45711
rect 13809 45665 13887 45711
rect 13933 45665 14011 45711
rect 14057 45665 14135 45711
rect 14181 45665 14259 45711
rect 14305 45665 14383 45711
rect 14429 45665 14507 45711
rect 14553 45665 14631 45711
rect 14677 45665 14755 45711
rect 14801 45665 14879 45711
rect 14925 45665 15003 45711
rect 15049 45665 15127 45711
rect 15173 45665 15251 45711
rect 15297 45665 15375 45711
rect 15421 45665 15499 45711
rect 15545 45665 15623 45711
rect 15669 45665 15747 45711
rect 15793 45665 15871 45711
rect 15917 45665 15995 45711
rect 16041 45665 16119 45711
rect 16165 45665 16243 45711
rect 16289 45665 16367 45711
rect 16413 45665 16491 45711
rect 16537 45665 16615 45711
rect 16661 45665 16739 45711
rect 16785 45665 16863 45711
rect 16909 45665 16987 45711
rect 17033 45665 17111 45711
rect 17157 45665 17235 45711
rect 17281 45665 17359 45711
rect 17405 45665 17483 45711
rect 17529 45665 17607 45711
rect 17653 45665 17731 45711
rect 17777 45665 17855 45711
rect 17901 45665 17979 45711
rect 18025 45665 18103 45711
rect 18149 45665 18227 45711
rect 18273 45665 18351 45711
rect 18397 45665 18475 45711
rect 18521 45665 18599 45711
rect 18645 45665 18723 45711
rect 18769 45665 18847 45711
rect 18893 45665 18971 45711
rect 19017 45665 19095 45711
rect 19141 45665 19219 45711
rect 19265 45665 19343 45711
rect 19389 45665 19467 45711
rect 19513 45665 19591 45711
rect 19637 45665 19715 45711
rect 19761 45665 19839 45711
rect 19885 45665 19963 45711
rect 20009 45665 20087 45711
rect 20133 45665 20211 45711
rect 20257 45665 20335 45711
rect 20381 45665 20459 45711
rect 20505 45665 20583 45711
rect 20629 45665 20707 45711
rect 20753 45665 20831 45711
rect 20877 45665 20955 45711
rect 21001 45665 21079 45711
rect 21125 45665 21203 45711
rect 21249 45665 21327 45711
rect 21373 45665 21451 45711
rect 21497 45665 21575 45711
rect 21621 45665 21699 45711
rect 21745 45665 21823 45711
rect 21869 45665 21947 45711
rect 21993 45665 22071 45711
rect 22117 45665 22195 45711
rect 22241 45665 22319 45711
rect 22365 45665 22443 45711
rect 22489 45665 22567 45711
rect 22613 45665 22691 45711
rect 22737 45665 22815 45711
rect 22861 45665 22939 45711
rect 22985 45665 23063 45711
rect 23109 45665 23187 45711
rect 23233 45665 23311 45711
rect 23357 45665 23435 45711
rect 23481 45665 23559 45711
rect 23605 45665 23683 45711
rect 23729 45665 23807 45711
rect 23853 45665 23931 45711
rect 23977 45665 24055 45711
rect 24101 45665 24179 45711
rect 24225 45665 24303 45711
rect 24349 45665 24427 45711
rect 24473 45665 24551 45711
rect 24597 45665 24675 45711
rect 24721 45665 24799 45711
rect 24845 45665 24923 45711
rect 24969 45665 25047 45711
rect 25093 45665 25171 45711
rect 25217 45665 25295 45711
rect 25341 45665 25419 45711
rect 25465 45665 25543 45711
rect 25589 45665 25667 45711
rect 25713 45665 25791 45711
rect 25837 45665 25915 45711
rect 25961 45665 26039 45711
rect 26085 45665 26163 45711
rect 26209 45665 26287 45711
rect 26333 45665 26411 45711
rect 26457 45665 26535 45711
rect 26581 45665 26659 45711
rect 26705 45665 26783 45711
rect 26829 45665 26907 45711
rect 26953 45665 27031 45711
rect 27077 45665 27155 45711
rect 27201 45665 27279 45711
rect 27325 45665 27403 45711
rect 27449 45665 27527 45711
rect 27573 45665 27651 45711
rect 27697 45665 27775 45711
rect 27821 45665 27899 45711
rect 27945 45665 28023 45711
rect 28069 45665 28147 45711
rect 28193 45665 28271 45711
rect 28317 45665 28395 45711
rect 28441 45665 28519 45711
rect 28565 45665 28643 45711
rect 28689 45665 28767 45711
rect 28813 45665 28891 45711
rect 28937 45665 29015 45711
rect 29061 45665 29139 45711
rect 29185 45665 29263 45711
rect 29309 45665 29387 45711
rect 29433 45665 29511 45711
rect 29557 45665 29635 45711
rect 29681 45665 29759 45711
rect 29805 45665 29883 45711
rect 29929 45665 30007 45711
rect 30053 45665 30131 45711
rect 30177 45665 30255 45711
rect 30301 45665 30379 45711
rect 30425 45665 30503 45711
rect 30549 45665 30627 45711
rect 30673 45665 30751 45711
rect 30797 45665 30875 45711
rect 30921 45665 30999 45711
rect 31045 45665 31123 45711
rect 31169 45665 31247 45711
rect 31293 45665 31371 45711
rect 31417 45665 31495 45711
rect 31541 45665 31619 45711
rect 31665 45665 31743 45711
rect 31789 45665 31867 45711
rect 31913 45665 31991 45711
rect 32037 45665 32115 45711
rect 32161 45665 32239 45711
rect 32285 45665 32363 45711
rect 32409 45665 32487 45711
rect 32533 45665 32611 45711
rect 32657 45665 32735 45711
rect 32781 45665 32859 45711
rect 32905 45665 32983 45711
rect 33029 45665 33107 45711
rect 33153 45665 33231 45711
rect 33277 45665 33355 45711
rect 33401 45665 33479 45711
rect 33525 45665 33603 45711
rect 33649 45665 33727 45711
rect 33773 45665 33851 45711
rect 33897 45665 33975 45711
rect 34021 45665 34099 45711
rect 34145 45665 34223 45711
rect 34269 45665 34347 45711
rect 34393 45665 34471 45711
rect 34517 45665 34595 45711
rect 34641 45665 34719 45711
rect 34765 45665 34843 45711
rect 34889 45665 34967 45711
rect 35013 45665 35091 45711
rect 35137 45665 35215 45711
rect 35261 45665 35339 45711
rect 35385 45665 35463 45711
rect 35509 45665 35587 45711
rect 35633 45665 35711 45711
rect 35757 45665 35835 45711
rect 35881 45665 35959 45711
rect 36005 45665 36083 45711
rect 36129 45665 36207 45711
rect 36253 45665 36331 45711
rect 36377 45665 36455 45711
rect 36501 45665 36579 45711
rect 36625 45665 36703 45711
rect 36749 45665 36827 45711
rect 36873 45665 36951 45711
rect 36997 45665 37075 45711
rect 37121 45665 37199 45711
rect 37245 45665 37323 45711
rect 37369 45665 37447 45711
rect 37493 45665 37571 45711
rect 37617 45665 37695 45711
rect 37741 45665 37819 45711
rect 37865 45665 37943 45711
rect 37989 45665 38067 45711
rect 38113 45665 38191 45711
rect 38237 45665 38315 45711
rect 38361 45665 38439 45711
rect 38485 45665 38563 45711
rect 38609 45665 38687 45711
rect 38733 45665 38811 45711
rect 38857 45665 38935 45711
rect 38981 45665 39059 45711
rect 39105 45665 39183 45711
rect 39229 45665 39307 45711
rect 39353 45665 39431 45711
rect 39477 45665 39555 45711
rect 39601 45665 39679 45711
rect 39725 45665 39803 45711
rect 39849 45665 39927 45711
rect 39973 45665 40051 45711
rect 40097 45665 40175 45711
rect 40221 45665 40299 45711
rect 40345 45665 40423 45711
rect 40469 45665 40547 45711
rect 40593 45665 40671 45711
rect 40717 45665 40795 45711
rect 40841 45665 40919 45711
rect 40965 45665 41043 45711
rect 41089 45665 41167 45711
rect 41213 45665 41291 45711
rect 41337 45665 41415 45711
rect 41461 45665 41539 45711
rect 41585 45665 41663 45711
rect 41709 45665 41787 45711
rect 41833 45665 41911 45711
rect 41957 45665 42035 45711
rect 42081 45665 42159 45711
rect 42205 45665 42283 45711
rect 42329 45665 42407 45711
rect 42453 45665 42531 45711
rect 42577 45665 42655 45711
rect 42701 45665 42779 45711
rect 42825 45665 42903 45711
rect 42949 45665 43027 45711
rect 43073 45665 43151 45711
rect 43197 45665 43275 45711
rect 43321 45665 43399 45711
rect 43445 45665 43523 45711
rect 43569 45665 43647 45711
rect 43693 45665 43771 45711
rect 43817 45665 43895 45711
rect 43941 45665 44019 45711
rect 44065 45665 44143 45711
rect 44189 45665 44267 45711
rect 44313 45665 44391 45711
rect 44437 45665 44515 45711
rect 44561 45665 44639 45711
rect 44685 45665 44763 45711
rect 44809 45665 44887 45711
rect 44933 45665 45011 45711
rect 45057 45665 45135 45711
rect 45181 45665 45259 45711
rect 45305 45665 45383 45711
rect 45429 45665 45507 45711
rect 45553 45665 45631 45711
rect 45677 45665 45755 45711
rect 45801 45665 45879 45711
rect 45925 45665 46003 45711
rect 46049 45665 46127 45711
rect 46173 45665 46251 45711
rect 46297 45665 46375 45711
rect 46421 45665 46499 45711
rect 46545 45665 46623 45711
rect 46669 45665 46747 45711
rect 46793 45665 46871 45711
rect 46917 45665 46995 45711
rect 47041 45665 47119 45711
rect 47165 45665 47243 45711
rect 47289 45665 47367 45711
rect 47413 45665 47491 45711
rect 47537 45665 47615 45711
rect 47661 45665 47739 45711
rect 47785 45665 47863 45711
rect 47909 45665 47987 45711
rect 48033 45665 48111 45711
rect 48157 45665 48235 45711
rect 48281 45665 48359 45711
rect 48405 45665 48483 45711
rect 48529 45665 48607 45711
rect 48653 45665 48731 45711
rect 48777 45665 48855 45711
rect 48901 45665 48979 45711
rect 49025 45665 49103 45711
rect 49149 45665 49227 45711
rect 49273 45665 49351 45711
rect 49397 45665 49475 45711
rect 49521 45665 49599 45711
rect 49645 45665 49723 45711
rect 49769 45665 49847 45711
rect 49893 45665 49971 45711
rect 50017 45665 50095 45711
rect 50141 45665 50219 45711
rect 50265 45665 50343 45711
rect 50389 45665 50467 45711
rect 50513 45665 50591 45711
rect 50637 45665 50715 45711
rect 50761 45665 50839 45711
rect 50885 45665 50963 45711
rect 51009 45665 51087 45711
rect 51133 45665 51211 45711
rect 51257 45665 51335 45711
rect 51381 45665 51459 45711
rect 51505 45665 51583 45711
rect 51629 45665 51707 45711
rect 51753 45665 51831 45711
rect 51877 45665 51955 45711
rect 52001 45665 52079 45711
rect 52125 45665 52203 45711
rect 52249 45665 52327 45711
rect 52373 45665 52451 45711
rect 52497 45665 52575 45711
rect 52621 45665 52699 45711
rect 52745 45665 52823 45711
rect 52869 45665 52947 45711
rect 52993 45665 53071 45711
rect 53117 45665 53195 45711
rect 53241 45665 53319 45711
rect 53365 45665 53443 45711
rect 53489 45665 53567 45711
rect 53613 45665 53691 45711
rect 53737 45665 53815 45711
rect 53861 45665 53939 45711
rect 53985 45665 54063 45711
rect 54109 45665 54187 45711
rect 54233 45665 54311 45711
rect 54357 45665 54435 45711
rect 54481 45665 54559 45711
rect 54605 45665 54683 45711
rect 54729 45665 54807 45711
rect 54853 45665 54931 45711
rect 54977 45665 55055 45711
rect 55101 45665 55179 45711
rect 55225 45665 55303 45711
rect 55349 45665 55427 45711
rect 55473 45665 55551 45711
rect 55597 45665 55675 45711
rect 55721 45665 55799 45711
rect 55845 45665 55923 45711
rect 55969 45665 56047 45711
rect 56093 45665 56171 45711
rect 56217 45665 56295 45711
rect 56341 45665 56419 45711
rect 56465 45665 56543 45711
rect 56589 45665 56667 45711
rect 56713 45665 56791 45711
rect 56837 45665 56915 45711
rect 56961 45665 57039 45711
rect 57085 45665 57163 45711
rect 57209 45665 57287 45711
rect 57333 45665 57411 45711
rect 57457 45665 57535 45711
rect 57581 45665 57659 45711
rect 57705 45665 57783 45711
rect 57829 45665 57907 45711
rect 57953 45665 58031 45711
rect 58077 45665 58155 45711
rect 58201 45665 58279 45711
rect 58325 45665 58403 45711
rect 58449 45665 58527 45711
rect 58573 45665 58651 45711
rect 58697 45665 58775 45711
rect 58821 45665 58899 45711
rect 58945 45665 59023 45711
rect 59069 45665 59147 45711
rect 59193 45665 59271 45711
rect 59317 45665 59395 45711
rect 59441 45665 59519 45711
rect 59565 45665 59643 45711
rect 59689 45665 59767 45711
rect 59813 45665 59891 45711
rect 59937 45665 60015 45711
rect 60061 45665 60139 45711
rect 60185 45665 60263 45711
rect 60309 45665 60387 45711
rect 60433 45665 60511 45711
rect 60557 45665 60635 45711
rect 60681 45665 60759 45711
rect 60805 45665 60883 45711
rect 60929 45665 61007 45711
rect 61053 45665 61131 45711
rect 61177 45665 61255 45711
rect 61301 45665 61379 45711
rect 61425 45665 61503 45711
rect 61549 45665 61627 45711
rect 61673 45665 61751 45711
rect 61797 45665 61875 45711
rect 61921 45665 61999 45711
rect 62045 45665 62123 45711
rect 62169 45665 62247 45711
rect 62293 45665 62371 45711
rect 62417 45665 62495 45711
rect 62541 45665 62619 45711
rect 62665 45665 62743 45711
rect 62789 45665 62867 45711
rect 62913 45665 62991 45711
rect 63037 45665 63115 45711
rect 63161 45665 63239 45711
rect 63285 45665 63363 45711
rect 63409 45665 63487 45711
rect 63533 45665 63611 45711
rect 63657 45665 63735 45711
rect 63781 45665 63859 45711
rect 63905 45665 63983 45711
rect 64029 45665 64107 45711
rect 64153 45665 64231 45711
rect 64277 45665 64355 45711
rect 64401 45665 64479 45711
rect 64525 45665 64603 45711
rect 64649 45665 64727 45711
rect 64773 45665 64851 45711
rect 64897 45665 64975 45711
rect 65021 45665 65099 45711
rect 65145 45665 65223 45711
rect 65269 45665 65347 45711
rect 65393 45665 65471 45711
rect 65517 45665 65595 45711
rect 65641 45665 65719 45711
rect 65765 45665 65843 45711
rect 65889 45665 65967 45711
rect 66013 45665 66091 45711
rect 66137 45665 66215 45711
rect 66261 45665 66339 45711
rect 66385 45665 66463 45711
rect 66509 45665 66587 45711
rect 66633 45665 66711 45711
rect 66757 45665 66835 45711
rect 66881 45665 66959 45711
rect 67005 45665 67083 45711
rect 67129 45665 67207 45711
rect 67253 45665 67331 45711
rect 67377 45665 67455 45711
rect 67501 45665 67579 45711
rect 67625 45665 67703 45711
rect 67749 45665 67827 45711
rect 67873 45665 67951 45711
rect 67997 45665 68075 45711
rect 68121 45665 68199 45711
rect 68245 45665 68323 45711
rect 68369 45665 68447 45711
rect 68493 45665 68571 45711
rect 68617 45665 68695 45711
rect 68741 45665 68819 45711
rect 68865 45665 68943 45711
rect 68989 45665 69067 45711
rect 69113 45665 69191 45711
rect 69237 45665 69315 45711
rect 69361 45665 69439 45711
rect 69485 45665 69563 45711
rect 69609 45665 69687 45711
rect 69733 45665 69811 45711
rect 69857 45665 69935 45711
rect 69981 45665 70059 45711
rect 70105 45665 70183 45711
rect 70229 45665 70307 45711
rect 70353 45665 70431 45711
rect 70477 45665 70555 45711
rect 70601 45665 70679 45711
rect 70725 45665 70803 45711
rect 70849 45665 70927 45711
rect 70973 45665 71051 45711
rect 71097 45665 71175 45711
rect 71221 45665 71299 45711
rect 71345 45665 71423 45711
rect 71469 45665 71547 45711
rect 71593 45665 71671 45711
rect 71717 45665 71795 45711
rect 71841 45665 71919 45711
rect 71965 45665 72043 45711
rect 72089 45665 72167 45711
rect 72213 45665 72291 45711
rect 72337 45665 72415 45711
rect 72461 45665 72539 45711
rect 72585 45665 72663 45711
rect 72709 45665 72787 45711
rect 72833 45665 72911 45711
rect 72957 45665 73035 45711
rect 73081 45665 73159 45711
rect 73205 45665 73283 45711
rect 73329 45665 73407 45711
rect 73453 45665 73531 45711
rect 73577 45665 73655 45711
rect 73701 45665 73779 45711
rect 73825 45665 73903 45711
rect 73949 45665 74027 45711
rect 74073 45665 74151 45711
rect 74197 45665 74275 45711
rect 74321 45665 74399 45711
rect 74445 45665 74523 45711
rect 74569 45665 74647 45711
rect 74693 45665 74771 45711
rect 74817 45665 74895 45711
rect 74941 45665 75019 45711
rect 75065 45665 75143 45711
rect 75189 45665 75267 45711
rect 75313 45665 75391 45711
rect 75437 45665 75515 45711
rect 75561 45665 75639 45711
rect 75685 45665 75763 45711
rect 75809 45665 75887 45711
rect 75933 45665 76011 45711
rect 76057 45665 76135 45711
rect 76181 45665 76259 45711
rect 76305 45665 76383 45711
rect 76429 45665 76507 45711
rect 76553 45665 76631 45711
rect 76677 45665 76755 45711
rect 76801 45665 76879 45711
rect 76925 45665 77003 45711
rect 77049 45665 77127 45711
rect 77173 45665 77251 45711
rect 77297 45665 77375 45711
rect 77421 45665 77499 45711
rect 77545 45665 77623 45711
rect 77669 45665 77747 45711
rect 77793 45665 77871 45711
rect 77917 45665 77995 45711
rect 78041 45665 78119 45711
rect 78165 45665 78243 45711
rect 78289 45665 78367 45711
rect 78413 45665 78491 45711
rect 78537 45665 78615 45711
rect 78661 45665 78739 45711
rect 78785 45665 78863 45711
rect 78909 45665 78987 45711
rect 79033 45665 79111 45711
rect 79157 45665 79235 45711
rect 79281 45665 79359 45711
rect 79405 45665 79483 45711
rect 79529 45665 79607 45711
rect 79653 45665 79731 45711
rect 79777 45665 79855 45711
rect 79901 45665 79979 45711
rect 80025 45665 80103 45711
rect 80149 45665 80227 45711
rect 80273 45665 80351 45711
rect 80397 45665 80475 45711
rect 80521 45665 80599 45711
rect 80645 45665 80723 45711
rect 80769 45665 80847 45711
rect 80893 45665 80971 45711
rect 81017 45665 81095 45711
rect 81141 45665 81219 45711
rect 81265 45665 81343 45711
rect 81389 45665 81467 45711
rect 81513 45665 81591 45711
rect 81637 45665 81715 45711
rect 81761 45665 81839 45711
rect 81885 45665 81963 45711
rect 82009 45665 82087 45711
rect 82133 45665 82211 45711
rect 82257 45665 82335 45711
rect 82381 45665 82459 45711
rect 82505 45665 82583 45711
rect 82629 45665 82707 45711
rect 82753 45665 82831 45711
rect 82877 45665 82955 45711
rect 83001 45665 83079 45711
rect 83125 45665 83203 45711
rect 83249 45665 83327 45711
rect 83373 45665 83451 45711
rect 83497 45665 83575 45711
rect 83621 45665 83699 45711
rect 83745 45665 83823 45711
rect 83869 45665 83947 45711
rect 83993 45665 84071 45711
rect 84117 45665 84195 45711
rect 84241 45665 84319 45711
rect 84365 45665 84443 45711
rect 84489 45665 84567 45711
rect 84613 45665 84691 45711
rect 84737 45665 84815 45711
rect 84861 45665 84939 45711
rect 84985 45665 85063 45711
rect 85109 45665 85187 45711
rect 85233 45665 85311 45711
rect 85357 45665 85435 45711
rect 85481 45665 85559 45711
rect 85605 45665 85683 45711
rect 85729 45665 85807 45711
rect 85853 45665 85931 45711
rect 85977 45665 86098 45711
rect 352 45646 86098 45665
rect 352 45563 736 45646
rect 352 1117 371 45563
rect 717 1117 736 45563
rect 352 1034 736 1117
rect 27479 45563 28911 45646
rect 27479 1117 27498 45563
rect 27744 45442 28911 45563
rect 27744 35996 27846 45442
rect 28492 44122 28911 45442
rect 56212 45463 57645 45646
rect 56212 45442 57380 45463
rect 32989 44309 34884 44366
rect 32989 44263 33044 44309
rect 33090 44263 33202 44309
rect 33248 44263 33360 44309
rect 33406 44263 33518 44309
rect 33564 44263 33677 44309
rect 33723 44263 33835 44309
rect 33881 44263 33993 44309
rect 34039 44263 34151 44309
rect 34197 44263 34309 44309
rect 34355 44263 34467 44309
rect 34513 44263 34625 44309
rect 34671 44263 34783 44309
rect 34829 44263 34884 44309
rect 32989 44206 34884 44263
rect 40062 44309 41957 44366
rect 40062 44263 40117 44309
rect 40163 44263 40275 44309
rect 40321 44263 40433 44309
rect 40479 44263 40591 44309
rect 40637 44263 40750 44309
rect 40796 44263 40908 44309
rect 40954 44263 41066 44309
rect 41112 44263 41224 44309
rect 41270 44263 41382 44309
rect 41428 44263 41540 44309
rect 41586 44263 41698 44309
rect 41744 44263 41856 44309
rect 41902 44263 41957 44309
rect 28492 44076 28810 44122
rect 28856 44076 28911 44122
rect 28492 43958 28911 44076
rect 28492 43912 28810 43958
rect 28856 43912 28911 43958
rect 28492 43795 28911 43912
rect 28492 43749 28810 43795
rect 28856 43749 28911 43795
rect 28492 43632 28911 43749
rect 28492 43586 28810 43632
rect 28856 43586 28911 43632
rect 28492 43468 28911 43586
rect 28492 43422 28810 43468
rect 28856 43422 28911 43468
rect 28492 43266 28911 43422
rect 40062 44206 41957 44263
rect 44459 44309 44931 44366
rect 44459 44263 44514 44309
rect 44560 44263 44672 44309
rect 44718 44263 44830 44309
rect 44876 44263 44931 44309
rect 44459 44206 44931 44263
rect 50074 44309 51969 44366
rect 50074 44263 50129 44309
rect 50175 44263 50287 44309
rect 50333 44263 50445 44309
rect 50491 44263 50603 44309
rect 50649 44263 50762 44309
rect 50808 44263 50920 44309
rect 50966 44263 51078 44309
rect 51124 44263 51236 44309
rect 51282 44263 51394 44309
rect 51440 44263 51552 44309
rect 51598 44263 51710 44309
rect 51756 44263 51868 44309
rect 51914 44263 51969 44309
rect 50074 44206 51969 44263
rect 28492 43220 28810 43266
rect 28856 43220 28911 43266
rect 28492 43103 28911 43220
rect 28492 43057 28810 43103
rect 28856 43057 28911 43103
rect 28492 42940 28911 43057
rect 28492 42894 28810 42940
rect 28856 42894 28911 42940
rect 28492 42777 28911 42894
rect 28492 42731 28810 42777
rect 28856 42731 28911 42777
rect 28492 42613 28911 42731
rect 28492 42567 28810 42613
rect 28856 42567 28911 42613
rect 28492 42450 28911 42567
rect 37938 43350 38492 43369
rect 37938 43304 37957 43350
rect 38473 43304 38492 43350
rect 37938 43285 38492 43304
rect 40779 43350 42995 43410
rect 40779 43304 40836 43350
rect 40882 43304 40994 43350
rect 41040 43304 41152 43350
rect 41198 43304 41310 43350
rect 41356 43304 41469 43350
rect 41515 43304 41627 43350
rect 41673 43304 41785 43350
rect 41831 43304 41943 43350
rect 41989 43304 42101 43350
rect 42147 43304 42259 43350
rect 42305 43304 42418 43350
rect 42464 43304 42576 43350
rect 42622 43304 42734 43350
rect 42780 43304 42892 43350
rect 42938 43304 42995 43350
rect 40779 43244 42995 43304
rect 56212 44122 56632 45442
rect 56212 44076 56267 44122
rect 56313 44076 56632 44122
rect 56212 43958 56632 44076
rect 56212 43912 56267 43958
rect 56313 43912 56632 43958
rect 56212 43795 56632 43912
rect 56212 43749 56267 43795
rect 56313 43749 56632 43795
rect 56212 43632 56632 43749
rect 56212 43586 56267 43632
rect 56313 43586 56632 43632
rect 56212 43468 56632 43586
rect 56212 43422 56267 43468
rect 56313 43422 56632 43468
rect 28492 42404 28810 42450
rect 28856 42404 28911 42450
rect 28492 42287 28911 42404
rect 28492 42241 28810 42287
rect 28856 42241 28911 42287
rect 28492 42123 28911 42241
rect 28492 42077 28810 42123
rect 28856 42077 28911 42123
rect 28492 41960 28911 42077
rect 28492 41914 28810 41960
rect 28856 41914 28911 41960
rect 28492 41797 28911 41914
rect 28492 41751 28810 41797
rect 28856 41751 28911 41797
rect 28492 41634 28911 41751
rect 28492 41588 28810 41634
rect 28856 41588 28911 41634
rect 28492 41466 28911 41588
rect 34861 42450 35017 42507
rect 34861 42404 34916 42450
rect 34962 42404 35017 42450
rect 34861 42347 35017 42404
rect 50103 42450 50263 42510
rect 50103 42404 50160 42450
rect 50206 42404 50263 42450
rect 50103 42344 50263 42404
rect 56212 43266 56632 43422
rect 56212 43220 56267 43266
rect 56313 43220 56632 43266
rect 56212 43103 56632 43220
rect 56212 43057 56267 43103
rect 56313 43057 56632 43103
rect 56212 42940 56632 43057
rect 56212 42894 56267 42940
rect 56313 42894 56632 42940
rect 56212 42777 56632 42894
rect 56212 42731 56267 42777
rect 56313 42731 56632 42777
rect 56212 42613 56632 42731
rect 56212 42567 56267 42613
rect 56313 42567 56632 42613
rect 56212 42450 56632 42567
rect 56212 42404 56267 42450
rect 56313 42404 56632 42450
rect 28492 41420 28810 41466
rect 28856 41420 28911 41466
rect 28492 41303 28911 41420
rect 28492 41257 28810 41303
rect 28856 41257 28911 41303
rect 28492 41140 28911 41257
rect 28492 41094 28810 41140
rect 28856 41094 28911 41140
rect 28492 40977 28911 41094
rect 28492 40931 28810 40977
rect 28856 40931 28911 40977
rect 28492 40813 28911 40931
rect 28492 40767 28810 40813
rect 28856 40767 28911 40813
rect 28492 40650 28911 40767
rect 37938 41550 38492 41569
rect 37938 41504 37957 41550
rect 38473 41504 38492 41550
rect 37938 41485 38492 41504
rect 40779 41550 42995 41610
rect 40779 41504 40836 41550
rect 40882 41504 40994 41550
rect 41040 41504 41152 41550
rect 41198 41504 41310 41550
rect 41356 41504 41469 41550
rect 41515 41504 41627 41550
rect 41673 41504 41785 41550
rect 41831 41504 41943 41550
rect 41989 41504 42101 41550
rect 42147 41504 42259 41550
rect 42305 41504 42418 41550
rect 42464 41504 42576 41550
rect 42622 41504 42734 41550
rect 42780 41504 42892 41550
rect 42938 41504 42995 41550
rect 40779 41444 42995 41504
rect 56212 42287 56632 42404
rect 56212 42241 56267 42287
rect 56313 42241 56632 42287
rect 56212 42123 56632 42241
rect 56212 42077 56267 42123
rect 56313 42077 56632 42123
rect 56212 41960 56632 42077
rect 56212 41914 56267 41960
rect 56313 41914 56632 41960
rect 56212 41797 56632 41914
rect 56212 41751 56267 41797
rect 56313 41751 56632 41797
rect 56212 41634 56632 41751
rect 56212 41588 56267 41634
rect 56313 41588 56632 41634
rect 28492 40604 28810 40650
rect 28856 40604 28911 40650
rect 28492 40487 28911 40604
rect 28492 40441 28810 40487
rect 28856 40441 28911 40487
rect 28492 40323 28911 40441
rect 28492 40277 28810 40323
rect 28856 40277 28911 40323
rect 28492 40160 28911 40277
rect 28492 40114 28810 40160
rect 28856 40114 28911 40160
rect 28492 39997 28911 40114
rect 28492 39951 28810 39997
rect 28856 39951 28911 39997
rect 28492 39834 28911 39951
rect 28492 39788 28810 39834
rect 28856 39788 28911 39834
rect 28492 39666 28911 39788
rect 34861 40650 35017 40707
rect 34861 40604 34916 40650
rect 34962 40604 35017 40650
rect 34861 40547 35017 40604
rect 50103 40650 50263 40710
rect 50103 40604 50160 40650
rect 50206 40604 50263 40650
rect 50103 40544 50263 40604
rect 56212 41466 56632 41588
rect 56212 41420 56267 41466
rect 56313 41420 56632 41466
rect 56212 41303 56632 41420
rect 56212 41257 56267 41303
rect 56313 41257 56632 41303
rect 56212 41140 56632 41257
rect 56212 41094 56267 41140
rect 56313 41094 56632 41140
rect 56212 40977 56632 41094
rect 56212 40931 56267 40977
rect 56313 40931 56632 40977
rect 56212 40813 56632 40931
rect 56212 40767 56267 40813
rect 56313 40767 56632 40813
rect 56212 40650 56632 40767
rect 56212 40604 56267 40650
rect 56313 40604 56632 40650
rect 28492 39620 28810 39666
rect 28856 39620 28911 39666
rect 28492 39503 28911 39620
rect 28492 39457 28810 39503
rect 28856 39457 28911 39503
rect 28492 39340 28911 39457
rect 28492 39294 28810 39340
rect 28856 39294 28911 39340
rect 28492 39177 28911 39294
rect 28492 39131 28810 39177
rect 28856 39131 28911 39177
rect 28492 39013 28911 39131
rect 28492 38967 28810 39013
rect 28856 38967 28911 39013
rect 28492 38850 28911 38967
rect 37938 39750 38492 39769
rect 37938 39704 37957 39750
rect 38473 39704 38492 39750
rect 37938 39685 38492 39704
rect 40779 39750 42995 39810
rect 40779 39704 40836 39750
rect 40882 39704 40994 39750
rect 41040 39704 41152 39750
rect 41198 39704 41310 39750
rect 41356 39704 41469 39750
rect 41515 39704 41627 39750
rect 41673 39704 41785 39750
rect 41831 39704 41943 39750
rect 41989 39704 42101 39750
rect 42147 39704 42259 39750
rect 42305 39704 42418 39750
rect 42464 39704 42576 39750
rect 42622 39704 42734 39750
rect 42780 39704 42892 39750
rect 42938 39704 42995 39750
rect 40779 39644 42995 39704
rect 56212 40487 56632 40604
rect 56212 40441 56267 40487
rect 56313 40441 56632 40487
rect 56212 40323 56632 40441
rect 56212 40277 56267 40323
rect 56313 40277 56632 40323
rect 56212 40160 56632 40277
rect 56212 40114 56267 40160
rect 56313 40114 56632 40160
rect 56212 39997 56632 40114
rect 56212 39951 56267 39997
rect 56313 39951 56632 39997
rect 56212 39834 56632 39951
rect 56212 39788 56267 39834
rect 56313 39788 56632 39834
rect 28492 38804 28810 38850
rect 28856 38804 28911 38850
rect 28492 38687 28911 38804
rect 28492 38641 28810 38687
rect 28856 38641 28911 38687
rect 28492 38523 28911 38641
rect 28492 38477 28810 38523
rect 28856 38477 28911 38523
rect 28492 38360 28911 38477
rect 28492 38314 28810 38360
rect 28856 38314 28911 38360
rect 28492 38197 28911 38314
rect 28492 38151 28810 38197
rect 28856 38151 28911 38197
rect 28492 38034 28911 38151
rect 28492 37988 28810 38034
rect 28856 37988 28911 38034
rect 28492 37866 28911 37988
rect 34861 38850 35017 38907
rect 34861 38804 34916 38850
rect 34962 38804 35017 38850
rect 34861 38747 35017 38804
rect 50103 38850 50263 38910
rect 50103 38804 50160 38850
rect 50206 38804 50263 38850
rect 50103 38744 50263 38804
rect 56212 39666 56632 39788
rect 56212 39620 56267 39666
rect 56313 39620 56632 39666
rect 56212 39503 56632 39620
rect 56212 39457 56267 39503
rect 56313 39457 56632 39503
rect 56212 39340 56632 39457
rect 56212 39294 56267 39340
rect 56313 39294 56632 39340
rect 56212 39177 56632 39294
rect 56212 39131 56267 39177
rect 56313 39131 56632 39177
rect 56212 39013 56632 39131
rect 56212 38967 56267 39013
rect 56313 38967 56632 39013
rect 56212 38850 56632 38967
rect 56212 38804 56267 38850
rect 56313 38804 56632 38850
rect 28492 37820 28810 37866
rect 28856 37820 28911 37866
rect 28492 37703 28911 37820
rect 28492 37657 28810 37703
rect 28856 37657 28911 37703
rect 28492 37540 28911 37657
rect 28492 37494 28810 37540
rect 28856 37494 28911 37540
rect 28492 37377 28911 37494
rect 28492 37331 28810 37377
rect 28856 37331 28911 37377
rect 28492 37213 28911 37331
rect 28492 37167 28810 37213
rect 28856 37167 28911 37213
rect 28492 37050 28911 37167
rect 37938 37950 38492 37969
rect 37938 37904 37957 37950
rect 38473 37904 38492 37950
rect 37938 37885 38492 37904
rect 40779 37950 42995 38010
rect 40779 37904 40836 37950
rect 40882 37904 40994 37950
rect 41040 37904 41152 37950
rect 41198 37904 41310 37950
rect 41356 37904 41469 37950
rect 41515 37904 41627 37950
rect 41673 37904 41785 37950
rect 41831 37904 41943 37950
rect 41989 37904 42101 37950
rect 42147 37904 42259 37950
rect 42305 37904 42418 37950
rect 42464 37904 42576 37950
rect 42622 37904 42734 37950
rect 42780 37904 42892 37950
rect 42938 37904 42995 37950
rect 40779 37844 42995 37904
rect 56212 38687 56632 38804
rect 56212 38641 56267 38687
rect 56313 38641 56632 38687
rect 56212 38523 56632 38641
rect 56212 38477 56267 38523
rect 56313 38477 56632 38523
rect 56212 38360 56632 38477
rect 56212 38314 56267 38360
rect 56313 38314 56632 38360
rect 56212 38197 56632 38314
rect 56212 38151 56267 38197
rect 56313 38151 56632 38197
rect 56212 38034 56632 38151
rect 56212 37988 56267 38034
rect 56313 37988 56632 38034
rect 28492 37004 28810 37050
rect 28856 37004 28911 37050
rect 28492 36887 28911 37004
rect 28492 36841 28810 36887
rect 28856 36841 28911 36887
rect 28492 36723 28911 36841
rect 28492 36677 28810 36723
rect 28856 36677 28911 36723
rect 28492 36560 28911 36677
rect 28492 36514 28810 36560
rect 28856 36514 28911 36560
rect 28492 36397 28911 36514
rect 28492 36351 28810 36397
rect 28856 36351 28911 36397
rect 28492 36234 28911 36351
rect 28492 36188 28810 36234
rect 28856 36188 28911 36234
rect 28492 35996 28911 36188
rect 34861 37050 35017 37107
rect 34861 37004 34916 37050
rect 34962 37004 35017 37050
rect 34861 36947 35017 37004
rect 50103 37050 50263 37110
rect 50103 37004 50160 37050
rect 50206 37004 50263 37050
rect 50103 36944 50263 37004
rect 56212 37866 56632 37988
rect 56212 37820 56267 37866
rect 56313 37820 56632 37866
rect 56212 37703 56632 37820
rect 56212 37657 56267 37703
rect 56313 37657 56632 37703
rect 56212 37540 56632 37657
rect 56212 37494 56267 37540
rect 56313 37494 56632 37540
rect 56212 37377 56632 37494
rect 56212 37331 56267 37377
rect 56313 37331 56632 37377
rect 56212 37213 56632 37331
rect 56212 37167 56267 37213
rect 56313 37167 56632 37213
rect 56212 37050 56632 37167
rect 56212 37004 56267 37050
rect 56313 37004 56632 37050
rect 37938 36150 38492 36169
rect 37938 36104 37957 36150
rect 38473 36104 38492 36150
rect 37938 36085 38492 36104
rect 40779 36150 42995 36210
rect 40779 36104 40836 36150
rect 40882 36104 40994 36150
rect 41040 36104 41152 36150
rect 41198 36104 41310 36150
rect 41356 36104 41469 36150
rect 41515 36104 41627 36150
rect 41673 36104 41785 36150
rect 41831 36104 41943 36150
rect 41989 36104 42101 36150
rect 42147 36104 42259 36150
rect 42305 36104 42418 36150
rect 42464 36104 42576 36150
rect 42622 36104 42734 36150
rect 42780 36104 42892 36150
rect 42938 36104 42995 36150
rect 40779 36044 42995 36104
rect 56212 36887 56632 37004
rect 56212 36841 56267 36887
rect 56313 36841 56632 36887
rect 56212 36723 56632 36841
rect 56212 36677 56267 36723
rect 56313 36677 56632 36723
rect 56212 36560 56632 36677
rect 56212 36514 56267 36560
rect 56313 36514 56632 36560
rect 56212 36397 56632 36514
rect 56212 36351 56267 36397
rect 56313 36351 56632 36397
rect 56212 36234 56632 36351
rect 56212 36188 56267 36234
rect 56313 36188 56632 36234
rect 27744 35977 28911 35996
rect 56212 35996 56632 36188
rect 57278 35996 57380 45442
rect 56212 35977 57380 35996
rect 27744 34621 27763 35977
rect 57361 34621 57380 35977
rect 27744 34602 57380 34621
rect 27744 34256 27846 34602
rect 57292 34256 57380 34602
rect 27744 34237 57380 34256
rect 27744 1117 27763 34237
rect 50826 3890 56594 3909
rect 27479 1034 27763 1117
rect 28620 3869 40188 3888
rect 28620 3823 28639 3869
rect 28685 3823 28755 3869
rect 28801 3823 28871 3869
rect 28917 3823 28987 3869
rect 29033 3823 29103 3869
rect 29149 3823 29219 3869
rect 29265 3823 29335 3869
rect 29381 3823 29451 3869
rect 29497 3823 29567 3869
rect 29613 3823 29683 3869
rect 29729 3823 29799 3869
rect 29845 3823 29915 3869
rect 29961 3823 30031 3869
rect 30077 3823 30147 3869
rect 30193 3823 30263 3869
rect 30309 3823 30379 3869
rect 30425 3823 30495 3869
rect 30541 3823 30611 3869
rect 30657 3823 30727 3869
rect 30773 3823 30843 3869
rect 30889 3823 30959 3869
rect 31005 3823 31075 3869
rect 31121 3823 31191 3869
rect 31237 3823 31307 3869
rect 31353 3823 31423 3869
rect 31469 3823 31539 3869
rect 31585 3823 31655 3869
rect 31701 3823 31771 3869
rect 31817 3823 31887 3869
rect 31933 3823 32003 3869
rect 32049 3823 32119 3869
rect 32165 3823 32235 3869
rect 32281 3823 32351 3869
rect 32397 3823 32467 3869
rect 32513 3823 32583 3869
rect 32629 3823 32699 3869
rect 32745 3823 32815 3869
rect 32861 3823 32931 3869
rect 32977 3823 33047 3869
rect 33093 3823 33163 3869
rect 33209 3823 33279 3869
rect 33325 3823 33395 3869
rect 33441 3823 33511 3869
rect 33557 3823 33627 3869
rect 33673 3823 33743 3869
rect 33789 3823 33859 3869
rect 33905 3823 33975 3869
rect 34021 3823 34091 3869
rect 34137 3823 34207 3869
rect 34253 3823 34323 3869
rect 34369 3823 34439 3869
rect 34485 3823 34555 3869
rect 34601 3823 34671 3869
rect 34717 3823 34787 3869
rect 34833 3823 34903 3869
rect 34949 3823 35019 3869
rect 35065 3823 35135 3869
rect 35181 3823 35251 3869
rect 35297 3823 35367 3869
rect 35413 3823 35483 3869
rect 35529 3823 35599 3869
rect 35645 3823 35715 3869
rect 35761 3823 35831 3869
rect 35877 3823 35947 3869
rect 35993 3823 36063 3869
rect 36109 3823 36179 3869
rect 36225 3823 36295 3869
rect 36341 3823 36411 3869
rect 36457 3823 36527 3869
rect 36573 3823 36643 3869
rect 36689 3823 36759 3869
rect 36805 3823 36875 3869
rect 36921 3823 36991 3869
rect 37037 3823 37107 3869
rect 37153 3823 37223 3869
rect 37269 3823 37339 3869
rect 37385 3823 37455 3869
rect 37501 3823 37571 3869
rect 37617 3823 37687 3869
rect 37733 3823 37803 3869
rect 37849 3823 37919 3869
rect 37965 3823 38035 3869
rect 38081 3823 38151 3869
rect 38197 3823 38267 3869
rect 38313 3823 38383 3869
rect 38429 3823 38499 3869
rect 38545 3823 38615 3869
rect 38661 3823 38731 3869
rect 38777 3823 38847 3869
rect 38893 3823 38963 3869
rect 39009 3823 39079 3869
rect 39125 3823 39195 3869
rect 39241 3823 39311 3869
rect 39357 3823 39427 3869
rect 39473 3823 39543 3869
rect 39589 3823 39659 3869
rect 39705 3823 39775 3869
rect 39821 3823 39891 3869
rect 39937 3823 40007 3869
rect 40053 3823 40123 3869
rect 40169 3823 40188 3869
rect 28620 3753 40188 3823
rect 28620 3707 28639 3753
rect 28685 3707 28755 3753
rect 28801 3707 28871 3753
rect 28917 3707 28987 3753
rect 29033 3707 29103 3753
rect 29149 3707 29219 3753
rect 29265 3707 29335 3753
rect 29381 3707 29451 3753
rect 29497 3707 29567 3753
rect 29613 3707 29683 3753
rect 29729 3707 29799 3753
rect 29845 3707 29915 3753
rect 29961 3707 30031 3753
rect 30077 3707 30147 3753
rect 30193 3707 30263 3753
rect 30309 3707 30379 3753
rect 30425 3707 30495 3753
rect 30541 3707 30611 3753
rect 30657 3707 30727 3753
rect 30773 3707 30843 3753
rect 30889 3707 30959 3753
rect 31005 3707 31075 3753
rect 31121 3707 31191 3753
rect 31237 3707 31307 3753
rect 31353 3707 31423 3753
rect 31469 3707 31539 3753
rect 31585 3707 31655 3753
rect 31701 3707 31771 3753
rect 31817 3707 31887 3753
rect 31933 3707 32003 3753
rect 32049 3707 32119 3753
rect 32165 3707 32235 3753
rect 32281 3707 32351 3753
rect 32397 3707 32467 3753
rect 32513 3707 32583 3753
rect 32629 3707 32699 3753
rect 32745 3707 32815 3753
rect 32861 3707 32931 3753
rect 32977 3707 33047 3753
rect 33093 3707 33163 3753
rect 33209 3707 33279 3753
rect 33325 3707 33395 3753
rect 33441 3707 33511 3753
rect 33557 3707 33627 3753
rect 33673 3707 33743 3753
rect 33789 3707 33859 3753
rect 33905 3707 33975 3753
rect 34021 3707 34091 3753
rect 34137 3707 34207 3753
rect 34253 3707 34323 3753
rect 34369 3707 34439 3753
rect 34485 3707 34555 3753
rect 34601 3707 34671 3753
rect 34717 3707 34787 3753
rect 34833 3707 34903 3753
rect 34949 3707 35019 3753
rect 35065 3707 35135 3753
rect 35181 3707 35251 3753
rect 35297 3707 35367 3753
rect 35413 3707 35483 3753
rect 35529 3707 35599 3753
rect 35645 3707 35715 3753
rect 35761 3707 35831 3753
rect 35877 3707 35947 3753
rect 35993 3707 36063 3753
rect 36109 3707 36179 3753
rect 36225 3707 36295 3753
rect 36341 3707 36411 3753
rect 36457 3707 36527 3753
rect 36573 3707 36643 3753
rect 36689 3707 36759 3753
rect 36805 3707 36875 3753
rect 36921 3707 36991 3753
rect 37037 3707 37107 3753
rect 37153 3707 37223 3753
rect 37269 3707 37339 3753
rect 37385 3707 37455 3753
rect 37501 3707 37571 3753
rect 37617 3707 37687 3753
rect 37733 3707 37803 3753
rect 37849 3707 37919 3753
rect 37965 3707 38035 3753
rect 38081 3707 38151 3753
rect 38197 3707 38267 3753
rect 38313 3707 38383 3753
rect 38429 3707 38499 3753
rect 38545 3707 38615 3753
rect 38661 3707 38731 3753
rect 38777 3707 38847 3753
rect 38893 3707 38963 3753
rect 39009 3707 39079 3753
rect 39125 3707 39195 3753
rect 39241 3707 39311 3753
rect 39357 3707 39427 3753
rect 39473 3707 39543 3753
rect 39589 3707 39659 3753
rect 39705 3707 39775 3753
rect 39821 3707 39891 3753
rect 39937 3707 40007 3753
rect 40053 3707 40123 3753
rect 40169 3707 40188 3753
rect 28620 3637 40188 3707
rect 28620 3591 28639 3637
rect 28685 3591 28755 3637
rect 28801 3591 28871 3637
rect 28917 3591 28987 3637
rect 29033 3591 29103 3637
rect 29149 3591 29219 3637
rect 29265 3591 29335 3637
rect 29381 3591 29451 3637
rect 29497 3591 29567 3637
rect 29613 3591 29683 3637
rect 29729 3591 29799 3637
rect 29845 3591 29915 3637
rect 29961 3591 30031 3637
rect 30077 3591 30147 3637
rect 30193 3591 30263 3637
rect 30309 3591 30379 3637
rect 30425 3591 30495 3637
rect 30541 3591 30611 3637
rect 30657 3591 30727 3637
rect 30773 3591 30843 3637
rect 30889 3591 30959 3637
rect 31005 3591 31075 3637
rect 31121 3591 31191 3637
rect 31237 3591 31307 3637
rect 31353 3591 31423 3637
rect 31469 3591 31539 3637
rect 31585 3591 31655 3637
rect 31701 3591 31771 3637
rect 31817 3591 31887 3637
rect 31933 3591 32003 3637
rect 32049 3591 32119 3637
rect 32165 3591 32235 3637
rect 32281 3591 32351 3637
rect 32397 3591 32467 3637
rect 32513 3591 32583 3637
rect 32629 3591 32699 3637
rect 32745 3591 32815 3637
rect 32861 3591 32931 3637
rect 32977 3591 33047 3637
rect 33093 3591 33163 3637
rect 33209 3591 33279 3637
rect 33325 3591 33395 3637
rect 33441 3591 33511 3637
rect 33557 3591 33627 3637
rect 33673 3591 33743 3637
rect 33789 3591 33859 3637
rect 33905 3591 33975 3637
rect 34021 3591 34091 3637
rect 34137 3591 34207 3637
rect 34253 3591 34323 3637
rect 34369 3591 34439 3637
rect 34485 3591 34555 3637
rect 34601 3591 34671 3637
rect 34717 3591 34787 3637
rect 34833 3591 34903 3637
rect 34949 3591 35019 3637
rect 35065 3591 35135 3637
rect 35181 3591 35251 3637
rect 35297 3591 35367 3637
rect 35413 3591 35483 3637
rect 35529 3591 35599 3637
rect 35645 3591 35715 3637
rect 35761 3591 35831 3637
rect 35877 3591 35947 3637
rect 35993 3591 36063 3637
rect 36109 3591 36179 3637
rect 36225 3591 36295 3637
rect 36341 3591 36411 3637
rect 36457 3591 36527 3637
rect 36573 3591 36643 3637
rect 36689 3591 36759 3637
rect 36805 3591 36875 3637
rect 36921 3591 36991 3637
rect 37037 3591 37107 3637
rect 37153 3591 37223 3637
rect 37269 3591 37339 3637
rect 37385 3591 37455 3637
rect 37501 3591 37571 3637
rect 37617 3591 37687 3637
rect 37733 3591 37803 3637
rect 37849 3591 37919 3637
rect 37965 3591 38035 3637
rect 38081 3591 38151 3637
rect 38197 3591 38267 3637
rect 38313 3591 38383 3637
rect 38429 3591 38499 3637
rect 38545 3591 38615 3637
rect 38661 3591 38731 3637
rect 38777 3591 38847 3637
rect 38893 3591 38963 3637
rect 39009 3591 39079 3637
rect 39125 3591 39195 3637
rect 39241 3591 39311 3637
rect 39357 3591 39427 3637
rect 39473 3591 39543 3637
rect 39589 3591 39659 3637
rect 39705 3591 39775 3637
rect 39821 3591 39891 3637
rect 39937 3591 40007 3637
rect 40053 3591 40123 3637
rect 40169 3591 40188 3637
rect 28620 3521 40188 3591
rect 28620 3475 28639 3521
rect 28685 3475 28755 3521
rect 28801 3475 28871 3521
rect 28917 3475 28987 3521
rect 29033 3475 29103 3521
rect 29149 3475 29219 3521
rect 29265 3475 29335 3521
rect 29381 3475 29451 3521
rect 29497 3475 29567 3521
rect 29613 3475 29683 3521
rect 29729 3475 29799 3521
rect 29845 3475 29915 3521
rect 29961 3475 30031 3521
rect 30077 3475 30147 3521
rect 30193 3475 30263 3521
rect 30309 3475 30379 3521
rect 30425 3475 30495 3521
rect 30541 3475 30611 3521
rect 30657 3475 30727 3521
rect 30773 3475 30843 3521
rect 30889 3475 30959 3521
rect 31005 3475 31075 3521
rect 31121 3475 31191 3521
rect 31237 3475 31307 3521
rect 31353 3475 31423 3521
rect 31469 3475 31539 3521
rect 31585 3475 31655 3521
rect 31701 3475 31771 3521
rect 31817 3475 31887 3521
rect 31933 3475 32003 3521
rect 32049 3475 32119 3521
rect 32165 3475 32235 3521
rect 32281 3475 32351 3521
rect 32397 3475 32467 3521
rect 32513 3475 32583 3521
rect 32629 3475 32699 3521
rect 32745 3475 32815 3521
rect 32861 3475 32931 3521
rect 32977 3475 33047 3521
rect 33093 3475 33163 3521
rect 33209 3475 33279 3521
rect 33325 3475 33395 3521
rect 33441 3475 33511 3521
rect 33557 3475 33627 3521
rect 33673 3475 33743 3521
rect 33789 3475 33859 3521
rect 33905 3475 33975 3521
rect 34021 3475 34091 3521
rect 34137 3475 34207 3521
rect 34253 3475 34323 3521
rect 34369 3475 34439 3521
rect 34485 3475 34555 3521
rect 34601 3475 34671 3521
rect 34717 3475 34787 3521
rect 34833 3475 34903 3521
rect 34949 3475 35019 3521
rect 35065 3475 35135 3521
rect 35181 3475 35251 3521
rect 35297 3475 35367 3521
rect 35413 3475 35483 3521
rect 35529 3475 35599 3521
rect 35645 3475 35715 3521
rect 35761 3475 35831 3521
rect 35877 3475 35947 3521
rect 35993 3475 36063 3521
rect 36109 3475 36179 3521
rect 36225 3475 36295 3521
rect 36341 3475 36411 3521
rect 36457 3475 36527 3521
rect 36573 3475 36643 3521
rect 36689 3475 36759 3521
rect 36805 3475 36875 3521
rect 36921 3475 36991 3521
rect 37037 3475 37107 3521
rect 37153 3475 37223 3521
rect 37269 3475 37339 3521
rect 37385 3475 37455 3521
rect 37501 3475 37571 3521
rect 37617 3475 37687 3521
rect 37733 3475 37803 3521
rect 37849 3475 37919 3521
rect 37965 3475 38035 3521
rect 38081 3475 38151 3521
rect 38197 3475 38267 3521
rect 38313 3475 38383 3521
rect 38429 3475 38499 3521
rect 38545 3475 38615 3521
rect 38661 3475 38731 3521
rect 38777 3475 38847 3521
rect 38893 3475 38963 3521
rect 39009 3475 39079 3521
rect 39125 3475 39195 3521
rect 39241 3475 39311 3521
rect 39357 3475 39427 3521
rect 39473 3475 39543 3521
rect 39589 3475 39659 3521
rect 39705 3475 39775 3521
rect 39821 3475 39891 3521
rect 39937 3475 40007 3521
rect 40053 3475 40123 3521
rect 40169 3475 40188 3521
rect 28620 3405 40188 3475
rect 28620 3359 28639 3405
rect 28685 3359 28755 3405
rect 28801 3359 28871 3405
rect 28917 3359 28987 3405
rect 29033 3359 29103 3405
rect 29149 3359 29219 3405
rect 29265 3359 29335 3405
rect 29381 3359 29451 3405
rect 29497 3359 29567 3405
rect 29613 3359 29683 3405
rect 29729 3359 29799 3405
rect 29845 3359 29915 3405
rect 29961 3359 30031 3405
rect 30077 3359 30147 3405
rect 30193 3359 30263 3405
rect 30309 3359 30379 3405
rect 30425 3359 30495 3405
rect 30541 3359 30611 3405
rect 30657 3359 30727 3405
rect 30773 3359 30843 3405
rect 30889 3359 30959 3405
rect 31005 3359 31075 3405
rect 31121 3359 31191 3405
rect 31237 3359 31307 3405
rect 31353 3359 31423 3405
rect 31469 3359 31539 3405
rect 31585 3359 31655 3405
rect 31701 3359 31771 3405
rect 31817 3359 31887 3405
rect 31933 3359 32003 3405
rect 32049 3359 32119 3405
rect 32165 3359 32235 3405
rect 32281 3359 32351 3405
rect 32397 3359 32467 3405
rect 32513 3359 32583 3405
rect 32629 3359 32699 3405
rect 32745 3359 32815 3405
rect 32861 3359 32931 3405
rect 32977 3359 33047 3405
rect 33093 3359 33163 3405
rect 33209 3359 33279 3405
rect 33325 3359 33395 3405
rect 33441 3359 33511 3405
rect 33557 3359 33627 3405
rect 33673 3359 33743 3405
rect 33789 3359 33859 3405
rect 33905 3359 33975 3405
rect 34021 3359 34091 3405
rect 34137 3359 34207 3405
rect 34253 3359 34323 3405
rect 34369 3359 34439 3405
rect 34485 3359 34555 3405
rect 34601 3359 34671 3405
rect 34717 3359 34787 3405
rect 34833 3359 34903 3405
rect 34949 3359 35019 3405
rect 35065 3359 35135 3405
rect 35181 3359 35251 3405
rect 35297 3359 35367 3405
rect 35413 3359 35483 3405
rect 35529 3359 35599 3405
rect 35645 3359 35715 3405
rect 35761 3359 35831 3405
rect 35877 3359 35947 3405
rect 35993 3359 36063 3405
rect 36109 3359 36179 3405
rect 36225 3359 36295 3405
rect 36341 3359 36411 3405
rect 36457 3359 36527 3405
rect 36573 3359 36643 3405
rect 36689 3359 36759 3405
rect 36805 3359 36875 3405
rect 36921 3359 36991 3405
rect 37037 3359 37107 3405
rect 37153 3359 37223 3405
rect 37269 3359 37339 3405
rect 37385 3359 37455 3405
rect 37501 3359 37571 3405
rect 37617 3359 37687 3405
rect 37733 3359 37803 3405
rect 37849 3359 37919 3405
rect 37965 3359 38035 3405
rect 38081 3359 38151 3405
rect 38197 3359 38267 3405
rect 38313 3359 38383 3405
rect 38429 3359 38499 3405
rect 38545 3359 38615 3405
rect 38661 3359 38731 3405
rect 38777 3359 38847 3405
rect 38893 3359 38963 3405
rect 39009 3359 39079 3405
rect 39125 3359 39195 3405
rect 39241 3359 39311 3405
rect 39357 3359 39427 3405
rect 39473 3359 39543 3405
rect 39589 3359 39659 3405
rect 39705 3359 39775 3405
rect 39821 3359 39891 3405
rect 39937 3359 40007 3405
rect 40053 3359 40123 3405
rect 40169 3359 40188 3405
rect 28620 3289 40188 3359
rect 28620 3243 28639 3289
rect 28685 3243 28755 3289
rect 28801 3243 28871 3289
rect 28917 3243 28987 3289
rect 29033 3243 29103 3289
rect 29149 3243 29219 3289
rect 29265 3243 29335 3289
rect 29381 3243 29451 3289
rect 29497 3243 29567 3289
rect 29613 3243 29683 3289
rect 29729 3243 29799 3289
rect 29845 3243 29915 3289
rect 29961 3243 30031 3289
rect 30077 3243 30147 3289
rect 30193 3243 30263 3289
rect 30309 3243 30379 3289
rect 30425 3243 30495 3289
rect 30541 3243 30611 3289
rect 30657 3243 30727 3289
rect 30773 3243 30843 3289
rect 30889 3243 30959 3289
rect 31005 3243 31075 3289
rect 31121 3243 31191 3289
rect 31237 3243 31307 3289
rect 31353 3243 31423 3289
rect 31469 3243 31539 3289
rect 31585 3243 31655 3289
rect 31701 3243 31771 3289
rect 31817 3243 31887 3289
rect 31933 3243 32003 3289
rect 32049 3243 32119 3289
rect 32165 3243 32235 3289
rect 32281 3243 32351 3289
rect 32397 3243 32467 3289
rect 32513 3243 32583 3289
rect 32629 3243 32699 3289
rect 32745 3243 32815 3289
rect 32861 3243 32931 3289
rect 32977 3243 33047 3289
rect 33093 3243 33163 3289
rect 33209 3243 33279 3289
rect 33325 3243 33395 3289
rect 33441 3243 33511 3289
rect 33557 3243 33627 3289
rect 33673 3243 33743 3289
rect 33789 3243 33859 3289
rect 33905 3243 33975 3289
rect 34021 3243 34091 3289
rect 34137 3243 34207 3289
rect 34253 3243 34323 3289
rect 34369 3243 34439 3289
rect 34485 3243 34555 3289
rect 34601 3243 34671 3289
rect 34717 3243 34787 3289
rect 34833 3243 34903 3289
rect 34949 3243 35019 3289
rect 35065 3243 35135 3289
rect 35181 3243 35251 3289
rect 35297 3243 35367 3289
rect 35413 3243 35483 3289
rect 35529 3243 35599 3289
rect 35645 3243 35715 3289
rect 35761 3243 35831 3289
rect 35877 3243 35947 3289
rect 35993 3243 36063 3289
rect 36109 3243 36179 3289
rect 36225 3243 36295 3289
rect 36341 3243 36411 3289
rect 36457 3243 36527 3289
rect 36573 3243 36643 3289
rect 36689 3243 36759 3289
rect 36805 3243 36875 3289
rect 36921 3243 36991 3289
rect 37037 3243 37107 3289
rect 37153 3243 37223 3289
rect 37269 3243 37339 3289
rect 37385 3243 37455 3289
rect 37501 3243 37571 3289
rect 37617 3243 37687 3289
rect 37733 3243 37803 3289
rect 37849 3243 37919 3289
rect 37965 3243 38035 3289
rect 38081 3243 38151 3289
rect 38197 3243 38267 3289
rect 38313 3243 38383 3289
rect 38429 3243 38499 3289
rect 38545 3243 38615 3289
rect 38661 3243 38731 3289
rect 38777 3243 38847 3289
rect 38893 3243 38963 3289
rect 39009 3243 39079 3289
rect 39125 3243 39195 3289
rect 39241 3243 39311 3289
rect 39357 3243 39427 3289
rect 39473 3243 39543 3289
rect 39589 3243 39659 3289
rect 39705 3243 39775 3289
rect 39821 3243 39891 3289
rect 39937 3243 40007 3289
rect 40053 3243 40123 3289
rect 40169 3243 40188 3289
rect 28620 3173 40188 3243
rect 28620 3127 28639 3173
rect 28685 3127 28755 3173
rect 28801 3127 28871 3173
rect 28917 3127 28987 3173
rect 29033 3127 29103 3173
rect 29149 3127 29219 3173
rect 29265 3127 29335 3173
rect 29381 3127 29451 3173
rect 29497 3127 29567 3173
rect 29613 3127 29683 3173
rect 29729 3127 29799 3173
rect 29845 3127 29915 3173
rect 29961 3127 30031 3173
rect 30077 3127 30147 3173
rect 30193 3127 30263 3173
rect 30309 3127 30379 3173
rect 30425 3127 30495 3173
rect 30541 3127 30611 3173
rect 30657 3127 30727 3173
rect 30773 3127 30843 3173
rect 30889 3127 30959 3173
rect 31005 3127 31075 3173
rect 31121 3127 31191 3173
rect 31237 3127 31307 3173
rect 31353 3127 31423 3173
rect 31469 3127 31539 3173
rect 31585 3127 31655 3173
rect 31701 3127 31771 3173
rect 31817 3127 31887 3173
rect 31933 3127 32003 3173
rect 32049 3127 32119 3173
rect 32165 3127 32235 3173
rect 32281 3127 32351 3173
rect 32397 3127 32467 3173
rect 32513 3127 32583 3173
rect 32629 3127 32699 3173
rect 32745 3127 32815 3173
rect 32861 3127 32931 3173
rect 32977 3127 33047 3173
rect 33093 3127 33163 3173
rect 33209 3127 33279 3173
rect 33325 3127 33395 3173
rect 33441 3127 33511 3173
rect 33557 3127 33627 3173
rect 33673 3127 33743 3173
rect 33789 3127 33859 3173
rect 33905 3127 33975 3173
rect 34021 3127 34091 3173
rect 34137 3127 34207 3173
rect 34253 3127 34323 3173
rect 34369 3127 34439 3173
rect 34485 3127 34555 3173
rect 34601 3127 34671 3173
rect 34717 3127 34787 3173
rect 34833 3127 34903 3173
rect 34949 3127 35019 3173
rect 35065 3127 35135 3173
rect 35181 3127 35251 3173
rect 35297 3127 35367 3173
rect 35413 3127 35483 3173
rect 35529 3127 35599 3173
rect 35645 3127 35715 3173
rect 35761 3127 35831 3173
rect 35877 3127 35947 3173
rect 35993 3127 36063 3173
rect 36109 3127 36179 3173
rect 36225 3127 36295 3173
rect 36341 3127 36411 3173
rect 36457 3127 36527 3173
rect 36573 3127 36643 3173
rect 36689 3127 36759 3173
rect 36805 3127 36875 3173
rect 36921 3127 36991 3173
rect 37037 3127 37107 3173
rect 37153 3127 37223 3173
rect 37269 3127 37339 3173
rect 37385 3127 37455 3173
rect 37501 3127 37571 3173
rect 37617 3127 37687 3173
rect 37733 3127 37803 3173
rect 37849 3127 37919 3173
rect 37965 3127 38035 3173
rect 38081 3127 38151 3173
rect 38197 3127 38267 3173
rect 38313 3127 38383 3173
rect 38429 3127 38499 3173
rect 38545 3127 38615 3173
rect 38661 3127 38731 3173
rect 38777 3127 38847 3173
rect 38893 3127 38963 3173
rect 39009 3127 39079 3173
rect 39125 3127 39195 3173
rect 39241 3127 39311 3173
rect 39357 3127 39427 3173
rect 39473 3127 39543 3173
rect 39589 3127 39659 3173
rect 39705 3127 39775 3173
rect 39821 3127 39891 3173
rect 39937 3127 40007 3173
rect 40053 3127 40123 3173
rect 40169 3127 40188 3173
rect 28620 3057 40188 3127
rect 28620 3011 28639 3057
rect 28685 3011 28755 3057
rect 28801 3011 28871 3057
rect 28917 3011 28987 3057
rect 29033 3011 29103 3057
rect 29149 3011 29219 3057
rect 29265 3011 29335 3057
rect 29381 3011 29451 3057
rect 29497 3011 29567 3057
rect 29613 3011 29683 3057
rect 29729 3011 29799 3057
rect 29845 3011 29915 3057
rect 29961 3011 30031 3057
rect 30077 3011 30147 3057
rect 30193 3011 30263 3057
rect 30309 3011 30379 3057
rect 30425 3011 30495 3057
rect 30541 3011 30611 3057
rect 30657 3011 30727 3057
rect 30773 3011 30843 3057
rect 30889 3011 30959 3057
rect 31005 3011 31075 3057
rect 31121 3011 31191 3057
rect 31237 3011 31307 3057
rect 31353 3011 31423 3057
rect 31469 3011 31539 3057
rect 31585 3011 31655 3057
rect 31701 3011 31771 3057
rect 31817 3011 31887 3057
rect 31933 3011 32003 3057
rect 32049 3011 32119 3057
rect 32165 3011 32235 3057
rect 32281 3011 32351 3057
rect 32397 3011 32467 3057
rect 32513 3011 32583 3057
rect 32629 3011 32699 3057
rect 32745 3011 32815 3057
rect 32861 3011 32931 3057
rect 32977 3011 33047 3057
rect 33093 3011 33163 3057
rect 33209 3011 33279 3057
rect 33325 3011 33395 3057
rect 33441 3011 33511 3057
rect 33557 3011 33627 3057
rect 33673 3011 33743 3057
rect 33789 3011 33859 3057
rect 33905 3011 33975 3057
rect 34021 3011 34091 3057
rect 34137 3011 34207 3057
rect 34253 3011 34323 3057
rect 34369 3011 34439 3057
rect 34485 3011 34555 3057
rect 34601 3011 34671 3057
rect 34717 3011 34787 3057
rect 34833 3011 34903 3057
rect 34949 3011 35019 3057
rect 35065 3011 35135 3057
rect 35181 3011 35251 3057
rect 35297 3011 35367 3057
rect 35413 3011 35483 3057
rect 35529 3011 35599 3057
rect 35645 3011 35715 3057
rect 35761 3011 35831 3057
rect 35877 3011 35947 3057
rect 35993 3011 36063 3057
rect 36109 3011 36179 3057
rect 36225 3011 36295 3057
rect 36341 3011 36411 3057
rect 36457 3011 36527 3057
rect 36573 3011 36643 3057
rect 36689 3011 36759 3057
rect 36805 3011 36875 3057
rect 36921 3011 36991 3057
rect 37037 3011 37107 3057
rect 37153 3011 37223 3057
rect 37269 3011 37339 3057
rect 37385 3011 37455 3057
rect 37501 3011 37571 3057
rect 37617 3011 37687 3057
rect 37733 3011 37803 3057
rect 37849 3011 37919 3057
rect 37965 3011 38035 3057
rect 38081 3011 38151 3057
rect 38197 3011 38267 3057
rect 38313 3011 38383 3057
rect 38429 3011 38499 3057
rect 38545 3011 38615 3057
rect 38661 3011 38731 3057
rect 38777 3011 38847 3057
rect 38893 3011 38963 3057
rect 39009 3011 39079 3057
rect 39125 3011 39195 3057
rect 39241 3011 39311 3057
rect 39357 3011 39427 3057
rect 39473 3011 39543 3057
rect 39589 3011 39659 3057
rect 39705 3011 39775 3057
rect 39821 3011 39891 3057
rect 39937 3011 40007 3057
rect 40053 3011 40123 3057
rect 40169 3011 40188 3057
rect 28620 2941 40188 3011
rect 28620 2895 28639 2941
rect 28685 2895 28755 2941
rect 28801 2895 28871 2941
rect 28917 2895 28987 2941
rect 29033 2895 29103 2941
rect 29149 2895 29219 2941
rect 29265 2895 29335 2941
rect 29381 2895 29451 2941
rect 29497 2895 29567 2941
rect 29613 2895 29683 2941
rect 29729 2895 29799 2941
rect 29845 2895 29915 2941
rect 29961 2895 30031 2941
rect 30077 2895 30147 2941
rect 30193 2895 30263 2941
rect 30309 2895 30379 2941
rect 30425 2895 30495 2941
rect 30541 2895 30611 2941
rect 30657 2895 30727 2941
rect 30773 2895 30843 2941
rect 30889 2895 30959 2941
rect 31005 2895 31075 2941
rect 31121 2895 31191 2941
rect 31237 2895 31307 2941
rect 31353 2895 31423 2941
rect 31469 2895 31539 2941
rect 31585 2895 31655 2941
rect 31701 2895 31771 2941
rect 31817 2895 31887 2941
rect 31933 2895 32003 2941
rect 32049 2895 32119 2941
rect 32165 2895 32235 2941
rect 32281 2895 32351 2941
rect 32397 2895 32467 2941
rect 32513 2895 32583 2941
rect 32629 2895 32699 2941
rect 32745 2895 32815 2941
rect 32861 2895 32931 2941
rect 32977 2895 33047 2941
rect 33093 2895 33163 2941
rect 33209 2895 33279 2941
rect 33325 2895 33395 2941
rect 33441 2895 33511 2941
rect 33557 2895 33627 2941
rect 33673 2895 33743 2941
rect 33789 2895 33859 2941
rect 33905 2895 33975 2941
rect 34021 2895 34091 2941
rect 34137 2895 34207 2941
rect 34253 2895 34323 2941
rect 34369 2895 34439 2941
rect 34485 2895 34555 2941
rect 34601 2895 34671 2941
rect 34717 2895 34787 2941
rect 34833 2895 34903 2941
rect 34949 2895 35019 2941
rect 35065 2895 35135 2941
rect 35181 2895 35251 2941
rect 35297 2895 35367 2941
rect 35413 2895 35483 2941
rect 35529 2895 35599 2941
rect 35645 2895 35715 2941
rect 35761 2895 35831 2941
rect 35877 2895 35947 2941
rect 35993 2895 36063 2941
rect 36109 2895 36179 2941
rect 36225 2895 36295 2941
rect 36341 2895 36411 2941
rect 36457 2895 36527 2941
rect 36573 2895 36643 2941
rect 36689 2895 36759 2941
rect 36805 2895 36875 2941
rect 36921 2895 36991 2941
rect 37037 2895 37107 2941
rect 37153 2895 37223 2941
rect 37269 2895 37339 2941
rect 37385 2895 37455 2941
rect 37501 2895 37571 2941
rect 37617 2895 37687 2941
rect 37733 2895 37803 2941
rect 37849 2895 37919 2941
rect 37965 2895 38035 2941
rect 38081 2895 38151 2941
rect 38197 2895 38267 2941
rect 38313 2895 38383 2941
rect 38429 2895 38499 2941
rect 38545 2895 38615 2941
rect 38661 2895 38731 2941
rect 38777 2895 38847 2941
rect 38893 2895 38963 2941
rect 39009 2895 39079 2941
rect 39125 2895 39195 2941
rect 39241 2895 39311 2941
rect 39357 2895 39427 2941
rect 39473 2895 39543 2941
rect 39589 2895 39659 2941
rect 39705 2895 39775 2941
rect 39821 2895 39891 2941
rect 39937 2895 40007 2941
rect 40053 2895 40123 2941
rect 40169 2895 40188 2941
rect 28620 2825 40188 2895
rect 28620 2779 28639 2825
rect 28685 2779 28755 2825
rect 28801 2779 28871 2825
rect 28917 2779 28987 2825
rect 29033 2779 29103 2825
rect 29149 2779 29219 2825
rect 29265 2779 29335 2825
rect 29381 2779 29451 2825
rect 29497 2779 29567 2825
rect 29613 2779 29683 2825
rect 29729 2779 29799 2825
rect 29845 2779 29915 2825
rect 29961 2779 30031 2825
rect 30077 2779 30147 2825
rect 30193 2779 30263 2825
rect 30309 2779 30379 2825
rect 30425 2779 30495 2825
rect 30541 2779 30611 2825
rect 30657 2779 30727 2825
rect 30773 2779 30843 2825
rect 30889 2779 30959 2825
rect 31005 2779 31075 2825
rect 31121 2779 31191 2825
rect 31237 2779 31307 2825
rect 31353 2779 31423 2825
rect 31469 2779 31539 2825
rect 31585 2779 31655 2825
rect 31701 2779 31771 2825
rect 31817 2779 31887 2825
rect 31933 2779 32003 2825
rect 32049 2779 32119 2825
rect 32165 2779 32235 2825
rect 32281 2779 32351 2825
rect 32397 2779 32467 2825
rect 32513 2779 32583 2825
rect 32629 2779 32699 2825
rect 32745 2779 32815 2825
rect 32861 2779 32931 2825
rect 32977 2779 33047 2825
rect 33093 2779 33163 2825
rect 33209 2779 33279 2825
rect 33325 2779 33395 2825
rect 33441 2779 33511 2825
rect 33557 2779 33627 2825
rect 33673 2779 33743 2825
rect 33789 2779 33859 2825
rect 33905 2779 33975 2825
rect 34021 2779 34091 2825
rect 34137 2779 34207 2825
rect 34253 2779 34323 2825
rect 34369 2779 34439 2825
rect 34485 2779 34555 2825
rect 34601 2779 34671 2825
rect 34717 2779 34787 2825
rect 34833 2779 34903 2825
rect 34949 2779 35019 2825
rect 35065 2779 35135 2825
rect 35181 2779 35251 2825
rect 35297 2779 35367 2825
rect 35413 2779 35483 2825
rect 35529 2779 35599 2825
rect 35645 2779 35715 2825
rect 35761 2779 35831 2825
rect 35877 2779 35947 2825
rect 35993 2779 36063 2825
rect 36109 2779 36179 2825
rect 36225 2779 36295 2825
rect 36341 2779 36411 2825
rect 36457 2779 36527 2825
rect 36573 2779 36643 2825
rect 36689 2779 36759 2825
rect 36805 2779 36875 2825
rect 36921 2779 36991 2825
rect 37037 2779 37107 2825
rect 37153 2779 37223 2825
rect 37269 2779 37339 2825
rect 37385 2779 37455 2825
rect 37501 2779 37571 2825
rect 37617 2779 37687 2825
rect 37733 2779 37803 2825
rect 37849 2779 37919 2825
rect 37965 2779 38035 2825
rect 38081 2779 38151 2825
rect 38197 2779 38267 2825
rect 38313 2779 38383 2825
rect 38429 2779 38499 2825
rect 38545 2779 38615 2825
rect 38661 2779 38731 2825
rect 38777 2779 38847 2825
rect 38893 2779 38963 2825
rect 39009 2779 39079 2825
rect 39125 2779 39195 2825
rect 39241 2779 39311 2825
rect 39357 2779 39427 2825
rect 39473 2779 39543 2825
rect 39589 2779 39659 2825
rect 39705 2779 39775 2825
rect 39821 2779 39891 2825
rect 39937 2779 40007 2825
rect 40053 2779 40123 2825
rect 40169 2779 40188 2825
rect 28620 2709 40188 2779
rect 28620 2663 28639 2709
rect 28685 2663 28755 2709
rect 28801 2663 28871 2709
rect 28917 2663 28987 2709
rect 29033 2663 29103 2709
rect 29149 2663 29219 2709
rect 29265 2663 29335 2709
rect 29381 2663 29451 2709
rect 29497 2663 29567 2709
rect 29613 2663 29683 2709
rect 29729 2663 29799 2709
rect 29845 2663 29915 2709
rect 29961 2663 30031 2709
rect 30077 2663 30147 2709
rect 30193 2663 30263 2709
rect 30309 2663 30379 2709
rect 30425 2663 30495 2709
rect 30541 2663 30611 2709
rect 30657 2663 30727 2709
rect 30773 2663 30843 2709
rect 30889 2663 30959 2709
rect 31005 2663 31075 2709
rect 31121 2663 31191 2709
rect 31237 2663 31307 2709
rect 31353 2663 31423 2709
rect 31469 2663 31539 2709
rect 31585 2663 31655 2709
rect 31701 2663 31771 2709
rect 31817 2663 31887 2709
rect 31933 2663 32003 2709
rect 32049 2663 32119 2709
rect 32165 2663 32235 2709
rect 32281 2663 32351 2709
rect 32397 2663 32467 2709
rect 32513 2663 32583 2709
rect 32629 2663 32699 2709
rect 32745 2663 32815 2709
rect 32861 2663 32931 2709
rect 32977 2663 33047 2709
rect 33093 2663 33163 2709
rect 33209 2663 33279 2709
rect 33325 2663 33395 2709
rect 33441 2663 33511 2709
rect 33557 2663 33627 2709
rect 33673 2663 33743 2709
rect 33789 2663 33859 2709
rect 33905 2663 33975 2709
rect 34021 2663 34091 2709
rect 34137 2663 34207 2709
rect 34253 2663 34323 2709
rect 34369 2663 34439 2709
rect 34485 2663 34555 2709
rect 34601 2663 34671 2709
rect 34717 2663 34787 2709
rect 34833 2663 34903 2709
rect 34949 2663 35019 2709
rect 35065 2663 35135 2709
rect 35181 2663 35251 2709
rect 35297 2663 35367 2709
rect 35413 2663 35483 2709
rect 35529 2663 35599 2709
rect 35645 2663 35715 2709
rect 35761 2663 35831 2709
rect 35877 2663 35947 2709
rect 35993 2663 36063 2709
rect 36109 2663 36179 2709
rect 36225 2663 36295 2709
rect 36341 2663 36411 2709
rect 36457 2663 36527 2709
rect 36573 2663 36643 2709
rect 36689 2663 36759 2709
rect 36805 2663 36875 2709
rect 36921 2663 36991 2709
rect 37037 2663 37107 2709
rect 37153 2663 37223 2709
rect 37269 2663 37339 2709
rect 37385 2663 37455 2709
rect 37501 2663 37571 2709
rect 37617 2663 37687 2709
rect 37733 2663 37803 2709
rect 37849 2663 37919 2709
rect 37965 2663 38035 2709
rect 38081 2663 38151 2709
rect 38197 2663 38267 2709
rect 38313 2663 38383 2709
rect 38429 2663 38499 2709
rect 38545 2663 38615 2709
rect 38661 2663 38731 2709
rect 38777 2663 38847 2709
rect 38893 2663 38963 2709
rect 39009 2663 39079 2709
rect 39125 2663 39195 2709
rect 39241 2663 39311 2709
rect 39357 2663 39427 2709
rect 39473 2663 39543 2709
rect 39589 2663 39659 2709
rect 39705 2663 39775 2709
rect 39821 2663 39891 2709
rect 39937 2663 40007 2709
rect 40053 2663 40123 2709
rect 40169 2663 40188 2709
rect 28620 2593 40188 2663
rect 28620 2547 28639 2593
rect 28685 2547 28755 2593
rect 28801 2547 28871 2593
rect 28917 2547 28987 2593
rect 29033 2547 29103 2593
rect 29149 2547 29219 2593
rect 29265 2547 29335 2593
rect 29381 2547 29451 2593
rect 29497 2547 29567 2593
rect 29613 2547 29683 2593
rect 29729 2547 29799 2593
rect 29845 2547 29915 2593
rect 29961 2547 30031 2593
rect 30077 2547 30147 2593
rect 30193 2547 30263 2593
rect 30309 2547 30379 2593
rect 30425 2547 30495 2593
rect 30541 2547 30611 2593
rect 30657 2547 30727 2593
rect 30773 2547 30843 2593
rect 30889 2547 30959 2593
rect 31005 2547 31075 2593
rect 31121 2547 31191 2593
rect 31237 2547 31307 2593
rect 31353 2547 31423 2593
rect 31469 2547 31539 2593
rect 31585 2547 31655 2593
rect 31701 2547 31771 2593
rect 31817 2547 31887 2593
rect 31933 2547 32003 2593
rect 32049 2547 32119 2593
rect 32165 2547 32235 2593
rect 32281 2547 32351 2593
rect 32397 2547 32467 2593
rect 32513 2547 32583 2593
rect 32629 2547 32699 2593
rect 32745 2547 32815 2593
rect 32861 2547 32931 2593
rect 32977 2547 33047 2593
rect 33093 2547 33163 2593
rect 33209 2547 33279 2593
rect 33325 2547 33395 2593
rect 33441 2547 33511 2593
rect 33557 2547 33627 2593
rect 33673 2547 33743 2593
rect 33789 2547 33859 2593
rect 33905 2547 33975 2593
rect 34021 2547 34091 2593
rect 34137 2547 34207 2593
rect 34253 2547 34323 2593
rect 34369 2547 34439 2593
rect 34485 2547 34555 2593
rect 34601 2547 34671 2593
rect 34717 2547 34787 2593
rect 34833 2547 34903 2593
rect 34949 2547 35019 2593
rect 35065 2547 35135 2593
rect 35181 2547 35251 2593
rect 35297 2547 35367 2593
rect 35413 2547 35483 2593
rect 35529 2547 35599 2593
rect 35645 2547 35715 2593
rect 35761 2547 35831 2593
rect 35877 2547 35947 2593
rect 35993 2547 36063 2593
rect 36109 2547 36179 2593
rect 36225 2547 36295 2593
rect 36341 2547 36411 2593
rect 36457 2547 36527 2593
rect 36573 2547 36643 2593
rect 36689 2547 36759 2593
rect 36805 2547 36875 2593
rect 36921 2547 36991 2593
rect 37037 2547 37107 2593
rect 37153 2547 37223 2593
rect 37269 2547 37339 2593
rect 37385 2547 37455 2593
rect 37501 2547 37571 2593
rect 37617 2547 37687 2593
rect 37733 2547 37803 2593
rect 37849 2547 37919 2593
rect 37965 2547 38035 2593
rect 38081 2547 38151 2593
rect 38197 2547 38267 2593
rect 38313 2547 38383 2593
rect 38429 2547 38499 2593
rect 38545 2547 38615 2593
rect 38661 2547 38731 2593
rect 38777 2547 38847 2593
rect 38893 2547 38963 2593
rect 39009 2547 39079 2593
rect 39125 2547 39195 2593
rect 39241 2547 39311 2593
rect 39357 2547 39427 2593
rect 39473 2547 39543 2593
rect 39589 2547 39659 2593
rect 39705 2547 39775 2593
rect 39821 2547 39891 2593
rect 39937 2547 40007 2593
rect 40053 2547 40123 2593
rect 40169 2547 40188 2593
rect 28620 2477 40188 2547
rect 28620 2431 28639 2477
rect 28685 2431 28755 2477
rect 28801 2431 28871 2477
rect 28917 2431 28987 2477
rect 29033 2431 29103 2477
rect 29149 2431 29219 2477
rect 29265 2431 29335 2477
rect 29381 2431 29451 2477
rect 29497 2431 29567 2477
rect 29613 2431 29683 2477
rect 29729 2431 29799 2477
rect 29845 2431 29915 2477
rect 29961 2431 30031 2477
rect 30077 2431 30147 2477
rect 30193 2431 30263 2477
rect 30309 2431 30379 2477
rect 30425 2431 30495 2477
rect 30541 2431 30611 2477
rect 30657 2431 30727 2477
rect 30773 2431 30843 2477
rect 30889 2431 30959 2477
rect 31005 2431 31075 2477
rect 31121 2431 31191 2477
rect 31237 2431 31307 2477
rect 31353 2431 31423 2477
rect 31469 2431 31539 2477
rect 31585 2431 31655 2477
rect 31701 2431 31771 2477
rect 31817 2431 31887 2477
rect 31933 2431 32003 2477
rect 32049 2431 32119 2477
rect 32165 2431 32235 2477
rect 32281 2431 32351 2477
rect 32397 2431 32467 2477
rect 32513 2431 32583 2477
rect 32629 2431 32699 2477
rect 32745 2431 32815 2477
rect 32861 2431 32931 2477
rect 32977 2431 33047 2477
rect 33093 2431 33163 2477
rect 33209 2431 33279 2477
rect 33325 2431 33395 2477
rect 33441 2431 33511 2477
rect 33557 2431 33627 2477
rect 33673 2431 33743 2477
rect 33789 2431 33859 2477
rect 33905 2431 33975 2477
rect 34021 2431 34091 2477
rect 34137 2431 34207 2477
rect 34253 2431 34323 2477
rect 34369 2431 34439 2477
rect 34485 2431 34555 2477
rect 34601 2431 34671 2477
rect 34717 2431 34787 2477
rect 34833 2431 34903 2477
rect 34949 2431 35019 2477
rect 35065 2431 35135 2477
rect 35181 2431 35251 2477
rect 35297 2431 35367 2477
rect 35413 2431 35483 2477
rect 35529 2431 35599 2477
rect 35645 2431 35715 2477
rect 35761 2431 35831 2477
rect 35877 2431 35947 2477
rect 35993 2431 36063 2477
rect 36109 2431 36179 2477
rect 36225 2431 36295 2477
rect 36341 2431 36411 2477
rect 36457 2431 36527 2477
rect 36573 2431 36643 2477
rect 36689 2431 36759 2477
rect 36805 2431 36875 2477
rect 36921 2431 36991 2477
rect 37037 2431 37107 2477
rect 37153 2431 37223 2477
rect 37269 2431 37339 2477
rect 37385 2431 37455 2477
rect 37501 2431 37571 2477
rect 37617 2431 37687 2477
rect 37733 2431 37803 2477
rect 37849 2431 37919 2477
rect 37965 2431 38035 2477
rect 38081 2431 38151 2477
rect 38197 2431 38267 2477
rect 38313 2431 38383 2477
rect 38429 2431 38499 2477
rect 38545 2431 38615 2477
rect 38661 2431 38731 2477
rect 38777 2431 38847 2477
rect 38893 2431 38963 2477
rect 39009 2431 39079 2477
rect 39125 2431 39195 2477
rect 39241 2431 39311 2477
rect 39357 2431 39427 2477
rect 39473 2431 39543 2477
rect 39589 2431 39659 2477
rect 39705 2431 39775 2477
rect 39821 2431 39891 2477
rect 39937 2431 40007 2477
rect 40053 2431 40123 2477
rect 40169 2431 40188 2477
rect 28620 2361 40188 2431
rect 28620 2315 28639 2361
rect 28685 2315 28755 2361
rect 28801 2315 28871 2361
rect 28917 2315 28987 2361
rect 29033 2315 29103 2361
rect 29149 2315 29219 2361
rect 29265 2315 29335 2361
rect 29381 2315 29451 2361
rect 29497 2315 29567 2361
rect 29613 2315 29683 2361
rect 29729 2315 29799 2361
rect 29845 2315 29915 2361
rect 29961 2315 30031 2361
rect 30077 2315 30147 2361
rect 30193 2315 30263 2361
rect 30309 2315 30379 2361
rect 30425 2315 30495 2361
rect 30541 2315 30611 2361
rect 30657 2315 30727 2361
rect 30773 2315 30843 2361
rect 30889 2315 30959 2361
rect 31005 2315 31075 2361
rect 31121 2315 31191 2361
rect 31237 2315 31307 2361
rect 31353 2315 31423 2361
rect 31469 2315 31539 2361
rect 31585 2315 31655 2361
rect 31701 2315 31771 2361
rect 31817 2315 31887 2361
rect 31933 2315 32003 2361
rect 32049 2315 32119 2361
rect 32165 2315 32235 2361
rect 32281 2315 32351 2361
rect 32397 2315 32467 2361
rect 32513 2315 32583 2361
rect 32629 2315 32699 2361
rect 32745 2315 32815 2361
rect 32861 2315 32931 2361
rect 32977 2315 33047 2361
rect 33093 2315 33163 2361
rect 33209 2315 33279 2361
rect 33325 2315 33395 2361
rect 33441 2315 33511 2361
rect 33557 2315 33627 2361
rect 33673 2315 33743 2361
rect 33789 2315 33859 2361
rect 33905 2315 33975 2361
rect 34021 2315 34091 2361
rect 34137 2315 34207 2361
rect 34253 2315 34323 2361
rect 34369 2315 34439 2361
rect 34485 2315 34555 2361
rect 34601 2315 34671 2361
rect 34717 2315 34787 2361
rect 34833 2315 34903 2361
rect 34949 2315 35019 2361
rect 35065 2315 35135 2361
rect 35181 2315 35251 2361
rect 35297 2315 35367 2361
rect 35413 2315 35483 2361
rect 35529 2315 35599 2361
rect 35645 2315 35715 2361
rect 35761 2315 35831 2361
rect 35877 2315 35947 2361
rect 35993 2315 36063 2361
rect 36109 2315 36179 2361
rect 36225 2315 36295 2361
rect 36341 2315 36411 2361
rect 36457 2315 36527 2361
rect 36573 2315 36643 2361
rect 36689 2315 36759 2361
rect 36805 2315 36875 2361
rect 36921 2315 36991 2361
rect 37037 2315 37107 2361
rect 37153 2315 37223 2361
rect 37269 2315 37339 2361
rect 37385 2315 37455 2361
rect 37501 2315 37571 2361
rect 37617 2315 37687 2361
rect 37733 2315 37803 2361
rect 37849 2315 37919 2361
rect 37965 2315 38035 2361
rect 38081 2315 38151 2361
rect 38197 2315 38267 2361
rect 38313 2315 38383 2361
rect 38429 2315 38499 2361
rect 38545 2315 38615 2361
rect 38661 2315 38731 2361
rect 38777 2315 38847 2361
rect 38893 2315 38963 2361
rect 39009 2315 39079 2361
rect 39125 2315 39195 2361
rect 39241 2315 39311 2361
rect 39357 2315 39427 2361
rect 39473 2315 39543 2361
rect 39589 2315 39659 2361
rect 39705 2315 39775 2361
rect 39821 2315 39891 2361
rect 39937 2315 40007 2361
rect 40053 2315 40123 2361
rect 40169 2315 40188 2361
rect 28620 2245 40188 2315
rect 28620 2199 28639 2245
rect 28685 2199 28755 2245
rect 28801 2199 28871 2245
rect 28917 2199 28987 2245
rect 29033 2199 29103 2245
rect 29149 2199 29219 2245
rect 29265 2199 29335 2245
rect 29381 2199 29451 2245
rect 29497 2199 29567 2245
rect 29613 2199 29683 2245
rect 29729 2199 29799 2245
rect 29845 2199 29915 2245
rect 29961 2199 30031 2245
rect 30077 2199 30147 2245
rect 30193 2199 30263 2245
rect 30309 2199 30379 2245
rect 30425 2199 30495 2245
rect 30541 2199 30611 2245
rect 30657 2199 30727 2245
rect 30773 2199 30843 2245
rect 30889 2199 30959 2245
rect 31005 2199 31075 2245
rect 31121 2199 31191 2245
rect 31237 2199 31307 2245
rect 31353 2199 31423 2245
rect 31469 2199 31539 2245
rect 31585 2199 31655 2245
rect 31701 2199 31771 2245
rect 31817 2199 31887 2245
rect 31933 2199 32003 2245
rect 32049 2199 32119 2245
rect 32165 2199 32235 2245
rect 32281 2199 32351 2245
rect 32397 2199 32467 2245
rect 32513 2199 32583 2245
rect 32629 2199 32699 2245
rect 32745 2199 32815 2245
rect 32861 2199 32931 2245
rect 32977 2199 33047 2245
rect 33093 2199 33163 2245
rect 33209 2199 33279 2245
rect 33325 2199 33395 2245
rect 33441 2199 33511 2245
rect 33557 2199 33627 2245
rect 33673 2199 33743 2245
rect 33789 2199 33859 2245
rect 33905 2199 33975 2245
rect 34021 2199 34091 2245
rect 34137 2199 34207 2245
rect 34253 2199 34323 2245
rect 34369 2199 34439 2245
rect 34485 2199 34555 2245
rect 34601 2199 34671 2245
rect 34717 2199 34787 2245
rect 34833 2199 34903 2245
rect 34949 2199 35019 2245
rect 35065 2199 35135 2245
rect 35181 2199 35251 2245
rect 35297 2199 35367 2245
rect 35413 2199 35483 2245
rect 35529 2199 35599 2245
rect 35645 2199 35715 2245
rect 35761 2199 35831 2245
rect 35877 2199 35947 2245
rect 35993 2199 36063 2245
rect 36109 2199 36179 2245
rect 36225 2199 36295 2245
rect 36341 2199 36411 2245
rect 36457 2199 36527 2245
rect 36573 2199 36643 2245
rect 36689 2199 36759 2245
rect 36805 2199 36875 2245
rect 36921 2199 36991 2245
rect 37037 2199 37107 2245
rect 37153 2199 37223 2245
rect 37269 2199 37339 2245
rect 37385 2199 37455 2245
rect 37501 2199 37571 2245
rect 37617 2199 37687 2245
rect 37733 2199 37803 2245
rect 37849 2199 37919 2245
rect 37965 2199 38035 2245
rect 38081 2199 38151 2245
rect 38197 2199 38267 2245
rect 38313 2199 38383 2245
rect 38429 2199 38499 2245
rect 38545 2199 38615 2245
rect 38661 2199 38731 2245
rect 38777 2199 38847 2245
rect 38893 2199 38963 2245
rect 39009 2199 39079 2245
rect 39125 2199 39195 2245
rect 39241 2199 39311 2245
rect 39357 2199 39427 2245
rect 39473 2199 39543 2245
rect 39589 2199 39659 2245
rect 39705 2199 39775 2245
rect 39821 2199 39891 2245
rect 39937 2199 40007 2245
rect 40053 2199 40123 2245
rect 40169 2199 40188 2245
rect 28620 2129 40188 2199
rect 28620 2083 28639 2129
rect 28685 2083 28755 2129
rect 28801 2083 28871 2129
rect 28917 2083 28987 2129
rect 29033 2083 29103 2129
rect 29149 2083 29219 2129
rect 29265 2083 29335 2129
rect 29381 2083 29451 2129
rect 29497 2083 29567 2129
rect 29613 2083 29683 2129
rect 29729 2083 29799 2129
rect 29845 2083 29915 2129
rect 29961 2083 30031 2129
rect 30077 2083 30147 2129
rect 30193 2083 30263 2129
rect 30309 2083 30379 2129
rect 30425 2083 30495 2129
rect 30541 2083 30611 2129
rect 30657 2083 30727 2129
rect 30773 2083 30843 2129
rect 30889 2083 30959 2129
rect 31005 2083 31075 2129
rect 31121 2083 31191 2129
rect 31237 2083 31307 2129
rect 31353 2083 31423 2129
rect 31469 2083 31539 2129
rect 31585 2083 31655 2129
rect 31701 2083 31771 2129
rect 31817 2083 31887 2129
rect 31933 2083 32003 2129
rect 32049 2083 32119 2129
rect 32165 2083 32235 2129
rect 32281 2083 32351 2129
rect 32397 2083 32467 2129
rect 32513 2083 32583 2129
rect 32629 2083 32699 2129
rect 32745 2083 32815 2129
rect 32861 2083 32931 2129
rect 32977 2083 33047 2129
rect 33093 2083 33163 2129
rect 33209 2083 33279 2129
rect 33325 2083 33395 2129
rect 33441 2083 33511 2129
rect 33557 2083 33627 2129
rect 33673 2083 33743 2129
rect 33789 2083 33859 2129
rect 33905 2083 33975 2129
rect 34021 2083 34091 2129
rect 34137 2083 34207 2129
rect 34253 2083 34323 2129
rect 34369 2083 34439 2129
rect 34485 2083 34555 2129
rect 34601 2083 34671 2129
rect 34717 2083 34787 2129
rect 34833 2083 34903 2129
rect 34949 2083 35019 2129
rect 35065 2083 35135 2129
rect 35181 2083 35251 2129
rect 35297 2083 35367 2129
rect 35413 2083 35483 2129
rect 35529 2083 35599 2129
rect 35645 2083 35715 2129
rect 35761 2083 35831 2129
rect 35877 2083 35947 2129
rect 35993 2083 36063 2129
rect 36109 2083 36179 2129
rect 36225 2083 36295 2129
rect 36341 2083 36411 2129
rect 36457 2083 36527 2129
rect 36573 2083 36643 2129
rect 36689 2083 36759 2129
rect 36805 2083 36875 2129
rect 36921 2083 36991 2129
rect 37037 2083 37107 2129
rect 37153 2083 37223 2129
rect 37269 2083 37339 2129
rect 37385 2083 37455 2129
rect 37501 2083 37571 2129
rect 37617 2083 37687 2129
rect 37733 2083 37803 2129
rect 37849 2083 37919 2129
rect 37965 2083 38035 2129
rect 38081 2083 38151 2129
rect 38197 2083 38267 2129
rect 38313 2083 38383 2129
rect 38429 2083 38499 2129
rect 38545 2083 38615 2129
rect 38661 2083 38731 2129
rect 38777 2083 38847 2129
rect 38893 2083 38963 2129
rect 39009 2083 39079 2129
rect 39125 2083 39195 2129
rect 39241 2083 39311 2129
rect 39357 2083 39427 2129
rect 39473 2083 39543 2129
rect 39589 2083 39659 2129
rect 39705 2083 39775 2129
rect 39821 2083 39891 2129
rect 39937 2083 40007 2129
rect 40053 2083 40123 2129
rect 40169 2083 40188 2129
rect 28620 2013 40188 2083
rect 28620 1967 28639 2013
rect 28685 1967 28755 2013
rect 28801 1967 28871 2013
rect 28917 1967 28987 2013
rect 29033 1967 29103 2013
rect 29149 1967 29219 2013
rect 29265 1967 29335 2013
rect 29381 1967 29451 2013
rect 29497 1967 29567 2013
rect 29613 1967 29683 2013
rect 29729 1967 29799 2013
rect 29845 1967 29915 2013
rect 29961 1967 30031 2013
rect 30077 1967 30147 2013
rect 30193 1967 30263 2013
rect 30309 1967 30379 2013
rect 30425 1967 30495 2013
rect 30541 1967 30611 2013
rect 30657 1967 30727 2013
rect 30773 1967 30843 2013
rect 30889 1967 30959 2013
rect 31005 1967 31075 2013
rect 31121 1967 31191 2013
rect 31237 1967 31307 2013
rect 31353 1967 31423 2013
rect 31469 1967 31539 2013
rect 31585 1967 31655 2013
rect 31701 1967 31771 2013
rect 31817 1967 31887 2013
rect 31933 1967 32003 2013
rect 32049 1967 32119 2013
rect 32165 1967 32235 2013
rect 32281 1967 32351 2013
rect 32397 1967 32467 2013
rect 32513 1967 32583 2013
rect 32629 1967 32699 2013
rect 32745 1967 32815 2013
rect 32861 1967 32931 2013
rect 32977 1967 33047 2013
rect 33093 1967 33163 2013
rect 33209 1967 33279 2013
rect 33325 1967 33395 2013
rect 33441 1967 33511 2013
rect 33557 1967 33627 2013
rect 33673 1967 33743 2013
rect 33789 1967 33859 2013
rect 33905 1967 33975 2013
rect 34021 1967 34091 2013
rect 34137 1967 34207 2013
rect 34253 1967 34323 2013
rect 34369 1967 34439 2013
rect 34485 1967 34555 2013
rect 34601 1967 34671 2013
rect 34717 1967 34787 2013
rect 34833 1967 34903 2013
rect 34949 1967 35019 2013
rect 35065 1967 35135 2013
rect 35181 1967 35251 2013
rect 35297 1967 35367 2013
rect 35413 1967 35483 2013
rect 35529 1967 35599 2013
rect 35645 1967 35715 2013
rect 35761 1967 35831 2013
rect 35877 1967 35947 2013
rect 35993 1967 36063 2013
rect 36109 1967 36179 2013
rect 36225 1967 36295 2013
rect 36341 1967 36411 2013
rect 36457 1967 36527 2013
rect 36573 1967 36643 2013
rect 36689 1967 36759 2013
rect 36805 1967 36875 2013
rect 36921 1967 36991 2013
rect 37037 1967 37107 2013
rect 37153 1967 37223 2013
rect 37269 1967 37339 2013
rect 37385 1967 37455 2013
rect 37501 1967 37571 2013
rect 37617 1967 37687 2013
rect 37733 1967 37803 2013
rect 37849 1967 37919 2013
rect 37965 1967 38035 2013
rect 38081 1967 38151 2013
rect 38197 1967 38267 2013
rect 38313 1967 38383 2013
rect 38429 1967 38499 2013
rect 38545 1967 38615 2013
rect 38661 1967 38731 2013
rect 38777 1967 38847 2013
rect 38893 1967 38963 2013
rect 39009 1967 39079 2013
rect 39125 1967 39195 2013
rect 39241 1967 39311 2013
rect 39357 1967 39427 2013
rect 39473 1967 39543 2013
rect 39589 1967 39659 2013
rect 39705 1967 39775 2013
rect 39821 1967 39891 2013
rect 39937 1967 40007 2013
rect 40053 1967 40123 2013
rect 40169 1967 40188 2013
rect 28620 1897 40188 1967
rect 28620 1851 28639 1897
rect 28685 1851 28755 1897
rect 28801 1851 28871 1897
rect 28917 1851 28987 1897
rect 29033 1851 29103 1897
rect 29149 1851 29219 1897
rect 29265 1851 29335 1897
rect 29381 1851 29451 1897
rect 29497 1851 29567 1897
rect 29613 1851 29683 1897
rect 29729 1851 29799 1897
rect 29845 1851 29915 1897
rect 29961 1851 30031 1897
rect 30077 1851 30147 1897
rect 30193 1851 30263 1897
rect 30309 1851 30379 1897
rect 30425 1851 30495 1897
rect 30541 1851 30611 1897
rect 30657 1851 30727 1897
rect 30773 1851 30843 1897
rect 30889 1851 30959 1897
rect 31005 1851 31075 1897
rect 31121 1851 31191 1897
rect 31237 1851 31307 1897
rect 31353 1851 31423 1897
rect 31469 1851 31539 1897
rect 31585 1851 31655 1897
rect 31701 1851 31771 1897
rect 31817 1851 31887 1897
rect 31933 1851 32003 1897
rect 32049 1851 32119 1897
rect 32165 1851 32235 1897
rect 32281 1851 32351 1897
rect 32397 1851 32467 1897
rect 32513 1851 32583 1897
rect 32629 1851 32699 1897
rect 32745 1851 32815 1897
rect 32861 1851 32931 1897
rect 32977 1851 33047 1897
rect 33093 1851 33163 1897
rect 33209 1851 33279 1897
rect 33325 1851 33395 1897
rect 33441 1851 33511 1897
rect 33557 1851 33627 1897
rect 33673 1851 33743 1897
rect 33789 1851 33859 1897
rect 33905 1851 33975 1897
rect 34021 1851 34091 1897
rect 34137 1851 34207 1897
rect 34253 1851 34323 1897
rect 34369 1851 34439 1897
rect 34485 1851 34555 1897
rect 34601 1851 34671 1897
rect 34717 1851 34787 1897
rect 34833 1851 34903 1897
rect 34949 1851 35019 1897
rect 35065 1851 35135 1897
rect 35181 1851 35251 1897
rect 35297 1851 35367 1897
rect 35413 1851 35483 1897
rect 35529 1851 35599 1897
rect 35645 1851 35715 1897
rect 35761 1851 35831 1897
rect 35877 1851 35947 1897
rect 35993 1851 36063 1897
rect 36109 1851 36179 1897
rect 36225 1851 36295 1897
rect 36341 1851 36411 1897
rect 36457 1851 36527 1897
rect 36573 1851 36643 1897
rect 36689 1851 36759 1897
rect 36805 1851 36875 1897
rect 36921 1851 36991 1897
rect 37037 1851 37107 1897
rect 37153 1851 37223 1897
rect 37269 1851 37339 1897
rect 37385 1851 37455 1897
rect 37501 1851 37571 1897
rect 37617 1851 37687 1897
rect 37733 1851 37803 1897
rect 37849 1851 37919 1897
rect 37965 1851 38035 1897
rect 38081 1851 38151 1897
rect 38197 1851 38267 1897
rect 38313 1851 38383 1897
rect 38429 1851 38499 1897
rect 38545 1851 38615 1897
rect 38661 1851 38731 1897
rect 38777 1851 38847 1897
rect 38893 1851 38963 1897
rect 39009 1851 39079 1897
rect 39125 1851 39195 1897
rect 39241 1851 39311 1897
rect 39357 1851 39427 1897
rect 39473 1851 39543 1897
rect 39589 1851 39659 1897
rect 39705 1851 39775 1897
rect 39821 1851 39891 1897
rect 39937 1851 40007 1897
rect 40053 1851 40123 1897
rect 40169 1851 40188 1897
rect 28620 1781 40188 1851
rect 28620 1735 28639 1781
rect 28685 1735 28755 1781
rect 28801 1735 28871 1781
rect 28917 1735 28987 1781
rect 29033 1735 29103 1781
rect 29149 1735 29219 1781
rect 29265 1735 29335 1781
rect 29381 1735 29451 1781
rect 29497 1735 29567 1781
rect 29613 1735 29683 1781
rect 29729 1735 29799 1781
rect 29845 1735 29915 1781
rect 29961 1735 30031 1781
rect 30077 1735 30147 1781
rect 30193 1735 30263 1781
rect 30309 1735 30379 1781
rect 30425 1735 30495 1781
rect 30541 1735 30611 1781
rect 30657 1735 30727 1781
rect 30773 1735 30843 1781
rect 30889 1735 30959 1781
rect 31005 1735 31075 1781
rect 31121 1735 31191 1781
rect 31237 1735 31307 1781
rect 31353 1735 31423 1781
rect 31469 1735 31539 1781
rect 31585 1735 31655 1781
rect 31701 1735 31771 1781
rect 31817 1735 31887 1781
rect 31933 1735 32003 1781
rect 32049 1735 32119 1781
rect 32165 1735 32235 1781
rect 32281 1735 32351 1781
rect 32397 1735 32467 1781
rect 32513 1735 32583 1781
rect 32629 1735 32699 1781
rect 32745 1735 32815 1781
rect 32861 1735 32931 1781
rect 32977 1735 33047 1781
rect 33093 1735 33163 1781
rect 33209 1735 33279 1781
rect 33325 1735 33395 1781
rect 33441 1735 33511 1781
rect 33557 1735 33627 1781
rect 33673 1735 33743 1781
rect 33789 1735 33859 1781
rect 33905 1735 33975 1781
rect 34021 1735 34091 1781
rect 34137 1735 34207 1781
rect 34253 1735 34323 1781
rect 34369 1735 34439 1781
rect 34485 1735 34555 1781
rect 34601 1735 34671 1781
rect 34717 1735 34787 1781
rect 34833 1735 34903 1781
rect 34949 1735 35019 1781
rect 35065 1735 35135 1781
rect 35181 1735 35251 1781
rect 35297 1735 35367 1781
rect 35413 1735 35483 1781
rect 35529 1735 35599 1781
rect 35645 1735 35715 1781
rect 35761 1735 35831 1781
rect 35877 1735 35947 1781
rect 35993 1735 36063 1781
rect 36109 1735 36179 1781
rect 36225 1735 36295 1781
rect 36341 1735 36411 1781
rect 36457 1735 36527 1781
rect 36573 1735 36643 1781
rect 36689 1735 36759 1781
rect 36805 1735 36875 1781
rect 36921 1735 36991 1781
rect 37037 1735 37107 1781
rect 37153 1735 37223 1781
rect 37269 1735 37339 1781
rect 37385 1735 37455 1781
rect 37501 1735 37571 1781
rect 37617 1735 37687 1781
rect 37733 1735 37803 1781
rect 37849 1735 37919 1781
rect 37965 1735 38035 1781
rect 38081 1735 38151 1781
rect 38197 1735 38267 1781
rect 38313 1735 38383 1781
rect 38429 1735 38499 1781
rect 38545 1735 38615 1781
rect 38661 1735 38731 1781
rect 38777 1735 38847 1781
rect 38893 1735 38963 1781
rect 39009 1735 39079 1781
rect 39125 1735 39195 1781
rect 39241 1735 39311 1781
rect 39357 1735 39427 1781
rect 39473 1735 39543 1781
rect 39589 1735 39659 1781
rect 39705 1735 39775 1781
rect 39821 1735 39891 1781
rect 39937 1735 40007 1781
rect 40053 1735 40123 1781
rect 40169 1735 40188 1781
rect 28620 1665 40188 1735
rect 28620 1619 28639 1665
rect 28685 1619 28755 1665
rect 28801 1619 28871 1665
rect 28917 1619 28987 1665
rect 29033 1619 29103 1665
rect 29149 1619 29219 1665
rect 29265 1619 29335 1665
rect 29381 1619 29451 1665
rect 29497 1619 29567 1665
rect 29613 1619 29683 1665
rect 29729 1619 29799 1665
rect 29845 1619 29915 1665
rect 29961 1619 30031 1665
rect 30077 1619 30147 1665
rect 30193 1619 30263 1665
rect 30309 1619 30379 1665
rect 30425 1619 30495 1665
rect 30541 1619 30611 1665
rect 30657 1619 30727 1665
rect 30773 1619 30843 1665
rect 30889 1619 30959 1665
rect 31005 1619 31075 1665
rect 31121 1619 31191 1665
rect 31237 1619 31307 1665
rect 31353 1619 31423 1665
rect 31469 1619 31539 1665
rect 31585 1619 31655 1665
rect 31701 1619 31771 1665
rect 31817 1619 31887 1665
rect 31933 1619 32003 1665
rect 32049 1619 32119 1665
rect 32165 1619 32235 1665
rect 32281 1619 32351 1665
rect 32397 1619 32467 1665
rect 32513 1619 32583 1665
rect 32629 1619 32699 1665
rect 32745 1619 32815 1665
rect 32861 1619 32931 1665
rect 32977 1619 33047 1665
rect 33093 1619 33163 1665
rect 33209 1619 33279 1665
rect 33325 1619 33395 1665
rect 33441 1619 33511 1665
rect 33557 1619 33627 1665
rect 33673 1619 33743 1665
rect 33789 1619 33859 1665
rect 33905 1619 33975 1665
rect 34021 1619 34091 1665
rect 34137 1619 34207 1665
rect 34253 1619 34323 1665
rect 34369 1619 34439 1665
rect 34485 1619 34555 1665
rect 34601 1619 34671 1665
rect 34717 1619 34787 1665
rect 34833 1619 34903 1665
rect 34949 1619 35019 1665
rect 35065 1619 35135 1665
rect 35181 1619 35251 1665
rect 35297 1619 35367 1665
rect 35413 1619 35483 1665
rect 35529 1619 35599 1665
rect 35645 1619 35715 1665
rect 35761 1619 35831 1665
rect 35877 1619 35947 1665
rect 35993 1619 36063 1665
rect 36109 1619 36179 1665
rect 36225 1619 36295 1665
rect 36341 1619 36411 1665
rect 36457 1619 36527 1665
rect 36573 1619 36643 1665
rect 36689 1619 36759 1665
rect 36805 1619 36875 1665
rect 36921 1619 36991 1665
rect 37037 1619 37107 1665
rect 37153 1619 37223 1665
rect 37269 1619 37339 1665
rect 37385 1619 37455 1665
rect 37501 1619 37571 1665
rect 37617 1619 37687 1665
rect 37733 1619 37803 1665
rect 37849 1619 37919 1665
rect 37965 1619 38035 1665
rect 38081 1619 38151 1665
rect 38197 1619 38267 1665
rect 38313 1619 38383 1665
rect 38429 1619 38499 1665
rect 38545 1619 38615 1665
rect 38661 1619 38731 1665
rect 38777 1619 38847 1665
rect 38893 1619 38963 1665
rect 39009 1619 39079 1665
rect 39125 1619 39195 1665
rect 39241 1619 39311 1665
rect 39357 1619 39427 1665
rect 39473 1619 39543 1665
rect 39589 1619 39659 1665
rect 39705 1619 39775 1665
rect 39821 1619 39891 1665
rect 39937 1619 40007 1665
rect 40053 1619 40123 1665
rect 40169 1619 40188 1665
rect 28620 1549 40188 1619
rect 28620 1503 28639 1549
rect 28685 1503 28755 1549
rect 28801 1503 28871 1549
rect 28917 1503 28987 1549
rect 29033 1503 29103 1549
rect 29149 1503 29219 1549
rect 29265 1503 29335 1549
rect 29381 1503 29451 1549
rect 29497 1503 29567 1549
rect 29613 1503 29683 1549
rect 29729 1503 29799 1549
rect 29845 1503 29915 1549
rect 29961 1503 30031 1549
rect 30077 1503 30147 1549
rect 30193 1503 30263 1549
rect 30309 1503 30379 1549
rect 30425 1503 30495 1549
rect 30541 1503 30611 1549
rect 30657 1503 30727 1549
rect 30773 1503 30843 1549
rect 30889 1503 30959 1549
rect 31005 1503 31075 1549
rect 31121 1503 31191 1549
rect 31237 1503 31307 1549
rect 31353 1503 31423 1549
rect 31469 1503 31539 1549
rect 31585 1503 31655 1549
rect 31701 1503 31771 1549
rect 31817 1503 31887 1549
rect 31933 1503 32003 1549
rect 32049 1503 32119 1549
rect 32165 1503 32235 1549
rect 32281 1503 32351 1549
rect 32397 1503 32467 1549
rect 32513 1503 32583 1549
rect 32629 1503 32699 1549
rect 32745 1503 32815 1549
rect 32861 1503 32931 1549
rect 32977 1503 33047 1549
rect 33093 1503 33163 1549
rect 33209 1503 33279 1549
rect 33325 1503 33395 1549
rect 33441 1503 33511 1549
rect 33557 1503 33627 1549
rect 33673 1503 33743 1549
rect 33789 1503 33859 1549
rect 33905 1503 33975 1549
rect 34021 1503 34091 1549
rect 34137 1503 34207 1549
rect 34253 1503 34323 1549
rect 34369 1503 34439 1549
rect 34485 1503 34555 1549
rect 34601 1503 34671 1549
rect 34717 1503 34787 1549
rect 34833 1503 34903 1549
rect 34949 1503 35019 1549
rect 35065 1503 35135 1549
rect 35181 1503 35251 1549
rect 35297 1503 35367 1549
rect 35413 1503 35483 1549
rect 35529 1503 35599 1549
rect 35645 1503 35715 1549
rect 35761 1503 35831 1549
rect 35877 1503 35947 1549
rect 35993 1503 36063 1549
rect 36109 1503 36179 1549
rect 36225 1503 36295 1549
rect 36341 1503 36411 1549
rect 36457 1503 36527 1549
rect 36573 1503 36643 1549
rect 36689 1503 36759 1549
rect 36805 1503 36875 1549
rect 36921 1503 36991 1549
rect 37037 1503 37107 1549
rect 37153 1503 37223 1549
rect 37269 1503 37339 1549
rect 37385 1503 37455 1549
rect 37501 1503 37571 1549
rect 37617 1503 37687 1549
rect 37733 1503 37803 1549
rect 37849 1503 37919 1549
rect 37965 1503 38035 1549
rect 38081 1503 38151 1549
rect 38197 1503 38267 1549
rect 38313 1503 38383 1549
rect 38429 1503 38499 1549
rect 38545 1503 38615 1549
rect 38661 1503 38731 1549
rect 38777 1503 38847 1549
rect 38893 1503 38963 1549
rect 39009 1503 39079 1549
rect 39125 1503 39195 1549
rect 39241 1503 39311 1549
rect 39357 1503 39427 1549
rect 39473 1503 39543 1549
rect 39589 1503 39659 1549
rect 39705 1503 39775 1549
rect 39821 1503 39891 1549
rect 39937 1503 40007 1549
rect 40053 1503 40123 1549
rect 40169 1503 40188 1549
rect 28620 1433 40188 1503
rect 28620 1387 28639 1433
rect 28685 1387 28755 1433
rect 28801 1387 28871 1433
rect 28917 1387 28987 1433
rect 29033 1387 29103 1433
rect 29149 1387 29219 1433
rect 29265 1387 29335 1433
rect 29381 1387 29451 1433
rect 29497 1387 29567 1433
rect 29613 1387 29683 1433
rect 29729 1387 29799 1433
rect 29845 1387 29915 1433
rect 29961 1387 30031 1433
rect 30077 1387 30147 1433
rect 30193 1387 30263 1433
rect 30309 1387 30379 1433
rect 30425 1387 30495 1433
rect 30541 1387 30611 1433
rect 30657 1387 30727 1433
rect 30773 1387 30843 1433
rect 30889 1387 30959 1433
rect 31005 1387 31075 1433
rect 31121 1387 31191 1433
rect 31237 1387 31307 1433
rect 31353 1387 31423 1433
rect 31469 1387 31539 1433
rect 31585 1387 31655 1433
rect 31701 1387 31771 1433
rect 31817 1387 31887 1433
rect 31933 1387 32003 1433
rect 32049 1387 32119 1433
rect 32165 1387 32235 1433
rect 32281 1387 32351 1433
rect 32397 1387 32467 1433
rect 32513 1387 32583 1433
rect 32629 1387 32699 1433
rect 32745 1387 32815 1433
rect 32861 1387 32931 1433
rect 32977 1387 33047 1433
rect 33093 1387 33163 1433
rect 33209 1387 33279 1433
rect 33325 1387 33395 1433
rect 33441 1387 33511 1433
rect 33557 1387 33627 1433
rect 33673 1387 33743 1433
rect 33789 1387 33859 1433
rect 33905 1387 33975 1433
rect 34021 1387 34091 1433
rect 34137 1387 34207 1433
rect 34253 1387 34323 1433
rect 34369 1387 34439 1433
rect 34485 1387 34555 1433
rect 34601 1387 34671 1433
rect 34717 1387 34787 1433
rect 34833 1387 34903 1433
rect 34949 1387 35019 1433
rect 35065 1387 35135 1433
rect 35181 1387 35251 1433
rect 35297 1387 35367 1433
rect 35413 1387 35483 1433
rect 35529 1387 35599 1433
rect 35645 1387 35715 1433
rect 35761 1387 35831 1433
rect 35877 1387 35947 1433
rect 35993 1387 36063 1433
rect 36109 1387 36179 1433
rect 36225 1387 36295 1433
rect 36341 1387 36411 1433
rect 36457 1387 36527 1433
rect 36573 1387 36643 1433
rect 36689 1387 36759 1433
rect 36805 1387 36875 1433
rect 36921 1387 36991 1433
rect 37037 1387 37107 1433
rect 37153 1387 37223 1433
rect 37269 1387 37339 1433
rect 37385 1387 37455 1433
rect 37501 1387 37571 1433
rect 37617 1387 37687 1433
rect 37733 1387 37803 1433
rect 37849 1387 37919 1433
rect 37965 1387 38035 1433
rect 38081 1387 38151 1433
rect 38197 1387 38267 1433
rect 38313 1387 38383 1433
rect 38429 1387 38499 1433
rect 38545 1387 38615 1433
rect 38661 1387 38731 1433
rect 38777 1387 38847 1433
rect 38893 1387 38963 1433
rect 39009 1387 39079 1433
rect 39125 1387 39195 1433
rect 39241 1387 39311 1433
rect 39357 1387 39427 1433
rect 39473 1387 39543 1433
rect 39589 1387 39659 1433
rect 39705 1387 39775 1433
rect 39821 1387 39891 1433
rect 39937 1387 40007 1433
rect 40053 1387 40123 1433
rect 40169 1387 40188 1433
rect 28620 1317 40188 1387
rect 28620 1271 28639 1317
rect 28685 1271 28755 1317
rect 28801 1271 28871 1317
rect 28917 1271 28987 1317
rect 29033 1271 29103 1317
rect 29149 1271 29219 1317
rect 29265 1271 29335 1317
rect 29381 1271 29451 1317
rect 29497 1271 29567 1317
rect 29613 1271 29683 1317
rect 29729 1271 29799 1317
rect 29845 1271 29915 1317
rect 29961 1271 30031 1317
rect 30077 1271 30147 1317
rect 30193 1271 30263 1317
rect 30309 1271 30379 1317
rect 30425 1271 30495 1317
rect 30541 1271 30611 1317
rect 30657 1271 30727 1317
rect 30773 1271 30843 1317
rect 30889 1271 30959 1317
rect 31005 1271 31075 1317
rect 31121 1271 31191 1317
rect 31237 1271 31307 1317
rect 31353 1271 31423 1317
rect 31469 1271 31539 1317
rect 31585 1271 31655 1317
rect 31701 1271 31771 1317
rect 31817 1271 31887 1317
rect 31933 1271 32003 1317
rect 32049 1271 32119 1317
rect 32165 1271 32235 1317
rect 32281 1271 32351 1317
rect 32397 1271 32467 1317
rect 32513 1271 32583 1317
rect 32629 1271 32699 1317
rect 32745 1271 32815 1317
rect 32861 1271 32931 1317
rect 32977 1271 33047 1317
rect 33093 1271 33163 1317
rect 33209 1271 33279 1317
rect 33325 1271 33395 1317
rect 33441 1271 33511 1317
rect 33557 1271 33627 1317
rect 33673 1271 33743 1317
rect 33789 1271 33859 1317
rect 33905 1271 33975 1317
rect 34021 1271 34091 1317
rect 34137 1271 34207 1317
rect 34253 1271 34323 1317
rect 34369 1271 34439 1317
rect 34485 1271 34555 1317
rect 34601 1271 34671 1317
rect 34717 1271 34787 1317
rect 34833 1271 34903 1317
rect 34949 1271 35019 1317
rect 35065 1271 35135 1317
rect 35181 1271 35251 1317
rect 35297 1271 35367 1317
rect 35413 1271 35483 1317
rect 35529 1271 35599 1317
rect 35645 1271 35715 1317
rect 35761 1271 35831 1317
rect 35877 1271 35947 1317
rect 35993 1271 36063 1317
rect 36109 1271 36179 1317
rect 36225 1271 36295 1317
rect 36341 1271 36411 1317
rect 36457 1271 36527 1317
rect 36573 1271 36643 1317
rect 36689 1271 36759 1317
rect 36805 1271 36875 1317
rect 36921 1271 36991 1317
rect 37037 1271 37107 1317
rect 37153 1271 37223 1317
rect 37269 1271 37339 1317
rect 37385 1271 37455 1317
rect 37501 1271 37571 1317
rect 37617 1271 37687 1317
rect 37733 1271 37803 1317
rect 37849 1271 37919 1317
rect 37965 1271 38035 1317
rect 38081 1271 38151 1317
rect 38197 1271 38267 1317
rect 38313 1271 38383 1317
rect 38429 1271 38499 1317
rect 38545 1271 38615 1317
rect 38661 1271 38731 1317
rect 38777 1271 38847 1317
rect 38893 1271 38963 1317
rect 39009 1271 39079 1317
rect 39125 1271 39195 1317
rect 39241 1271 39311 1317
rect 39357 1271 39427 1317
rect 39473 1271 39543 1317
rect 39589 1271 39659 1317
rect 39705 1271 39775 1317
rect 39821 1271 39891 1317
rect 39937 1271 40007 1317
rect 40053 1271 40123 1317
rect 40169 1271 40188 1317
rect 28620 1201 40188 1271
rect 28620 1155 28639 1201
rect 28685 1155 28755 1201
rect 28801 1155 28871 1201
rect 28917 1155 28987 1201
rect 29033 1155 29103 1201
rect 29149 1155 29219 1201
rect 29265 1155 29335 1201
rect 29381 1155 29451 1201
rect 29497 1155 29567 1201
rect 29613 1155 29683 1201
rect 29729 1155 29799 1201
rect 29845 1155 29915 1201
rect 29961 1155 30031 1201
rect 30077 1155 30147 1201
rect 30193 1155 30263 1201
rect 30309 1155 30379 1201
rect 30425 1155 30495 1201
rect 30541 1155 30611 1201
rect 30657 1155 30727 1201
rect 30773 1155 30843 1201
rect 30889 1155 30959 1201
rect 31005 1155 31075 1201
rect 31121 1155 31191 1201
rect 31237 1155 31307 1201
rect 31353 1155 31423 1201
rect 31469 1155 31539 1201
rect 31585 1155 31655 1201
rect 31701 1155 31771 1201
rect 31817 1155 31887 1201
rect 31933 1155 32003 1201
rect 32049 1155 32119 1201
rect 32165 1155 32235 1201
rect 32281 1155 32351 1201
rect 32397 1155 32467 1201
rect 32513 1155 32583 1201
rect 32629 1155 32699 1201
rect 32745 1155 32815 1201
rect 32861 1155 32931 1201
rect 32977 1155 33047 1201
rect 33093 1155 33163 1201
rect 33209 1155 33279 1201
rect 33325 1155 33395 1201
rect 33441 1155 33511 1201
rect 33557 1155 33627 1201
rect 33673 1155 33743 1201
rect 33789 1155 33859 1201
rect 33905 1155 33975 1201
rect 34021 1155 34091 1201
rect 34137 1155 34207 1201
rect 34253 1155 34323 1201
rect 34369 1155 34439 1201
rect 34485 1155 34555 1201
rect 34601 1155 34671 1201
rect 34717 1155 34787 1201
rect 34833 1155 34903 1201
rect 34949 1155 35019 1201
rect 35065 1155 35135 1201
rect 35181 1155 35251 1201
rect 35297 1155 35367 1201
rect 35413 1155 35483 1201
rect 35529 1155 35599 1201
rect 35645 1155 35715 1201
rect 35761 1155 35831 1201
rect 35877 1155 35947 1201
rect 35993 1155 36063 1201
rect 36109 1155 36179 1201
rect 36225 1155 36295 1201
rect 36341 1155 36411 1201
rect 36457 1155 36527 1201
rect 36573 1155 36643 1201
rect 36689 1155 36759 1201
rect 36805 1155 36875 1201
rect 36921 1155 36991 1201
rect 37037 1155 37107 1201
rect 37153 1155 37223 1201
rect 37269 1155 37339 1201
rect 37385 1155 37455 1201
rect 37501 1155 37571 1201
rect 37617 1155 37687 1201
rect 37733 1155 37803 1201
rect 37849 1155 37919 1201
rect 37965 1155 38035 1201
rect 38081 1155 38151 1201
rect 38197 1155 38267 1201
rect 38313 1155 38383 1201
rect 38429 1155 38499 1201
rect 38545 1155 38615 1201
rect 38661 1155 38731 1201
rect 38777 1155 38847 1201
rect 38893 1155 38963 1201
rect 39009 1155 39079 1201
rect 39125 1155 39195 1201
rect 39241 1155 39311 1201
rect 39357 1155 39427 1201
rect 39473 1155 39543 1201
rect 39589 1155 39659 1201
rect 39705 1155 39775 1201
rect 39821 1155 39891 1201
rect 39937 1155 40007 1201
rect 40053 1155 40123 1201
rect 40169 1155 40188 1201
rect 28620 1034 40188 1155
rect 50826 3844 50845 3890
rect 50891 3844 50961 3890
rect 51007 3844 51077 3890
rect 51123 3844 51193 3890
rect 51239 3844 51309 3890
rect 51355 3844 51425 3890
rect 51471 3844 51541 3890
rect 51587 3844 51657 3890
rect 51703 3844 51773 3890
rect 51819 3844 51889 3890
rect 51935 3844 52005 3890
rect 52051 3844 52121 3890
rect 52167 3844 52237 3890
rect 52283 3844 52353 3890
rect 52399 3844 52469 3890
rect 52515 3844 52585 3890
rect 52631 3844 52701 3890
rect 52747 3844 52817 3890
rect 52863 3844 52933 3890
rect 52979 3844 53049 3890
rect 53095 3844 53165 3890
rect 53211 3844 53281 3890
rect 53327 3844 53397 3890
rect 53443 3844 53513 3890
rect 53559 3844 53629 3890
rect 53675 3844 53745 3890
rect 53791 3844 53861 3890
rect 53907 3844 53977 3890
rect 54023 3844 54093 3890
rect 54139 3844 54209 3890
rect 54255 3844 54325 3890
rect 54371 3844 54441 3890
rect 54487 3844 54557 3890
rect 54603 3844 54673 3890
rect 54719 3844 54789 3890
rect 54835 3844 54905 3890
rect 54951 3844 55021 3890
rect 55067 3844 55137 3890
rect 55183 3844 55253 3890
rect 55299 3844 55369 3890
rect 55415 3844 55485 3890
rect 55531 3844 55601 3890
rect 55647 3844 55717 3890
rect 55763 3844 55833 3890
rect 55879 3844 55949 3890
rect 55995 3844 56065 3890
rect 56111 3844 56181 3890
rect 56227 3844 56297 3890
rect 56343 3844 56413 3890
rect 56459 3844 56529 3890
rect 56575 3844 56594 3890
rect 50826 3774 56594 3844
rect 50826 3728 50845 3774
rect 50891 3728 50961 3774
rect 51007 3728 51077 3774
rect 51123 3728 51193 3774
rect 51239 3728 51309 3774
rect 51355 3728 51425 3774
rect 51471 3728 51541 3774
rect 51587 3728 51657 3774
rect 51703 3728 51773 3774
rect 51819 3728 51889 3774
rect 51935 3728 52005 3774
rect 52051 3728 52121 3774
rect 52167 3728 52237 3774
rect 52283 3728 52353 3774
rect 52399 3728 52469 3774
rect 52515 3728 52585 3774
rect 52631 3728 52701 3774
rect 52747 3728 52817 3774
rect 52863 3728 52933 3774
rect 52979 3728 53049 3774
rect 53095 3728 53165 3774
rect 53211 3728 53281 3774
rect 53327 3728 53397 3774
rect 53443 3728 53513 3774
rect 53559 3728 53629 3774
rect 53675 3728 53745 3774
rect 53791 3728 53861 3774
rect 53907 3728 53977 3774
rect 54023 3728 54093 3774
rect 54139 3728 54209 3774
rect 54255 3728 54325 3774
rect 54371 3728 54441 3774
rect 54487 3728 54557 3774
rect 54603 3728 54673 3774
rect 54719 3728 54789 3774
rect 54835 3728 54905 3774
rect 54951 3728 55021 3774
rect 55067 3728 55137 3774
rect 55183 3728 55253 3774
rect 55299 3728 55369 3774
rect 55415 3728 55485 3774
rect 55531 3728 55601 3774
rect 55647 3728 55717 3774
rect 55763 3728 55833 3774
rect 55879 3728 55949 3774
rect 55995 3728 56065 3774
rect 56111 3728 56181 3774
rect 56227 3728 56297 3774
rect 56343 3728 56413 3774
rect 56459 3728 56529 3774
rect 56575 3728 56594 3774
rect 50826 3658 56594 3728
rect 50826 3612 50845 3658
rect 50891 3612 50961 3658
rect 51007 3612 51077 3658
rect 51123 3612 51193 3658
rect 51239 3612 51309 3658
rect 51355 3612 51425 3658
rect 51471 3612 51541 3658
rect 51587 3612 51657 3658
rect 51703 3612 51773 3658
rect 51819 3612 51889 3658
rect 51935 3612 52005 3658
rect 52051 3612 52121 3658
rect 52167 3612 52237 3658
rect 52283 3612 52353 3658
rect 52399 3612 52469 3658
rect 52515 3612 52585 3658
rect 52631 3612 52701 3658
rect 52747 3612 52817 3658
rect 52863 3612 52933 3658
rect 52979 3612 53049 3658
rect 53095 3612 53165 3658
rect 53211 3612 53281 3658
rect 53327 3612 53397 3658
rect 53443 3612 53513 3658
rect 53559 3612 53629 3658
rect 53675 3612 53745 3658
rect 53791 3612 53861 3658
rect 53907 3612 53977 3658
rect 54023 3612 54093 3658
rect 54139 3612 54209 3658
rect 54255 3612 54325 3658
rect 54371 3612 54441 3658
rect 54487 3612 54557 3658
rect 54603 3612 54673 3658
rect 54719 3612 54789 3658
rect 54835 3612 54905 3658
rect 54951 3612 55021 3658
rect 55067 3612 55137 3658
rect 55183 3612 55253 3658
rect 55299 3612 55369 3658
rect 55415 3612 55485 3658
rect 55531 3612 55601 3658
rect 55647 3612 55717 3658
rect 55763 3612 55833 3658
rect 55879 3612 55949 3658
rect 55995 3612 56065 3658
rect 56111 3612 56181 3658
rect 56227 3612 56297 3658
rect 56343 3612 56413 3658
rect 56459 3612 56529 3658
rect 56575 3612 56594 3658
rect 50826 3542 56594 3612
rect 50826 3496 50845 3542
rect 50891 3496 50961 3542
rect 51007 3496 51077 3542
rect 51123 3496 51193 3542
rect 51239 3496 51309 3542
rect 51355 3496 51425 3542
rect 51471 3496 51541 3542
rect 51587 3496 51657 3542
rect 51703 3496 51773 3542
rect 51819 3496 51889 3542
rect 51935 3496 52005 3542
rect 52051 3496 52121 3542
rect 52167 3496 52237 3542
rect 52283 3496 52353 3542
rect 52399 3496 52469 3542
rect 52515 3496 52585 3542
rect 52631 3496 52701 3542
rect 52747 3496 52817 3542
rect 52863 3496 52933 3542
rect 52979 3496 53049 3542
rect 53095 3496 53165 3542
rect 53211 3496 53281 3542
rect 53327 3496 53397 3542
rect 53443 3496 53513 3542
rect 53559 3496 53629 3542
rect 53675 3496 53745 3542
rect 53791 3496 53861 3542
rect 53907 3496 53977 3542
rect 54023 3496 54093 3542
rect 54139 3496 54209 3542
rect 54255 3496 54325 3542
rect 54371 3496 54441 3542
rect 54487 3496 54557 3542
rect 54603 3496 54673 3542
rect 54719 3496 54789 3542
rect 54835 3496 54905 3542
rect 54951 3496 55021 3542
rect 55067 3496 55137 3542
rect 55183 3496 55253 3542
rect 55299 3496 55369 3542
rect 55415 3496 55485 3542
rect 55531 3496 55601 3542
rect 55647 3496 55717 3542
rect 55763 3496 55833 3542
rect 55879 3496 55949 3542
rect 55995 3496 56065 3542
rect 56111 3496 56181 3542
rect 56227 3496 56297 3542
rect 56343 3496 56413 3542
rect 56459 3496 56529 3542
rect 56575 3496 56594 3542
rect 50826 3426 56594 3496
rect 50826 3380 50845 3426
rect 50891 3380 50961 3426
rect 51007 3380 51077 3426
rect 51123 3380 51193 3426
rect 51239 3380 51309 3426
rect 51355 3380 51425 3426
rect 51471 3380 51541 3426
rect 51587 3380 51657 3426
rect 51703 3380 51773 3426
rect 51819 3380 51889 3426
rect 51935 3380 52005 3426
rect 52051 3380 52121 3426
rect 52167 3380 52237 3426
rect 52283 3380 52353 3426
rect 52399 3380 52469 3426
rect 52515 3380 52585 3426
rect 52631 3380 52701 3426
rect 52747 3380 52817 3426
rect 52863 3380 52933 3426
rect 52979 3380 53049 3426
rect 53095 3380 53165 3426
rect 53211 3380 53281 3426
rect 53327 3380 53397 3426
rect 53443 3380 53513 3426
rect 53559 3380 53629 3426
rect 53675 3380 53745 3426
rect 53791 3380 53861 3426
rect 53907 3380 53977 3426
rect 54023 3380 54093 3426
rect 54139 3380 54209 3426
rect 54255 3380 54325 3426
rect 54371 3380 54441 3426
rect 54487 3380 54557 3426
rect 54603 3380 54673 3426
rect 54719 3380 54789 3426
rect 54835 3380 54905 3426
rect 54951 3380 55021 3426
rect 55067 3380 55137 3426
rect 55183 3380 55253 3426
rect 55299 3380 55369 3426
rect 55415 3380 55485 3426
rect 55531 3380 55601 3426
rect 55647 3380 55717 3426
rect 55763 3380 55833 3426
rect 55879 3380 55949 3426
rect 55995 3380 56065 3426
rect 56111 3380 56181 3426
rect 56227 3380 56297 3426
rect 56343 3380 56413 3426
rect 56459 3380 56529 3426
rect 56575 3380 56594 3426
rect 50826 3310 56594 3380
rect 50826 3264 50845 3310
rect 50891 3264 50961 3310
rect 51007 3264 51077 3310
rect 51123 3264 51193 3310
rect 51239 3264 51309 3310
rect 51355 3264 51425 3310
rect 51471 3264 51541 3310
rect 51587 3264 51657 3310
rect 51703 3264 51773 3310
rect 51819 3264 51889 3310
rect 51935 3264 52005 3310
rect 52051 3264 52121 3310
rect 52167 3264 52237 3310
rect 52283 3264 52353 3310
rect 52399 3264 52469 3310
rect 52515 3264 52585 3310
rect 52631 3264 52701 3310
rect 52747 3264 52817 3310
rect 52863 3264 52933 3310
rect 52979 3264 53049 3310
rect 53095 3264 53165 3310
rect 53211 3264 53281 3310
rect 53327 3264 53397 3310
rect 53443 3264 53513 3310
rect 53559 3264 53629 3310
rect 53675 3264 53745 3310
rect 53791 3264 53861 3310
rect 53907 3264 53977 3310
rect 54023 3264 54093 3310
rect 54139 3264 54209 3310
rect 54255 3264 54325 3310
rect 54371 3264 54441 3310
rect 54487 3264 54557 3310
rect 54603 3264 54673 3310
rect 54719 3264 54789 3310
rect 54835 3264 54905 3310
rect 54951 3264 55021 3310
rect 55067 3264 55137 3310
rect 55183 3264 55253 3310
rect 55299 3264 55369 3310
rect 55415 3264 55485 3310
rect 55531 3264 55601 3310
rect 55647 3264 55717 3310
rect 55763 3264 55833 3310
rect 55879 3264 55949 3310
rect 55995 3264 56065 3310
rect 56111 3264 56181 3310
rect 56227 3264 56297 3310
rect 56343 3264 56413 3310
rect 56459 3264 56529 3310
rect 56575 3264 56594 3310
rect 50826 3194 56594 3264
rect 50826 3148 50845 3194
rect 50891 3148 50961 3194
rect 51007 3148 51077 3194
rect 51123 3148 51193 3194
rect 51239 3148 51309 3194
rect 51355 3148 51425 3194
rect 51471 3148 51541 3194
rect 51587 3148 51657 3194
rect 51703 3148 51773 3194
rect 51819 3148 51889 3194
rect 51935 3148 52005 3194
rect 52051 3148 52121 3194
rect 52167 3148 52237 3194
rect 52283 3148 52353 3194
rect 52399 3148 52469 3194
rect 52515 3148 52585 3194
rect 52631 3148 52701 3194
rect 52747 3148 52817 3194
rect 52863 3148 52933 3194
rect 52979 3148 53049 3194
rect 53095 3148 53165 3194
rect 53211 3148 53281 3194
rect 53327 3148 53397 3194
rect 53443 3148 53513 3194
rect 53559 3148 53629 3194
rect 53675 3148 53745 3194
rect 53791 3148 53861 3194
rect 53907 3148 53977 3194
rect 54023 3148 54093 3194
rect 54139 3148 54209 3194
rect 54255 3148 54325 3194
rect 54371 3148 54441 3194
rect 54487 3148 54557 3194
rect 54603 3148 54673 3194
rect 54719 3148 54789 3194
rect 54835 3148 54905 3194
rect 54951 3148 55021 3194
rect 55067 3148 55137 3194
rect 55183 3148 55253 3194
rect 55299 3148 55369 3194
rect 55415 3148 55485 3194
rect 55531 3148 55601 3194
rect 55647 3148 55717 3194
rect 55763 3148 55833 3194
rect 55879 3148 55949 3194
rect 55995 3148 56065 3194
rect 56111 3148 56181 3194
rect 56227 3148 56297 3194
rect 56343 3148 56413 3194
rect 56459 3148 56529 3194
rect 56575 3148 56594 3194
rect 50826 3078 56594 3148
rect 50826 3032 50845 3078
rect 50891 3032 50961 3078
rect 51007 3032 51077 3078
rect 51123 3032 51193 3078
rect 51239 3032 51309 3078
rect 51355 3032 51425 3078
rect 51471 3032 51541 3078
rect 51587 3032 51657 3078
rect 51703 3032 51773 3078
rect 51819 3032 51889 3078
rect 51935 3032 52005 3078
rect 52051 3032 52121 3078
rect 52167 3032 52237 3078
rect 52283 3032 52353 3078
rect 52399 3032 52469 3078
rect 52515 3032 52585 3078
rect 52631 3032 52701 3078
rect 52747 3032 52817 3078
rect 52863 3032 52933 3078
rect 52979 3032 53049 3078
rect 53095 3032 53165 3078
rect 53211 3032 53281 3078
rect 53327 3032 53397 3078
rect 53443 3032 53513 3078
rect 53559 3032 53629 3078
rect 53675 3032 53745 3078
rect 53791 3032 53861 3078
rect 53907 3032 53977 3078
rect 54023 3032 54093 3078
rect 54139 3032 54209 3078
rect 54255 3032 54325 3078
rect 54371 3032 54441 3078
rect 54487 3032 54557 3078
rect 54603 3032 54673 3078
rect 54719 3032 54789 3078
rect 54835 3032 54905 3078
rect 54951 3032 55021 3078
rect 55067 3032 55137 3078
rect 55183 3032 55253 3078
rect 55299 3032 55369 3078
rect 55415 3032 55485 3078
rect 55531 3032 55601 3078
rect 55647 3032 55717 3078
rect 55763 3032 55833 3078
rect 55879 3032 55949 3078
rect 55995 3032 56065 3078
rect 56111 3032 56181 3078
rect 56227 3032 56297 3078
rect 56343 3032 56413 3078
rect 56459 3032 56529 3078
rect 56575 3032 56594 3078
rect 50826 2962 56594 3032
rect 50826 2916 50845 2962
rect 50891 2916 50961 2962
rect 51007 2916 51077 2962
rect 51123 2916 51193 2962
rect 51239 2916 51309 2962
rect 51355 2916 51425 2962
rect 51471 2916 51541 2962
rect 51587 2916 51657 2962
rect 51703 2916 51773 2962
rect 51819 2916 51889 2962
rect 51935 2916 52005 2962
rect 52051 2916 52121 2962
rect 52167 2916 52237 2962
rect 52283 2916 52353 2962
rect 52399 2916 52469 2962
rect 52515 2916 52585 2962
rect 52631 2916 52701 2962
rect 52747 2916 52817 2962
rect 52863 2916 52933 2962
rect 52979 2916 53049 2962
rect 53095 2916 53165 2962
rect 53211 2916 53281 2962
rect 53327 2916 53397 2962
rect 53443 2916 53513 2962
rect 53559 2916 53629 2962
rect 53675 2916 53745 2962
rect 53791 2916 53861 2962
rect 53907 2916 53977 2962
rect 54023 2916 54093 2962
rect 54139 2916 54209 2962
rect 54255 2916 54325 2962
rect 54371 2916 54441 2962
rect 54487 2916 54557 2962
rect 54603 2916 54673 2962
rect 54719 2916 54789 2962
rect 54835 2916 54905 2962
rect 54951 2916 55021 2962
rect 55067 2916 55137 2962
rect 55183 2916 55253 2962
rect 55299 2916 55369 2962
rect 55415 2916 55485 2962
rect 55531 2916 55601 2962
rect 55647 2916 55717 2962
rect 55763 2916 55833 2962
rect 55879 2916 55949 2962
rect 55995 2916 56065 2962
rect 56111 2916 56181 2962
rect 56227 2916 56297 2962
rect 56343 2916 56413 2962
rect 56459 2916 56529 2962
rect 56575 2916 56594 2962
rect 50826 2846 56594 2916
rect 50826 2800 50845 2846
rect 50891 2800 50961 2846
rect 51007 2800 51077 2846
rect 51123 2800 51193 2846
rect 51239 2800 51309 2846
rect 51355 2800 51425 2846
rect 51471 2800 51541 2846
rect 51587 2800 51657 2846
rect 51703 2800 51773 2846
rect 51819 2800 51889 2846
rect 51935 2800 52005 2846
rect 52051 2800 52121 2846
rect 52167 2800 52237 2846
rect 52283 2800 52353 2846
rect 52399 2800 52469 2846
rect 52515 2800 52585 2846
rect 52631 2800 52701 2846
rect 52747 2800 52817 2846
rect 52863 2800 52933 2846
rect 52979 2800 53049 2846
rect 53095 2800 53165 2846
rect 53211 2800 53281 2846
rect 53327 2800 53397 2846
rect 53443 2800 53513 2846
rect 53559 2800 53629 2846
rect 53675 2800 53745 2846
rect 53791 2800 53861 2846
rect 53907 2800 53977 2846
rect 54023 2800 54093 2846
rect 54139 2800 54209 2846
rect 54255 2800 54325 2846
rect 54371 2800 54441 2846
rect 54487 2800 54557 2846
rect 54603 2800 54673 2846
rect 54719 2800 54789 2846
rect 54835 2800 54905 2846
rect 54951 2800 55021 2846
rect 55067 2800 55137 2846
rect 55183 2800 55253 2846
rect 55299 2800 55369 2846
rect 55415 2800 55485 2846
rect 55531 2800 55601 2846
rect 55647 2800 55717 2846
rect 55763 2800 55833 2846
rect 55879 2800 55949 2846
rect 55995 2800 56065 2846
rect 56111 2800 56181 2846
rect 56227 2800 56297 2846
rect 56343 2800 56413 2846
rect 56459 2800 56529 2846
rect 56575 2800 56594 2846
rect 50826 2730 56594 2800
rect 50826 2684 50845 2730
rect 50891 2684 50961 2730
rect 51007 2684 51077 2730
rect 51123 2684 51193 2730
rect 51239 2684 51309 2730
rect 51355 2684 51425 2730
rect 51471 2684 51541 2730
rect 51587 2684 51657 2730
rect 51703 2684 51773 2730
rect 51819 2684 51889 2730
rect 51935 2684 52005 2730
rect 52051 2684 52121 2730
rect 52167 2684 52237 2730
rect 52283 2684 52353 2730
rect 52399 2684 52469 2730
rect 52515 2684 52585 2730
rect 52631 2684 52701 2730
rect 52747 2684 52817 2730
rect 52863 2684 52933 2730
rect 52979 2684 53049 2730
rect 53095 2684 53165 2730
rect 53211 2684 53281 2730
rect 53327 2684 53397 2730
rect 53443 2684 53513 2730
rect 53559 2684 53629 2730
rect 53675 2684 53745 2730
rect 53791 2684 53861 2730
rect 53907 2684 53977 2730
rect 54023 2684 54093 2730
rect 54139 2684 54209 2730
rect 54255 2684 54325 2730
rect 54371 2684 54441 2730
rect 54487 2684 54557 2730
rect 54603 2684 54673 2730
rect 54719 2684 54789 2730
rect 54835 2684 54905 2730
rect 54951 2684 55021 2730
rect 55067 2684 55137 2730
rect 55183 2684 55253 2730
rect 55299 2684 55369 2730
rect 55415 2684 55485 2730
rect 55531 2684 55601 2730
rect 55647 2684 55717 2730
rect 55763 2684 55833 2730
rect 55879 2684 55949 2730
rect 55995 2684 56065 2730
rect 56111 2684 56181 2730
rect 56227 2684 56297 2730
rect 56343 2684 56413 2730
rect 56459 2684 56529 2730
rect 56575 2684 56594 2730
rect 50826 2614 56594 2684
rect 50826 2568 50845 2614
rect 50891 2568 50961 2614
rect 51007 2568 51077 2614
rect 51123 2568 51193 2614
rect 51239 2568 51309 2614
rect 51355 2568 51425 2614
rect 51471 2568 51541 2614
rect 51587 2568 51657 2614
rect 51703 2568 51773 2614
rect 51819 2568 51889 2614
rect 51935 2568 52005 2614
rect 52051 2568 52121 2614
rect 52167 2568 52237 2614
rect 52283 2568 52353 2614
rect 52399 2568 52469 2614
rect 52515 2568 52585 2614
rect 52631 2568 52701 2614
rect 52747 2568 52817 2614
rect 52863 2568 52933 2614
rect 52979 2568 53049 2614
rect 53095 2568 53165 2614
rect 53211 2568 53281 2614
rect 53327 2568 53397 2614
rect 53443 2568 53513 2614
rect 53559 2568 53629 2614
rect 53675 2568 53745 2614
rect 53791 2568 53861 2614
rect 53907 2568 53977 2614
rect 54023 2568 54093 2614
rect 54139 2568 54209 2614
rect 54255 2568 54325 2614
rect 54371 2568 54441 2614
rect 54487 2568 54557 2614
rect 54603 2568 54673 2614
rect 54719 2568 54789 2614
rect 54835 2568 54905 2614
rect 54951 2568 55021 2614
rect 55067 2568 55137 2614
rect 55183 2568 55253 2614
rect 55299 2568 55369 2614
rect 55415 2568 55485 2614
rect 55531 2568 55601 2614
rect 55647 2568 55717 2614
rect 55763 2568 55833 2614
rect 55879 2568 55949 2614
rect 55995 2568 56065 2614
rect 56111 2568 56181 2614
rect 56227 2568 56297 2614
rect 56343 2568 56413 2614
rect 56459 2568 56529 2614
rect 56575 2568 56594 2614
rect 50826 2498 56594 2568
rect 50826 2452 50845 2498
rect 50891 2452 50961 2498
rect 51007 2452 51077 2498
rect 51123 2452 51193 2498
rect 51239 2452 51309 2498
rect 51355 2452 51425 2498
rect 51471 2452 51541 2498
rect 51587 2452 51657 2498
rect 51703 2452 51773 2498
rect 51819 2452 51889 2498
rect 51935 2452 52005 2498
rect 52051 2452 52121 2498
rect 52167 2452 52237 2498
rect 52283 2452 52353 2498
rect 52399 2452 52469 2498
rect 52515 2452 52585 2498
rect 52631 2452 52701 2498
rect 52747 2452 52817 2498
rect 52863 2452 52933 2498
rect 52979 2452 53049 2498
rect 53095 2452 53165 2498
rect 53211 2452 53281 2498
rect 53327 2452 53397 2498
rect 53443 2452 53513 2498
rect 53559 2452 53629 2498
rect 53675 2452 53745 2498
rect 53791 2452 53861 2498
rect 53907 2452 53977 2498
rect 54023 2452 54093 2498
rect 54139 2452 54209 2498
rect 54255 2452 54325 2498
rect 54371 2452 54441 2498
rect 54487 2452 54557 2498
rect 54603 2452 54673 2498
rect 54719 2452 54789 2498
rect 54835 2452 54905 2498
rect 54951 2452 55021 2498
rect 55067 2452 55137 2498
rect 55183 2452 55253 2498
rect 55299 2452 55369 2498
rect 55415 2452 55485 2498
rect 55531 2452 55601 2498
rect 55647 2452 55717 2498
rect 55763 2452 55833 2498
rect 55879 2452 55949 2498
rect 55995 2452 56065 2498
rect 56111 2452 56181 2498
rect 56227 2452 56297 2498
rect 56343 2452 56413 2498
rect 56459 2452 56529 2498
rect 56575 2452 56594 2498
rect 50826 2382 56594 2452
rect 50826 2336 50845 2382
rect 50891 2336 50961 2382
rect 51007 2336 51077 2382
rect 51123 2336 51193 2382
rect 51239 2336 51309 2382
rect 51355 2336 51425 2382
rect 51471 2336 51541 2382
rect 51587 2336 51657 2382
rect 51703 2336 51773 2382
rect 51819 2336 51889 2382
rect 51935 2336 52005 2382
rect 52051 2336 52121 2382
rect 52167 2336 52237 2382
rect 52283 2336 52353 2382
rect 52399 2336 52469 2382
rect 52515 2336 52585 2382
rect 52631 2336 52701 2382
rect 52747 2336 52817 2382
rect 52863 2336 52933 2382
rect 52979 2336 53049 2382
rect 53095 2336 53165 2382
rect 53211 2336 53281 2382
rect 53327 2336 53397 2382
rect 53443 2336 53513 2382
rect 53559 2336 53629 2382
rect 53675 2336 53745 2382
rect 53791 2336 53861 2382
rect 53907 2336 53977 2382
rect 54023 2336 54093 2382
rect 54139 2336 54209 2382
rect 54255 2336 54325 2382
rect 54371 2336 54441 2382
rect 54487 2336 54557 2382
rect 54603 2336 54673 2382
rect 54719 2336 54789 2382
rect 54835 2336 54905 2382
rect 54951 2336 55021 2382
rect 55067 2336 55137 2382
rect 55183 2336 55253 2382
rect 55299 2336 55369 2382
rect 55415 2336 55485 2382
rect 55531 2336 55601 2382
rect 55647 2336 55717 2382
rect 55763 2336 55833 2382
rect 55879 2336 55949 2382
rect 55995 2336 56065 2382
rect 56111 2336 56181 2382
rect 56227 2336 56297 2382
rect 56343 2336 56413 2382
rect 56459 2336 56529 2382
rect 56575 2336 56594 2382
rect 50826 2266 56594 2336
rect 50826 2220 50845 2266
rect 50891 2220 50961 2266
rect 51007 2220 51077 2266
rect 51123 2220 51193 2266
rect 51239 2220 51309 2266
rect 51355 2220 51425 2266
rect 51471 2220 51541 2266
rect 51587 2220 51657 2266
rect 51703 2220 51773 2266
rect 51819 2220 51889 2266
rect 51935 2220 52005 2266
rect 52051 2220 52121 2266
rect 52167 2220 52237 2266
rect 52283 2220 52353 2266
rect 52399 2220 52469 2266
rect 52515 2220 52585 2266
rect 52631 2220 52701 2266
rect 52747 2220 52817 2266
rect 52863 2220 52933 2266
rect 52979 2220 53049 2266
rect 53095 2220 53165 2266
rect 53211 2220 53281 2266
rect 53327 2220 53397 2266
rect 53443 2220 53513 2266
rect 53559 2220 53629 2266
rect 53675 2220 53745 2266
rect 53791 2220 53861 2266
rect 53907 2220 53977 2266
rect 54023 2220 54093 2266
rect 54139 2220 54209 2266
rect 54255 2220 54325 2266
rect 54371 2220 54441 2266
rect 54487 2220 54557 2266
rect 54603 2220 54673 2266
rect 54719 2220 54789 2266
rect 54835 2220 54905 2266
rect 54951 2220 55021 2266
rect 55067 2220 55137 2266
rect 55183 2220 55253 2266
rect 55299 2220 55369 2266
rect 55415 2220 55485 2266
rect 55531 2220 55601 2266
rect 55647 2220 55717 2266
rect 55763 2220 55833 2266
rect 55879 2220 55949 2266
rect 55995 2220 56065 2266
rect 56111 2220 56181 2266
rect 56227 2220 56297 2266
rect 56343 2220 56413 2266
rect 56459 2220 56529 2266
rect 56575 2220 56594 2266
rect 50826 2150 56594 2220
rect 50826 2104 50845 2150
rect 50891 2104 50961 2150
rect 51007 2104 51077 2150
rect 51123 2104 51193 2150
rect 51239 2104 51309 2150
rect 51355 2104 51425 2150
rect 51471 2104 51541 2150
rect 51587 2104 51657 2150
rect 51703 2104 51773 2150
rect 51819 2104 51889 2150
rect 51935 2104 52005 2150
rect 52051 2104 52121 2150
rect 52167 2104 52237 2150
rect 52283 2104 52353 2150
rect 52399 2104 52469 2150
rect 52515 2104 52585 2150
rect 52631 2104 52701 2150
rect 52747 2104 52817 2150
rect 52863 2104 52933 2150
rect 52979 2104 53049 2150
rect 53095 2104 53165 2150
rect 53211 2104 53281 2150
rect 53327 2104 53397 2150
rect 53443 2104 53513 2150
rect 53559 2104 53629 2150
rect 53675 2104 53745 2150
rect 53791 2104 53861 2150
rect 53907 2104 53977 2150
rect 54023 2104 54093 2150
rect 54139 2104 54209 2150
rect 54255 2104 54325 2150
rect 54371 2104 54441 2150
rect 54487 2104 54557 2150
rect 54603 2104 54673 2150
rect 54719 2104 54789 2150
rect 54835 2104 54905 2150
rect 54951 2104 55021 2150
rect 55067 2104 55137 2150
rect 55183 2104 55253 2150
rect 55299 2104 55369 2150
rect 55415 2104 55485 2150
rect 55531 2104 55601 2150
rect 55647 2104 55717 2150
rect 55763 2104 55833 2150
rect 55879 2104 55949 2150
rect 55995 2104 56065 2150
rect 56111 2104 56181 2150
rect 56227 2104 56297 2150
rect 56343 2104 56413 2150
rect 56459 2104 56529 2150
rect 56575 2104 56594 2150
rect 50826 2034 56594 2104
rect 50826 1988 50845 2034
rect 50891 1988 50961 2034
rect 51007 1988 51077 2034
rect 51123 1988 51193 2034
rect 51239 1988 51309 2034
rect 51355 1988 51425 2034
rect 51471 1988 51541 2034
rect 51587 1988 51657 2034
rect 51703 1988 51773 2034
rect 51819 1988 51889 2034
rect 51935 1988 52005 2034
rect 52051 1988 52121 2034
rect 52167 1988 52237 2034
rect 52283 1988 52353 2034
rect 52399 1988 52469 2034
rect 52515 1988 52585 2034
rect 52631 1988 52701 2034
rect 52747 1988 52817 2034
rect 52863 1988 52933 2034
rect 52979 1988 53049 2034
rect 53095 1988 53165 2034
rect 53211 1988 53281 2034
rect 53327 1988 53397 2034
rect 53443 1988 53513 2034
rect 53559 1988 53629 2034
rect 53675 1988 53745 2034
rect 53791 1988 53861 2034
rect 53907 1988 53977 2034
rect 54023 1988 54093 2034
rect 54139 1988 54209 2034
rect 54255 1988 54325 2034
rect 54371 1988 54441 2034
rect 54487 1988 54557 2034
rect 54603 1988 54673 2034
rect 54719 1988 54789 2034
rect 54835 1988 54905 2034
rect 54951 1988 55021 2034
rect 55067 1988 55137 2034
rect 55183 1988 55253 2034
rect 55299 1988 55369 2034
rect 55415 1988 55485 2034
rect 55531 1988 55601 2034
rect 55647 1988 55717 2034
rect 55763 1988 55833 2034
rect 55879 1988 55949 2034
rect 55995 1988 56065 2034
rect 56111 1988 56181 2034
rect 56227 1988 56297 2034
rect 56343 1988 56413 2034
rect 56459 1988 56529 2034
rect 56575 1988 56594 2034
rect 50826 1918 56594 1988
rect 50826 1872 50845 1918
rect 50891 1872 50961 1918
rect 51007 1872 51077 1918
rect 51123 1872 51193 1918
rect 51239 1872 51309 1918
rect 51355 1872 51425 1918
rect 51471 1872 51541 1918
rect 51587 1872 51657 1918
rect 51703 1872 51773 1918
rect 51819 1872 51889 1918
rect 51935 1872 52005 1918
rect 52051 1872 52121 1918
rect 52167 1872 52237 1918
rect 52283 1872 52353 1918
rect 52399 1872 52469 1918
rect 52515 1872 52585 1918
rect 52631 1872 52701 1918
rect 52747 1872 52817 1918
rect 52863 1872 52933 1918
rect 52979 1872 53049 1918
rect 53095 1872 53165 1918
rect 53211 1872 53281 1918
rect 53327 1872 53397 1918
rect 53443 1872 53513 1918
rect 53559 1872 53629 1918
rect 53675 1872 53745 1918
rect 53791 1872 53861 1918
rect 53907 1872 53977 1918
rect 54023 1872 54093 1918
rect 54139 1872 54209 1918
rect 54255 1872 54325 1918
rect 54371 1872 54441 1918
rect 54487 1872 54557 1918
rect 54603 1872 54673 1918
rect 54719 1872 54789 1918
rect 54835 1872 54905 1918
rect 54951 1872 55021 1918
rect 55067 1872 55137 1918
rect 55183 1872 55253 1918
rect 55299 1872 55369 1918
rect 55415 1872 55485 1918
rect 55531 1872 55601 1918
rect 55647 1872 55717 1918
rect 55763 1872 55833 1918
rect 55879 1872 55949 1918
rect 55995 1872 56065 1918
rect 56111 1872 56181 1918
rect 56227 1872 56297 1918
rect 56343 1872 56413 1918
rect 56459 1872 56529 1918
rect 56575 1872 56594 1918
rect 50826 1802 56594 1872
rect 50826 1756 50845 1802
rect 50891 1756 50961 1802
rect 51007 1756 51077 1802
rect 51123 1756 51193 1802
rect 51239 1756 51309 1802
rect 51355 1756 51425 1802
rect 51471 1756 51541 1802
rect 51587 1756 51657 1802
rect 51703 1756 51773 1802
rect 51819 1756 51889 1802
rect 51935 1756 52005 1802
rect 52051 1756 52121 1802
rect 52167 1756 52237 1802
rect 52283 1756 52353 1802
rect 52399 1756 52469 1802
rect 52515 1756 52585 1802
rect 52631 1756 52701 1802
rect 52747 1756 52817 1802
rect 52863 1756 52933 1802
rect 52979 1756 53049 1802
rect 53095 1756 53165 1802
rect 53211 1756 53281 1802
rect 53327 1756 53397 1802
rect 53443 1756 53513 1802
rect 53559 1756 53629 1802
rect 53675 1756 53745 1802
rect 53791 1756 53861 1802
rect 53907 1756 53977 1802
rect 54023 1756 54093 1802
rect 54139 1756 54209 1802
rect 54255 1756 54325 1802
rect 54371 1756 54441 1802
rect 54487 1756 54557 1802
rect 54603 1756 54673 1802
rect 54719 1756 54789 1802
rect 54835 1756 54905 1802
rect 54951 1756 55021 1802
rect 55067 1756 55137 1802
rect 55183 1756 55253 1802
rect 55299 1756 55369 1802
rect 55415 1756 55485 1802
rect 55531 1756 55601 1802
rect 55647 1756 55717 1802
rect 55763 1756 55833 1802
rect 55879 1756 55949 1802
rect 55995 1756 56065 1802
rect 56111 1756 56181 1802
rect 56227 1756 56297 1802
rect 56343 1756 56413 1802
rect 56459 1756 56529 1802
rect 56575 1756 56594 1802
rect 50826 1686 56594 1756
rect 50826 1640 50845 1686
rect 50891 1640 50961 1686
rect 51007 1640 51077 1686
rect 51123 1640 51193 1686
rect 51239 1640 51309 1686
rect 51355 1640 51425 1686
rect 51471 1640 51541 1686
rect 51587 1640 51657 1686
rect 51703 1640 51773 1686
rect 51819 1640 51889 1686
rect 51935 1640 52005 1686
rect 52051 1640 52121 1686
rect 52167 1640 52237 1686
rect 52283 1640 52353 1686
rect 52399 1640 52469 1686
rect 52515 1640 52585 1686
rect 52631 1640 52701 1686
rect 52747 1640 52817 1686
rect 52863 1640 52933 1686
rect 52979 1640 53049 1686
rect 53095 1640 53165 1686
rect 53211 1640 53281 1686
rect 53327 1640 53397 1686
rect 53443 1640 53513 1686
rect 53559 1640 53629 1686
rect 53675 1640 53745 1686
rect 53791 1640 53861 1686
rect 53907 1640 53977 1686
rect 54023 1640 54093 1686
rect 54139 1640 54209 1686
rect 54255 1640 54325 1686
rect 54371 1640 54441 1686
rect 54487 1640 54557 1686
rect 54603 1640 54673 1686
rect 54719 1640 54789 1686
rect 54835 1640 54905 1686
rect 54951 1640 55021 1686
rect 55067 1640 55137 1686
rect 55183 1640 55253 1686
rect 55299 1640 55369 1686
rect 55415 1640 55485 1686
rect 55531 1640 55601 1686
rect 55647 1640 55717 1686
rect 55763 1640 55833 1686
rect 55879 1640 55949 1686
rect 55995 1640 56065 1686
rect 56111 1640 56181 1686
rect 56227 1640 56297 1686
rect 56343 1640 56413 1686
rect 56459 1640 56529 1686
rect 56575 1640 56594 1686
rect 50826 1570 56594 1640
rect 50826 1524 50845 1570
rect 50891 1524 50961 1570
rect 51007 1524 51077 1570
rect 51123 1524 51193 1570
rect 51239 1524 51309 1570
rect 51355 1524 51425 1570
rect 51471 1524 51541 1570
rect 51587 1524 51657 1570
rect 51703 1524 51773 1570
rect 51819 1524 51889 1570
rect 51935 1524 52005 1570
rect 52051 1524 52121 1570
rect 52167 1524 52237 1570
rect 52283 1524 52353 1570
rect 52399 1524 52469 1570
rect 52515 1524 52585 1570
rect 52631 1524 52701 1570
rect 52747 1524 52817 1570
rect 52863 1524 52933 1570
rect 52979 1524 53049 1570
rect 53095 1524 53165 1570
rect 53211 1524 53281 1570
rect 53327 1524 53397 1570
rect 53443 1524 53513 1570
rect 53559 1524 53629 1570
rect 53675 1524 53745 1570
rect 53791 1524 53861 1570
rect 53907 1524 53977 1570
rect 54023 1524 54093 1570
rect 54139 1524 54209 1570
rect 54255 1524 54325 1570
rect 54371 1524 54441 1570
rect 54487 1524 54557 1570
rect 54603 1524 54673 1570
rect 54719 1524 54789 1570
rect 54835 1524 54905 1570
rect 54951 1524 55021 1570
rect 55067 1524 55137 1570
rect 55183 1524 55253 1570
rect 55299 1524 55369 1570
rect 55415 1524 55485 1570
rect 55531 1524 55601 1570
rect 55647 1524 55717 1570
rect 55763 1524 55833 1570
rect 55879 1524 55949 1570
rect 55995 1524 56065 1570
rect 56111 1524 56181 1570
rect 56227 1524 56297 1570
rect 56343 1524 56413 1570
rect 56459 1524 56529 1570
rect 56575 1524 56594 1570
rect 50826 1454 56594 1524
rect 50826 1408 50845 1454
rect 50891 1408 50961 1454
rect 51007 1408 51077 1454
rect 51123 1408 51193 1454
rect 51239 1408 51309 1454
rect 51355 1408 51425 1454
rect 51471 1408 51541 1454
rect 51587 1408 51657 1454
rect 51703 1408 51773 1454
rect 51819 1408 51889 1454
rect 51935 1408 52005 1454
rect 52051 1408 52121 1454
rect 52167 1408 52237 1454
rect 52283 1408 52353 1454
rect 52399 1408 52469 1454
rect 52515 1408 52585 1454
rect 52631 1408 52701 1454
rect 52747 1408 52817 1454
rect 52863 1408 52933 1454
rect 52979 1408 53049 1454
rect 53095 1408 53165 1454
rect 53211 1408 53281 1454
rect 53327 1408 53397 1454
rect 53443 1408 53513 1454
rect 53559 1408 53629 1454
rect 53675 1408 53745 1454
rect 53791 1408 53861 1454
rect 53907 1408 53977 1454
rect 54023 1408 54093 1454
rect 54139 1408 54209 1454
rect 54255 1408 54325 1454
rect 54371 1408 54441 1454
rect 54487 1408 54557 1454
rect 54603 1408 54673 1454
rect 54719 1408 54789 1454
rect 54835 1408 54905 1454
rect 54951 1408 55021 1454
rect 55067 1408 55137 1454
rect 55183 1408 55253 1454
rect 55299 1408 55369 1454
rect 55415 1408 55485 1454
rect 55531 1408 55601 1454
rect 55647 1408 55717 1454
rect 55763 1408 55833 1454
rect 55879 1408 55949 1454
rect 55995 1408 56065 1454
rect 56111 1408 56181 1454
rect 56227 1408 56297 1454
rect 56343 1408 56413 1454
rect 56459 1408 56529 1454
rect 56575 1408 56594 1454
rect 50826 1338 56594 1408
rect 50826 1292 50845 1338
rect 50891 1292 50961 1338
rect 51007 1292 51077 1338
rect 51123 1292 51193 1338
rect 51239 1292 51309 1338
rect 51355 1292 51425 1338
rect 51471 1292 51541 1338
rect 51587 1292 51657 1338
rect 51703 1292 51773 1338
rect 51819 1292 51889 1338
rect 51935 1292 52005 1338
rect 52051 1292 52121 1338
rect 52167 1292 52237 1338
rect 52283 1292 52353 1338
rect 52399 1292 52469 1338
rect 52515 1292 52585 1338
rect 52631 1292 52701 1338
rect 52747 1292 52817 1338
rect 52863 1292 52933 1338
rect 52979 1292 53049 1338
rect 53095 1292 53165 1338
rect 53211 1292 53281 1338
rect 53327 1292 53397 1338
rect 53443 1292 53513 1338
rect 53559 1292 53629 1338
rect 53675 1292 53745 1338
rect 53791 1292 53861 1338
rect 53907 1292 53977 1338
rect 54023 1292 54093 1338
rect 54139 1292 54209 1338
rect 54255 1292 54325 1338
rect 54371 1292 54441 1338
rect 54487 1292 54557 1338
rect 54603 1292 54673 1338
rect 54719 1292 54789 1338
rect 54835 1292 54905 1338
rect 54951 1292 55021 1338
rect 55067 1292 55137 1338
rect 55183 1292 55253 1338
rect 55299 1292 55369 1338
rect 55415 1292 55485 1338
rect 55531 1292 55601 1338
rect 55647 1292 55717 1338
rect 55763 1292 55833 1338
rect 55879 1292 55949 1338
rect 55995 1292 56065 1338
rect 56111 1292 56181 1338
rect 56227 1292 56297 1338
rect 56343 1292 56413 1338
rect 56459 1292 56529 1338
rect 56575 1292 56594 1338
rect 50826 1222 56594 1292
rect 50826 1176 50845 1222
rect 50891 1176 50961 1222
rect 51007 1176 51077 1222
rect 51123 1176 51193 1222
rect 51239 1176 51309 1222
rect 51355 1176 51425 1222
rect 51471 1176 51541 1222
rect 51587 1176 51657 1222
rect 51703 1176 51773 1222
rect 51819 1176 51889 1222
rect 51935 1176 52005 1222
rect 52051 1176 52121 1222
rect 52167 1176 52237 1222
rect 52283 1176 52353 1222
rect 52399 1176 52469 1222
rect 52515 1176 52585 1222
rect 52631 1176 52701 1222
rect 52747 1176 52817 1222
rect 52863 1176 52933 1222
rect 52979 1176 53049 1222
rect 53095 1176 53165 1222
rect 53211 1176 53281 1222
rect 53327 1176 53397 1222
rect 53443 1176 53513 1222
rect 53559 1176 53629 1222
rect 53675 1176 53745 1222
rect 53791 1176 53861 1222
rect 53907 1176 53977 1222
rect 54023 1176 54093 1222
rect 54139 1176 54209 1222
rect 54255 1176 54325 1222
rect 54371 1176 54441 1222
rect 54487 1176 54557 1222
rect 54603 1176 54673 1222
rect 54719 1176 54789 1222
rect 54835 1176 54905 1222
rect 54951 1176 55021 1222
rect 55067 1176 55137 1222
rect 55183 1176 55253 1222
rect 55299 1176 55369 1222
rect 55415 1176 55485 1222
rect 55531 1176 55601 1222
rect 55647 1176 55717 1222
rect 55763 1176 55833 1222
rect 55879 1176 55949 1222
rect 55995 1176 56065 1222
rect 56111 1176 56181 1222
rect 56227 1176 56297 1222
rect 56343 1176 56413 1222
rect 56459 1176 56529 1222
rect 56575 1176 56594 1222
rect 50826 1034 56594 1176
rect 57361 1117 57380 34237
rect 57626 1117 57645 45463
rect 57361 1034 57645 1117
rect 85714 45563 86098 45646
rect 85714 1117 85733 45563
rect 86079 1117 86098 45563
rect 85714 1034 86098 1117
rect 352 1015 86098 1034
rect 352 969 371 1015
rect 417 969 495 1015
rect 541 969 619 1015
rect 665 969 743 1015
rect 789 969 867 1015
rect 913 969 991 1015
rect 1037 969 1115 1015
rect 1161 969 1239 1015
rect 1285 969 1363 1015
rect 1409 969 1487 1015
rect 1533 969 1611 1015
rect 1657 969 1735 1015
rect 1781 969 1859 1015
rect 1905 969 1983 1015
rect 2029 969 2107 1015
rect 2153 969 2231 1015
rect 2277 969 2355 1015
rect 2401 969 2479 1015
rect 2525 969 2603 1015
rect 2649 969 2727 1015
rect 2773 969 2851 1015
rect 2897 969 2975 1015
rect 3021 969 3099 1015
rect 3145 969 3223 1015
rect 3269 969 3347 1015
rect 3393 969 3471 1015
rect 3517 969 3595 1015
rect 3641 969 3719 1015
rect 3765 969 3843 1015
rect 3889 969 3967 1015
rect 4013 969 4091 1015
rect 4137 969 4215 1015
rect 4261 969 4339 1015
rect 4385 969 4463 1015
rect 4509 969 4587 1015
rect 4633 969 4711 1015
rect 4757 969 4835 1015
rect 4881 969 4959 1015
rect 5005 969 5083 1015
rect 5129 969 5207 1015
rect 5253 969 5331 1015
rect 5377 969 5455 1015
rect 5501 969 5579 1015
rect 5625 969 5703 1015
rect 5749 969 5827 1015
rect 5873 969 5951 1015
rect 5997 969 6075 1015
rect 6121 969 6199 1015
rect 6245 969 6323 1015
rect 6369 969 6447 1015
rect 6493 969 6571 1015
rect 6617 969 6695 1015
rect 6741 969 6819 1015
rect 6865 969 6943 1015
rect 6989 969 7067 1015
rect 7113 969 7191 1015
rect 7237 969 7315 1015
rect 7361 969 7439 1015
rect 7485 969 7563 1015
rect 7609 969 7687 1015
rect 7733 969 7811 1015
rect 7857 969 7935 1015
rect 7981 969 8059 1015
rect 8105 969 8183 1015
rect 8229 969 8307 1015
rect 8353 969 8431 1015
rect 8477 969 8555 1015
rect 8601 969 8679 1015
rect 8725 969 8803 1015
rect 8849 969 8927 1015
rect 8973 969 9051 1015
rect 9097 969 9175 1015
rect 9221 969 9299 1015
rect 9345 969 9423 1015
rect 9469 969 9547 1015
rect 9593 969 9671 1015
rect 9717 969 9795 1015
rect 9841 969 9919 1015
rect 9965 969 10043 1015
rect 10089 969 10167 1015
rect 10213 969 10291 1015
rect 10337 969 10415 1015
rect 10461 969 10539 1015
rect 10585 969 10663 1015
rect 10709 969 10787 1015
rect 10833 969 10911 1015
rect 10957 969 11035 1015
rect 11081 969 11159 1015
rect 11205 969 11283 1015
rect 11329 969 11407 1015
rect 11453 969 11531 1015
rect 11577 969 11655 1015
rect 11701 969 11779 1015
rect 11825 969 11903 1015
rect 11949 969 12027 1015
rect 12073 969 12151 1015
rect 12197 969 12275 1015
rect 12321 969 12399 1015
rect 12445 969 12523 1015
rect 12569 969 12647 1015
rect 12693 969 12771 1015
rect 12817 969 12895 1015
rect 12941 969 13019 1015
rect 13065 969 13143 1015
rect 13189 969 13267 1015
rect 13313 969 13391 1015
rect 13437 969 13515 1015
rect 13561 969 13639 1015
rect 13685 969 13763 1015
rect 13809 969 13887 1015
rect 13933 969 14011 1015
rect 14057 969 14135 1015
rect 14181 969 14259 1015
rect 14305 969 14383 1015
rect 14429 969 14507 1015
rect 14553 969 14631 1015
rect 14677 969 14755 1015
rect 14801 969 14879 1015
rect 14925 969 15003 1015
rect 15049 969 15127 1015
rect 15173 969 15251 1015
rect 15297 969 15375 1015
rect 15421 969 15499 1015
rect 15545 969 15623 1015
rect 15669 969 15747 1015
rect 15793 969 15871 1015
rect 15917 969 15995 1015
rect 16041 969 16119 1015
rect 16165 969 16243 1015
rect 16289 969 16367 1015
rect 16413 969 16491 1015
rect 16537 969 16615 1015
rect 16661 969 16739 1015
rect 16785 969 16863 1015
rect 16909 969 16987 1015
rect 17033 969 17111 1015
rect 17157 969 17235 1015
rect 17281 969 17359 1015
rect 17405 969 17483 1015
rect 17529 969 17607 1015
rect 17653 969 17731 1015
rect 17777 969 17855 1015
rect 17901 969 17979 1015
rect 18025 969 18103 1015
rect 18149 969 18227 1015
rect 18273 969 18351 1015
rect 18397 969 18475 1015
rect 18521 969 18599 1015
rect 18645 969 18723 1015
rect 18769 969 18847 1015
rect 18893 969 18971 1015
rect 19017 969 19095 1015
rect 19141 969 19219 1015
rect 19265 969 19343 1015
rect 19389 969 19467 1015
rect 19513 969 19591 1015
rect 19637 969 19715 1015
rect 19761 969 19839 1015
rect 19885 969 19963 1015
rect 20009 969 20087 1015
rect 20133 969 20211 1015
rect 20257 969 20335 1015
rect 20381 969 20459 1015
rect 20505 969 20583 1015
rect 20629 969 20707 1015
rect 20753 969 20831 1015
rect 20877 969 20955 1015
rect 21001 969 21079 1015
rect 21125 969 21203 1015
rect 21249 969 21327 1015
rect 21373 969 21451 1015
rect 21497 969 21575 1015
rect 21621 969 21699 1015
rect 21745 969 21823 1015
rect 21869 969 21947 1015
rect 21993 969 22071 1015
rect 22117 969 22195 1015
rect 22241 969 22319 1015
rect 22365 969 22443 1015
rect 22489 969 22567 1015
rect 22613 969 22691 1015
rect 22737 969 22815 1015
rect 22861 969 22939 1015
rect 22985 969 23063 1015
rect 23109 969 23187 1015
rect 23233 969 23311 1015
rect 23357 969 23435 1015
rect 23481 969 23559 1015
rect 23605 969 23683 1015
rect 23729 969 23807 1015
rect 23853 969 23931 1015
rect 23977 969 24055 1015
rect 24101 969 24179 1015
rect 24225 969 24303 1015
rect 24349 969 24427 1015
rect 24473 969 24551 1015
rect 24597 969 24675 1015
rect 24721 969 24799 1015
rect 24845 969 24923 1015
rect 24969 969 25047 1015
rect 25093 969 25171 1015
rect 25217 969 25295 1015
rect 25341 969 25419 1015
rect 25465 969 25543 1015
rect 25589 969 25667 1015
rect 25713 969 25791 1015
rect 25837 969 25915 1015
rect 25961 969 26039 1015
rect 26085 969 26163 1015
rect 26209 969 26287 1015
rect 26333 969 26411 1015
rect 26457 969 26535 1015
rect 26581 969 26659 1015
rect 26705 969 26783 1015
rect 26829 969 26907 1015
rect 26953 969 27031 1015
rect 27077 969 27155 1015
rect 27201 969 27279 1015
rect 27325 969 27403 1015
rect 27449 969 27527 1015
rect 27573 969 27651 1015
rect 27697 969 27775 1015
rect 27821 969 27899 1015
rect 27945 969 28023 1015
rect 28069 969 28147 1015
rect 28193 969 28271 1015
rect 28317 969 28395 1015
rect 28441 969 28519 1015
rect 28565 969 28643 1015
rect 28689 969 28767 1015
rect 28813 969 28891 1015
rect 28937 969 29015 1015
rect 29061 969 29139 1015
rect 29185 969 29263 1015
rect 29309 969 29387 1015
rect 29433 969 29511 1015
rect 29557 969 29635 1015
rect 29681 969 29759 1015
rect 29805 969 29883 1015
rect 29929 969 30007 1015
rect 30053 969 30131 1015
rect 30177 969 30255 1015
rect 30301 969 30379 1015
rect 30425 969 30503 1015
rect 30549 969 30627 1015
rect 30673 969 30751 1015
rect 30797 969 30875 1015
rect 30921 969 30999 1015
rect 31045 969 31123 1015
rect 31169 969 31247 1015
rect 31293 969 31371 1015
rect 31417 969 31495 1015
rect 31541 969 31619 1015
rect 31665 969 31743 1015
rect 31789 969 31867 1015
rect 31913 969 31991 1015
rect 32037 969 32115 1015
rect 32161 969 32239 1015
rect 32285 969 32363 1015
rect 32409 969 32487 1015
rect 32533 969 32611 1015
rect 32657 969 32735 1015
rect 32781 969 32859 1015
rect 32905 969 32983 1015
rect 33029 969 33107 1015
rect 33153 969 33231 1015
rect 33277 969 33355 1015
rect 33401 969 33479 1015
rect 33525 969 33603 1015
rect 33649 969 33727 1015
rect 33773 969 33851 1015
rect 33897 969 33975 1015
rect 34021 969 34099 1015
rect 34145 969 34223 1015
rect 34269 969 34347 1015
rect 34393 969 34471 1015
rect 34517 969 34595 1015
rect 34641 969 34719 1015
rect 34765 969 34843 1015
rect 34889 969 34967 1015
rect 35013 969 35091 1015
rect 35137 969 35215 1015
rect 35261 969 35339 1015
rect 35385 969 35463 1015
rect 35509 969 35587 1015
rect 35633 969 35711 1015
rect 35757 969 35835 1015
rect 35881 969 35959 1015
rect 36005 969 36083 1015
rect 36129 969 36207 1015
rect 36253 969 36331 1015
rect 36377 969 36455 1015
rect 36501 969 36579 1015
rect 36625 969 36703 1015
rect 36749 969 36827 1015
rect 36873 969 36951 1015
rect 36997 969 37075 1015
rect 37121 969 37199 1015
rect 37245 969 37323 1015
rect 37369 969 37447 1015
rect 37493 969 37571 1015
rect 37617 969 37695 1015
rect 37741 969 37819 1015
rect 37865 969 37943 1015
rect 37989 969 38067 1015
rect 38113 969 38191 1015
rect 38237 969 38315 1015
rect 38361 969 38439 1015
rect 38485 969 38563 1015
rect 38609 969 38687 1015
rect 38733 969 38811 1015
rect 38857 969 38935 1015
rect 38981 969 39059 1015
rect 39105 969 39183 1015
rect 39229 969 39307 1015
rect 39353 969 39431 1015
rect 39477 969 39555 1015
rect 39601 969 39679 1015
rect 39725 969 39803 1015
rect 39849 969 39927 1015
rect 39973 969 40051 1015
rect 40097 969 40175 1015
rect 40221 969 40299 1015
rect 40345 969 40423 1015
rect 40469 969 40547 1015
rect 40593 969 40671 1015
rect 40717 969 40795 1015
rect 40841 969 40919 1015
rect 40965 969 41043 1015
rect 41089 969 41167 1015
rect 41213 969 41291 1015
rect 41337 969 41415 1015
rect 41461 969 41539 1015
rect 41585 969 41663 1015
rect 41709 969 41787 1015
rect 41833 969 41911 1015
rect 41957 969 42035 1015
rect 42081 969 42159 1015
rect 42205 969 42283 1015
rect 42329 969 42407 1015
rect 42453 969 42531 1015
rect 42577 969 42655 1015
rect 42701 969 42779 1015
rect 42825 969 42903 1015
rect 42949 969 43027 1015
rect 43073 969 43151 1015
rect 43197 969 43275 1015
rect 43321 969 43399 1015
rect 43445 969 43523 1015
rect 43569 969 43647 1015
rect 43693 969 43771 1015
rect 43817 969 43895 1015
rect 43941 969 44019 1015
rect 44065 969 44143 1015
rect 44189 969 44267 1015
rect 44313 969 44391 1015
rect 44437 969 44515 1015
rect 44561 969 44639 1015
rect 44685 969 44763 1015
rect 44809 969 44887 1015
rect 44933 969 45011 1015
rect 45057 969 45135 1015
rect 45181 969 45259 1015
rect 45305 969 45383 1015
rect 45429 969 45507 1015
rect 45553 969 45631 1015
rect 45677 969 45755 1015
rect 45801 969 45879 1015
rect 45925 969 46003 1015
rect 46049 969 46127 1015
rect 46173 969 46251 1015
rect 46297 969 46375 1015
rect 46421 969 46499 1015
rect 46545 969 46623 1015
rect 46669 969 46747 1015
rect 46793 969 46871 1015
rect 46917 969 46995 1015
rect 47041 969 47119 1015
rect 47165 969 47243 1015
rect 47289 969 47367 1015
rect 47413 969 47491 1015
rect 47537 969 47615 1015
rect 47661 969 47739 1015
rect 47785 969 47863 1015
rect 47909 969 47987 1015
rect 48033 969 48111 1015
rect 48157 969 48235 1015
rect 48281 969 48359 1015
rect 48405 969 48483 1015
rect 48529 969 48607 1015
rect 48653 969 48731 1015
rect 48777 969 48855 1015
rect 48901 969 48979 1015
rect 49025 969 49103 1015
rect 49149 969 49227 1015
rect 49273 969 49351 1015
rect 49397 969 49475 1015
rect 49521 969 49599 1015
rect 49645 969 49723 1015
rect 49769 969 49847 1015
rect 49893 969 49971 1015
rect 50017 969 50095 1015
rect 50141 969 50219 1015
rect 50265 969 50343 1015
rect 50389 969 50467 1015
rect 50513 969 50591 1015
rect 50637 969 50715 1015
rect 50761 969 50839 1015
rect 50885 969 50963 1015
rect 51009 969 51087 1015
rect 51133 969 51211 1015
rect 51257 969 51335 1015
rect 51381 969 51459 1015
rect 51505 969 51583 1015
rect 51629 969 51707 1015
rect 51753 969 51831 1015
rect 51877 969 51955 1015
rect 52001 969 52079 1015
rect 52125 969 52203 1015
rect 52249 969 52327 1015
rect 52373 969 52451 1015
rect 52497 969 52575 1015
rect 52621 969 52699 1015
rect 52745 969 52823 1015
rect 52869 969 52947 1015
rect 52993 969 53071 1015
rect 53117 969 53195 1015
rect 53241 969 53319 1015
rect 53365 969 53443 1015
rect 53489 969 53567 1015
rect 53613 969 53691 1015
rect 53737 969 53815 1015
rect 53861 969 53939 1015
rect 53985 969 54063 1015
rect 54109 969 54187 1015
rect 54233 969 54311 1015
rect 54357 969 54435 1015
rect 54481 969 54559 1015
rect 54605 969 54683 1015
rect 54729 969 54807 1015
rect 54853 969 54931 1015
rect 54977 969 55055 1015
rect 55101 969 55179 1015
rect 55225 969 55303 1015
rect 55349 969 55427 1015
rect 55473 969 55551 1015
rect 55597 969 55675 1015
rect 55721 969 55799 1015
rect 55845 969 55923 1015
rect 55969 969 56047 1015
rect 56093 969 56171 1015
rect 56217 969 56295 1015
rect 56341 969 56419 1015
rect 56465 969 56543 1015
rect 56589 969 56667 1015
rect 56713 969 56791 1015
rect 56837 969 56915 1015
rect 56961 969 57039 1015
rect 57085 969 57163 1015
rect 57209 969 57287 1015
rect 57333 969 57411 1015
rect 57457 969 57535 1015
rect 57581 969 57659 1015
rect 57705 969 57783 1015
rect 57829 969 57907 1015
rect 57953 969 58031 1015
rect 58077 969 58155 1015
rect 58201 969 58279 1015
rect 58325 969 58403 1015
rect 58449 969 58527 1015
rect 58573 969 58651 1015
rect 58697 969 58775 1015
rect 58821 969 58899 1015
rect 58945 969 59023 1015
rect 59069 969 59147 1015
rect 59193 969 59271 1015
rect 59317 969 59395 1015
rect 59441 969 59519 1015
rect 59565 969 59643 1015
rect 59689 969 59767 1015
rect 59813 969 59891 1015
rect 59937 969 60015 1015
rect 60061 969 60139 1015
rect 60185 969 60263 1015
rect 60309 969 60387 1015
rect 60433 969 60511 1015
rect 60557 969 60635 1015
rect 60681 969 60759 1015
rect 60805 969 60883 1015
rect 60929 969 61007 1015
rect 61053 969 61131 1015
rect 61177 969 61255 1015
rect 61301 969 61379 1015
rect 61425 969 61503 1015
rect 61549 969 61627 1015
rect 61673 969 61751 1015
rect 61797 969 61875 1015
rect 61921 969 61999 1015
rect 62045 969 62123 1015
rect 62169 969 62247 1015
rect 62293 969 62371 1015
rect 62417 969 62495 1015
rect 62541 969 62619 1015
rect 62665 969 62743 1015
rect 62789 969 62867 1015
rect 62913 969 62991 1015
rect 63037 969 63115 1015
rect 63161 969 63239 1015
rect 63285 969 63363 1015
rect 63409 969 63487 1015
rect 63533 969 63611 1015
rect 63657 969 63735 1015
rect 63781 969 63859 1015
rect 63905 969 63983 1015
rect 64029 969 64107 1015
rect 64153 969 64231 1015
rect 64277 969 64355 1015
rect 64401 969 64479 1015
rect 64525 969 64603 1015
rect 64649 969 64727 1015
rect 64773 969 64851 1015
rect 64897 969 64975 1015
rect 65021 969 65099 1015
rect 65145 969 65223 1015
rect 65269 969 65347 1015
rect 65393 969 65471 1015
rect 65517 969 65595 1015
rect 65641 969 65719 1015
rect 65765 969 65843 1015
rect 65889 969 65967 1015
rect 66013 969 66091 1015
rect 66137 969 66215 1015
rect 66261 969 66339 1015
rect 66385 969 66463 1015
rect 66509 969 66587 1015
rect 66633 969 66711 1015
rect 66757 969 66835 1015
rect 66881 969 66959 1015
rect 67005 969 67083 1015
rect 67129 969 67207 1015
rect 67253 969 67331 1015
rect 67377 969 67455 1015
rect 67501 969 67579 1015
rect 67625 969 67703 1015
rect 67749 969 67827 1015
rect 67873 969 67951 1015
rect 67997 969 68075 1015
rect 68121 969 68199 1015
rect 68245 969 68323 1015
rect 68369 969 68447 1015
rect 68493 969 68571 1015
rect 68617 969 68695 1015
rect 68741 969 68819 1015
rect 68865 969 68943 1015
rect 68989 969 69067 1015
rect 69113 969 69191 1015
rect 69237 969 69315 1015
rect 69361 969 69439 1015
rect 69485 969 69563 1015
rect 69609 969 69687 1015
rect 69733 969 69811 1015
rect 69857 969 69935 1015
rect 69981 969 70059 1015
rect 70105 969 70183 1015
rect 70229 969 70307 1015
rect 70353 969 70431 1015
rect 70477 969 70555 1015
rect 70601 969 70679 1015
rect 70725 969 70803 1015
rect 70849 969 70927 1015
rect 70973 969 71051 1015
rect 71097 969 71175 1015
rect 71221 969 71299 1015
rect 71345 969 71423 1015
rect 71469 969 71547 1015
rect 71593 969 71671 1015
rect 71717 969 71795 1015
rect 71841 969 71919 1015
rect 71965 969 72043 1015
rect 72089 969 72167 1015
rect 72213 969 72291 1015
rect 72337 969 72415 1015
rect 72461 969 72539 1015
rect 72585 969 72663 1015
rect 72709 969 72787 1015
rect 72833 969 72911 1015
rect 72957 969 73035 1015
rect 73081 969 73159 1015
rect 73205 969 73283 1015
rect 73329 969 73407 1015
rect 73453 969 73531 1015
rect 73577 969 73655 1015
rect 73701 969 73779 1015
rect 73825 969 73903 1015
rect 73949 969 74027 1015
rect 74073 969 74151 1015
rect 74197 969 74275 1015
rect 74321 969 74399 1015
rect 74445 969 74523 1015
rect 74569 969 74647 1015
rect 74693 969 74771 1015
rect 74817 969 74895 1015
rect 74941 969 75019 1015
rect 75065 969 75143 1015
rect 75189 969 75267 1015
rect 75313 969 75391 1015
rect 75437 969 75515 1015
rect 75561 969 75639 1015
rect 75685 969 75763 1015
rect 75809 969 75887 1015
rect 75933 969 76011 1015
rect 76057 969 76135 1015
rect 76181 969 76259 1015
rect 76305 969 76383 1015
rect 76429 969 76507 1015
rect 76553 969 76631 1015
rect 76677 969 76755 1015
rect 76801 969 76879 1015
rect 76925 969 77003 1015
rect 77049 969 77127 1015
rect 77173 969 77251 1015
rect 77297 969 77375 1015
rect 77421 969 77499 1015
rect 77545 969 77623 1015
rect 77669 969 77747 1015
rect 77793 969 77871 1015
rect 77917 969 77995 1015
rect 78041 969 78119 1015
rect 78165 969 78243 1015
rect 78289 969 78367 1015
rect 78413 969 78491 1015
rect 78537 969 78615 1015
rect 78661 969 78739 1015
rect 78785 969 78863 1015
rect 78909 969 78987 1015
rect 79033 969 79111 1015
rect 79157 969 79235 1015
rect 79281 969 79359 1015
rect 79405 969 79483 1015
rect 79529 969 79607 1015
rect 79653 969 79731 1015
rect 79777 969 79855 1015
rect 79901 969 79979 1015
rect 80025 969 80103 1015
rect 80149 969 80227 1015
rect 80273 969 80351 1015
rect 80397 969 80475 1015
rect 80521 969 80599 1015
rect 80645 969 80723 1015
rect 80769 969 80847 1015
rect 80893 969 80971 1015
rect 81017 969 81095 1015
rect 81141 969 81219 1015
rect 81265 969 81343 1015
rect 81389 969 81467 1015
rect 81513 969 81591 1015
rect 81637 969 81715 1015
rect 81761 969 81839 1015
rect 81885 969 81963 1015
rect 82009 969 82087 1015
rect 82133 969 82211 1015
rect 82257 969 82335 1015
rect 82381 969 82459 1015
rect 82505 969 82583 1015
rect 82629 969 82707 1015
rect 82753 969 82831 1015
rect 82877 969 82955 1015
rect 83001 969 83079 1015
rect 83125 969 83203 1015
rect 83249 969 83327 1015
rect 83373 969 83451 1015
rect 83497 969 83575 1015
rect 83621 969 83699 1015
rect 83745 969 83823 1015
rect 83869 969 83947 1015
rect 83993 969 84071 1015
rect 84117 969 84195 1015
rect 84241 969 84319 1015
rect 84365 969 84443 1015
rect 84489 969 84567 1015
rect 84613 969 84691 1015
rect 84737 969 84815 1015
rect 84861 969 84939 1015
rect 84985 969 85063 1015
rect 85109 969 85187 1015
rect 85233 969 85311 1015
rect 85357 969 85435 1015
rect 85481 969 85559 1015
rect 85605 969 85683 1015
rect 85729 969 85807 1015
rect 85853 969 85931 1015
rect 85977 969 86098 1015
rect 352 891 86098 969
rect 352 845 371 891
rect 417 845 495 891
rect 541 845 619 891
rect 665 845 743 891
rect 789 845 867 891
rect 913 845 991 891
rect 1037 845 1115 891
rect 1161 845 1239 891
rect 1285 845 1363 891
rect 1409 845 1487 891
rect 1533 845 1611 891
rect 1657 845 1735 891
rect 1781 845 1859 891
rect 1905 845 1983 891
rect 2029 845 2107 891
rect 2153 845 2231 891
rect 2277 845 2355 891
rect 2401 845 2479 891
rect 2525 845 2603 891
rect 2649 845 2727 891
rect 2773 845 2851 891
rect 2897 845 2975 891
rect 3021 845 3099 891
rect 3145 845 3223 891
rect 3269 845 3347 891
rect 3393 845 3471 891
rect 3517 845 3595 891
rect 3641 845 3719 891
rect 3765 845 3843 891
rect 3889 845 3967 891
rect 4013 845 4091 891
rect 4137 845 4215 891
rect 4261 845 4339 891
rect 4385 845 4463 891
rect 4509 845 4587 891
rect 4633 845 4711 891
rect 4757 845 4835 891
rect 4881 845 4959 891
rect 5005 845 5083 891
rect 5129 845 5207 891
rect 5253 845 5331 891
rect 5377 845 5455 891
rect 5501 845 5579 891
rect 5625 845 5703 891
rect 5749 845 5827 891
rect 5873 845 5951 891
rect 5997 845 6075 891
rect 6121 845 6199 891
rect 6245 845 6323 891
rect 6369 845 6447 891
rect 6493 845 6571 891
rect 6617 845 6695 891
rect 6741 845 6819 891
rect 6865 845 6943 891
rect 6989 845 7067 891
rect 7113 845 7191 891
rect 7237 845 7315 891
rect 7361 845 7439 891
rect 7485 845 7563 891
rect 7609 845 7687 891
rect 7733 845 7811 891
rect 7857 845 7935 891
rect 7981 845 8059 891
rect 8105 845 8183 891
rect 8229 845 8307 891
rect 8353 845 8431 891
rect 8477 845 8555 891
rect 8601 845 8679 891
rect 8725 845 8803 891
rect 8849 845 8927 891
rect 8973 845 9051 891
rect 9097 845 9175 891
rect 9221 845 9299 891
rect 9345 845 9423 891
rect 9469 845 9547 891
rect 9593 845 9671 891
rect 9717 845 9795 891
rect 9841 845 9919 891
rect 9965 845 10043 891
rect 10089 845 10167 891
rect 10213 845 10291 891
rect 10337 845 10415 891
rect 10461 845 10539 891
rect 10585 845 10663 891
rect 10709 845 10787 891
rect 10833 845 10911 891
rect 10957 845 11035 891
rect 11081 845 11159 891
rect 11205 845 11283 891
rect 11329 845 11407 891
rect 11453 845 11531 891
rect 11577 845 11655 891
rect 11701 845 11779 891
rect 11825 845 11903 891
rect 11949 845 12027 891
rect 12073 845 12151 891
rect 12197 845 12275 891
rect 12321 845 12399 891
rect 12445 845 12523 891
rect 12569 845 12647 891
rect 12693 845 12771 891
rect 12817 845 12895 891
rect 12941 845 13019 891
rect 13065 845 13143 891
rect 13189 845 13267 891
rect 13313 845 13391 891
rect 13437 845 13515 891
rect 13561 845 13639 891
rect 13685 845 13763 891
rect 13809 845 13887 891
rect 13933 845 14011 891
rect 14057 845 14135 891
rect 14181 845 14259 891
rect 14305 845 14383 891
rect 14429 845 14507 891
rect 14553 845 14631 891
rect 14677 845 14755 891
rect 14801 845 14879 891
rect 14925 845 15003 891
rect 15049 845 15127 891
rect 15173 845 15251 891
rect 15297 845 15375 891
rect 15421 845 15499 891
rect 15545 845 15623 891
rect 15669 845 15747 891
rect 15793 845 15871 891
rect 15917 845 15995 891
rect 16041 845 16119 891
rect 16165 845 16243 891
rect 16289 845 16367 891
rect 16413 845 16491 891
rect 16537 845 16615 891
rect 16661 845 16739 891
rect 16785 845 16863 891
rect 16909 845 16987 891
rect 17033 845 17111 891
rect 17157 845 17235 891
rect 17281 845 17359 891
rect 17405 845 17483 891
rect 17529 845 17607 891
rect 17653 845 17731 891
rect 17777 845 17855 891
rect 17901 845 17979 891
rect 18025 845 18103 891
rect 18149 845 18227 891
rect 18273 845 18351 891
rect 18397 845 18475 891
rect 18521 845 18599 891
rect 18645 845 18723 891
rect 18769 845 18847 891
rect 18893 845 18971 891
rect 19017 845 19095 891
rect 19141 845 19219 891
rect 19265 845 19343 891
rect 19389 845 19467 891
rect 19513 845 19591 891
rect 19637 845 19715 891
rect 19761 845 19839 891
rect 19885 845 19963 891
rect 20009 845 20087 891
rect 20133 845 20211 891
rect 20257 845 20335 891
rect 20381 845 20459 891
rect 20505 845 20583 891
rect 20629 845 20707 891
rect 20753 845 20831 891
rect 20877 845 20955 891
rect 21001 845 21079 891
rect 21125 845 21203 891
rect 21249 845 21327 891
rect 21373 845 21451 891
rect 21497 845 21575 891
rect 21621 845 21699 891
rect 21745 845 21823 891
rect 21869 845 21947 891
rect 21993 845 22071 891
rect 22117 845 22195 891
rect 22241 845 22319 891
rect 22365 845 22443 891
rect 22489 845 22567 891
rect 22613 845 22691 891
rect 22737 845 22815 891
rect 22861 845 22939 891
rect 22985 845 23063 891
rect 23109 845 23187 891
rect 23233 845 23311 891
rect 23357 845 23435 891
rect 23481 845 23559 891
rect 23605 845 23683 891
rect 23729 845 23807 891
rect 23853 845 23931 891
rect 23977 845 24055 891
rect 24101 845 24179 891
rect 24225 845 24303 891
rect 24349 845 24427 891
rect 24473 845 24551 891
rect 24597 845 24675 891
rect 24721 845 24799 891
rect 24845 845 24923 891
rect 24969 845 25047 891
rect 25093 845 25171 891
rect 25217 845 25295 891
rect 25341 845 25419 891
rect 25465 845 25543 891
rect 25589 845 25667 891
rect 25713 845 25791 891
rect 25837 845 25915 891
rect 25961 845 26039 891
rect 26085 845 26163 891
rect 26209 845 26287 891
rect 26333 845 26411 891
rect 26457 845 26535 891
rect 26581 845 26659 891
rect 26705 845 26783 891
rect 26829 845 26907 891
rect 26953 845 27031 891
rect 27077 845 27155 891
rect 27201 845 27279 891
rect 27325 845 27403 891
rect 27449 845 27527 891
rect 27573 845 27651 891
rect 27697 845 27775 891
rect 27821 845 27899 891
rect 27945 845 28023 891
rect 28069 845 28147 891
rect 28193 845 28271 891
rect 28317 845 28395 891
rect 28441 845 28519 891
rect 28565 845 28643 891
rect 28689 845 28767 891
rect 28813 845 28891 891
rect 28937 845 29015 891
rect 29061 845 29139 891
rect 29185 845 29263 891
rect 29309 845 29387 891
rect 29433 845 29511 891
rect 29557 845 29635 891
rect 29681 845 29759 891
rect 29805 845 29883 891
rect 29929 845 30007 891
rect 30053 845 30131 891
rect 30177 845 30255 891
rect 30301 845 30379 891
rect 30425 845 30503 891
rect 30549 845 30627 891
rect 30673 845 30751 891
rect 30797 845 30875 891
rect 30921 845 30999 891
rect 31045 845 31123 891
rect 31169 845 31247 891
rect 31293 845 31371 891
rect 31417 845 31495 891
rect 31541 845 31619 891
rect 31665 845 31743 891
rect 31789 845 31867 891
rect 31913 845 31991 891
rect 32037 845 32115 891
rect 32161 845 32239 891
rect 32285 845 32363 891
rect 32409 845 32487 891
rect 32533 845 32611 891
rect 32657 845 32735 891
rect 32781 845 32859 891
rect 32905 845 32983 891
rect 33029 845 33107 891
rect 33153 845 33231 891
rect 33277 845 33355 891
rect 33401 845 33479 891
rect 33525 845 33603 891
rect 33649 845 33727 891
rect 33773 845 33851 891
rect 33897 845 33975 891
rect 34021 845 34099 891
rect 34145 845 34223 891
rect 34269 845 34347 891
rect 34393 845 34471 891
rect 34517 845 34595 891
rect 34641 845 34719 891
rect 34765 845 34843 891
rect 34889 845 34967 891
rect 35013 845 35091 891
rect 35137 845 35215 891
rect 35261 845 35339 891
rect 35385 845 35463 891
rect 35509 845 35587 891
rect 35633 845 35711 891
rect 35757 845 35835 891
rect 35881 845 35959 891
rect 36005 845 36083 891
rect 36129 845 36207 891
rect 36253 845 36331 891
rect 36377 845 36455 891
rect 36501 845 36579 891
rect 36625 845 36703 891
rect 36749 845 36827 891
rect 36873 845 36951 891
rect 36997 845 37075 891
rect 37121 845 37199 891
rect 37245 845 37323 891
rect 37369 845 37447 891
rect 37493 845 37571 891
rect 37617 845 37695 891
rect 37741 845 37819 891
rect 37865 845 37943 891
rect 37989 845 38067 891
rect 38113 845 38191 891
rect 38237 845 38315 891
rect 38361 845 38439 891
rect 38485 845 38563 891
rect 38609 845 38687 891
rect 38733 845 38811 891
rect 38857 845 38935 891
rect 38981 845 39059 891
rect 39105 845 39183 891
rect 39229 845 39307 891
rect 39353 845 39431 891
rect 39477 845 39555 891
rect 39601 845 39679 891
rect 39725 845 39803 891
rect 39849 845 39927 891
rect 39973 845 40051 891
rect 40097 845 40175 891
rect 40221 845 40299 891
rect 40345 845 40423 891
rect 40469 845 40547 891
rect 40593 845 40671 891
rect 40717 845 40795 891
rect 40841 845 40919 891
rect 40965 845 41043 891
rect 41089 845 41167 891
rect 41213 845 41291 891
rect 41337 845 41415 891
rect 41461 845 41539 891
rect 41585 845 41663 891
rect 41709 845 41787 891
rect 41833 845 41911 891
rect 41957 845 42035 891
rect 42081 845 42159 891
rect 42205 845 42283 891
rect 42329 845 42407 891
rect 42453 845 42531 891
rect 42577 845 42655 891
rect 42701 845 42779 891
rect 42825 845 42903 891
rect 42949 845 43027 891
rect 43073 845 43151 891
rect 43197 845 43275 891
rect 43321 845 43399 891
rect 43445 845 43523 891
rect 43569 845 43647 891
rect 43693 845 43771 891
rect 43817 845 43895 891
rect 43941 845 44019 891
rect 44065 845 44143 891
rect 44189 845 44267 891
rect 44313 845 44391 891
rect 44437 845 44515 891
rect 44561 845 44639 891
rect 44685 845 44763 891
rect 44809 845 44887 891
rect 44933 845 45011 891
rect 45057 845 45135 891
rect 45181 845 45259 891
rect 45305 845 45383 891
rect 45429 845 45507 891
rect 45553 845 45631 891
rect 45677 845 45755 891
rect 45801 845 45879 891
rect 45925 845 46003 891
rect 46049 845 46127 891
rect 46173 845 46251 891
rect 46297 845 46375 891
rect 46421 845 46499 891
rect 46545 845 46623 891
rect 46669 845 46747 891
rect 46793 845 46871 891
rect 46917 845 46995 891
rect 47041 845 47119 891
rect 47165 845 47243 891
rect 47289 845 47367 891
rect 47413 845 47491 891
rect 47537 845 47615 891
rect 47661 845 47739 891
rect 47785 845 47863 891
rect 47909 845 47987 891
rect 48033 845 48111 891
rect 48157 845 48235 891
rect 48281 845 48359 891
rect 48405 845 48483 891
rect 48529 845 48607 891
rect 48653 845 48731 891
rect 48777 845 48855 891
rect 48901 845 48979 891
rect 49025 845 49103 891
rect 49149 845 49227 891
rect 49273 845 49351 891
rect 49397 845 49475 891
rect 49521 845 49599 891
rect 49645 845 49723 891
rect 49769 845 49847 891
rect 49893 845 49971 891
rect 50017 845 50095 891
rect 50141 845 50219 891
rect 50265 845 50343 891
rect 50389 845 50467 891
rect 50513 845 50591 891
rect 50637 845 50715 891
rect 50761 845 50839 891
rect 50885 845 50963 891
rect 51009 845 51087 891
rect 51133 845 51211 891
rect 51257 845 51335 891
rect 51381 845 51459 891
rect 51505 845 51583 891
rect 51629 845 51707 891
rect 51753 845 51831 891
rect 51877 845 51955 891
rect 52001 845 52079 891
rect 52125 845 52203 891
rect 52249 845 52327 891
rect 52373 845 52451 891
rect 52497 845 52575 891
rect 52621 845 52699 891
rect 52745 845 52823 891
rect 52869 845 52947 891
rect 52993 845 53071 891
rect 53117 845 53195 891
rect 53241 845 53319 891
rect 53365 845 53443 891
rect 53489 845 53567 891
rect 53613 845 53691 891
rect 53737 845 53815 891
rect 53861 845 53939 891
rect 53985 845 54063 891
rect 54109 845 54187 891
rect 54233 845 54311 891
rect 54357 845 54435 891
rect 54481 845 54559 891
rect 54605 845 54683 891
rect 54729 845 54807 891
rect 54853 845 54931 891
rect 54977 845 55055 891
rect 55101 845 55179 891
rect 55225 845 55303 891
rect 55349 845 55427 891
rect 55473 845 55551 891
rect 55597 845 55675 891
rect 55721 845 55799 891
rect 55845 845 55923 891
rect 55969 845 56047 891
rect 56093 845 56171 891
rect 56217 845 56295 891
rect 56341 845 56419 891
rect 56465 845 56543 891
rect 56589 845 56667 891
rect 56713 845 56791 891
rect 56837 845 56915 891
rect 56961 845 57039 891
rect 57085 845 57163 891
rect 57209 845 57287 891
rect 57333 845 57411 891
rect 57457 845 57535 891
rect 57581 845 57659 891
rect 57705 845 57783 891
rect 57829 845 57907 891
rect 57953 845 58031 891
rect 58077 845 58155 891
rect 58201 845 58279 891
rect 58325 845 58403 891
rect 58449 845 58527 891
rect 58573 845 58651 891
rect 58697 845 58775 891
rect 58821 845 58899 891
rect 58945 845 59023 891
rect 59069 845 59147 891
rect 59193 845 59271 891
rect 59317 845 59395 891
rect 59441 845 59519 891
rect 59565 845 59643 891
rect 59689 845 59767 891
rect 59813 845 59891 891
rect 59937 845 60015 891
rect 60061 845 60139 891
rect 60185 845 60263 891
rect 60309 845 60387 891
rect 60433 845 60511 891
rect 60557 845 60635 891
rect 60681 845 60759 891
rect 60805 845 60883 891
rect 60929 845 61007 891
rect 61053 845 61131 891
rect 61177 845 61255 891
rect 61301 845 61379 891
rect 61425 845 61503 891
rect 61549 845 61627 891
rect 61673 845 61751 891
rect 61797 845 61875 891
rect 61921 845 61999 891
rect 62045 845 62123 891
rect 62169 845 62247 891
rect 62293 845 62371 891
rect 62417 845 62495 891
rect 62541 845 62619 891
rect 62665 845 62743 891
rect 62789 845 62867 891
rect 62913 845 62991 891
rect 63037 845 63115 891
rect 63161 845 63239 891
rect 63285 845 63363 891
rect 63409 845 63487 891
rect 63533 845 63611 891
rect 63657 845 63735 891
rect 63781 845 63859 891
rect 63905 845 63983 891
rect 64029 845 64107 891
rect 64153 845 64231 891
rect 64277 845 64355 891
rect 64401 845 64479 891
rect 64525 845 64603 891
rect 64649 845 64727 891
rect 64773 845 64851 891
rect 64897 845 64975 891
rect 65021 845 65099 891
rect 65145 845 65223 891
rect 65269 845 65347 891
rect 65393 845 65471 891
rect 65517 845 65595 891
rect 65641 845 65719 891
rect 65765 845 65843 891
rect 65889 845 65967 891
rect 66013 845 66091 891
rect 66137 845 66215 891
rect 66261 845 66339 891
rect 66385 845 66463 891
rect 66509 845 66587 891
rect 66633 845 66711 891
rect 66757 845 66835 891
rect 66881 845 66959 891
rect 67005 845 67083 891
rect 67129 845 67207 891
rect 67253 845 67331 891
rect 67377 845 67455 891
rect 67501 845 67579 891
rect 67625 845 67703 891
rect 67749 845 67827 891
rect 67873 845 67951 891
rect 67997 845 68075 891
rect 68121 845 68199 891
rect 68245 845 68323 891
rect 68369 845 68447 891
rect 68493 845 68571 891
rect 68617 845 68695 891
rect 68741 845 68819 891
rect 68865 845 68943 891
rect 68989 845 69067 891
rect 69113 845 69191 891
rect 69237 845 69315 891
rect 69361 845 69439 891
rect 69485 845 69563 891
rect 69609 845 69687 891
rect 69733 845 69811 891
rect 69857 845 69935 891
rect 69981 845 70059 891
rect 70105 845 70183 891
rect 70229 845 70307 891
rect 70353 845 70431 891
rect 70477 845 70555 891
rect 70601 845 70679 891
rect 70725 845 70803 891
rect 70849 845 70927 891
rect 70973 845 71051 891
rect 71097 845 71175 891
rect 71221 845 71299 891
rect 71345 845 71423 891
rect 71469 845 71547 891
rect 71593 845 71671 891
rect 71717 845 71795 891
rect 71841 845 71919 891
rect 71965 845 72043 891
rect 72089 845 72167 891
rect 72213 845 72291 891
rect 72337 845 72415 891
rect 72461 845 72539 891
rect 72585 845 72663 891
rect 72709 845 72787 891
rect 72833 845 72911 891
rect 72957 845 73035 891
rect 73081 845 73159 891
rect 73205 845 73283 891
rect 73329 845 73407 891
rect 73453 845 73531 891
rect 73577 845 73655 891
rect 73701 845 73779 891
rect 73825 845 73903 891
rect 73949 845 74027 891
rect 74073 845 74151 891
rect 74197 845 74275 891
rect 74321 845 74399 891
rect 74445 845 74523 891
rect 74569 845 74647 891
rect 74693 845 74771 891
rect 74817 845 74895 891
rect 74941 845 75019 891
rect 75065 845 75143 891
rect 75189 845 75267 891
rect 75313 845 75391 891
rect 75437 845 75515 891
rect 75561 845 75639 891
rect 75685 845 75763 891
rect 75809 845 75887 891
rect 75933 845 76011 891
rect 76057 845 76135 891
rect 76181 845 76259 891
rect 76305 845 76383 891
rect 76429 845 76507 891
rect 76553 845 76631 891
rect 76677 845 76755 891
rect 76801 845 76879 891
rect 76925 845 77003 891
rect 77049 845 77127 891
rect 77173 845 77251 891
rect 77297 845 77375 891
rect 77421 845 77499 891
rect 77545 845 77623 891
rect 77669 845 77747 891
rect 77793 845 77871 891
rect 77917 845 77995 891
rect 78041 845 78119 891
rect 78165 845 78243 891
rect 78289 845 78367 891
rect 78413 845 78491 891
rect 78537 845 78615 891
rect 78661 845 78739 891
rect 78785 845 78863 891
rect 78909 845 78987 891
rect 79033 845 79111 891
rect 79157 845 79235 891
rect 79281 845 79359 891
rect 79405 845 79483 891
rect 79529 845 79607 891
rect 79653 845 79731 891
rect 79777 845 79855 891
rect 79901 845 79979 891
rect 80025 845 80103 891
rect 80149 845 80227 891
rect 80273 845 80351 891
rect 80397 845 80475 891
rect 80521 845 80599 891
rect 80645 845 80723 891
rect 80769 845 80847 891
rect 80893 845 80971 891
rect 81017 845 81095 891
rect 81141 845 81219 891
rect 81265 845 81343 891
rect 81389 845 81467 891
rect 81513 845 81591 891
rect 81637 845 81715 891
rect 81761 845 81839 891
rect 81885 845 81963 891
rect 82009 845 82087 891
rect 82133 845 82211 891
rect 82257 845 82335 891
rect 82381 845 82459 891
rect 82505 845 82583 891
rect 82629 845 82707 891
rect 82753 845 82831 891
rect 82877 845 82955 891
rect 83001 845 83079 891
rect 83125 845 83203 891
rect 83249 845 83327 891
rect 83373 845 83451 891
rect 83497 845 83575 891
rect 83621 845 83699 891
rect 83745 845 83823 891
rect 83869 845 83947 891
rect 83993 845 84071 891
rect 84117 845 84195 891
rect 84241 845 84319 891
rect 84365 845 84443 891
rect 84489 845 84567 891
rect 84613 845 84691 891
rect 84737 845 84815 891
rect 84861 845 84939 891
rect 84985 845 85063 891
rect 85109 845 85187 891
rect 85233 845 85311 891
rect 85357 845 85435 891
rect 85481 845 85559 891
rect 85605 845 85683 891
rect 85729 845 85807 891
rect 85853 845 85931 891
rect 85977 845 86098 891
rect 352 767 86098 845
rect 352 721 371 767
rect 417 721 495 767
rect 541 721 619 767
rect 665 721 743 767
rect 789 721 867 767
rect 913 721 991 767
rect 1037 721 1115 767
rect 1161 721 1239 767
rect 1285 721 1363 767
rect 1409 721 1487 767
rect 1533 721 1611 767
rect 1657 721 1735 767
rect 1781 721 1859 767
rect 1905 721 1983 767
rect 2029 721 2107 767
rect 2153 721 2231 767
rect 2277 721 2355 767
rect 2401 721 2479 767
rect 2525 721 2603 767
rect 2649 721 2727 767
rect 2773 721 2851 767
rect 2897 721 2975 767
rect 3021 721 3099 767
rect 3145 721 3223 767
rect 3269 721 3347 767
rect 3393 721 3471 767
rect 3517 721 3595 767
rect 3641 721 3719 767
rect 3765 721 3843 767
rect 3889 721 3967 767
rect 4013 721 4091 767
rect 4137 721 4215 767
rect 4261 721 4339 767
rect 4385 721 4463 767
rect 4509 721 4587 767
rect 4633 721 4711 767
rect 4757 721 4835 767
rect 4881 721 4959 767
rect 5005 721 5083 767
rect 5129 721 5207 767
rect 5253 721 5331 767
rect 5377 721 5455 767
rect 5501 721 5579 767
rect 5625 721 5703 767
rect 5749 721 5827 767
rect 5873 721 5951 767
rect 5997 721 6075 767
rect 6121 721 6199 767
rect 6245 721 6323 767
rect 6369 721 6447 767
rect 6493 721 6571 767
rect 6617 721 6695 767
rect 6741 721 6819 767
rect 6865 721 6943 767
rect 6989 721 7067 767
rect 7113 721 7191 767
rect 7237 721 7315 767
rect 7361 721 7439 767
rect 7485 721 7563 767
rect 7609 721 7687 767
rect 7733 721 7811 767
rect 7857 721 7935 767
rect 7981 721 8059 767
rect 8105 721 8183 767
rect 8229 721 8307 767
rect 8353 721 8431 767
rect 8477 721 8555 767
rect 8601 721 8679 767
rect 8725 721 8803 767
rect 8849 721 8927 767
rect 8973 721 9051 767
rect 9097 721 9175 767
rect 9221 721 9299 767
rect 9345 721 9423 767
rect 9469 721 9547 767
rect 9593 721 9671 767
rect 9717 721 9795 767
rect 9841 721 9919 767
rect 9965 721 10043 767
rect 10089 721 10167 767
rect 10213 721 10291 767
rect 10337 721 10415 767
rect 10461 721 10539 767
rect 10585 721 10663 767
rect 10709 721 10787 767
rect 10833 721 10911 767
rect 10957 721 11035 767
rect 11081 721 11159 767
rect 11205 721 11283 767
rect 11329 721 11407 767
rect 11453 721 11531 767
rect 11577 721 11655 767
rect 11701 721 11779 767
rect 11825 721 11903 767
rect 11949 721 12027 767
rect 12073 721 12151 767
rect 12197 721 12275 767
rect 12321 721 12399 767
rect 12445 721 12523 767
rect 12569 721 12647 767
rect 12693 721 12771 767
rect 12817 721 12895 767
rect 12941 721 13019 767
rect 13065 721 13143 767
rect 13189 721 13267 767
rect 13313 721 13391 767
rect 13437 721 13515 767
rect 13561 721 13639 767
rect 13685 721 13763 767
rect 13809 721 13887 767
rect 13933 721 14011 767
rect 14057 721 14135 767
rect 14181 721 14259 767
rect 14305 721 14383 767
rect 14429 721 14507 767
rect 14553 721 14631 767
rect 14677 721 14755 767
rect 14801 721 14879 767
rect 14925 721 15003 767
rect 15049 721 15127 767
rect 15173 721 15251 767
rect 15297 721 15375 767
rect 15421 721 15499 767
rect 15545 721 15623 767
rect 15669 721 15747 767
rect 15793 721 15871 767
rect 15917 721 15995 767
rect 16041 721 16119 767
rect 16165 721 16243 767
rect 16289 721 16367 767
rect 16413 721 16491 767
rect 16537 721 16615 767
rect 16661 721 16739 767
rect 16785 721 16863 767
rect 16909 721 16987 767
rect 17033 721 17111 767
rect 17157 721 17235 767
rect 17281 721 17359 767
rect 17405 721 17483 767
rect 17529 721 17607 767
rect 17653 721 17731 767
rect 17777 721 17855 767
rect 17901 721 17979 767
rect 18025 721 18103 767
rect 18149 721 18227 767
rect 18273 721 18351 767
rect 18397 721 18475 767
rect 18521 721 18599 767
rect 18645 721 18723 767
rect 18769 721 18847 767
rect 18893 721 18971 767
rect 19017 721 19095 767
rect 19141 721 19219 767
rect 19265 721 19343 767
rect 19389 721 19467 767
rect 19513 721 19591 767
rect 19637 721 19715 767
rect 19761 721 19839 767
rect 19885 721 19963 767
rect 20009 721 20087 767
rect 20133 721 20211 767
rect 20257 721 20335 767
rect 20381 721 20459 767
rect 20505 721 20583 767
rect 20629 721 20707 767
rect 20753 721 20831 767
rect 20877 721 20955 767
rect 21001 721 21079 767
rect 21125 721 21203 767
rect 21249 721 21327 767
rect 21373 721 21451 767
rect 21497 721 21575 767
rect 21621 721 21699 767
rect 21745 721 21823 767
rect 21869 721 21947 767
rect 21993 721 22071 767
rect 22117 721 22195 767
rect 22241 721 22319 767
rect 22365 721 22443 767
rect 22489 721 22567 767
rect 22613 721 22691 767
rect 22737 721 22815 767
rect 22861 721 22939 767
rect 22985 721 23063 767
rect 23109 721 23187 767
rect 23233 721 23311 767
rect 23357 721 23435 767
rect 23481 721 23559 767
rect 23605 721 23683 767
rect 23729 721 23807 767
rect 23853 721 23931 767
rect 23977 721 24055 767
rect 24101 721 24179 767
rect 24225 721 24303 767
rect 24349 721 24427 767
rect 24473 721 24551 767
rect 24597 721 24675 767
rect 24721 721 24799 767
rect 24845 721 24923 767
rect 24969 721 25047 767
rect 25093 721 25171 767
rect 25217 721 25295 767
rect 25341 721 25419 767
rect 25465 721 25543 767
rect 25589 721 25667 767
rect 25713 721 25791 767
rect 25837 721 25915 767
rect 25961 721 26039 767
rect 26085 721 26163 767
rect 26209 721 26287 767
rect 26333 721 26411 767
rect 26457 721 26535 767
rect 26581 721 26659 767
rect 26705 721 26783 767
rect 26829 721 26907 767
rect 26953 721 27031 767
rect 27077 721 27155 767
rect 27201 721 27279 767
rect 27325 721 27403 767
rect 27449 721 27527 767
rect 27573 721 27651 767
rect 27697 721 27775 767
rect 27821 721 27899 767
rect 27945 721 28023 767
rect 28069 721 28147 767
rect 28193 721 28271 767
rect 28317 721 28395 767
rect 28441 721 28519 767
rect 28565 721 28643 767
rect 28689 721 28767 767
rect 28813 721 28891 767
rect 28937 721 29015 767
rect 29061 721 29139 767
rect 29185 721 29263 767
rect 29309 721 29387 767
rect 29433 721 29511 767
rect 29557 721 29635 767
rect 29681 721 29759 767
rect 29805 721 29883 767
rect 29929 721 30007 767
rect 30053 721 30131 767
rect 30177 721 30255 767
rect 30301 721 30379 767
rect 30425 721 30503 767
rect 30549 721 30627 767
rect 30673 721 30751 767
rect 30797 721 30875 767
rect 30921 721 30999 767
rect 31045 721 31123 767
rect 31169 721 31247 767
rect 31293 721 31371 767
rect 31417 721 31495 767
rect 31541 721 31619 767
rect 31665 721 31743 767
rect 31789 721 31867 767
rect 31913 721 31991 767
rect 32037 721 32115 767
rect 32161 721 32239 767
rect 32285 721 32363 767
rect 32409 721 32487 767
rect 32533 721 32611 767
rect 32657 721 32735 767
rect 32781 721 32859 767
rect 32905 721 32983 767
rect 33029 721 33107 767
rect 33153 721 33231 767
rect 33277 721 33355 767
rect 33401 721 33479 767
rect 33525 721 33603 767
rect 33649 721 33727 767
rect 33773 721 33851 767
rect 33897 721 33975 767
rect 34021 721 34099 767
rect 34145 721 34223 767
rect 34269 721 34347 767
rect 34393 721 34471 767
rect 34517 721 34595 767
rect 34641 721 34719 767
rect 34765 721 34843 767
rect 34889 721 34967 767
rect 35013 721 35091 767
rect 35137 721 35215 767
rect 35261 721 35339 767
rect 35385 721 35463 767
rect 35509 721 35587 767
rect 35633 721 35711 767
rect 35757 721 35835 767
rect 35881 721 35959 767
rect 36005 721 36083 767
rect 36129 721 36207 767
rect 36253 721 36331 767
rect 36377 721 36455 767
rect 36501 721 36579 767
rect 36625 721 36703 767
rect 36749 721 36827 767
rect 36873 721 36951 767
rect 36997 721 37075 767
rect 37121 721 37199 767
rect 37245 721 37323 767
rect 37369 721 37447 767
rect 37493 721 37571 767
rect 37617 721 37695 767
rect 37741 721 37819 767
rect 37865 721 37943 767
rect 37989 721 38067 767
rect 38113 721 38191 767
rect 38237 721 38315 767
rect 38361 721 38439 767
rect 38485 721 38563 767
rect 38609 721 38687 767
rect 38733 721 38811 767
rect 38857 721 38935 767
rect 38981 721 39059 767
rect 39105 721 39183 767
rect 39229 721 39307 767
rect 39353 721 39431 767
rect 39477 721 39555 767
rect 39601 721 39679 767
rect 39725 721 39803 767
rect 39849 721 39927 767
rect 39973 721 40051 767
rect 40097 721 40175 767
rect 40221 721 40299 767
rect 40345 721 40423 767
rect 40469 721 40547 767
rect 40593 721 40671 767
rect 40717 721 40795 767
rect 40841 721 40919 767
rect 40965 721 41043 767
rect 41089 721 41167 767
rect 41213 721 41291 767
rect 41337 721 41415 767
rect 41461 721 41539 767
rect 41585 721 41663 767
rect 41709 721 41787 767
rect 41833 721 41911 767
rect 41957 721 42035 767
rect 42081 721 42159 767
rect 42205 721 42283 767
rect 42329 721 42407 767
rect 42453 721 42531 767
rect 42577 721 42655 767
rect 42701 721 42779 767
rect 42825 721 42903 767
rect 42949 721 43027 767
rect 43073 721 43151 767
rect 43197 721 43275 767
rect 43321 721 43399 767
rect 43445 721 43523 767
rect 43569 721 43647 767
rect 43693 721 43771 767
rect 43817 721 43895 767
rect 43941 721 44019 767
rect 44065 721 44143 767
rect 44189 721 44267 767
rect 44313 721 44391 767
rect 44437 721 44515 767
rect 44561 721 44639 767
rect 44685 721 44763 767
rect 44809 721 44887 767
rect 44933 721 45011 767
rect 45057 721 45135 767
rect 45181 721 45259 767
rect 45305 721 45383 767
rect 45429 721 45507 767
rect 45553 721 45631 767
rect 45677 721 45755 767
rect 45801 721 45879 767
rect 45925 721 46003 767
rect 46049 721 46127 767
rect 46173 721 46251 767
rect 46297 721 46375 767
rect 46421 721 46499 767
rect 46545 721 46623 767
rect 46669 721 46747 767
rect 46793 721 46871 767
rect 46917 721 46995 767
rect 47041 721 47119 767
rect 47165 721 47243 767
rect 47289 721 47367 767
rect 47413 721 47491 767
rect 47537 721 47615 767
rect 47661 721 47739 767
rect 47785 721 47863 767
rect 47909 721 47987 767
rect 48033 721 48111 767
rect 48157 721 48235 767
rect 48281 721 48359 767
rect 48405 721 48483 767
rect 48529 721 48607 767
rect 48653 721 48731 767
rect 48777 721 48855 767
rect 48901 721 48979 767
rect 49025 721 49103 767
rect 49149 721 49227 767
rect 49273 721 49351 767
rect 49397 721 49475 767
rect 49521 721 49599 767
rect 49645 721 49723 767
rect 49769 721 49847 767
rect 49893 721 49971 767
rect 50017 721 50095 767
rect 50141 721 50219 767
rect 50265 721 50343 767
rect 50389 721 50467 767
rect 50513 721 50591 767
rect 50637 721 50715 767
rect 50761 721 50839 767
rect 50885 721 50963 767
rect 51009 721 51087 767
rect 51133 721 51211 767
rect 51257 721 51335 767
rect 51381 721 51459 767
rect 51505 721 51583 767
rect 51629 721 51707 767
rect 51753 721 51831 767
rect 51877 721 51955 767
rect 52001 721 52079 767
rect 52125 721 52203 767
rect 52249 721 52327 767
rect 52373 721 52451 767
rect 52497 721 52575 767
rect 52621 721 52699 767
rect 52745 721 52823 767
rect 52869 721 52947 767
rect 52993 721 53071 767
rect 53117 721 53195 767
rect 53241 721 53319 767
rect 53365 721 53443 767
rect 53489 721 53567 767
rect 53613 721 53691 767
rect 53737 721 53815 767
rect 53861 721 53939 767
rect 53985 721 54063 767
rect 54109 721 54187 767
rect 54233 721 54311 767
rect 54357 721 54435 767
rect 54481 721 54559 767
rect 54605 721 54683 767
rect 54729 721 54807 767
rect 54853 721 54931 767
rect 54977 721 55055 767
rect 55101 721 55179 767
rect 55225 721 55303 767
rect 55349 721 55427 767
rect 55473 721 55551 767
rect 55597 721 55675 767
rect 55721 721 55799 767
rect 55845 721 55923 767
rect 55969 721 56047 767
rect 56093 721 56171 767
rect 56217 721 56295 767
rect 56341 721 56419 767
rect 56465 721 56543 767
rect 56589 721 56667 767
rect 56713 721 56791 767
rect 56837 721 56915 767
rect 56961 721 57039 767
rect 57085 721 57163 767
rect 57209 721 57287 767
rect 57333 721 57411 767
rect 57457 721 57535 767
rect 57581 721 57659 767
rect 57705 721 57783 767
rect 57829 721 57907 767
rect 57953 721 58031 767
rect 58077 721 58155 767
rect 58201 721 58279 767
rect 58325 721 58403 767
rect 58449 721 58527 767
rect 58573 721 58651 767
rect 58697 721 58775 767
rect 58821 721 58899 767
rect 58945 721 59023 767
rect 59069 721 59147 767
rect 59193 721 59271 767
rect 59317 721 59395 767
rect 59441 721 59519 767
rect 59565 721 59643 767
rect 59689 721 59767 767
rect 59813 721 59891 767
rect 59937 721 60015 767
rect 60061 721 60139 767
rect 60185 721 60263 767
rect 60309 721 60387 767
rect 60433 721 60511 767
rect 60557 721 60635 767
rect 60681 721 60759 767
rect 60805 721 60883 767
rect 60929 721 61007 767
rect 61053 721 61131 767
rect 61177 721 61255 767
rect 61301 721 61379 767
rect 61425 721 61503 767
rect 61549 721 61627 767
rect 61673 721 61751 767
rect 61797 721 61875 767
rect 61921 721 61999 767
rect 62045 721 62123 767
rect 62169 721 62247 767
rect 62293 721 62371 767
rect 62417 721 62495 767
rect 62541 721 62619 767
rect 62665 721 62743 767
rect 62789 721 62867 767
rect 62913 721 62991 767
rect 63037 721 63115 767
rect 63161 721 63239 767
rect 63285 721 63363 767
rect 63409 721 63487 767
rect 63533 721 63611 767
rect 63657 721 63735 767
rect 63781 721 63859 767
rect 63905 721 63983 767
rect 64029 721 64107 767
rect 64153 721 64231 767
rect 64277 721 64355 767
rect 64401 721 64479 767
rect 64525 721 64603 767
rect 64649 721 64727 767
rect 64773 721 64851 767
rect 64897 721 64975 767
rect 65021 721 65099 767
rect 65145 721 65223 767
rect 65269 721 65347 767
rect 65393 721 65471 767
rect 65517 721 65595 767
rect 65641 721 65719 767
rect 65765 721 65843 767
rect 65889 721 65967 767
rect 66013 721 66091 767
rect 66137 721 66215 767
rect 66261 721 66339 767
rect 66385 721 66463 767
rect 66509 721 66587 767
rect 66633 721 66711 767
rect 66757 721 66835 767
rect 66881 721 66959 767
rect 67005 721 67083 767
rect 67129 721 67207 767
rect 67253 721 67331 767
rect 67377 721 67455 767
rect 67501 721 67579 767
rect 67625 721 67703 767
rect 67749 721 67827 767
rect 67873 721 67951 767
rect 67997 721 68075 767
rect 68121 721 68199 767
rect 68245 721 68323 767
rect 68369 721 68447 767
rect 68493 721 68571 767
rect 68617 721 68695 767
rect 68741 721 68819 767
rect 68865 721 68943 767
rect 68989 721 69067 767
rect 69113 721 69191 767
rect 69237 721 69315 767
rect 69361 721 69439 767
rect 69485 721 69563 767
rect 69609 721 69687 767
rect 69733 721 69811 767
rect 69857 721 69935 767
rect 69981 721 70059 767
rect 70105 721 70183 767
rect 70229 721 70307 767
rect 70353 721 70431 767
rect 70477 721 70555 767
rect 70601 721 70679 767
rect 70725 721 70803 767
rect 70849 721 70927 767
rect 70973 721 71051 767
rect 71097 721 71175 767
rect 71221 721 71299 767
rect 71345 721 71423 767
rect 71469 721 71547 767
rect 71593 721 71671 767
rect 71717 721 71795 767
rect 71841 721 71919 767
rect 71965 721 72043 767
rect 72089 721 72167 767
rect 72213 721 72291 767
rect 72337 721 72415 767
rect 72461 721 72539 767
rect 72585 721 72663 767
rect 72709 721 72787 767
rect 72833 721 72911 767
rect 72957 721 73035 767
rect 73081 721 73159 767
rect 73205 721 73283 767
rect 73329 721 73407 767
rect 73453 721 73531 767
rect 73577 721 73655 767
rect 73701 721 73779 767
rect 73825 721 73903 767
rect 73949 721 74027 767
rect 74073 721 74151 767
rect 74197 721 74275 767
rect 74321 721 74399 767
rect 74445 721 74523 767
rect 74569 721 74647 767
rect 74693 721 74771 767
rect 74817 721 74895 767
rect 74941 721 75019 767
rect 75065 721 75143 767
rect 75189 721 75267 767
rect 75313 721 75391 767
rect 75437 721 75515 767
rect 75561 721 75639 767
rect 75685 721 75763 767
rect 75809 721 75887 767
rect 75933 721 76011 767
rect 76057 721 76135 767
rect 76181 721 76259 767
rect 76305 721 76383 767
rect 76429 721 76507 767
rect 76553 721 76631 767
rect 76677 721 76755 767
rect 76801 721 76879 767
rect 76925 721 77003 767
rect 77049 721 77127 767
rect 77173 721 77251 767
rect 77297 721 77375 767
rect 77421 721 77499 767
rect 77545 721 77623 767
rect 77669 721 77747 767
rect 77793 721 77871 767
rect 77917 721 77995 767
rect 78041 721 78119 767
rect 78165 721 78243 767
rect 78289 721 78367 767
rect 78413 721 78491 767
rect 78537 721 78615 767
rect 78661 721 78739 767
rect 78785 721 78863 767
rect 78909 721 78987 767
rect 79033 721 79111 767
rect 79157 721 79235 767
rect 79281 721 79359 767
rect 79405 721 79483 767
rect 79529 721 79607 767
rect 79653 721 79731 767
rect 79777 721 79855 767
rect 79901 721 79979 767
rect 80025 721 80103 767
rect 80149 721 80227 767
rect 80273 721 80351 767
rect 80397 721 80475 767
rect 80521 721 80599 767
rect 80645 721 80723 767
rect 80769 721 80847 767
rect 80893 721 80971 767
rect 81017 721 81095 767
rect 81141 721 81219 767
rect 81265 721 81343 767
rect 81389 721 81467 767
rect 81513 721 81591 767
rect 81637 721 81715 767
rect 81761 721 81839 767
rect 81885 721 81963 767
rect 82009 721 82087 767
rect 82133 721 82211 767
rect 82257 721 82335 767
rect 82381 721 82459 767
rect 82505 721 82583 767
rect 82629 721 82707 767
rect 82753 721 82831 767
rect 82877 721 82955 767
rect 83001 721 83079 767
rect 83125 721 83203 767
rect 83249 721 83327 767
rect 83373 721 83451 767
rect 83497 721 83575 767
rect 83621 721 83699 767
rect 83745 721 83823 767
rect 83869 721 83947 767
rect 83993 721 84071 767
rect 84117 721 84195 767
rect 84241 721 84319 767
rect 84365 721 84443 767
rect 84489 721 84567 767
rect 84613 721 84691 767
rect 84737 721 84815 767
rect 84861 721 84939 767
rect 84985 721 85063 767
rect 85109 721 85187 767
rect 85233 721 85311 767
rect 85357 721 85435 767
rect 85481 721 85559 767
rect 85605 721 85683 767
rect 85729 721 85807 767
rect 85853 721 85931 767
rect 85977 721 86098 767
rect 352 643 86098 721
rect 352 597 371 643
rect 417 597 495 643
rect 541 597 619 643
rect 665 597 743 643
rect 789 597 867 643
rect 913 597 991 643
rect 1037 597 1115 643
rect 1161 597 1239 643
rect 1285 597 1363 643
rect 1409 597 1487 643
rect 1533 597 1611 643
rect 1657 597 1735 643
rect 1781 597 1859 643
rect 1905 597 1983 643
rect 2029 597 2107 643
rect 2153 597 2231 643
rect 2277 597 2355 643
rect 2401 597 2479 643
rect 2525 597 2603 643
rect 2649 597 2727 643
rect 2773 597 2851 643
rect 2897 597 2975 643
rect 3021 597 3099 643
rect 3145 597 3223 643
rect 3269 597 3347 643
rect 3393 597 3471 643
rect 3517 597 3595 643
rect 3641 597 3719 643
rect 3765 597 3843 643
rect 3889 597 3967 643
rect 4013 597 4091 643
rect 4137 597 4215 643
rect 4261 597 4339 643
rect 4385 597 4463 643
rect 4509 597 4587 643
rect 4633 597 4711 643
rect 4757 597 4835 643
rect 4881 597 4959 643
rect 5005 597 5083 643
rect 5129 597 5207 643
rect 5253 597 5331 643
rect 5377 597 5455 643
rect 5501 597 5579 643
rect 5625 597 5703 643
rect 5749 597 5827 643
rect 5873 597 5951 643
rect 5997 597 6075 643
rect 6121 597 6199 643
rect 6245 597 6323 643
rect 6369 597 6447 643
rect 6493 597 6571 643
rect 6617 597 6695 643
rect 6741 597 6819 643
rect 6865 597 6943 643
rect 6989 597 7067 643
rect 7113 597 7191 643
rect 7237 597 7315 643
rect 7361 597 7439 643
rect 7485 597 7563 643
rect 7609 597 7687 643
rect 7733 597 7811 643
rect 7857 597 7935 643
rect 7981 597 8059 643
rect 8105 597 8183 643
rect 8229 597 8307 643
rect 8353 597 8431 643
rect 8477 597 8555 643
rect 8601 597 8679 643
rect 8725 597 8803 643
rect 8849 597 8927 643
rect 8973 597 9051 643
rect 9097 597 9175 643
rect 9221 597 9299 643
rect 9345 597 9423 643
rect 9469 597 9547 643
rect 9593 597 9671 643
rect 9717 597 9795 643
rect 9841 597 9919 643
rect 9965 597 10043 643
rect 10089 597 10167 643
rect 10213 597 10291 643
rect 10337 597 10415 643
rect 10461 597 10539 643
rect 10585 597 10663 643
rect 10709 597 10787 643
rect 10833 597 10911 643
rect 10957 597 11035 643
rect 11081 597 11159 643
rect 11205 597 11283 643
rect 11329 597 11407 643
rect 11453 597 11531 643
rect 11577 597 11655 643
rect 11701 597 11779 643
rect 11825 597 11903 643
rect 11949 597 12027 643
rect 12073 597 12151 643
rect 12197 597 12275 643
rect 12321 597 12399 643
rect 12445 597 12523 643
rect 12569 597 12647 643
rect 12693 597 12771 643
rect 12817 597 12895 643
rect 12941 597 13019 643
rect 13065 597 13143 643
rect 13189 597 13267 643
rect 13313 597 13391 643
rect 13437 597 13515 643
rect 13561 597 13639 643
rect 13685 597 13763 643
rect 13809 597 13887 643
rect 13933 597 14011 643
rect 14057 597 14135 643
rect 14181 597 14259 643
rect 14305 597 14383 643
rect 14429 597 14507 643
rect 14553 597 14631 643
rect 14677 597 14755 643
rect 14801 597 14879 643
rect 14925 597 15003 643
rect 15049 597 15127 643
rect 15173 597 15251 643
rect 15297 597 15375 643
rect 15421 597 15499 643
rect 15545 597 15623 643
rect 15669 597 15747 643
rect 15793 597 15871 643
rect 15917 597 15995 643
rect 16041 597 16119 643
rect 16165 597 16243 643
rect 16289 597 16367 643
rect 16413 597 16491 643
rect 16537 597 16615 643
rect 16661 597 16739 643
rect 16785 597 16863 643
rect 16909 597 16987 643
rect 17033 597 17111 643
rect 17157 597 17235 643
rect 17281 597 17359 643
rect 17405 597 17483 643
rect 17529 597 17607 643
rect 17653 597 17731 643
rect 17777 597 17855 643
rect 17901 597 17979 643
rect 18025 597 18103 643
rect 18149 597 18227 643
rect 18273 597 18351 643
rect 18397 597 18475 643
rect 18521 597 18599 643
rect 18645 597 18723 643
rect 18769 597 18847 643
rect 18893 597 18971 643
rect 19017 597 19095 643
rect 19141 597 19219 643
rect 19265 597 19343 643
rect 19389 597 19467 643
rect 19513 597 19591 643
rect 19637 597 19715 643
rect 19761 597 19839 643
rect 19885 597 19963 643
rect 20009 597 20087 643
rect 20133 597 20211 643
rect 20257 597 20335 643
rect 20381 597 20459 643
rect 20505 597 20583 643
rect 20629 597 20707 643
rect 20753 597 20831 643
rect 20877 597 20955 643
rect 21001 597 21079 643
rect 21125 597 21203 643
rect 21249 597 21327 643
rect 21373 597 21451 643
rect 21497 597 21575 643
rect 21621 597 21699 643
rect 21745 597 21823 643
rect 21869 597 21947 643
rect 21993 597 22071 643
rect 22117 597 22195 643
rect 22241 597 22319 643
rect 22365 597 22443 643
rect 22489 597 22567 643
rect 22613 597 22691 643
rect 22737 597 22815 643
rect 22861 597 22939 643
rect 22985 597 23063 643
rect 23109 597 23187 643
rect 23233 597 23311 643
rect 23357 597 23435 643
rect 23481 597 23559 643
rect 23605 597 23683 643
rect 23729 597 23807 643
rect 23853 597 23931 643
rect 23977 597 24055 643
rect 24101 597 24179 643
rect 24225 597 24303 643
rect 24349 597 24427 643
rect 24473 597 24551 643
rect 24597 597 24675 643
rect 24721 597 24799 643
rect 24845 597 24923 643
rect 24969 597 25047 643
rect 25093 597 25171 643
rect 25217 597 25295 643
rect 25341 597 25419 643
rect 25465 597 25543 643
rect 25589 597 25667 643
rect 25713 597 25791 643
rect 25837 597 25915 643
rect 25961 597 26039 643
rect 26085 597 26163 643
rect 26209 597 26287 643
rect 26333 597 26411 643
rect 26457 597 26535 643
rect 26581 597 26659 643
rect 26705 597 26783 643
rect 26829 597 26907 643
rect 26953 597 27031 643
rect 27077 597 27155 643
rect 27201 597 27279 643
rect 27325 597 27403 643
rect 27449 597 27527 643
rect 27573 597 27651 643
rect 27697 597 27775 643
rect 27821 597 27899 643
rect 27945 597 28023 643
rect 28069 597 28147 643
rect 28193 597 28271 643
rect 28317 597 28395 643
rect 28441 597 28519 643
rect 28565 597 28643 643
rect 28689 597 28767 643
rect 28813 597 28891 643
rect 28937 597 29015 643
rect 29061 597 29139 643
rect 29185 597 29263 643
rect 29309 597 29387 643
rect 29433 597 29511 643
rect 29557 597 29635 643
rect 29681 597 29759 643
rect 29805 597 29883 643
rect 29929 597 30007 643
rect 30053 597 30131 643
rect 30177 597 30255 643
rect 30301 597 30379 643
rect 30425 597 30503 643
rect 30549 597 30627 643
rect 30673 597 30751 643
rect 30797 597 30875 643
rect 30921 597 30999 643
rect 31045 597 31123 643
rect 31169 597 31247 643
rect 31293 597 31371 643
rect 31417 597 31495 643
rect 31541 597 31619 643
rect 31665 597 31743 643
rect 31789 597 31867 643
rect 31913 597 31991 643
rect 32037 597 32115 643
rect 32161 597 32239 643
rect 32285 597 32363 643
rect 32409 597 32487 643
rect 32533 597 32611 643
rect 32657 597 32735 643
rect 32781 597 32859 643
rect 32905 597 32983 643
rect 33029 597 33107 643
rect 33153 597 33231 643
rect 33277 597 33355 643
rect 33401 597 33479 643
rect 33525 597 33603 643
rect 33649 597 33727 643
rect 33773 597 33851 643
rect 33897 597 33975 643
rect 34021 597 34099 643
rect 34145 597 34223 643
rect 34269 597 34347 643
rect 34393 597 34471 643
rect 34517 597 34595 643
rect 34641 597 34719 643
rect 34765 597 34843 643
rect 34889 597 34967 643
rect 35013 597 35091 643
rect 35137 597 35215 643
rect 35261 597 35339 643
rect 35385 597 35463 643
rect 35509 597 35587 643
rect 35633 597 35711 643
rect 35757 597 35835 643
rect 35881 597 35959 643
rect 36005 597 36083 643
rect 36129 597 36207 643
rect 36253 597 36331 643
rect 36377 597 36455 643
rect 36501 597 36579 643
rect 36625 597 36703 643
rect 36749 597 36827 643
rect 36873 597 36951 643
rect 36997 597 37075 643
rect 37121 597 37199 643
rect 37245 597 37323 643
rect 37369 597 37447 643
rect 37493 597 37571 643
rect 37617 597 37695 643
rect 37741 597 37819 643
rect 37865 597 37943 643
rect 37989 597 38067 643
rect 38113 597 38191 643
rect 38237 597 38315 643
rect 38361 597 38439 643
rect 38485 597 38563 643
rect 38609 597 38687 643
rect 38733 597 38811 643
rect 38857 597 38935 643
rect 38981 597 39059 643
rect 39105 597 39183 643
rect 39229 597 39307 643
rect 39353 597 39431 643
rect 39477 597 39555 643
rect 39601 597 39679 643
rect 39725 597 39803 643
rect 39849 597 39927 643
rect 39973 597 40051 643
rect 40097 597 40175 643
rect 40221 597 40299 643
rect 40345 597 40423 643
rect 40469 597 40547 643
rect 40593 597 40671 643
rect 40717 597 40795 643
rect 40841 597 40919 643
rect 40965 597 41043 643
rect 41089 597 41167 643
rect 41213 597 41291 643
rect 41337 597 41415 643
rect 41461 597 41539 643
rect 41585 597 41663 643
rect 41709 597 41787 643
rect 41833 597 41911 643
rect 41957 597 42035 643
rect 42081 597 42159 643
rect 42205 597 42283 643
rect 42329 597 42407 643
rect 42453 597 42531 643
rect 42577 597 42655 643
rect 42701 597 42779 643
rect 42825 597 42903 643
rect 42949 597 43027 643
rect 43073 597 43151 643
rect 43197 597 43275 643
rect 43321 597 43399 643
rect 43445 597 43523 643
rect 43569 597 43647 643
rect 43693 597 43771 643
rect 43817 597 43895 643
rect 43941 597 44019 643
rect 44065 597 44143 643
rect 44189 597 44267 643
rect 44313 597 44391 643
rect 44437 597 44515 643
rect 44561 597 44639 643
rect 44685 597 44763 643
rect 44809 597 44887 643
rect 44933 597 45011 643
rect 45057 597 45135 643
rect 45181 597 45259 643
rect 45305 597 45383 643
rect 45429 597 45507 643
rect 45553 597 45631 643
rect 45677 597 45755 643
rect 45801 597 45879 643
rect 45925 597 46003 643
rect 46049 597 46127 643
rect 46173 597 46251 643
rect 46297 597 46375 643
rect 46421 597 46499 643
rect 46545 597 46623 643
rect 46669 597 46747 643
rect 46793 597 46871 643
rect 46917 597 46995 643
rect 47041 597 47119 643
rect 47165 597 47243 643
rect 47289 597 47367 643
rect 47413 597 47491 643
rect 47537 597 47615 643
rect 47661 597 47739 643
rect 47785 597 47863 643
rect 47909 597 47987 643
rect 48033 597 48111 643
rect 48157 597 48235 643
rect 48281 597 48359 643
rect 48405 597 48483 643
rect 48529 597 48607 643
rect 48653 597 48731 643
rect 48777 597 48855 643
rect 48901 597 48979 643
rect 49025 597 49103 643
rect 49149 597 49227 643
rect 49273 597 49351 643
rect 49397 597 49475 643
rect 49521 597 49599 643
rect 49645 597 49723 643
rect 49769 597 49847 643
rect 49893 597 49971 643
rect 50017 597 50095 643
rect 50141 597 50219 643
rect 50265 597 50343 643
rect 50389 597 50467 643
rect 50513 597 50591 643
rect 50637 597 50715 643
rect 50761 597 50839 643
rect 50885 597 50963 643
rect 51009 597 51087 643
rect 51133 597 51211 643
rect 51257 597 51335 643
rect 51381 597 51459 643
rect 51505 597 51583 643
rect 51629 597 51707 643
rect 51753 597 51831 643
rect 51877 597 51955 643
rect 52001 597 52079 643
rect 52125 597 52203 643
rect 52249 597 52327 643
rect 52373 597 52451 643
rect 52497 597 52575 643
rect 52621 597 52699 643
rect 52745 597 52823 643
rect 52869 597 52947 643
rect 52993 597 53071 643
rect 53117 597 53195 643
rect 53241 597 53319 643
rect 53365 597 53443 643
rect 53489 597 53567 643
rect 53613 597 53691 643
rect 53737 597 53815 643
rect 53861 597 53939 643
rect 53985 597 54063 643
rect 54109 597 54187 643
rect 54233 597 54311 643
rect 54357 597 54435 643
rect 54481 597 54559 643
rect 54605 597 54683 643
rect 54729 597 54807 643
rect 54853 597 54931 643
rect 54977 597 55055 643
rect 55101 597 55179 643
rect 55225 597 55303 643
rect 55349 597 55427 643
rect 55473 597 55551 643
rect 55597 597 55675 643
rect 55721 597 55799 643
rect 55845 597 55923 643
rect 55969 597 56047 643
rect 56093 597 56171 643
rect 56217 597 56295 643
rect 56341 597 56419 643
rect 56465 597 56543 643
rect 56589 597 56667 643
rect 56713 597 56791 643
rect 56837 597 56915 643
rect 56961 597 57039 643
rect 57085 597 57163 643
rect 57209 597 57287 643
rect 57333 597 57411 643
rect 57457 597 57535 643
rect 57581 597 57659 643
rect 57705 597 57783 643
rect 57829 597 57907 643
rect 57953 597 58031 643
rect 58077 597 58155 643
rect 58201 597 58279 643
rect 58325 597 58403 643
rect 58449 597 58527 643
rect 58573 597 58651 643
rect 58697 597 58775 643
rect 58821 597 58899 643
rect 58945 597 59023 643
rect 59069 597 59147 643
rect 59193 597 59271 643
rect 59317 597 59395 643
rect 59441 597 59519 643
rect 59565 597 59643 643
rect 59689 597 59767 643
rect 59813 597 59891 643
rect 59937 597 60015 643
rect 60061 597 60139 643
rect 60185 597 60263 643
rect 60309 597 60387 643
rect 60433 597 60511 643
rect 60557 597 60635 643
rect 60681 597 60759 643
rect 60805 597 60883 643
rect 60929 597 61007 643
rect 61053 597 61131 643
rect 61177 597 61255 643
rect 61301 597 61379 643
rect 61425 597 61503 643
rect 61549 597 61627 643
rect 61673 597 61751 643
rect 61797 597 61875 643
rect 61921 597 61999 643
rect 62045 597 62123 643
rect 62169 597 62247 643
rect 62293 597 62371 643
rect 62417 597 62495 643
rect 62541 597 62619 643
rect 62665 597 62743 643
rect 62789 597 62867 643
rect 62913 597 62991 643
rect 63037 597 63115 643
rect 63161 597 63239 643
rect 63285 597 63363 643
rect 63409 597 63487 643
rect 63533 597 63611 643
rect 63657 597 63735 643
rect 63781 597 63859 643
rect 63905 597 63983 643
rect 64029 597 64107 643
rect 64153 597 64231 643
rect 64277 597 64355 643
rect 64401 597 64479 643
rect 64525 597 64603 643
rect 64649 597 64727 643
rect 64773 597 64851 643
rect 64897 597 64975 643
rect 65021 597 65099 643
rect 65145 597 65223 643
rect 65269 597 65347 643
rect 65393 597 65471 643
rect 65517 597 65595 643
rect 65641 597 65719 643
rect 65765 597 65843 643
rect 65889 597 65967 643
rect 66013 597 66091 643
rect 66137 597 66215 643
rect 66261 597 66339 643
rect 66385 597 66463 643
rect 66509 597 66587 643
rect 66633 597 66711 643
rect 66757 597 66835 643
rect 66881 597 66959 643
rect 67005 597 67083 643
rect 67129 597 67207 643
rect 67253 597 67331 643
rect 67377 597 67455 643
rect 67501 597 67579 643
rect 67625 597 67703 643
rect 67749 597 67827 643
rect 67873 597 67951 643
rect 67997 597 68075 643
rect 68121 597 68199 643
rect 68245 597 68323 643
rect 68369 597 68447 643
rect 68493 597 68571 643
rect 68617 597 68695 643
rect 68741 597 68819 643
rect 68865 597 68943 643
rect 68989 597 69067 643
rect 69113 597 69191 643
rect 69237 597 69315 643
rect 69361 597 69439 643
rect 69485 597 69563 643
rect 69609 597 69687 643
rect 69733 597 69811 643
rect 69857 597 69935 643
rect 69981 597 70059 643
rect 70105 597 70183 643
rect 70229 597 70307 643
rect 70353 597 70431 643
rect 70477 597 70555 643
rect 70601 597 70679 643
rect 70725 597 70803 643
rect 70849 597 70927 643
rect 70973 597 71051 643
rect 71097 597 71175 643
rect 71221 597 71299 643
rect 71345 597 71423 643
rect 71469 597 71547 643
rect 71593 597 71671 643
rect 71717 597 71795 643
rect 71841 597 71919 643
rect 71965 597 72043 643
rect 72089 597 72167 643
rect 72213 597 72291 643
rect 72337 597 72415 643
rect 72461 597 72539 643
rect 72585 597 72663 643
rect 72709 597 72787 643
rect 72833 597 72911 643
rect 72957 597 73035 643
rect 73081 597 73159 643
rect 73205 597 73283 643
rect 73329 597 73407 643
rect 73453 597 73531 643
rect 73577 597 73655 643
rect 73701 597 73779 643
rect 73825 597 73903 643
rect 73949 597 74027 643
rect 74073 597 74151 643
rect 74197 597 74275 643
rect 74321 597 74399 643
rect 74445 597 74523 643
rect 74569 597 74647 643
rect 74693 597 74771 643
rect 74817 597 74895 643
rect 74941 597 75019 643
rect 75065 597 75143 643
rect 75189 597 75267 643
rect 75313 597 75391 643
rect 75437 597 75515 643
rect 75561 597 75639 643
rect 75685 597 75763 643
rect 75809 597 75887 643
rect 75933 597 76011 643
rect 76057 597 76135 643
rect 76181 597 76259 643
rect 76305 597 76383 643
rect 76429 597 76507 643
rect 76553 597 76631 643
rect 76677 597 76755 643
rect 76801 597 76879 643
rect 76925 597 77003 643
rect 77049 597 77127 643
rect 77173 597 77251 643
rect 77297 597 77375 643
rect 77421 597 77499 643
rect 77545 597 77623 643
rect 77669 597 77747 643
rect 77793 597 77871 643
rect 77917 597 77995 643
rect 78041 597 78119 643
rect 78165 597 78243 643
rect 78289 597 78367 643
rect 78413 597 78491 643
rect 78537 597 78615 643
rect 78661 597 78739 643
rect 78785 597 78863 643
rect 78909 597 78987 643
rect 79033 597 79111 643
rect 79157 597 79235 643
rect 79281 597 79359 643
rect 79405 597 79483 643
rect 79529 597 79607 643
rect 79653 597 79731 643
rect 79777 597 79855 643
rect 79901 597 79979 643
rect 80025 597 80103 643
rect 80149 597 80227 643
rect 80273 597 80351 643
rect 80397 597 80475 643
rect 80521 597 80599 643
rect 80645 597 80723 643
rect 80769 597 80847 643
rect 80893 597 80971 643
rect 81017 597 81095 643
rect 81141 597 81219 643
rect 81265 597 81343 643
rect 81389 597 81467 643
rect 81513 597 81591 643
rect 81637 597 81715 643
rect 81761 597 81839 643
rect 81885 597 81963 643
rect 82009 597 82087 643
rect 82133 597 82211 643
rect 82257 597 82335 643
rect 82381 597 82459 643
rect 82505 597 82583 643
rect 82629 597 82707 643
rect 82753 597 82831 643
rect 82877 597 82955 643
rect 83001 597 83079 643
rect 83125 597 83203 643
rect 83249 597 83327 643
rect 83373 597 83451 643
rect 83497 597 83575 643
rect 83621 597 83699 643
rect 83745 597 83823 643
rect 83869 597 83947 643
rect 83993 597 84071 643
rect 84117 597 84195 643
rect 84241 597 84319 643
rect 84365 597 84443 643
rect 84489 597 84567 643
rect 84613 597 84691 643
rect 84737 597 84815 643
rect 84861 597 84939 643
rect 84985 597 85063 643
rect 85109 597 85187 643
rect 85233 597 85311 643
rect 85357 597 85435 643
rect 85481 597 85559 643
rect 85605 597 85683 643
rect 85729 597 85807 643
rect 85853 597 85931 643
rect 85977 597 86098 643
rect 352 578 86098 597
<< mvnsubdiff >>
rect 30583 44293 30802 44294
rect 30583 44236 32694 44293
rect 30583 44190 30854 44236
rect 30900 44190 31012 44236
rect 31058 44190 31170 44236
rect 31216 44190 31328 44236
rect 31374 44190 31487 44236
rect 31533 44190 31645 44236
rect 31691 44190 31803 44236
rect 31849 44190 31961 44236
rect 32007 44190 32119 44236
rect 32165 44190 32277 44236
rect 32323 44190 32435 44236
rect 32481 44190 32593 44236
rect 32639 44190 32694 44236
rect 30583 44122 32694 44190
rect 42662 44309 43608 44366
rect 42662 44263 42717 44309
rect 42763 44263 42875 44309
rect 42921 44263 43033 44309
rect 43079 44263 43191 44309
rect 43237 44263 43350 44309
rect 43396 44263 43508 44309
rect 43554 44263 43608 44309
rect 42662 44206 43608 44263
rect 30583 44076 30637 44122
rect 30683 44076 32694 44122
rect 30583 44073 32694 44076
rect 30583 44027 30854 44073
rect 30900 44027 31012 44073
rect 31058 44027 31170 44073
rect 31216 44027 31328 44073
rect 31374 44027 31487 44073
rect 31533 44027 31645 44073
rect 31691 44027 31803 44073
rect 31849 44027 31961 44073
rect 32007 44027 32119 44073
rect 32165 44027 32277 44073
rect 32323 44027 32435 44073
rect 32481 44027 32593 44073
rect 32639 44027 32694 44073
rect 30583 43958 32694 44027
rect 30583 43912 30637 43958
rect 30683 43912 32694 43958
rect 30583 43909 32694 43912
rect 30583 43863 30854 43909
rect 30900 43863 31012 43909
rect 31058 43863 31170 43909
rect 31216 43863 31328 43909
rect 31374 43863 31487 43909
rect 31533 43863 31645 43909
rect 31691 43863 31803 43909
rect 31849 43863 31961 43909
rect 32007 43863 32119 43909
rect 32165 43863 32277 43909
rect 32323 43863 32435 43909
rect 32481 43863 32593 43909
rect 32639 43863 32694 43909
rect 30583 43795 32694 43863
rect 54321 44293 54540 44294
rect 52428 44236 54540 44293
rect 52428 44190 52483 44236
rect 52529 44190 52641 44236
rect 52687 44190 52799 44236
rect 52845 44190 52957 44236
rect 53003 44190 53115 44236
rect 53161 44190 53273 44236
rect 53319 44190 53431 44236
rect 53477 44190 53589 44236
rect 53635 44190 53748 44236
rect 53794 44190 53906 44236
rect 53952 44190 54064 44236
rect 54110 44190 54222 44236
rect 54268 44190 54540 44236
rect 30583 43749 30637 43795
rect 30683 43749 32694 43795
rect 30583 43746 32694 43749
rect 30583 43700 30854 43746
rect 30900 43700 31012 43746
rect 31058 43700 31170 43746
rect 31216 43700 31328 43746
rect 31374 43700 31487 43746
rect 31533 43700 31645 43746
rect 31691 43700 31803 43746
rect 31849 43700 31961 43746
rect 32007 43700 32119 43746
rect 32165 43700 32277 43746
rect 32323 43700 32435 43746
rect 32481 43700 32593 43746
rect 32639 43700 32694 43746
rect 52428 44122 54540 44190
rect 52428 44076 54440 44122
rect 54486 44076 54540 44122
rect 52428 44073 54540 44076
rect 52428 44027 52483 44073
rect 52529 44027 52641 44073
rect 52687 44027 52799 44073
rect 52845 44027 52957 44073
rect 53003 44027 53115 44073
rect 53161 44027 53273 44073
rect 53319 44027 53431 44073
rect 53477 44027 53589 44073
rect 53635 44027 53748 44073
rect 53794 44027 53906 44073
rect 53952 44027 54064 44073
rect 54110 44027 54222 44073
rect 54268 44027 54540 44073
rect 52428 43958 54540 44027
rect 52428 43912 54440 43958
rect 54486 43912 54540 43958
rect 52428 43909 54540 43912
rect 52428 43863 52483 43909
rect 52529 43863 52641 43909
rect 52687 43863 52799 43909
rect 52845 43863 52957 43909
rect 53003 43863 53115 43909
rect 53161 43863 53273 43909
rect 53319 43863 53431 43909
rect 53477 43863 53589 43909
rect 53635 43863 53748 43909
rect 53794 43863 53906 43909
rect 53952 43863 54064 43909
rect 54110 43863 54222 43909
rect 54268 43863 54540 43909
rect 52428 43795 54540 43863
rect 52428 43749 54440 43795
rect 54486 43749 54540 43795
rect 52428 43746 54540 43749
rect 30583 43643 32694 43700
rect 52428 43700 52483 43746
rect 52529 43700 52641 43746
rect 52687 43700 52799 43746
rect 52845 43700 52957 43746
rect 53003 43700 53115 43746
rect 53161 43700 53273 43746
rect 53319 43700 53431 43746
rect 53477 43700 53589 43746
rect 53635 43700 53748 43746
rect 53794 43700 53906 43746
rect 53952 43700 54064 43746
rect 54110 43700 54222 43746
rect 54268 43700 54540 43746
rect 52428 43643 54540 43700
rect 30583 43632 30955 43643
rect 30583 43586 30637 43632
rect 30683 43586 30955 43632
rect 30583 43468 30955 43586
rect 30583 43422 30637 43468
rect 30683 43422 30955 43468
rect 30583 43389 30955 43422
rect 54167 43632 54540 43643
rect 54167 43586 54440 43632
rect 54486 43586 54540 43632
rect 54167 43468 54540 43586
rect 54167 43422 54440 43468
rect 54486 43422 54540 43468
rect 30583 43266 30956 43389
rect 36348 43350 36861 43396
rect 36348 43304 36489 43350
rect 36723 43304 36861 43350
rect 30583 43220 30637 43266
rect 30683 43226 30956 43266
rect 30683 43220 30855 43226
rect 30583 43180 30855 43220
rect 30901 43180 30956 43226
rect 30583 43103 30956 43180
rect 30583 43057 30637 43103
rect 30683 43062 30956 43103
rect 30683 43057 30855 43062
rect 30583 43016 30855 43057
rect 30901 43016 30956 43062
rect 30583 42940 30956 43016
rect 30583 42894 30637 42940
rect 30683 42899 30956 42940
rect 30683 42894 30855 42899
rect 30583 42853 30855 42894
rect 30901 42853 30956 42899
rect 30583 42777 30956 42853
rect 30583 42731 30637 42777
rect 30683 42736 30956 42777
rect 30683 42731 30855 42736
rect 30583 42690 30855 42731
rect 30901 42690 30956 42736
rect 36348 43258 36861 43304
rect 39007 43350 39321 43407
rect 39007 43304 39062 43350
rect 39108 43304 39220 43350
rect 39266 43304 39321 43350
rect 39007 43247 39321 43304
rect 45564 43396 48566 43407
rect 45564 43350 48766 43396
rect 54167 43387 54540 43422
rect 45564 43304 45619 43350
rect 45665 43304 45777 43350
rect 45823 43304 45935 43350
rect 45981 43304 46093 43350
rect 46139 43304 46251 43350
rect 46297 43304 46409 43350
rect 46455 43304 46568 43350
rect 46614 43304 46726 43350
rect 46772 43304 46884 43350
rect 46930 43304 47042 43350
rect 47088 43304 47200 43350
rect 47246 43304 47358 43350
rect 47404 43304 47516 43350
rect 47562 43304 47675 43350
rect 47721 43304 47833 43350
rect 47879 43304 47991 43350
rect 48037 43304 48149 43350
rect 48195 43304 48307 43350
rect 48353 43304 48465 43350
rect 48511 43304 48766 43350
rect 45564 43258 48766 43304
rect 45564 43186 48566 43258
rect 45564 43140 45619 43186
rect 45665 43140 45777 43186
rect 45823 43140 45935 43186
rect 45981 43140 46093 43186
rect 46139 43140 46251 43186
rect 46297 43140 46409 43186
rect 46455 43140 46568 43186
rect 46614 43140 46726 43186
rect 46772 43140 46884 43186
rect 46930 43140 47042 43186
rect 47088 43140 47200 43186
rect 47246 43140 47358 43186
rect 47404 43140 47516 43186
rect 47562 43140 47675 43186
rect 47721 43140 47833 43186
rect 47879 43140 47991 43186
rect 48037 43140 48149 43186
rect 48195 43140 48307 43186
rect 48353 43140 48465 43186
rect 48511 43140 48566 43186
rect 54168 43266 54540 43387
rect 54168 43226 54440 43266
rect 54168 43180 54223 43226
rect 54269 43220 54440 43226
rect 54486 43220 54540 43266
rect 54269 43180 54540 43220
rect 45564 43083 48566 43140
rect 30583 42613 30956 42690
rect 30583 42567 30637 42613
rect 30683 42573 30956 42613
rect 30683 42567 30855 42573
rect 30583 42527 30855 42567
rect 30901 42527 30956 42573
rect 54168 43103 54540 43180
rect 54168 43062 54440 43103
rect 54168 43016 54223 43062
rect 54269 43057 54440 43062
rect 54486 43057 54540 43103
rect 54269 43016 54540 43057
rect 54168 42940 54540 43016
rect 54168 42894 54440 42940
rect 54486 42894 54540 42940
rect 54168 42777 54540 42894
rect 54168 42731 54440 42777
rect 54486 42731 54540 42777
rect 54168 42613 54540 42731
rect 54168 42573 54440 42613
rect 30583 42450 30956 42527
rect 54168 42527 54223 42573
rect 54269 42567 54440 42573
rect 54486 42567 54540 42613
rect 54269 42527 54540 42567
rect 30583 42404 30637 42450
rect 30683 42404 30956 42450
rect 30583 42327 30956 42404
rect 54168 42450 54540 42527
rect 54168 42404 54440 42450
rect 54486 42404 54540 42450
rect 30583 42287 30855 42327
rect 30583 42241 30637 42287
rect 30683 42281 30855 42287
rect 30901 42281 30956 42327
rect 54168 42327 54540 42404
rect 30683 42241 30956 42281
rect 30583 42164 30956 42241
rect 30583 42123 30855 42164
rect 30583 42077 30637 42123
rect 30683 42118 30855 42123
rect 30901 42118 30956 42164
rect 30683 42077 30956 42118
rect 30583 42001 30956 42077
rect 30583 41960 30855 42001
rect 30583 41914 30637 41960
rect 30683 41955 30855 41960
rect 30901 41955 30956 42001
rect 30683 41914 30956 41955
rect 30583 41838 30956 41914
rect 30583 41797 30855 41838
rect 30583 41751 30637 41797
rect 30683 41792 30855 41797
rect 30901 41792 30956 41838
rect 30683 41751 30956 41792
rect 30583 41674 30956 41751
rect 30583 41634 30855 41674
rect 30583 41588 30637 41634
rect 30683 41628 30855 41634
rect 30901 41628 30956 41674
rect 30683 41588 30956 41628
rect 30583 41466 30956 41588
rect 54168 42281 54223 42327
rect 54269 42287 54540 42327
rect 54269 42281 54440 42287
rect 54168 42241 54440 42281
rect 54486 42241 54540 42287
rect 36348 41550 36861 41596
rect 36348 41504 36489 41550
rect 36723 41504 36861 41550
rect 30583 41420 30637 41466
rect 30683 41426 30956 41466
rect 30683 41420 30855 41426
rect 30583 41380 30855 41420
rect 30901 41380 30956 41426
rect 30583 41303 30956 41380
rect 30583 41257 30637 41303
rect 30683 41262 30956 41303
rect 30683 41257 30855 41262
rect 30583 41216 30855 41257
rect 30901 41216 30956 41262
rect 30583 41140 30956 41216
rect 30583 41094 30637 41140
rect 30683 41099 30956 41140
rect 30683 41094 30855 41099
rect 30583 41053 30855 41094
rect 30901 41053 30956 41099
rect 30583 40977 30956 41053
rect 30583 40931 30637 40977
rect 30683 40936 30956 40977
rect 30683 40931 30855 40936
rect 30583 40890 30855 40931
rect 30901 40890 30956 40936
rect 36348 41458 36861 41504
rect 39007 41550 39321 41607
rect 39007 41504 39062 41550
rect 39108 41504 39220 41550
rect 39266 41504 39321 41550
rect 39007 41447 39321 41504
rect 45564 41714 48566 41771
rect 45564 41668 45619 41714
rect 45665 41668 45777 41714
rect 45823 41668 45935 41714
rect 45981 41668 46093 41714
rect 46139 41668 46251 41714
rect 46297 41668 46409 41714
rect 46455 41668 46568 41714
rect 46614 41668 46726 41714
rect 46772 41668 46884 41714
rect 46930 41668 47042 41714
rect 47088 41668 47200 41714
rect 47246 41668 47358 41714
rect 47404 41668 47516 41714
rect 47562 41668 47675 41714
rect 47721 41668 47833 41714
rect 47879 41668 47991 41714
rect 48037 41668 48149 41714
rect 48195 41668 48307 41714
rect 48353 41668 48465 41714
rect 48511 41668 48566 41714
rect 54168 42123 54540 42241
rect 54168 42077 54440 42123
rect 54486 42077 54540 42123
rect 54168 41960 54540 42077
rect 54168 41914 54440 41960
rect 54486 41914 54540 41960
rect 54168 41838 54540 41914
rect 54168 41792 54223 41838
rect 54269 41797 54540 41838
rect 54269 41792 54440 41797
rect 54168 41751 54440 41792
rect 54486 41751 54540 41797
rect 45564 41596 48566 41668
rect 45564 41550 48766 41596
rect 54168 41674 54540 41751
rect 54168 41628 54223 41674
rect 54269 41634 54540 41674
rect 54269 41628 54440 41634
rect 54168 41588 54440 41628
rect 54486 41588 54540 41634
rect 45564 41504 45619 41550
rect 45665 41504 45777 41550
rect 45823 41504 45935 41550
rect 45981 41504 46093 41550
rect 46139 41504 46251 41550
rect 46297 41504 46409 41550
rect 46455 41504 46568 41550
rect 46614 41504 46726 41550
rect 46772 41504 46884 41550
rect 46930 41504 47042 41550
rect 47088 41504 47200 41550
rect 47246 41504 47358 41550
rect 47404 41504 47516 41550
rect 47562 41504 47675 41550
rect 47721 41504 47833 41550
rect 47879 41504 47991 41550
rect 48037 41504 48149 41550
rect 48195 41504 48307 41550
rect 48353 41504 48465 41550
rect 48511 41504 48766 41550
rect 45564 41458 48766 41504
rect 45564 41386 48566 41458
rect 45564 41340 45619 41386
rect 45665 41340 45777 41386
rect 45823 41340 45935 41386
rect 45981 41340 46093 41386
rect 46139 41340 46251 41386
rect 46297 41340 46409 41386
rect 46455 41340 46568 41386
rect 46614 41340 46726 41386
rect 46772 41340 46884 41386
rect 46930 41340 47042 41386
rect 47088 41340 47200 41386
rect 47246 41340 47358 41386
rect 47404 41340 47516 41386
rect 47562 41340 47675 41386
rect 47721 41340 47833 41386
rect 47879 41340 47991 41386
rect 48037 41340 48149 41386
rect 48195 41340 48307 41386
rect 48353 41340 48465 41386
rect 48511 41340 48566 41386
rect 54168 41466 54540 41588
rect 54168 41426 54440 41466
rect 54168 41380 54223 41426
rect 54269 41420 54440 41426
rect 54486 41420 54540 41466
rect 54269 41380 54540 41420
rect 45564 41283 48566 41340
rect 30583 40813 30956 40890
rect 30583 40767 30637 40813
rect 30683 40773 30956 40813
rect 30683 40767 30855 40773
rect 30583 40727 30855 40767
rect 30901 40727 30956 40773
rect 54168 41303 54540 41380
rect 54168 41262 54440 41303
rect 54168 41216 54223 41262
rect 54269 41257 54440 41262
rect 54486 41257 54540 41303
rect 54269 41216 54540 41257
rect 54168 41140 54540 41216
rect 54168 41094 54440 41140
rect 54486 41094 54540 41140
rect 54168 40977 54540 41094
rect 54168 40931 54440 40977
rect 54486 40931 54540 40977
rect 54168 40813 54540 40931
rect 54168 40773 54440 40813
rect 30583 40650 30956 40727
rect 54168 40727 54223 40773
rect 54269 40767 54440 40773
rect 54486 40767 54540 40813
rect 54269 40727 54540 40767
rect 30583 40604 30637 40650
rect 30683 40604 30956 40650
rect 30583 40527 30956 40604
rect 54168 40650 54540 40727
rect 54168 40604 54440 40650
rect 54486 40604 54540 40650
rect 30583 40487 30855 40527
rect 30583 40441 30637 40487
rect 30683 40481 30855 40487
rect 30901 40481 30956 40527
rect 54168 40527 54540 40604
rect 30683 40441 30956 40481
rect 30583 40364 30956 40441
rect 30583 40323 30855 40364
rect 30583 40277 30637 40323
rect 30683 40318 30855 40323
rect 30901 40318 30956 40364
rect 30683 40277 30956 40318
rect 30583 40201 30956 40277
rect 30583 40160 30855 40201
rect 30583 40114 30637 40160
rect 30683 40155 30855 40160
rect 30901 40155 30956 40201
rect 30683 40114 30956 40155
rect 30583 40038 30956 40114
rect 30583 39997 30855 40038
rect 30583 39951 30637 39997
rect 30683 39992 30855 39997
rect 30901 39992 30956 40038
rect 30683 39951 30956 39992
rect 30583 39874 30956 39951
rect 30583 39834 30855 39874
rect 30583 39788 30637 39834
rect 30683 39828 30855 39834
rect 30901 39828 30956 39874
rect 30683 39788 30956 39828
rect 30583 39666 30956 39788
rect 54168 40481 54223 40527
rect 54269 40487 54540 40527
rect 54269 40481 54440 40487
rect 54168 40441 54440 40481
rect 54486 40441 54540 40487
rect 36348 39750 36861 39796
rect 36348 39704 36489 39750
rect 36723 39704 36861 39750
rect 30583 39620 30637 39666
rect 30683 39626 30956 39666
rect 30683 39620 30855 39626
rect 30583 39580 30855 39620
rect 30901 39580 30956 39626
rect 30583 39503 30956 39580
rect 30583 39457 30637 39503
rect 30683 39462 30956 39503
rect 30683 39457 30855 39462
rect 30583 39416 30855 39457
rect 30901 39416 30956 39462
rect 30583 39340 30956 39416
rect 30583 39294 30637 39340
rect 30683 39299 30956 39340
rect 30683 39294 30855 39299
rect 30583 39253 30855 39294
rect 30901 39253 30956 39299
rect 30583 39177 30956 39253
rect 30583 39131 30637 39177
rect 30683 39136 30956 39177
rect 30683 39131 30855 39136
rect 30583 39090 30855 39131
rect 30901 39090 30956 39136
rect 36348 39658 36861 39704
rect 39007 39750 39321 39807
rect 39007 39704 39062 39750
rect 39108 39704 39220 39750
rect 39266 39704 39321 39750
rect 39007 39647 39321 39704
rect 45564 39914 48566 39971
rect 45564 39868 45619 39914
rect 45665 39868 45777 39914
rect 45823 39868 45935 39914
rect 45981 39868 46093 39914
rect 46139 39868 46251 39914
rect 46297 39868 46409 39914
rect 46455 39868 46568 39914
rect 46614 39868 46726 39914
rect 46772 39868 46884 39914
rect 46930 39868 47042 39914
rect 47088 39868 47200 39914
rect 47246 39868 47358 39914
rect 47404 39868 47516 39914
rect 47562 39868 47675 39914
rect 47721 39868 47833 39914
rect 47879 39868 47991 39914
rect 48037 39868 48149 39914
rect 48195 39868 48307 39914
rect 48353 39868 48465 39914
rect 48511 39868 48566 39914
rect 54168 40323 54540 40441
rect 54168 40277 54440 40323
rect 54486 40277 54540 40323
rect 54168 40160 54540 40277
rect 54168 40114 54440 40160
rect 54486 40114 54540 40160
rect 54168 40038 54540 40114
rect 54168 39992 54223 40038
rect 54269 39997 54540 40038
rect 54269 39992 54440 39997
rect 54168 39951 54440 39992
rect 54486 39951 54540 39997
rect 45564 39796 48566 39868
rect 45564 39750 48766 39796
rect 54168 39874 54540 39951
rect 54168 39828 54223 39874
rect 54269 39834 54540 39874
rect 54269 39828 54440 39834
rect 54168 39788 54440 39828
rect 54486 39788 54540 39834
rect 45564 39704 45619 39750
rect 45665 39704 45777 39750
rect 45823 39704 45935 39750
rect 45981 39704 46093 39750
rect 46139 39704 46251 39750
rect 46297 39704 46409 39750
rect 46455 39704 46568 39750
rect 46614 39704 46726 39750
rect 46772 39704 46884 39750
rect 46930 39704 47042 39750
rect 47088 39704 47200 39750
rect 47246 39704 47358 39750
rect 47404 39704 47516 39750
rect 47562 39704 47675 39750
rect 47721 39704 47833 39750
rect 47879 39704 47991 39750
rect 48037 39704 48149 39750
rect 48195 39704 48307 39750
rect 48353 39704 48465 39750
rect 48511 39704 48766 39750
rect 45564 39658 48766 39704
rect 45564 39586 48566 39658
rect 45564 39540 45619 39586
rect 45665 39540 45777 39586
rect 45823 39540 45935 39586
rect 45981 39540 46093 39586
rect 46139 39540 46251 39586
rect 46297 39540 46409 39586
rect 46455 39540 46568 39586
rect 46614 39540 46726 39586
rect 46772 39540 46884 39586
rect 46930 39540 47042 39586
rect 47088 39540 47200 39586
rect 47246 39540 47358 39586
rect 47404 39540 47516 39586
rect 47562 39540 47675 39586
rect 47721 39540 47833 39586
rect 47879 39540 47991 39586
rect 48037 39540 48149 39586
rect 48195 39540 48307 39586
rect 48353 39540 48465 39586
rect 48511 39540 48566 39586
rect 54168 39666 54540 39788
rect 54168 39626 54440 39666
rect 54168 39580 54223 39626
rect 54269 39620 54440 39626
rect 54486 39620 54540 39666
rect 54269 39580 54540 39620
rect 45564 39483 48566 39540
rect 30583 39013 30956 39090
rect 30583 38967 30637 39013
rect 30683 38973 30956 39013
rect 30683 38967 30855 38973
rect 30583 38927 30855 38967
rect 30901 38927 30956 38973
rect 54168 39503 54540 39580
rect 54168 39462 54440 39503
rect 54168 39416 54223 39462
rect 54269 39457 54440 39462
rect 54486 39457 54540 39503
rect 54269 39416 54540 39457
rect 54168 39340 54540 39416
rect 54168 39294 54440 39340
rect 54486 39294 54540 39340
rect 54168 39177 54540 39294
rect 54168 39131 54440 39177
rect 54486 39131 54540 39177
rect 54168 39013 54540 39131
rect 54168 38973 54440 39013
rect 30583 38850 30956 38927
rect 54168 38927 54223 38973
rect 54269 38967 54440 38973
rect 54486 38967 54540 39013
rect 54269 38927 54540 38967
rect 30583 38804 30637 38850
rect 30683 38804 30956 38850
rect 30583 38727 30956 38804
rect 54168 38850 54540 38927
rect 54168 38804 54440 38850
rect 54486 38804 54540 38850
rect 30583 38687 30855 38727
rect 30583 38641 30637 38687
rect 30683 38681 30855 38687
rect 30901 38681 30956 38727
rect 54168 38727 54540 38804
rect 30683 38641 30956 38681
rect 30583 38564 30956 38641
rect 30583 38523 30855 38564
rect 30583 38477 30637 38523
rect 30683 38518 30855 38523
rect 30901 38518 30956 38564
rect 30683 38477 30956 38518
rect 30583 38401 30956 38477
rect 30583 38360 30855 38401
rect 30583 38314 30637 38360
rect 30683 38355 30855 38360
rect 30901 38355 30956 38401
rect 30683 38314 30956 38355
rect 30583 38238 30956 38314
rect 30583 38197 30855 38238
rect 30583 38151 30637 38197
rect 30683 38192 30855 38197
rect 30901 38192 30956 38238
rect 30683 38151 30956 38192
rect 30583 38074 30956 38151
rect 30583 38034 30855 38074
rect 30583 37988 30637 38034
rect 30683 38028 30855 38034
rect 30901 38028 30956 38074
rect 30683 37988 30956 38028
rect 30583 37866 30956 37988
rect 54168 38681 54223 38727
rect 54269 38687 54540 38727
rect 54269 38681 54440 38687
rect 54168 38641 54440 38681
rect 54486 38641 54540 38687
rect 36348 37950 36861 37996
rect 36348 37904 36489 37950
rect 36723 37904 36861 37950
rect 30583 37820 30637 37866
rect 30683 37826 30956 37866
rect 30683 37820 30855 37826
rect 30583 37780 30855 37820
rect 30901 37780 30956 37826
rect 30583 37703 30956 37780
rect 30583 37657 30637 37703
rect 30683 37662 30956 37703
rect 30683 37657 30855 37662
rect 30583 37616 30855 37657
rect 30901 37616 30956 37662
rect 30583 37540 30956 37616
rect 30583 37494 30637 37540
rect 30683 37499 30956 37540
rect 30683 37494 30855 37499
rect 30583 37453 30855 37494
rect 30901 37453 30956 37499
rect 30583 37377 30956 37453
rect 30583 37331 30637 37377
rect 30683 37336 30956 37377
rect 30683 37331 30855 37336
rect 30583 37290 30855 37331
rect 30901 37290 30956 37336
rect 36348 37858 36861 37904
rect 39007 37950 39321 38007
rect 39007 37904 39062 37950
rect 39108 37904 39220 37950
rect 39266 37904 39321 37950
rect 39007 37847 39321 37904
rect 45564 38114 48566 38171
rect 45564 38068 45619 38114
rect 45665 38068 45777 38114
rect 45823 38068 45935 38114
rect 45981 38068 46093 38114
rect 46139 38068 46251 38114
rect 46297 38068 46409 38114
rect 46455 38068 46568 38114
rect 46614 38068 46726 38114
rect 46772 38068 46884 38114
rect 46930 38068 47042 38114
rect 47088 38068 47200 38114
rect 47246 38068 47358 38114
rect 47404 38068 47516 38114
rect 47562 38068 47675 38114
rect 47721 38068 47833 38114
rect 47879 38068 47991 38114
rect 48037 38068 48149 38114
rect 48195 38068 48307 38114
rect 48353 38068 48465 38114
rect 48511 38068 48566 38114
rect 54168 38523 54540 38641
rect 54168 38477 54440 38523
rect 54486 38477 54540 38523
rect 54168 38360 54540 38477
rect 54168 38314 54440 38360
rect 54486 38314 54540 38360
rect 54168 38238 54540 38314
rect 54168 38192 54223 38238
rect 54269 38197 54540 38238
rect 54269 38192 54440 38197
rect 54168 38151 54440 38192
rect 54486 38151 54540 38197
rect 45564 37996 48566 38068
rect 45564 37950 48766 37996
rect 54168 38074 54540 38151
rect 54168 38028 54223 38074
rect 54269 38034 54540 38074
rect 54269 38028 54440 38034
rect 54168 37988 54440 38028
rect 54486 37988 54540 38034
rect 45564 37904 45619 37950
rect 45665 37904 45777 37950
rect 45823 37904 45935 37950
rect 45981 37904 46093 37950
rect 46139 37904 46251 37950
rect 46297 37904 46409 37950
rect 46455 37904 46568 37950
rect 46614 37904 46726 37950
rect 46772 37904 46884 37950
rect 46930 37904 47042 37950
rect 47088 37904 47200 37950
rect 47246 37904 47358 37950
rect 47404 37904 47516 37950
rect 47562 37904 47675 37950
rect 47721 37904 47833 37950
rect 47879 37904 47991 37950
rect 48037 37904 48149 37950
rect 48195 37904 48307 37950
rect 48353 37904 48465 37950
rect 48511 37904 48766 37950
rect 45564 37858 48766 37904
rect 45564 37786 48566 37858
rect 45564 37740 45619 37786
rect 45665 37740 45777 37786
rect 45823 37740 45935 37786
rect 45981 37740 46093 37786
rect 46139 37740 46251 37786
rect 46297 37740 46409 37786
rect 46455 37740 46568 37786
rect 46614 37740 46726 37786
rect 46772 37740 46884 37786
rect 46930 37740 47042 37786
rect 47088 37740 47200 37786
rect 47246 37740 47358 37786
rect 47404 37740 47516 37786
rect 47562 37740 47675 37786
rect 47721 37740 47833 37786
rect 47879 37740 47991 37786
rect 48037 37740 48149 37786
rect 48195 37740 48307 37786
rect 48353 37740 48465 37786
rect 48511 37740 48566 37786
rect 54168 37866 54540 37988
rect 54168 37826 54440 37866
rect 54168 37780 54223 37826
rect 54269 37820 54440 37826
rect 54486 37820 54540 37866
rect 54269 37780 54540 37820
rect 45564 37683 48566 37740
rect 30583 37213 30956 37290
rect 30583 37167 30637 37213
rect 30683 37173 30956 37213
rect 30683 37167 30855 37173
rect 30583 37127 30855 37167
rect 30901 37127 30956 37173
rect 54168 37703 54540 37780
rect 54168 37662 54440 37703
rect 54168 37616 54223 37662
rect 54269 37657 54440 37662
rect 54486 37657 54540 37703
rect 54269 37616 54540 37657
rect 54168 37540 54540 37616
rect 54168 37494 54440 37540
rect 54486 37494 54540 37540
rect 54168 37377 54540 37494
rect 54168 37331 54440 37377
rect 54486 37331 54540 37377
rect 54168 37213 54540 37331
rect 54168 37173 54440 37213
rect 30583 37050 30956 37127
rect 54168 37127 54223 37173
rect 54269 37167 54440 37173
rect 54486 37167 54540 37213
rect 54269 37127 54540 37167
rect 30583 37004 30637 37050
rect 30683 37004 30956 37050
rect 30583 36927 30956 37004
rect 54168 37050 54540 37127
rect 54168 37004 54440 37050
rect 54486 37004 54540 37050
rect 30583 36887 30855 36927
rect 30583 36841 30637 36887
rect 30683 36881 30855 36887
rect 30901 36881 30956 36927
rect 54168 36927 54540 37004
rect 30683 36841 30956 36881
rect 30583 36764 30956 36841
rect 30583 36723 30855 36764
rect 30583 36677 30637 36723
rect 30683 36718 30855 36723
rect 30901 36718 30956 36764
rect 30683 36677 30956 36718
rect 30583 36601 30956 36677
rect 30583 36560 30855 36601
rect 30583 36514 30637 36560
rect 30683 36555 30855 36560
rect 30901 36555 30956 36601
rect 30683 36514 30956 36555
rect 30583 36438 30956 36514
rect 30583 36397 30855 36438
rect 30583 36351 30637 36397
rect 30683 36392 30855 36397
rect 30901 36392 30956 36438
rect 30683 36351 30956 36392
rect 30583 36274 30956 36351
rect 30583 36234 30855 36274
rect 30583 36188 30637 36234
rect 30683 36228 30855 36234
rect 30901 36228 30956 36274
rect 30683 36188 30956 36228
rect 30583 36065 30956 36188
rect 54168 36881 54223 36927
rect 54269 36887 54540 36927
rect 54269 36881 54440 36887
rect 54168 36841 54440 36881
rect 54486 36841 54540 36887
rect 36348 36150 36861 36196
rect 36348 36104 36489 36150
rect 36723 36104 36861 36150
rect 30583 36061 30802 36065
rect 36348 36058 36861 36104
rect 39007 36150 39321 36207
rect 39007 36104 39062 36150
rect 39108 36104 39220 36150
rect 39266 36104 39321 36150
rect 39007 36047 39321 36104
rect 45564 36314 48566 36371
rect 45564 36268 45619 36314
rect 45665 36268 45777 36314
rect 45823 36268 45935 36314
rect 45981 36268 46093 36314
rect 46139 36268 46251 36314
rect 46297 36268 46409 36314
rect 46455 36268 46568 36314
rect 46614 36268 46726 36314
rect 46772 36268 46884 36314
rect 46930 36268 47042 36314
rect 47088 36268 47200 36314
rect 47246 36268 47358 36314
rect 47404 36268 47516 36314
rect 47562 36268 47675 36314
rect 47721 36268 47833 36314
rect 47879 36268 47991 36314
rect 48037 36268 48149 36314
rect 48195 36268 48307 36314
rect 48353 36268 48465 36314
rect 48511 36268 48566 36314
rect 54168 36723 54540 36841
rect 54168 36677 54440 36723
rect 54486 36677 54540 36723
rect 54168 36560 54540 36677
rect 54168 36514 54440 36560
rect 54486 36514 54540 36560
rect 54168 36438 54540 36514
rect 54168 36392 54223 36438
rect 54269 36397 54540 36438
rect 54269 36392 54440 36397
rect 54168 36351 54440 36392
rect 54486 36351 54540 36397
rect 45564 36196 48566 36268
rect 45564 36150 48766 36196
rect 54168 36274 54540 36351
rect 54168 36228 54223 36274
rect 54269 36234 54540 36274
rect 54269 36228 54440 36234
rect 54168 36188 54440 36228
rect 54486 36188 54540 36234
rect 45564 36104 45619 36150
rect 45665 36104 45777 36150
rect 45823 36104 45935 36150
rect 45981 36104 46093 36150
rect 46139 36104 46251 36150
rect 46297 36104 46409 36150
rect 46455 36104 46568 36150
rect 46614 36104 46726 36150
rect 46772 36104 46884 36150
rect 46930 36104 47042 36150
rect 47088 36104 47200 36150
rect 47246 36104 47358 36150
rect 47404 36104 47516 36150
rect 47562 36104 47675 36150
rect 47721 36104 47833 36150
rect 47879 36104 47991 36150
rect 48037 36104 48149 36150
rect 48195 36104 48307 36150
rect 48353 36104 48465 36150
rect 48511 36104 48766 36150
rect 45564 36058 48766 36104
rect 54168 36065 54540 36188
rect 54321 36061 54540 36065
rect 45564 36047 48566 36058
<< mvpsubdiffcont >>
rect 371 46037 417 46083
rect 495 46037 541 46083
rect 619 46037 665 46083
rect 743 46037 789 46083
rect 867 46037 913 46083
rect 991 46037 1037 46083
rect 1115 46037 1161 46083
rect 1239 46037 1285 46083
rect 1363 46037 1409 46083
rect 1487 46037 1533 46083
rect 1611 46037 1657 46083
rect 1735 46037 1781 46083
rect 1859 46037 1905 46083
rect 1983 46037 2029 46083
rect 2107 46037 2153 46083
rect 2231 46037 2277 46083
rect 2355 46037 2401 46083
rect 2479 46037 2525 46083
rect 2603 46037 2649 46083
rect 2727 46037 2773 46083
rect 2851 46037 2897 46083
rect 2975 46037 3021 46083
rect 3099 46037 3145 46083
rect 3223 46037 3269 46083
rect 3347 46037 3393 46083
rect 3471 46037 3517 46083
rect 3595 46037 3641 46083
rect 3719 46037 3765 46083
rect 3843 46037 3889 46083
rect 3967 46037 4013 46083
rect 4091 46037 4137 46083
rect 4215 46037 4261 46083
rect 4339 46037 4385 46083
rect 4463 46037 4509 46083
rect 4587 46037 4633 46083
rect 4711 46037 4757 46083
rect 4835 46037 4881 46083
rect 4959 46037 5005 46083
rect 5083 46037 5129 46083
rect 5207 46037 5253 46083
rect 5331 46037 5377 46083
rect 5455 46037 5501 46083
rect 5579 46037 5625 46083
rect 5703 46037 5749 46083
rect 5827 46037 5873 46083
rect 5951 46037 5997 46083
rect 6075 46037 6121 46083
rect 6199 46037 6245 46083
rect 6323 46037 6369 46083
rect 6447 46037 6493 46083
rect 6571 46037 6617 46083
rect 6695 46037 6741 46083
rect 6819 46037 6865 46083
rect 6943 46037 6989 46083
rect 7067 46037 7113 46083
rect 7191 46037 7237 46083
rect 7315 46037 7361 46083
rect 7439 46037 7485 46083
rect 7563 46037 7609 46083
rect 7687 46037 7733 46083
rect 7811 46037 7857 46083
rect 7935 46037 7981 46083
rect 8059 46037 8105 46083
rect 8183 46037 8229 46083
rect 8307 46037 8353 46083
rect 8431 46037 8477 46083
rect 8555 46037 8601 46083
rect 8679 46037 8725 46083
rect 8803 46037 8849 46083
rect 8927 46037 8973 46083
rect 9051 46037 9097 46083
rect 9175 46037 9221 46083
rect 9299 46037 9345 46083
rect 9423 46037 9469 46083
rect 9547 46037 9593 46083
rect 9671 46037 9717 46083
rect 9795 46037 9841 46083
rect 9919 46037 9965 46083
rect 10043 46037 10089 46083
rect 10167 46037 10213 46083
rect 10291 46037 10337 46083
rect 10415 46037 10461 46083
rect 10539 46037 10585 46083
rect 10663 46037 10709 46083
rect 10787 46037 10833 46083
rect 10911 46037 10957 46083
rect 11035 46037 11081 46083
rect 11159 46037 11205 46083
rect 11283 46037 11329 46083
rect 11407 46037 11453 46083
rect 11531 46037 11577 46083
rect 11655 46037 11701 46083
rect 11779 46037 11825 46083
rect 11903 46037 11949 46083
rect 12027 46037 12073 46083
rect 12151 46037 12197 46083
rect 12275 46037 12321 46083
rect 12399 46037 12445 46083
rect 12523 46037 12569 46083
rect 12647 46037 12693 46083
rect 12771 46037 12817 46083
rect 12895 46037 12941 46083
rect 13019 46037 13065 46083
rect 13143 46037 13189 46083
rect 13267 46037 13313 46083
rect 13391 46037 13437 46083
rect 13515 46037 13561 46083
rect 13639 46037 13685 46083
rect 13763 46037 13809 46083
rect 13887 46037 13933 46083
rect 14011 46037 14057 46083
rect 14135 46037 14181 46083
rect 14259 46037 14305 46083
rect 14383 46037 14429 46083
rect 14507 46037 14553 46083
rect 14631 46037 14677 46083
rect 14755 46037 14801 46083
rect 14879 46037 14925 46083
rect 15003 46037 15049 46083
rect 15127 46037 15173 46083
rect 15251 46037 15297 46083
rect 15375 46037 15421 46083
rect 15499 46037 15545 46083
rect 15623 46037 15669 46083
rect 15747 46037 15793 46083
rect 15871 46037 15917 46083
rect 15995 46037 16041 46083
rect 16119 46037 16165 46083
rect 16243 46037 16289 46083
rect 16367 46037 16413 46083
rect 16491 46037 16537 46083
rect 16615 46037 16661 46083
rect 16739 46037 16785 46083
rect 16863 46037 16909 46083
rect 16987 46037 17033 46083
rect 17111 46037 17157 46083
rect 17235 46037 17281 46083
rect 17359 46037 17405 46083
rect 17483 46037 17529 46083
rect 17607 46037 17653 46083
rect 17731 46037 17777 46083
rect 17855 46037 17901 46083
rect 17979 46037 18025 46083
rect 18103 46037 18149 46083
rect 18227 46037 18273 46083
rect 18351 46037 18397 46083
rect 18475 46037 18521 46083
rect 18599 46037 18645 46083
rect 18723 46037 18769 46083
rect 18847 46037 18893 46083
rect 18971 46037 19017 46083
rect 19095 46037 19141 46083
rect 19219 46037 19265 46083
rect 19343 46037 19389 46083
rect 19467 46037 19513 46083
rect 19591 46037 19637 46083
rect 19715 46037 19761 46083
rect 19839 46037 19885 46083
rect 19963 46037 20009 46083
rect 20087 46037 20133 46083
rect 20211 46037 20257 46083
rect 20335 46037 20381 46083
rect 20459 46037 20505 46083
rect 20583 46037 20629 46083
rect 20707 46037 20753 46083
rect 20831 46037 20877 46083
rect 20955 46037 21001 46083
rect 21079 46037 21125 46083
rect 21203 46037 21249 46083
rect 21327 46037 21373 46083
rect 21451 46037 21497 46083
rect 21575 46037 21621 46083
rect 21699 46037 21745 46083
rect 21823 46037 21869 46083
rect 21947 46037 21993 46083
rect 22071 46037 22117 46083
rect 22195 46037 22241 46083
rect 22319 46037 22365 46083
rect 22443 46037 22489 46083
rect 22567 46037 22613 46083
rect 22691 46037 22737 46083
rect 22815 46037 22861 46083
rect 22939 46037 22985 46083
rect 23063 46037 23109 46083
rect 23187 46037 23233 46083
rect 23311 46037 23357 46083
rect 23435 46037 23481 46083
rect 23559 46037 23605 46083
rect 23683 46037 23729 46083
rect 23807 46037 23853 46083
rect 23931 46037 23977 46083
rect 24055 46037 24101 46083
rect 24179 46037 24225 46083
rect 24303 46037 24349 46083
rect 24427 46037 24473 46083
rect 24551 46037 24597 46083
rect 24675 46037 24721 46083
rect 24799 46037 24845 46083
rect 24923 46037 24969 46083
rect 25047 46037 25093 46083
rect 25171 46037 25217 46083
rect 25295 46037 25341 46083
rect 25419 46037 25465 46083
rect 25543 46037 25589 46083
rect 25667 46037 25713 46083
rect 25791 46037 25837 46083
rect 25915 46037 25961 46083
rect 26039 46037 26085 46083
rect 26163 46037 26209 46083
rect 26287 46037 26333 46083
rect 26411 46037 26457 46083
rect 26535 46037 26581 46083
rect 26659 46037 26705 46083
rect 26783 46037 26829 46083
rect 26907 46037 26953 46083
rect 27031 46037 27077 46083
rect 27155 46037 27201 46083
rect 27279 46037 27325 46083
rect 27403 46037 27449 46083
rect 27527 46037 27573 46083
rect 27651 46037 27697 46083
rect 27775 46037 27821 46083
rect 27899 46037 27945 46083
rect 28023 46037 28069 46083
rect 28147 46037 28193 46083
rect 28271 46037 28317 46083
rect 28395 46037 28441 46083
rect 28519 46037 28565 46083
rect 28643 46037 28689 46083
rect 28767 46037 28813 46083
rect 28891 46037 28937 46083
rect 29015 46037 29061 46083
rect 29139 46037 29185 46083
rect 29263 46037 29309 46083
rect 29387 46037 29433 46083
rect 29511 46037 29557 46083
rect 29635 46037 29681 46083
rect 29759 46037 29805 46083
rect 29883 46037 29929 46083
rect 30007 46037 30053 46083
rect 30131 46037 30177 46083
rect 30255 46037 30301 46083
rect 30379 46037 30425 46083
rect 30503 46037 30549 46083
rect 30627 46037 30673 46083
rect 30751 46037 30797 46083
rect 30875 46037 30921 46083
rect 30999 46037 31045 46083
rect 31123 46037 31169 46083
rect 31247 46037 31293 46083
rect 31371 46037 31417 46083
rect 31495 46037 31541 46083
rect 31619 46037 31665 46083
rect 31743 46037 31789 46083
rect 31867 46037 31913 46083
rect 31991 46037 32037 46083
rect 32115 46037 32161 46083
rect 32239 46037 32285 46083
rect 32363 46037 32409 46083
rect 32487 46037 32533 46083
rect 32611 46037 32657 46083
rect 32735 46037 32781 46083
rect 32859 46037 32905 46083
rect 32983 46037 33029 46083
rect 33107 46037 33153 46083
rect 33231 46037 33277 46083
rect 33355 46037 33401 46083
rect 33479 46037 33525 46083
rect 33603 46037 33649 46083
rect 33727 46037 33773 46083
rect 33851 46037 33897 46083
rect 33975 46037 34021 46083
rect 34099 46037 34145 46083
rect 34223 46037 34269 46083
rect 34347 46037 34393 46083
rect 34471 46037 34517 46083
rect 34595 46037 34641 46083
rect 34719 46037 34765 46083
rect 34843 46037 34889 46083
rect 34967 46037 35013 46083
rect 35091 46037 35137 46083
rect 35215 46037 35261 46083
rect 35339 46037 35385 46083
rect 35463 46037 35509 46083
rect 35587 46037 35633 46083
rect 35711 46037 35757 46083
rect 35835 46037 35881 46083
rect 35959 46037 36005 46083
rect 36083 46037 36129 46083
rect 36207 46037 36253 46083
rect 36331 46037 36377 46083
rect 36455 46037 36501 46083
rect 36579 46037 36625 46083
rect 36703 46037 36749 46083
rect 36827 46037 36873 46083
rect 36951 46037 36997 46083
rect 37075 46037 37121 46083
rect 37199 46037 37245 46083
rect 37323 46037 37369 46083
rect 37447 46037 37493 46083
rect 37571 46037 37617 46083
rect 37695 46037 37741 46083
rect 37819 46037 37865 46083
rect 37943 46037 37989 46083
rect 38067 46037 38113 46083
rect 38191 46037 38237 46083
rect 38315 46037 38361 46083
rect 38439 46037 38485 46083
rect 38563 46037 38609 46083
rect 38687 46037 38733 46083
rect 38811 46037 38857 46083
rect 38935 46037 38981 46083
rect 39059 46037 39105 46083
rect 39183 46037 39229 46083
rect 39307 46037 39353 46083
rect 39431 46037 39477 46083
rect 39555 46037 39601 46083
rect 39679 46037 39725 46083
rect 39803 46037 39849 46083
rect 39927 46037 39973 46083
rect 40051 46037 40097 46083
rect 40175 46037 40221 46083
rect 40299 46037 40345 46083
rect 40423 46037 40469 46083
rect 40547 46037 40593 46083
rect 40671 46037 40717 46083
rect 40795 46037 40841 46083
rect 40919 46037 40965 46083
rect 41043 46037 41089 46083
rect 41167 46037 41213 46083
rect 41291 46037 41337 46083
rect 41415 46037 41461 46083
rect 41539 46037 41585 46083
rect 41663 46037 41709 46083
rect 41787 46037 41833 46083
rect 41911 46037 41957 46083
rect 42035 46037 42081 46083
rect 42159 46037 42205 46083
rect 42283 46037 42329 46083
rect 42407 46037 42453 46083
rect 42531 46037 42577 46083
rect 42655 46037 42701 46083
rect 42779 46037 42825 46083
rect 42903 46037 42949 46083
rect 43027 46037 43073 46083
rect 43151 46037 43197 46083
rect 43275 46037 43321 46083
rect 43399 46037 43445 46083
rect 43523 46037 43569 46083
rect 43647 46037 43693 46083
rect 43771 46037 43817 46083
rect 43895 46037 43941 46083
rect 44019 46037 44065 46083
rect 44143 46037 44189 46083
rect 44267 46037 44313 46083
rect 44391 46037 44437 46083
rect 44515 46037 44561 46083
rect 44639 46037 44685 46083
rect 44763 46037 44809 46083
rect 44887 46037 44933 46083
rect 45011 46037 45057 46083
rect 45135 46037 45181 46083
rect 45259 46037 45305 46083
rect 45383 46037 45429 46083
rect 45507 46037 45553 46083
rect 45631 46037 45677 46083
rect 45755 46037 45801 46083
rect 45879 46037 45925 46083
rect 46003 46037 46049 46083
rect 46127 46037 46173 46083
rect 46251 46037 46297 46083
rect 46375 46037 46421 46083
rect 46499 46037 46545 46083
rect 46623 46037 46669 46083
rect 46747 46037 46793 46083
rect 46871 46037 46917 46083
rect 46995 46037 47041 46083
rect 47119 46037 47165 46083
rect 47243 46037 47289 46083
rect 47367 46037 47413 46083
rect 47491 46037 47537 46083
rect 47615 46037 47661 46083
rect 47739 46037 47785 46083
rect 47863 46037 47909 46083
rect 47987 46037 48033 46083
rect 48111 46037 48157 46083
rect 48235 46037 48281 46083
rect 48359 46037 48405 46083
rect 48483 46037 48529 46083
rect 48607 46037 48653 46083
rect 48731 46037 48777 46083
rect 48855 46037 48901 46083
rect 48979 46037 49025 46083
rect 49103 46037 49149 46083
rect 49227 46037 49273 46083
rect 49351 46037 49397 46083
rect 49475 46037 49521 46083
rect 49599 46037 49645 46083
rect 49723 46037 49769 46083
rect 49847 46037 49893 46083
rect 49971 46037 50017 46083
rect 50095 46037 50141 46083
rect 50219 46037 50265 46083
rect 50343 46037 50389 46083
rect 50467 46037 50513 46083
rect 50591 46037 50637 46083
rect 50715 46037 50761 46083
rect 50839 46037 50885 46083
rect 50963 46037 51009 46083
rect 51087 46037 51133 46083
rect 51211 46037 51257 46083
rect 51335 46037 51381 46083
rect 51459 46037 51505 46083
rect 51583 46037 51629 46083
rect 51707 46037 51753 46083
rect 51831 46037 51877 46083
rect 51955 46037 52001 46083
rect 52079 46037 52125 46083
rect 52203 46037 52249 46083
rect 52327 46037 52373 46083
rect 52451 46037 52497 46083
rect 52575 46037 52621 46083
rect 52699 46037 52745 46083
rect 52823 46037 52869 46083
rect 52947 46037 52993 46083
rect 53071 46037 53117 46083
rect 53195 46037 53241 46083
rect 53319 46037 53365 46083
rect 53443 46037 53489 46083
rect 53567 46037 53613 46083
rect 53691 46037 53737 46083
rect 53815 46037 53861 46083
rect 53939 46037 53985 46083
rect 54063 46037 54109 46083
rect 54187 46037 54233 46083
rect 54311 46037 54357 46083
rect 54435 46037 54481 46083
rect 54559 46037 54605 46083
rect 54683 46037 54729 46083
rect 54807 46037 54853 46083
rect 54931 46037 54977 46083
rect 55055 46037 55101 46083
rect 55179 46037 55225 46083
rect 55303 46037 55349 46083
rect 55427 46037 55473 46083
rect 55551 46037 55597 46083
rect 55675 46037 55721 46083
rect 55799 46037 55845 46083
rect 55923 46037 55969 46083
rect 56047 46037 56093 46083
rect 56171 46037 56217 46083
rect 56295 46037 56341 46083
rect 56419 46037 56465 46083
rect 56543 46037 56589 46083
rect 56667 46037 56713 46083
rect 56791 46037 56837 46083
rect 56915 46037 56961 46083
rect 57039 46037 57085 46083
rect 57163 46037 57209 46083
rect 57287 46037 57333 46083
rect 57411 46037 57457 46083
rect 57535 46037 57581 46083
rect 57659 46037 57705 46083
rect 57783 46037 57829 46083
rect 57907 46037 57953 46083
rect 58031 46037 58077 46083
rect 58155 46037 58201 46083
rect 58279 46037 58325 46083
rect 58403 46037 58449 46083
rect 58527 46037 58573 46083
rect 58651 46037 58697 46083
rect 58775 46037 58821 46083
rect 58899 46037 58945 46083
rect 59023 46037 59069 46083
rect 59147 46037 59193 46083
rect 59271 46037 59317 46083
rect 59395 46037 59441 46083
rect 59519 46037 59565 46083
rect 59643 46037 59689 46083
rect 59767 46037 59813 46083
rect 59891 46037 59937 46083
rect 60015 46037 60061 46083
rect 60139 46037 60185 46083
rect 60263 46037 60309 46083
rect 60387 46037 60433 46083
rect 60511 46037 60557 46083
rect 60635 46037 60681 46083
rect 60759 46037 60805 46083
rect 60883 46037 60929 46083
rect 61007 46037 61053 46083
rect 61131 46037 61177 46083
rect 61255 46037 61301 46083
rect 61379 46037 61425 46083
rect 61503 46037 61549 46083
rect 61627 46037 61673 46083
rect 61751 46037 61797 46083
rect 61875 46037 61921 46083
rect 61999 46037 62045 46083
rect 62123 46037 62169 46083
rect 62247 46037 62293 46083
rect 62371 46037 62417 46083
rect 62495 46037 62541 46083
rect 62619 46037 62665 46083
rect 62743 46037 62789 46083
rect 62867 46037 62913 46083
rect 62991 46037 63037 46083
rect 63115 46037 63161 46083
rect 63239 46037 63285 46083
rect 63363 46037 63409 46083
rect 63487 46037 63533 46083
rect 63611 46037 63657 46083
rect 63735 46037 63781 46083
rect 63859 46037 63905 46083
rect 63983 46037 64029 46083
rect 64107 46037 64153 46083
rect 64231 46037 64277 46083
rect 64355 46037 64401 46083
rect 64479 46037 64525 46083
rect 64603 46037 64649 46083
rect 64727 46037 64773 46083
rect 64851 46037 64897 46083
rect 64975 46037 65021 46083
rect 65099 46037 65145 46083
rect 65223 46037 65269 46083
rect 65347 46037 65393 46083
rect 65471 46037 65517 46083
rect 65595 46037 65641 46083
rect 65719 46037 65765 46083
rect 65843 46037 65889 46083
rect 65967 46037 66013 46083
rect 66091 46037 66137 46083
rect 66215 46037 66261 46083
rect 66339 46037 66385 46083
rect 66463 46037 66509 46083
rect 66587 46037 66633 46083
rect 66711 46037 66757 46083
rect 66835 46037 66881 46083
rect 66959 46037 67005 46083
rect 67083 46037 67129 46083
rect 67207 46037 67253 46083
rect 67331 46037 67377 46083
rect 67455 46037 67501 46083
rect 67579 46037 67625 46083
rect 67703 46037 67749 46083
rect 67827 46037 67873 46083
rect 67951 46037 67997 46083
rect 68075 46037 68121 46083
rect 68199 46037 68245 46083
rect 68323 46037 68369 46083
rect 68447 46037 68493 46083
rect 68571 46037 68617 46083
rect 68695 46037 68741 46083
rect 68819 46037 68865 46083
rect 68943 46037 68989 46083
rect 69067 46037 69113 46083
rect 69191 46037 69237 46083
rect 69315 46037 69361 46083
rect 69439 46037 69485 46083
rect 69563 46037 69609 46083
rect 69687 46037 69733 46083
rect 69811 46037 69857 46083
rect 69935 46037 69981 46083
rect 70059 46037 70105 46083
rect 70183 46037 70229 46083
rect 70307 46037 70353 46083
rect 70431 46037 70477 46083
rect 70555 46037 70601 46083
rect 70679 46037 70725 46083
rect 70803 46037 70849 46083
rect 70927 46037 70973 46083
rect 71051 46037 71097 46083
rect 71175 46037 71221 46083
rect 71299 46037 71345 46083
rect 71423 46037 71469 46083
rect 71547 46037 71593 46083
rect 71671 46037 71717 46083
rect 71795 46037 71841 46083
rect 71919 46037 71965 46083
rect 72043 46037 72089 46083
rect 72167 46037 72213 46083
rect 72291 46037 72337 46083
rect 72415 46037 72461 46083
rect 72539 46037 72585 46083
rect 72663 46037 72709 46083
rect 72787 46037 72833 46083
rect 72911 46037 72957 46083
rect 73035 46037 73081 46083
rect 73159 46037 73205 46083
rect 73283 46037 73329 46083
rect 73407 46037 73453 46083
rect 73531 46037 73577 46083
rect 73655 46037 73701 46083
rect 73779 46037 73825 46083
rect 73903 46037 73949 46083
rect 74027 46037 74073 46083
rect 74151 46037 74197 46083
rect 74275 46037 74321 46083
rect 74399 46037 74445 46083
rect 74523 46037 74569 46083
rect 74647 46037 74693 46083
rect 74771 46037 74817 46083
rect 74895 46037 74941 46083
rect 75019 46037 75065 46083
rect 75143 46037 75189 46083
rect 75267 46037 75313 46083
rect 75391 46037 75437 46083
rect 75515 46037 75561 46083
rect 75639 46037 75685 46083
rect 75763 46037 75809 46083
rect 75887 46037 75933 46083
rect 76011 46037 76057 46083
rect 76135 46037 76181 46083
rect 76259 46037 76305 46083
rect 76383 46037 76429 46083
rect 76507 46037 76553 46083
rect 76631 46037 76677 46083
rect 76755 46037 76801 46083
rect 76879 46037 76925 46083
rect 77003 46037 77049 46083
rect 77127 46037 77173 46083
rect 77251 46037 77297 46083
rect 77375 46037 77421 46083
rect 77499 46037 77545 46083
rect 77623 46037 77669 46083
rect 77747 46037 77793 46083
rect 77871 46037 77917 46083
rect 77995 46037 78041 46083
rect 78119 46037 78165 46083
rect 78243 46037 78289 46083
rect 78367 46037 78413 46083
rect 78491 46037 78537 46083
rect 78615 46037 78661 46083
rect 78739 46037 78785 46083
rect 78863 46037 78909 46083
rect 78987 46037 79033 46083
rect 79111 46037 79157 46083
rect 79235 46037 79281 46083
rect 79359 46037 79405 46083
rect 79483 46037 79529 46083
rect 79607 46037 79653 46083
rect 79731 46037 79777 46083
rect 79855 46037 79901 46083
rect 79979 46037 80025 46083
rect 80103 46037 80149 46083
rect 80227 46037 80273 46083
rect 80351 46037 80397 46083
rect 80475 46037 80521 46083
rect 80599 46037 80645 46083
rect 80723 46037 80769 46083
rect 80847 46037 80893 46083
rect 80971 46037 81017 46083
rect 81095 46037 81141 46083
rect 81219 46037 81265 46083
rect 81343 46037 81389 46083
rect 81467 46037 81513 46083
rect 81591 46037 81637 46083
rect 81715 46037 81761 46083
rect 81839 46037 81885 46083
rect 81963 46037 82009 46083
rect 82087 46037 82133 46083
rect 82211 46037 82257 46083
rect 82335 46037 82381 46083
rect 82459 46037 82505 46083
rect 82583 46037 82629 46083
rect 82707 46037 82753 46083
rect 82831 46037 82877 46083
rect 82955 46037 83001 46083
rect 83079 46037 83125 46083
rect 83203 46037 83249 46083
rect 83327 46037 83373 46083
rect 83451 46037 83497 46083
rect 83575 46037 83621 46083
rect 83699 46037 83745 46083
rect 83823 46037 83869 46083
rect 83947 46037 83993 46083
rect 84071 46037 84117 46083
rect 84195 46037 84241 46083
rect 84319 46037 84365 46083
rect 84443 46037 84489 46083
rect 84567 46037 84613 46083
rect 84691 46037 84737 46083
rect 84815 46037 84861 46083
rect 84939 46037 84985 46083
rect 85063 46037 85109 46083
rect 85187 46037 85233 46083
rect 85311 46037 85357 46083
rect 85435 46037 85481 46083
rect 85559 46037 85605 46083
rect 85683 46037 85729 46083
rect 85807 46037 85853 46083
rect 85931 46037 85977 46083
rect 371 45913 417 45959
rect 495 45913 541 45959
rect 619 45913 665 45959
rect 743 45913 789 45959
rect 867 45913 913 45959
rect 991 45913 1037 45959
rect 1115 45913 1161 45959
rect 1239 45913 1285 45959
rect 1363 45913 1409 45959
rect 1487 45913 1533 45959
rect 1611 45913 1657 45959
rect 1735 45913 1781 45959
rect 1859 45913 1905 45959
rect 1983 45913 2029 45959
rect 2107 45913 2153 45959
rect 2231 45913 2277 45959
rect 2355 45913 2401 45959
rect 2479 45913 2525 45959
rect 2603 45913 2649 45959
rect 2727 45913 2773 45959
rect 2851 45913 2897 45959
rect 2975 45913 3021 45959
rect 3099 45913 3145 45959
rect 3223 45913 3269 45959
rect 3347 45913 3393 45959
rect 3471 45913 3517 45959
rect 3595 45913 3641 45959
rect 3719 45913 3765 45959
rect 3843 45913 3889 45959
rect 3967 45913 4013 45959
rect 4091 45913 4137 45959
rect 4215 45913 4261 45959
rect 4339 45913 4385 45959
rect 4463 45913 4509 45959
rect 4587 45913 4633 45959
rect 4711 45913 4757 45959
rect 4835 45913 4881 45959
rect 4959 45913 5005 45959
rect 5083 45913 5129 45959
rect 5207 45913 5253 45959
rect 5331 45913 5377 45959
rect 5455 45913 5501 45959
rect 5579 45913 5625 45959
rect 5703 45913 5749 45959
rect 5827 45913 5873 45959
rect 5951 45913 5997 45959
rect 6075 45913 6121 45959
rect 6199 45913 6245 45959
rect 6323 45913 6369 45959
rect 6447 45913 6493 45959
rect 6571 45913 6617 45959
rect 6695 45913 6741 45959
rect 6819 45913 6865 45959
rect 6943 45913 6989 45959
rect 7067 45913 7113 45959
rect 7191 45913 7237 45959
rect 7315 45913 7361 45959
rect 7439 45913 7485 45959
rect 7563 45913 7609 45959
rect 7687 45913 7733 45959
rect 7811 45913 7857 45959
rect 7935 45913 7981 45959
rect 8059 45913 8105 45959
rect 8183 45913 8229 45959
rect 8307 45913 8353 45959
rect 8431 45913 8477 45959
rect 8555 45913 8601 45959
rect 8679 45913 8725 45959
rect 8803 45913 8849 45959
rect 8927 45913 8973 45959
rect 9051 45913 9097 45959
rect 9175 45913 9221 45959
rect 9299 45913 9345 45959
rect 9423 45913 9469 45959
rect 9547 45913 9593 45959
rect 9671 45913 9717 45959
rect 9795 45913 9841 45959
rect 9919 45913 9965 45959
rect 10043 45913 10089 45959
rect 10167 45913 10213 45959
rect 10291 45913 10337 45959
rect 10415 45913 10461 45959
rect 10539 45913 10585 45959
rect 10663 45913 10709 45959
rect 10787 45913 10833 45959
rect 10911 45913 10957 45959
rect 11035 45913 11081 45959
rect 11159 45913 11205 45959
rect 11283 45913 11329 45959
rect 11407 45913 11453 45959
rect 11531 45913 11577 45959
rect 11655 45913 11701 45959
rect 11779 45913 11825 45959
rect 11903 45913 11949 45959
rect 12027 45913 12073 45959
rect 12151 45913 12197 45959
rect 12275 45913 12321 45959
rect 12399 45913 12445 45959
rect 12523 45913 12569 45959
rect 12647 45913 12693 45959
rect 12771 45913 12817 45959
rect 12895 45913 12941 45959
rect 13019 45913 13065 45959
rect 13143 45913 13189 45959
rect 13267 45913 13313 45959
rect 13391 45913 13437 45959
rect 13515 45913 13561 45959
rect 13639 45913 13685 45959
rect 13763 45913 13809 45959
rect 13887 45913 13933 45959
rect 14011 45913 14057 45959
rect 14135 45913 14181 45959
rect 14259 45913 14305 45959
rect 14383 45913 14429 45959
rect 14507 45913 14553 45959
rect 14631 45913 14677 45959
rect 14755 45913 14801 45959
rect 14879 45913 14925 45959
rect 15003 45913 15049 45959
rect 15127 45913 15173 45959
rect 15251 45913 15297 45959
rect 15375 45913 15421 45959
rect 15499 45913 15545 45959
rect 15623 45913 15669 45959
rect 15747 45913 15793 45959
rect 15871 45913 15917 45959
rect 15995 45913 16041 45959
rect 16119 45913 16165 45959
rect 16243 45913 16289 45959
rect 16367 45913 16413 45959
rect 16491 45913 16537 45959
rect 16615 45913 16661 45959
rect 16739 45913 16785 45959
rect 16863 45913 16909 45959
rect 16987 45913 17033 45959
rect 17111 45913 17157 45959
rect 17235 45913 17281 45959
rect 17359 45913 17405 45959
rect 17483 45913 17529 45959
rect 17607 45913 17653 45959
rect 17731 45913 17777 45959
rect 17855 45913 17901 45959
rect 17979 45913 18025 45959
rect 18103 45913 18149 45959
rect 18227 45913 18273 45959
rect 18351 45913 18397 45959
rect 18475 45913 18521 45959
rect 18599 45913 18645 45959
rect 18723 45913 18769 45959
rect 18847 45913 18893 45959
rect 18971 45913 19017 45959
rect 19095 45913 19141 45959
rect 19219 45913 19265 45959
rect 19343 45913 19389 45959
rect 19467 45913 19513 45959
rect 19591 45913 19637 45959
rect 19715 45913 19761 45959
rect 19839 45913 19885 45959
rect 19963 45913 20009 45959
rect 20087 45913 20133 45959
rect 20211 45913 20257 45959
rect 20335 45913 20381 45959
rect 20459 45913 20505 45959
rect 20583 45913 20629 45959
rect 20707 45913 20753 45959
rect 20831 45913 20877 45959
rect 20955 45913 21001 45959
rect 21079 45913 21125 45959
rect 21203 45913 21249 45959
rect 21327 45913 21373 45959
rect 21451 45913 21497 45959
rect 21575 45913 21621 45959
rect 21699 45913 21745 45959
rect 21823 45913 21869 45959
rect 21947 45913 21993 45959
rect 22071 45913 22117 45959
rect 22195 45913 22241 45959
rect 22319 45913 22365 45959
rect 22443 45913 22489 45959
rect 22567 45913 22613 45959
rect 22691 45913 22737 45959
rect 22815 45913 22861 45959
rect 22939 45913 22985 45959
rect 23063 45913 23109 45959
rect 23187 45913 23233 45959
rect 23311 45913 23357 45959
rect 23435 45913 23481 45959
rect 23559 45913 23605 45959
rect 23683 45913 23729 45959
rect 23807 45913 23853 45959
rect 23931 45913 23977 45959
rect 24055 45913 24101 45959
rect 24179 45913 24225 45959
rect 24303 45913 24349 45959
rect 24427 45913 24473 45959
rect 24551 45913 24597 45959
rect 24675 45913 24721 45959
rect 24799 45913 24845 45959
rect 24923 45913 24969 45959
rect 25047 45913 25093 45959
rect 25171 45913 25217 45959
rect 25295 45913 25341 45959
rect 25419 45913 25465 45959
rect 25543 45913 25589 45959
rect 25667 45913 25713 45959
rect 25791 45913 25837 45959
rect 25915 45913 25961 45959
rect 26039 45913 26085 45959
rect 26163 45913 26209 45959
rect 26287 45913 26333 45959
rect 26411 45913 26457 45959
rect 26535 45913 26581 45959
rect 26659 45913 26705 45959
rect 26783 45913 26829 45959
rect 26907 45913 26953 45959
rect 27031 45913 27077 45959
rect 27155 45913 27201 45959
rect 27279 45913 27325 45959
rect 27403 45913 27449 45959
rect 27527 45913 27573 45959
rect 27651 45913 27697 45959
rect 27775 45913 27821 45959
rect 27899 45913 27945 45959
rect 28023 45913 28069 45959
rect 28147 45913 28193 45959
rect 28271 45913 28317 45959
rect 28395 45913 28441 45959
rect 28519 45913 28565 45959
rect 28643 45913 28689 45959
rect 28767 45913 28813 45959
rect 28891 45913 28937 45959
rect 29015 45913 29061 45959
rect 29139 45913 29185 45959
rect 29263 45913 29309 45959
rect 29387 45913 29433 45959
rect 29511 45913 29557 45959
rect 29635 45913 29681 45959
rect 29759 45913 29805 45959
rect 29883 45913 29929 45959
rect 30007 45913 30053 45959
rect 30131 45913 30177 45959
rect 30255 45913 30301 45959
rect 30379 45913 30425 45959
rect 30503 45913 30549 45959
rect 30627 45913 30673 45959
rect 30751 45913 30797 45959
rect 30875 45913 30921 45959
rect 30999 45913 31045 45959
rect 31123 45913 31169 45959
rect 31247 45913 31293 45959
rect 31371 45913 31417 45959
rect 31495 45913 31541 45959
rect 31619 45913 31665 45959
rect 31743 45913 31789 45959
rect 31867 45913 31913 45959
rect 31991 45913 32037 45959
rect 32115 45913 32161 45959
rect 32239 45913 32285 45959
rect 32363 45913 32409 45959
rect 32487 45913 32533 45959
rect 32611 45913 32657 45959
rect 32735 45913 32781 45959
rect 32859 45913 32905 45959
rect 32983 45913 33029 45959
rect 33107 45913 33153 45959
rect 33231 45913 33277 45959
rect 33355 45913 33401 45959
rect 33479 45913 33525 45959
rect 33603 45913 33649 45959
rect 33727 45913 33773 45959
rect 33851 45913 33897 45959
rect 33975 45913 34021 45959
rect 34099 45913 34145 45959
rect 34223 45913 34269 45959
rect 34347 45913 34393 45959
rect 34471 45913 34517 45959
rect 34595 45913 34641 45959
rect 34719 45913 34765 45959
rect 34843 45913 34889 45959
rect 34967 45913 35013 45959
rect 35091 45913 35137 45959
rect 35215 45913 35261 45959
rect 35339 45913 35385 45959
rect 35463 45913 35509 45959
rect 35587 45913 35633 45959
rect 35711 45913 35757 45959
rect 35835 45913 35881 45959
rect 35959 45913 36005 45959
rect 36083 45913 36129 45959
rect 36207 45913 36253 45959
rect 36331 45913 36377 45959
rect 36455 45913 36501 45959
rect 36579 45913 36625 45959
rect 36703 45913 36749 45959
rect 36827 45913 36873 45959
rect 36951 45913 36997 45959
rect 37075 45913 37121 45959
rect 37199 45913 37245 45959
rect 37323 45913 37369 45959
rect 37447 45913 37493 45959
rect 37571 45913 37617 45959
rect 37695 45913 37741 45959
rect 37819 45913 37865 45959
rect 37943 45913 37989 45959
rect 38067 45913 38113 45959
rect 38191 45913 38237 45959
rect 38315 45913 38361 45959
rect 38439 45913 38485 45959
rect 38563 45913 38609 45959
rect 38687 45913 38733 45959
rect 38811 45913 38857 45959
rect 38935 45913 38981 45959
rect 39059 45913 39105 45959
rect 39183 45913 39229 45959
rect 39307 45913 39353 45959
rect 39431 45913 39477 45959
rect 39555 45913 39601 45959
rect 39679 45913 39725 45959
rect 39803 45913 39849 45959
rect 39927 45913 39973 45959
rect 40051 45913 40097 45959
rect 40175 45913 40221 45959
rect 40299 45913 40345 45959
rect 40423 45913 40469 45959
rect 40547 45913 40593 45959
rect 40671 45913 40717 45959
rect 40795 45913 40841 45959
rect 40919 45913 40965 45959
rect 41043 45913 41089 45959
rect 41167 45913 41213 45959
rect 41291 45913 41337 45959
rect 41415 45913 41461 45959
rect 41539 45913 41585 45959
rect 41663 45913 41709 45959
rect 41787 45913 41833 45959
rect 41911 45913 41957 45959
rect 42035 45913 42081 45959
rect 42159 45913 42205 45959
rect 42283 45913 42329 45959
rect 42407 45913 42453 45959
rect 42531 45913 42577 45959
rect 42655 45913 42701 45959
rect 42779 45913 42825 45959
rect 42903 45913 42949 45959
rect 43027 45913 43073 45959
rect 43151 45913 43197 45959
rect 43275 45913 43321 45959
rect 43399 45913 43445 45959
rect 43523 45913 43569 45959
rect 43647 45913 43693 45959
rect 43771 45913 43817 45959
rect 43895 45913 43941 45959
rect 44019 45913 44065 45959
rect 44143 45913 44189 45959
rect 44267 45913 44313 45959
rect 44391 45913 44437 45959
rect 44515 45913 44561 45959
rect 44639 45913 44685 45959
rect 44763 45913 44809 45959
rect 44887 45913 44933 45959
rect 45011 45913 45057 45959
rect 45135 45913 45181 45959
rect 45259 45913 45305 45959
rect 45383 45913 45429 45959
rect 45507 45913 45553 45959
rect 45631 45913 45677 45959
rect 45755 45913 45801 45959
rect 45879 45913 45925 45959
rect 46003 45913 46049 45959
rect 46127 45913 46173 45959
rect 46251 45913 46297 45959
rect 46375 45913 46421 45959
rect 46499 45913 46545 45959
rect 46623 45913 46669 45959
rect 46747 45913 46793 45959
rect 46871 45913 46917 45959
rect 46995 45913 47041 45959
rect 47119 45913 47165 45959
rect 47243 45913 47289 45959
rect 47367 45913 47413 45959
rect 47491 45913 47537 45959
rect 47615 45913 47661 45959
rect 47739 45913 47785 45959
rect 47863 45913 47909 45959
rect 47987 45913 48033 45959
rect 48111 45913 48157 45959
rect 48235 45913 48281 45959
rect 48359 45913 48405 45959
rect 48483 45913 48529 45959
rect 48607 45913 48653 45959
rect 48731 45913 48777 45959
rect 48855 45913 48901 45959
rect 48979 45913 49025 45959
rect 49103 45913 49149 45959
rect 49227 45913 49273 45959
rect 49351 45913 49397 45959
rect 49475 45913 49521 45959
rect 49599 45913 49645 45959
rect 49723 45913 49769 45959
rect 49847 45913 49893 45959
rect 49971 45913 50017 45959
rect 50095 45913 50141 45959
rect 50219 45913 50265 45959
rect 50343 45913 50389 45959
rect 50467 45913 50513 45959
rect 50591 45913 50637 45959
rect 50715 45913 50761 45959
rect 50839 45913 50885 45959
rect 50963 45913 51009 45959
rect 51087 45913 51133 45959
rect 51211 45913 51257 45959
rect 51335 45913 51381 45959
rect 51459 45913 51505 45959
rect 51583 45913 51629 45959
rect 51707 45913 51753 45959
rect 51831 45913 51877 45959
rect 51955 45913 52001 45959
rect 52079 45913 52125 45959
rect 52203 45913 52249 45959
rect 52327 45913 52373 45959
rect 52451 45913 52497 45959
rect 52575 45913 52621 45959
rect 52699 45913 52745 45959
rect 52823 45913 52869 45959
rect 52947 45913 52993 45959
rect 53071 45913 53117 45959
rect 53195 45913 53241 45959
rect 53319 45913 53365 45959
rect 53443 45913 53489 45959
rect 53567 45913 53613 45959
rect 53691 45913 53737 45959
rect 53815 45913 53861 45959
rect 53939 45913 53985 45959
rect 54063 45913 54109 45959
rect 54187 45913 54233 45959
rect 54311 45913 54357 45959
rect 54435 45913 54481 45959
rect 54559 45913 54605 45959
rect 54683 45913 54729 45959
rect 54807 45913 54853 45959
rect 54931 45913 54977 45959
rect 55055 45913 55101 45959
rect 55179 45913 55225 45959
rect 55303 45913 55349 45959
rect 55427 45913 55473 45959
rect 55551 45913 55597 45959
rect 55675 45913 55721 45959
rect 55799 45913 55845 45959
rect 55923 45913 55969 45959
rect 56047 45913 56093 45959
rect 56171 45913 56217 45959
rect 56295 45913 56341 45959
rect 56419 45913 56465 45959
rect 56543 45913 56589 45959
rect 56667 45913 56713 45959
rect 56791 45913 56837 45959
rect 56915 45913 56961 45959
rect 57039 45913 57085 45959
rect 57163 45913 57209 45959
rect 57287 45913 57333 45959
rect 57411 45913 57457 45959
rect 57535 45913 57581 45959
rect 57659 45913 57705 45959
rect 57783 45913 57829 45959
rect 57907 45913 57953 45959
rect 58031 45913 58077 45959
rect 58155 45913 58201 45959
rect 58279 45913 58325 45959
rect 58403 45913 58449 45959
rect 58527 45913 58573 45959
rect 58651 45913 58697 45959
rect 58775 45913 58821 45959
rect 58899 45913 58945 45959
rect 59023 45913 59069 45959
rect 59147 45913 59193 45959
rect 59271 45913 59317 45959
rect 59395 45913 59441 45959
rect 59519 45913 59565 45959
rect 59643 45913 59689 45959
rect 59767 45913 59813 45959
rect 59891 45913 59937 45959
rect 60015 45913 60061 45959
rect 60139 45913 60185 45959
rect 60263 45913 60309 45959
rect 60387 45913 60433 45959
rect 60511 45913 60557 45959
rect 60635 45913 60681 45959
rect 60759 45913 60805 45959
rect 60883 45913 60929 45959
rect 61007 45913 61053 45959
rect 61131 45913 61177 45959
rect 61255 45913 61301 45959
rect 61379 45913 61425 45959
rect 61503 45913 61549 45959
rect 61627 45913 61673 45959
rect 61751 45913 61797 45959
rect 61875 45913 61921 45959
rect 61999 45913 62045 45959
rect 62123 45913 62169 45959
rect 62247 45913 62293 45959
rect 62371 45913 62417 45959
rect 62495 45913 62541 45959
rect 62619 45913 62665 45959
rect 62743 45913 62789 45959
rect 62867 45913 62913 45959
rect 62991 45913 63037 45959
rect 63115 45913 63161 45959
rect 63239 45913 63285 45959
rect 63363 45913 63409 45959
rect 63487 45913 63533 45959
rect 63611 45913 63657 45959
rect 63735 45913 63781 45959
rect 63859 45913 63905 45959
rect 63983 45913 64029 45959
rect 64107 45913 64153 45959
rect 64231 45913 64277 45959
rect 64355 45913 64401 45959
rect 64479 45913 64525 45959
rect 64603 45913 64649 45959
rect 64727 45913 64773 45959
rect 64851 45913 64897 45959
rect 64975 45913 65021 45959
rect 65099 45913 65145 45959
rect 65223 45913 65269 45959
rect 65347 45913 65393 45959
rect 65471 45913 65517 45959
rect 65595 45913 65641 45959
rect 65719 45913 65765 45959
rect 65843 45913 65889 45959
rect 65967 45913 66013 45959
rect 66091 45913 66137 45959
rect 66215 45913 66261 45959
rect 66339 45913 66385 45959
rect 66463 45913 66509 45959
rect 66587 45913 66633 45959
rect 66711 45913 66757 45959
rect 66835 45913 66881 45959
rect 66959 45913 67005 45959
rect 67083 45913 67129 45959
rect 67207 45913 67253 45959
rect 67331 45913 67377 45959
rect 67455 45913 67501 45959
rect 67579 45913 67625 45959
rect 67703 45913 67749 45959
rect 67827 45913 67873 45959
rect 67951 45913 67997 45959
rect 68075 45913 68121 45959
rect 68199 45913 68245 45959
rect 68323 45913 68369 45959
rect 68447 45913 68493 45959
rect 68571 45913 68617 45959
rect 68695 45913 68741 45959
rect 68819 45913 68865 45959
rect 68943 45913 68989 45959
rect 69067 45913 69113 45959
rect 69191 45913 69237 45959
rect 69315 45913 69361 45959
rect 69439 45913 69485 45959
rect 69563 45913 69609 45959
rect 69687 45913 69733 45959
rect 69811 45913 69857 45959
rect 69935 45913 69981 45959
rect 70059 45913 70105 45959
rect 70183 45913 70229 45959
rect 70307 45913 70353 45959
rect 70431 45913 70477 45959
rect 70555 45913 70601 45959
rect 70679 45913 70725 45959
rect 70803 45913 70849 45959
rect 70927 45913 70973 45959
rect 71051 45913 71097 45959
rect 71175 45913 71221 45959
rect 71299 45913 71345 45959
rect 71423 45913 71469 45959
rect 71547 45913 71593 45959
rect 71671 45913 71717 45959
rect 71795 45913 71841 45959
rect 71919 45913 71965 45959
rect 72043 45913 72089 45959
rect 72167 45913 72213 45959
rect 72291 45913 72337 45959
rect 72415 45913 72461 45959
rect 72539 45913 72585 45959
rect 72663 45913 72709 45959
rect 72787 45913 72833 45959
rect 72911 45913 72957 45959
rect 73035 45913 73081 45959
rect 73159 45913 73205 45959
rect 73283 45913 73329 45959
rect 73407 45913 73453 45959
rect 73531 45913 73577 45959
rect 73655 45913 73701 45959
rect 73779 45913 73825 45959
rect 73903 45913 73949 45959
rect 74027 45913 74073 45959
rect 74151 45913 74197 45959
rect 74275 45913 74321 45959
rect 74399 45913 74445 45959
rect 74523 45913 74569 45959
rect 74647 45913 74693 45959
rect 74771 45913 74817 45959
rect 74895 45913 74941 45959
rect 75019 45913 75065 45959
rect 75143 45913 75189 45959
rect 75267 45913 75313 45959
rect 75391 45913 75437 45959
rect 75515 45913 75561 45959
rect 75639 45913 75685 45959
rect 75763 45913 75809 45959
rect 75887 45913 75933 45959
rect 76011 45913 76057 45959
rect 76135 45913 76181 45959
rect 76259 45913 76305 45959
rect 76383 45913 76429 45959
rect 76507 45913 76553 45959
rect 76631 45913 76677 45959
rect 76755 45913 76801 45959
rect 76879 45913 76925 45959
rect 77003 45913 77049 45959
rect 77127 45913 77173 45959
rect 77251 45913 77297 45959
rect 77375 45913 77421 45959
rect 77499 45913 77545 45959
rect 77623 45913 77669 45959
rect 77747 45913 77793 45959
rect 77871 45913 77917 45959
rect 77995 45913 78041 45959
rect 78119 45913 78165 45959
rect 78243 45913 78289 45959
rect 78367 45913 78413 45959
rect 78491 45913 78537 45959
rect 78615 45913 78661 45959
rect 78739 45913 78785 45959
rect 78863 45913 78909 45959
rect 78987 45913 79033 45959
rect 79111 45913 79157 45959
rect 79235 45913 79281 45959
rect 79359 45913 79405 45959
rect 79483 45913 79529 45959
rect 79607 45913 79653 45959
rect 79731 45913 79777 45959
rect 79855 45913 79901 45959
rect 79979 45913 80025 45959
rect 80103 45913 80149 45959
rect 80227 45913 80273 45959
rect 80351 45913 80397 45959
rect 80475 45913 80521 45959
rect 80599 45913 80645 45959
rect 80723 45913 80769 45959
rect 80847 45913 80893 45959
rect 80971 45913 81017 45959
rect 81095 45913 81141 45959
rect 81219 45913 81265 45959
rect 81343 45913 81389 45959
rect 81467 45913 81513 45959
rect 81591 45913 81637 45959
rect 81715 45913 81761 45959
rect 81839 45913 81885 45959
rect 81963 45913 82009 45959
rect 82087 45913 82133 45959
rect 82211 45913 82257 45959
rect 82335 45913 82381 45959
rect 82459 45913 82505 45959
rect 82583 45913 82629 45959
rect 82707 45913 82753 45959
rect 82831 45913 82877 45959
rect 82955 45913 83001 45959
rect 83079 45913 83125 45959
rect 83203 45913 83249 45959
rect 83327 45913 83373 45959
rect 83451 45913 83497 45959
rect 83575 45913 83621 45959
rect 83699 45913 83745 45959
rect 83823 45913 83869 45959
rect 83947 45913 83993 45959
rect 84071 45913 84117 45959
rect 84195 45913 84241 45959
rect 84319 45913 84365 45959
rect 84443 45913 84489 45959
rect 84567 45913 84613 45959
rect 84691 45913 84737 45959
rect 84815 45913 84861 45959
rect 84939 45913 84985 45959
rect 85063 45913 85109 45959
rect 85187 45913 85233 45959
rect 85311 45913 85357 45959
rect 85435 45913 85481 45959
rect 85559 45913 85605 45959
rect 85683 45913 85729 45959
rect 85807 45913 85853 45959
rect 85931 45913 85977 45959
rect 371 45789 417 45835
rect 495 45789 541 45835
rect 619 45789 665 45835
rect 743 45789 789 45835
rect 867 45789 913 45835
rect 991 45789 1037 45835
rect 1115 45789 1161 45835
rect 1239 45789 1285 45835
rect 1363 45789 1409 45835
rect 1487 45789 1533 45835
rect 1611 45789 1657 45835
rect 1735 45789 1781 45835
rect 1859 45789 1905 45835
rect 1983 45789 2029 45835
rect 2107 45789 2153 45835
rect 2231 45789 2277 45835
rect 2355 45789 2401 45835
rect 2479 45789 2525 45835
rect 2603 45789 2649 45835
rect 2727 45789 2773 45835
rect 2851 45789 2897 45835
rect 2975 45789 3021 45835
rect 3099 45789 3145 45835
rect 3223 45789 3269 45835
rect 3347 45789 3393 45835
rect 3471 45789 3517 45835
rect 3595 45789 3641 45835
rect 3719 45789 3765 45835
rect 3843 45789 3889 45835
rect 3967 45789 4013 45835
rect 4091 45789 4137 45835
rect 4215 45789 4261 45835
rect 4339 45789 4385 45835
rect 4463 45789 4509 45835
rect 4587 45789 4633 45835
rect 4711 45789 4757 45835
rect 4835 45789 4881 45835
rect 4959 45789 5005 45835
rect 5083 45789 5129 45835
rect 5207 45789 5253 45835
rect 5331 45789 5377 45835
rect 5455 45789 5501 45835
rect 5579 45789 5625 45835
rect 5703 45789 5749 45835
rect 5827 45789 5873 45835
rect 5951 45789 5997 45835
rect 6075 45789 6121 45835
rect 6199 45789 6245 45835
rect 6323 45789 6369 45835
rect 6447 45789 6493 45835
rect 6571 45789 6617 45835
rect 6695 45789 6741 45835
rect 6819 45789 6865 45835
rect 6943 45789 6989 45835
rect 7067 45789 7113 45835
rect 7191 45789 7237 45835
rect 7315 45789 7361 45835
rect 7439 45789 7485 45835
rect 7563 45789 7609 45835
rect 7687 45789 7733 45835
rect 7811 45789 7857 45835
rect 7935 45789 7981 45835
rect 8059 45789 8105 45835
rect 8183 45789 8229 45835
rect 8307 45789 8353 45835
rect 8431 45789 8477 45835
rect 8555 45789 8601 45835
rect 8679 45789 8725 45835
rect 8803 45789 8849 45835
rect 8927 45789 8973 45835
rect 9051 45789 9097 45835
rect 9175 45789 9221 45835
rect 9299 45789 9345 45835
rect 9423 45789 9469 45835
rect 9547 45789 9593 45835
rect 9671 45789 9717 45835
rect 9795 45789 9841 45835
rect 9919 45789 9965 45835
rect 10043 45789 10089 45835
rect 10167 45789 10213 45835
rect 10291 45789 10337 45835
rect 10415 45789 10461 45835
rect 10539 45789 10585 45835
rect 10663 45789 10709 45835
rect 10787 45789 10833 45835
rect 10911 45789 10957 45835
rect 11035 45789 11081 45835
rect 11159 45789 11205 45835
rect 11283 45789 11329 45835
rect 11407 45789 11453 45835
rect 11531 45789 11577 45835
rect 11655 45789 11701 45835
rect 11779 45789 11825 45835
rect 11903 45789 11949 45835
rect 12027 45789 12073 45835
rect 12151 45789 12197 45835
rect 12275 45789 12321 45835
rect 12399 45789 12445 45835
rect 12523 45789 12569 45835
rect 12647 45789 12693 45835
rect 12771 45789 12817 45835
rect 12895 45789 12941 45835
rect 13019 45789 13065 45835
rect 13143 45789 13189 45835
rect 13267 45789 13313 45835
rect 13391 45789 13437 45835
rect 13515 45789 13561 45835
rect 13639 45789 13685 45835
rect 13763 45789 13809 45835
rect 13887 45789 13933 45835
rect 14011 45789 14057 45835
rect 14135 45789 14181 45835
rect 14259 45789 14305 45835
rect 14383 45789 14429 45835
rect 14507 45789 14553 45835
rect 14631 45789 14677 45835
rect 14755 45789 14801 45835
rect 14879 45789 14925 45835
rect 15003 45789 15049 45835
rect 15127 45789 15173 45835
rect 15251 45789 15297 45835
rect 15375 45789 15421 45835
rect 15499 45789 15545 45835
rect 15623 45789 15669 45835
rect 15747 45789 15793 45835
rect 15871 45789 15917 45835
rect 15995 45789 16041 45835
rect 16119 45789 16165 45835
rect 16243 45789 16289 45835
rect 16367 45789 16413 45835
rect 16491 45789 16537 45835
rect 16615 45789 16661 45835
rect 16739 45789 16785 45835
rect 16863 45789 16909 45835
rect 16987 45789 17033 45835
rect 17111 45789 17157 45835
rect 17235 45789 17281 45835
rect 17359 45789 17405 45835
rect 17483 45789 17529 45835
rect 17607 45789 17653 45835
rect 17731 45789 17777 45835
rect 17855 45789 17901 45835
rect 17979 45789 18025 45835
rect 18103 45789 18149 45835
rect 18227 45789 18273 45835
rect 18351 45789 18397 45835
rect 18475 45789 18521 45835
rect 18599 45789 18645 45835
rect 18723 45789 18769 45835
rect 18847 45789 18893 45835
rect 18971 45789 19017 45835
rect 19095 45789 19141 45835
rect 19219 45789 19265 45835
rect 19343 45789 19389 45835
rect 19467 45789 19513 45835
rect 19591 45789 19637 45835
rect 19715 45789 19761 45835
rect 19839 45789 19885 45835
rect 19963 45789 20009 45835
rect 20087 45789 20133 45835
rect 20211 45789 20257 45835
rect 20335 45789 20381 45835
rect 20459 45789 20505 45835
rect 20583 45789 20629 45835
rect 20707 45789 20753 45835
rect 20831 45789 20877 45835
rect 20955 45789 21001 45835
rect 21079 45789 21125 45835
rect 21203 45789 21249 45835
rect 21327 45789 21373 45835
rect 21451 45789 21497 45835
rect 21575 45789 21621 45835
rect 21699 45789 21745 45835
rect 21823 45789 21869 45835
rect 21947 45789 21993 45835
rect 22071 45789 22117 45835
rect 22195 45789 22241 45835
rect 22319 45789 22365 45835
rect 22443 45789 22489 45835
rect 22567 45789 22613 45835
rect 22691 45789 22737 45835
rect 22815 45789 22861 45835
rect 22939 45789 22985 45835
rect 23063 45789 23109 45835
rect 23187 45789 23233 45835
rect 23311 45789 23357 45835
rect 23435 45789 23481 45835
rect 23559 45789 23605 45835
rect 23683 45789 23729 45835
rect 23807 45789 23853 45835
rect 23931 45789 23977 45835
rect 24055 45789 24101 45835
rect 24179 45789 24225 45835
rect 24303 45789 24349 45835
rect 24427 45789 24473 45835
rect 24551 45789 24597 45835
rect 24675 45789 24721 45835
rect 24799 45789 24845 45835
rect 24923 45789 24969 45835
rect 25047 45789 25093 45835
rect 25171 45789 25217 45835
rect 25295 45789 25341 45835
rect 25419 45789 25465 45835
rect 25543 45789 25589 45835
rect 25667 45789 25713 45835
rect 25791 45789 25837 45835
rect 25915 45789 25961 45835
rect 26039 45789 26085 45835
rect 26163 45789 26209 45835
rect 26287 45789 26333 45835
rect 26411 45789 26457 45835
rect 26535 45789 26581 45835
rect 26659 45789 26705 45835
rect 26783 45789 26829 45835
rect 26907 45789 26953 45835
rect 27031 45789 27077 45835
rect 27155 45789 27201 45835
rect 27279 45789 27325 45835
rect 27403 45789 27449 45835
rect 27527 45789 27573 45835
rect 27651 45789 27697 45835
rect 27775 45789 27821 45835
rect 27899 45789 27945 45835
rect 28023 45789 28069 45835
rect 28147 45789 28193 45835
rect 28271 45789 28317 45835
rect 28395 45789 28441 45835
rect 28519 45789 28565 45835
rect 28643 45789 28689 45835
rect 28767 45789 28813 45835
rect 28891 45789 28937 45835
rect 29015 45789 29061 45835
rect 29139 45789 29185 45835
rect 29263 45789 29309 45835
rect 29387 45789 29433 45835
rect 29511 45789 29557 45835
rect 29635 45789 29681 45835
rect 29759 45789 29805 45835
rect 29883 45789 29929 45835
rect 30007 45789 30053 45835
rect 30131 45789 30177 45835
rect 30255 45789 30301 45835
rect 30379 45789 30425 45835
rect 30503 45789 30549 45835
rect 30627 45789 30673 45835
rect 30751 45789 30797 45835
rect 30875 45789 30921 45835
rect 30999 45789 31045 45835
rect 31123 45789 31169 45835
rect 31247 45789 31293 45835
rect 31371 45789 31417 45835
rect 31495 45789 31541 45835
rect 31619 45789 31665 45835
rect 31743 45789 31789 45835
rect 31867 45789 31913 45835
rect 31991 45789 32037 45835
rect 32115 45789 32161 45835
rect 32239 45789 32285 45835
rect 32363 45789 32409 45835
rect 32487 45789 32533 45835
rect 32611 45789 32657 45835
rect 32735 45789 32781 45835
rect 32859 45789 32905 45835
rect 32983 45789 33029 45835
rect 33107 45789 33153 45835
rect 33231 45789 33277 45835
rect 33355 45789 33401 45835
rect 33479 45789 33525 45835
rect 33603 45789 33649 45835
rect 33727 45789 33773 45835
rect 33851 45789 33897 45835
rect 33975 45789 34021 45835
rect 34099 45789 34145 45835
rect 34223 45789 34269 45835
rect 34347 45789 34393 45835
rect 34471 45789 34517 45835
rect 34595 45789 34641 45835
rect 34719 45789 34765 45835
rect 34843 45789 34889 45835
rect 34967 45789 35013 45835
rect 35091 45789 35137 45835
rect 35215 45789 35261 45835
rect 35339 45789 35385 45835
rect 35463 45789 35509 45835
rect 35587 45789 35633 45835
rect 35711 45789 35757 45835
rect 35835 45789 35881 45835
rect 35959 45789 36005 45835
rect 36083 45789 36129 45835
rect 36207 45789 36253 45835
rect 36331 45789 36377 45835
rect 36455 45789 36501 45835
rect 36579 45789 36625 45835
rect 36703 45789 36749 45835
rect 36827 45789 36873 45835
rect 36951 45789 36997 45835
rect 37075 45789 37121 45835
rect 37199 45789 37245 45835
rect 37323 45789 37369 45835
rect 37447 45789 37493 45835
rect 37571 45789 37617 45835
rect 37695 45789 37741 45835
rect 37819 45789 37865 45835
rect 37943 45789 37989 45835
rect 38067 45789 38113 45835
rect 38191 45789 38237 45835
rect 38315 45789 38361 45835
rect 38439 45789 38485 45835
rect 38563 45789 38609 45835
rect 38687 45789 38733 45835
rect 38811 45789 38857 45835
rect 38935 45789 38981 45835
rect 39059 45789 39105 45835
rect 39183 45789 39229 45835
rect 39307 45789 39353 45835
rect 39431 45789 39477 45835
rect 39555 45789 39601 45835
rect 39679 45789 39725 45835
rect 39803 45789 39849 45835
rect 39927 45789 39973 45835
rect 40051 45789 40097 45835
rect 40175 45789 40221 45835
rect 40299 45789 40345 45835
rect 40423 45789 40469 45835
rect 40547 45789 40593 45835
rect 40671 45789 40717 45835
rect 40795 45789 40841 45835
rect 40919 45789 40965 45835
rect 41043 45789 41089 45835
rect 41167 45789 41213 45835
rect 41291 45789 41337 45835
rect 41415 45789 41461 45835
rect 41539 45789 41585 45835
rect 41663 45789 41709 45835
rect 41787 45789 41833 45835
rect 41911 45789 41957 45835
rect 42035 45789 42081 45835
rect 42159 45789 42205 45835
rect 42283 45789 42329 45835
rect 42407 45789 42453 45835
rect 42531 45789 42577 45835
rect 42655 45789 42701 45835
rect 42779 45789 42825 45835
rect 42903 45789 42949 45835
rect 43027 45789 43073 45835
rect 43151 45789 43197 45835
rect 43275 45789 43321 45835
rect 43399 45789 43445 45835
rect 43523 45789 43569 45835
rect 43647 45789 43693 45835
rect 43771 45789 43817 45835
rect 43895 45789 43941 45835
rect 44019 45789 44065 45835
rect 44143 45789 44189 45835
rect 44267 45789 44313 45835
rect 44391 45789 44437 45835
rect 44515 45789 44561 45835
rect 44639 45789 44685 45835
rect 44763 45789 44809 45835
rect 44887 45789 44933 45835
rect 45011 45789 45057 45835
rect 45135 45789 45181 45835
rect 45259 45789 45305 45835
rect 45383 45789 45429 45835
rect 45507 45789 45553 45835
rect 45631 45789 45677 45835
rect 45755 45789 45801 45835
rect 45879 45789 45925 45835
rect 46003 45789 46049 45835
rect 46127 45789 46173 45835
rect 46251 45789 46297 45835
rect 46375 45789 46421 45835
rect 46499 45789 46545 45835
rect 46623 45789 46669 45835
rect 46747 45789 46793 45835
rect 46871 45789 46917 45835
rect 46995 45789 47041 45835
rect 47119 45789 47165 45835
rect 47243 45789 47289 45835
rect 47367 45789 47413 45835
rect 47491 45789 47537 45835
rect 47615 45789 47661 45835
rect 47739 45789 47785 45835
rect 47863 45789 47909 45835
rect 47987 45789 48033 45835
rect 48111 45789 48157 45835
rect 48235 45789 48281 45835
rect 48359 45789 48405 45835
rect 48483 45789 48529 45835
rect 48607 45789 48653 45835
rect 48731 45789 48777 45835
rect 48855 45789 48901 45835
rect 48979 45789 49025 45835
rect 49103 45789 49149 45835
rect 49227 45789 49273 45835
rect 49351 45789 49397 45835
rect 49475 45789 49521 45835
rect 49599 45789 49645 45835
rect 49723 45789 49769 45835
rect 49847 45789 49893 45835
rect 49971 45789 50017 45835
rect 50095 45789 50141 45835
rect 50219 45789 50265 45835
rect 50343 45789 50389 45835
rect 50467 45789 50513 45835
rect 50591 45789 50637 45835
rect 50715 45789 50761 45835
rect 50839 45789 50885 45835
rect 50963 45789 51009 45835
rect 51087 45789 51133 45835
rect 51211 45789 51257 45835
rect 51335 45789 51381 45835
rect 51459 45789 51505 45835
rect 51583 45789 51629 45835
rect 51707 45789 51753 45835
rect 51831 45789 51877 45835
rect 51955 45789 52001 45835
rect 52079 45789 52125 45835
rect 52203 45789 52249 45835
rect 52327 45789 52373 45835
rect 52451 45789 52497 45835
rect 52575 45789 52621 45835
rect 52699 45789 52745 45835
rect 52823 45789 52869 45835
rect 52947 45789 52993 45835
rect 53071 45789 53117 45835
rect 53195 45789 53241 45835
rect 53319 45789 53365 45835
rect 53443 45789 53489 45835
rect 53567 45789 53613 45835
rect 53691 45789 53737 45835
rect 53815 45789 53861 45835
rect 53939 45789 53985 45835
rect 54063 45789 54109 45835
rect 54187 45789 54233 45835
rect 54311 45789 54357 45835
rect 54435 45789 54481 45835
rect 54559 45789 54605 45835
rect 54683 45789 54729 45835
rect 54807 45789 54853 45835
rect 54931 45789 54977 45835
rect 55055 45789 55101 45835
rect 55179 45789 55225 45835
rect 55303 45789 55349 45835
rect 55427 45789 55473 45835
rect 55551 45789 55597 45835
rect 55675 45789 55721 45835
rect 55799 45789 55845 45835
rect 55923 45789 55969 45835
rect 56047 45789 56093 45835
rect 56171 45789 56217 45835
rect 56295 45789 56341 45835
rect 56419 45789 56465 45835
rect 56543 45789 56589 45835
rect 56667 45789 56713 45835
rect 56791 45789 56837 45835
rect 56915 45789 56961 45835
rect 57039 45789 57085 45835
rect 57163 45789 57209 45835
rect 57287 45789 57333 45835
rect 57411 45789 57457 45835
rect 57535 45789 57581 45835
rect 57659 45789 57705 45835
rect 57783 45789 57829 45835
rect 57907 45789 57953 45835
rect 58031 45789 58077 45835
rect 58155 45789 58201 45835
rect 58279 45789 58325 45835
rect 58403 45789 58449 45835
rect 58527 45789 58573 45835
rect 58651 45789 58697 45835
rect 58775 45789 58821 45835
rect 58899 45789 58945 45835
rect 59023 45789 59069 45835
rect 59147 45789 59193 45835
rect 59271 45789 59317 45835
rect 59395 45789 59441 45835
rect 59519 45789 59565 45835
rect 59643 45789 59689 45835
rect 59767 45789 59813 45835
rect 59891 45789 59937 45835
rect 60015 45789 60061 45835
rect 60139 45789 60185 45835
rect 60263 45789 60309 45835
rect 60387 45789 60433 45835
rect 60511 45789 60557 45835
rect 60635 45789 60681 45835
rect 60759 45789 60805 45835
rect 60883 45789 60929 45835
rect 61007 45789 61053 45835
rect 61131 45789 61177 45835
rect 61255 45789 61301 45835
rect 61379 45789 61425 45835
rect 61503 45789 61549 45835
rect 61627 45789 61673 45835
rect 61751 45789 61797 45835
rect 61875 45789 61921 45835
rect 61999 45789 62045 45835
rect 62123 45789 62169 45835
rect 62247 45789 62293 45835
rect 62371 45789 62417 45835
rect 62495 45789 62541 45835
rect 62619 45789 62665 45835
rect 62743 45789 62789 45835
rect 62867 45789 62913 45835
rect 62991 45789 63037 45835
rect 63115 45789 63161 45835
rect 63239 45789 63285 45835
rect 63363 45789 63409 45835
rect 63487 45789 63533 45835
rect 63611 45789 63657 45835
rect 63735 45789 63781 45835
rect 63859 45789 63905 45835
rect 63983 45789 64029 45835
rect 64107 45789 64153 45835
rect 64231 45789 64277 45835
rect 64355 45789 64401 45835
rect 64479 45789 64525 45835
rect 64603 45789 64649 45835
rect 64727 45789 64773 45835
rect 64851 45789 64897 45835
rect 64975 45789 65021 45835
rect 65099 45789 65145 45835
rect 65223 45789 65269 45835
rect 65347 45789 65393 45835
rect 65471 45789 65517 45835
rect 65595 45789 65641 45835
rect 65719 45789 65765 45835
rect 65843 45789 65889 45835
rect 65967 45789 66013 45835
rect 66091 45789 66137 45835
rect 66215 45789 66261 45835
rect 66339 45789 66385 45835
rect 66463 45789 66509 45835
rect 66587 45789 66633 45835
rect 66711 45789 66757 45835
rect 66835 45789 66881 45835
rect 66959 45789 67005 45835
rect 67083 45789 67129 45835
rect 67207 45789 67253 45835
rect 67331 45789 67377 45835
rect 67455 45789 67501 45835
rect 67579 45789 67625 45835
rect 67703 45789 67749 45835
rect 67827 45789 67873 45835
rect 67951 45789 67997 45835
rect 68075 45789 68121 45835
rect 68199 45789 68245 45835
rect 68323 45789 68369 45835
rect 68447 45789 68493 45835
rect 68571 45789 68617 45835
rect 68695 45789 68741 45835
rect 68819 45789 68865 45835
rect 68943 45789 68989 45835
rect 69067 45789 69113 45835
rect 69191 45789 69237 45835
rect 69315 45789 69361 45835
rect 69439 45789 69485 45835
rect 69563 45789 69609 45835
rect 69687 45789 69733 45835
rect 69811 45789 69857 45835
rect 69935 45789 69981 45835
rect 70059 45789 70105 45835
rect 70183 45789 70229 45835
rect 70307 45789 70353 45835
rect 70431 45789 70477 45835
rect 70555 45789 70601 45835
rect 70679 45789 70725 45835
rect 70803 45789 70849 45835
rect 70927 45789 70973 45835
rect 71051 45789 71097 45835
rect 71175 45789 71221 45835
rect 71299 45789 71345 45835
rect 71423 45789 71469 45835
rect 71547 45789 71593 45835
rect 71671 45789 71717 45835
rect 71795 45789 71841 45835
rect 71919 45789 71965 45835
rect 72043 45789 72089 45835
rect 72167 45789 72213 45835
rect 72291 45789 72337 45835
rect 72415 45789 72461 45835
rect 72539 45789 72585 45835
rect 72663 45789 72709 45835
rect 72787 45789 72833 45835
rect 72911 45789 72957 45835
rect 73035 45789 73081 45835
rect 73159 45789 73205 45835
rect 73283 45789 73329 45835
rect 73407 45789 73453 45835
rect 73531 45789 73577 45835
rect 73655 45789 73701 45835
rect 73779 45789 73825 45835
rect 73903 45789 73949 45835
rect 74027 45789 74073 45835
rect 74151 45789 74197 45835
rect 74275 45789 74321 45835
rect 74399 45789 74445 45835
rect 74523 45789 74569 45835
rect 74647 45789 74693 45835
rect 74771 45789 74817 45835
rect 74895 45789 74941 45835
rect 75019 45789 75065 45835
rect 75143 45789 75189 45835
rect 75267 45789 75313 45835
rect 75391 45789 75437 45835
rect 75515 45789 75561 45835
rect 75639 45789 75685 45835
rect 75763 45789 75809 45835
rect 75887 45789 75933 45835
rect 76011 45789 76057 45835
rect 76135 45789 76181 45835
rect 76259 45789 76305 45835
rect 76383 45789 76429 45835
rect 76507 45789 76553 45835
rect 76631 45789 76677 45835
rect 76755 45789 76801 45835
rect 76879 45789 76925 45835
rect 77003 45789 77049 45835
rect 77127 45789 77173 45835
rect 77251 45789 77297 45835
rect 77375 45789 77421 45835
rect 77499 45789 77545 45835
rect 77623 45789 77669 45835
rect 77747 45789 77793 45835
rect 77871 45789 77917 45835
rect 77995 45789 78041 45835
rect 78119 45789 78165 45835
rect 78243 45789 78289 45835
rect 78367 45789 78413 45835
rect 78491 45789 78537 45835
rect 78615 45789 78661 45835
rect 78739 45789 78785 45835
rect 78863 45789 78909 45835
rect 78987 45789 79033 45835
rect 79111 45789 79157 45835
rect 79235 45789 79281 45835
rect 79359 45789 79405 45835
rect 79483 45789 79529 45835
rect 79607 45789 79653 45835
rect 79731 45789 79777 45835
rect 79855 45789 79901 45835
rect 79979 45789 80025 45835
rect 80103 45789 80149 45835
rect 80227 45789 80273 45835
rect 80351 45789 80397 45835
rect 80475 45789 80521 45835
rect 80599 45789 80645 45835
rect 80723 45789 80769 45835
rect 80847 45789 80893 45835
rect 80971 45789 81017 45835
rect 81095 45789 81141 45835
rect 81219 45789 81265 45835
rect 81343 45789 81389 45835
rect 81467 45789 81513 45835
rect 81591 45789 81637 45835
rect 81715 45789 81761 45835
rect 81839 45789 81885 45835
rect 81963 45789 82009 45835
rect 82087 45789 82133 45835
rect 82211 45789 82257 45835
rect 82335 45789 82381 45835
rect 82459 45789 82505 45835
rect 82583 45789 82629 45835
rect 82707 45789 82753 45835
rect 82831 45789 82877 45835
rect 82955 45789 83001 45835
rect 83079 45789 83125 45835
rect 83203 45789 83249 45835
rect 83327 45789 83373 45835
rect 83451 45789 83497 45835
rect 83575 45789 83621 45835
rect 83699 45789 83745 45835
rect 83823 45789 83869 45835
rect 83947 45789 83993 45835
rect 84071 45789 84117 45835
rect 84195 45789 84241 45835
rect 84319 45789 84365 45835
rect 84443 45789 84489 45835
rect 84567 45789 84613 45835
rect 84691 45789 84737 45835
rect 84815 45789 84861 45835
rect 84939 45789 84985 45835
rect 85063 45789 85109 45835
rect 85187 45789 85233 45835
rect 85311 45789 85357 45835
rect 85435 45789 85481 45835
rect 85559 45789 85605 45835
rect 85683 45789 85729 45835
rect 85807 45789 85853 45835
rect 85931 45789 85977 45835
rect 371 45665 417 45711
rect 495 45665 541 45711
rect 619 45665 665 45711
rect 743 45665 789 45711
rect 867 45665 913 45711
rect 991 45665 1037 45711
rect 1115 45665 1161 45711
rect 1239 45665 1285 45711
rect 1363 45665 1409 45711
rect 1487 45665 1533 45711
rect 1611 45665 1657 45711
rect 1735 45665 1781 45711
rect 1859 45665 1905 45711
rect 1983 45665 2029 45711
rect 2107 45665 2153 45711
rect 2231 45665 2277 45711
rect 2355 45665 2401 45711
rect 2479 45665 2525 45711
rect 2603 45665 2649 45711
rect 2727 45665 2773 45711
rect 2851 45665 2897 45711
rect 2975 45665 3021 45711
rect 3099 45665 3145 45711
rect 3223 45665 3269 45711
rect 3347 45665 3393 45711
rect 3471 45665 3517 45711
rect 3595 45665 3641 45711
rect 3719 45665 3765 45711
rect 3843 45665 3889 45711
rect 3967 45665 4013 45711
rect 4091 45665 4137 45711
rect 4215 45665 4261 45711
rect 4339 45665 4385 45711
rect 4463 45665 4509 45711
rect 4587 45665 4633 45711
rect 4711 45665 4757 45711
rect 4835 45665 4881 45711
rect 4959 45665 5005 45711
rect 5083 45665 5129 45711
rect 5207 45665 5253 45711
rect 5331 45665 5377 45711
rect 5455 45665 5501 45711
rect 5579 45665 5625 45711
rect 5703 45665 5749 45711
rect 5827 45665 5873 45711
rect 5951 45665 5997 45711
rect 6075 45665 6121 45711
rect 6199 45665 6245 45711
rect 6323 45665 6369 45711
rect 6447 45665 6493 45711
rect 6571 45665 6617 45711
rect 6695 45665 6741 45711
rect 6819 45665 6865 45711
rect 6943 45665 6989 45711
rect 7067 45665 7113 45711
rect 7191 45665 7237 45711
rect 7315 45665 7361 45711
rect 7439 45665 7485 45711
rect 7563 45665 7609 45711
rect 7687 45665 7733 45711
rect 7811 45665 7857 45711
rect 7935 45665 7981 45711
rect 8059 45665 8105 45711
rect 8183 45665 8229 45711
rect 8307 45665 8353 45711
rect 8431 45665 8477 45711
rect 8555 45665 8601 45711
rect 8679 45665 8725 45711
rect 8803 45665 8849 45711
rect 8927 45665 8973 45711
rect 9051 45665 9097 45711
rect 9175 45665 9221 45711
rect 9299 45665 9345 45711
rect 9423 45665 9469 45711
rect 9547 45665 9593 45711
rect 9671 45665 9717 45711
rect 9795 45665 9841 45711
rect 9919 45665 9965 45711
rect 10043 45665 10089 45711
rect 10167 45665 10213 45711
rect 10291 45665 10337 45711
rect 10415 45665 10461 45711
rect 10539 45665 10585 45711
rect 10663 45665 10709 45711
rect 10787 45665 10833 45711
rect 10911 45665 10957 45711
rect 11035 45665 11081 45711
rect 11159 45665 11205 45711
rect 11283 45665 11329 45711
rect 11407 45665 11453 45711
rect 11531 45665 11577 45711
rect 11655 45665 11701 45711
rect 11779 45665 11825 45711
rect 11903 45665 11949 45711
rect 12027 45665 12073 45711
rect 12151 45665 12197 45711
rect 12275 45665 12321 45711
rect 12399 45665 12445 45711
rect 12523 45665 12569 45711
rect 12647 45665 12693 45711
rect 12771 45665 12817 45711
rect 12895 45665 12941 45711
rect 13019 45665 13065 45711
rect 13143 45665 13189 45711
rect 13267 45665 13313 45711
rect 13391 45665 13437 45711
rect 13515 45665 13561 45711
rect 13639 45665 13685 45711
rect 13763 45665 13809 45711
rect 13887 45665 13933 45711
rect 14011 45665 14057 45711
rect 14135 45665 14181 45711
rect 14259 45665 14305 45711
rect 14383 45665 14429 45711
rect 14507 45665 14553 45711
rect 14631 45665 14677 45711
rect 14755 45665 14801 45711
rect 14879 45665 14925 45711
rect 15003 45665 15049 45711
rect 15127 45665 15173 45711
rect 15251 45665 15297 45711
rect 15375 45665 15421 45711
rect 15499 45665 15545 45711
rect 15623 45665 15669 45711
rect 15747 45665 15793 45711
rect 15871 45665 15917 45711
rect 15995 45665 16041 45711
rect 16119 45665 16165 45711
rect 16243 45665 16289 45711
rect 16367 45665 16413 45711
rect 16491 45665 16537 45711
rect 16615 45665 16661 45711
rect 16739 45665 16785 45711
rect 16863 45665 16909 45711
rect 16987 45665 17033 45711
rect 17111 45665 17157 45711
rect 17235 45665 17281 45711
rect 17359 45665 17405 45711
rect 17483 45665 17529 45711
rect 17607 45665 17653 45711
rect 17731 45665 17777 45711
rect 17855 45665 17901 45711
rect 17979 45665 18025 45711
rect 18103 45665 18149 45711
rect 18227 45665 18273 45711
rect 18351 45665 18397 45711
rect 18475 45665 18521 45711
rect 18599 45665 18645 45711
rect 18723 45665 18769 45711
rect 18847 45665 18893 45711
rect 18971 45665 19017 45711
rect 19095 45665 19141 45711
rect 19219 45665 19265 45711
rect 19343 45665 19389 45711
rect 19467 45665 19513 45711
rect 19591 45665 19637 45711
rect 19715 45665 19761 45711
rect 19839 45665 19885 45711
rect 19963 45665 20009 45711
rect 20087 45665 20133 45711
rect 20211 45665 20257 45711
rect 20335 45665 20381 45711
rect 20459 45665 20505 45711
rect 20583 45665 20629 45711
rect 20707 45665 20753 45711
rect 20831 45665 20877 45711
rect 20955 45665 21001 45711
rect 21079 45665 21125 45711
rect 21203 45665 21249 45711
rect 21327 45665 21373 45711
rect 21451 45665 21497 45711
rect 21575 45665 21621 45711
rect 21699 45665 21745 45711
rect 21823 45665 21869 45711
rect 21947 45665 21993 45711
rect 22071 45665 22117 45711
rect 22195 45665 22241 45711
rect 22319 45665 22365 45711
rect 22443 45665 22489 45711
rect 22567 45665 22613 45711
rect 22691 45665 22737 45711
rect 22815 45665 22861 45711
rect 22939 45665 22985 45711
rect 23063 45665 23109 45711
rect 23187 45665 23233 45711
rect 23311 45665 23357 45711
rect 23435 45665 23481 45711
rect 23559 45665 23605 45711
rect 23683 45665 23729 45711
rect 23807 45665 23853 45711
rect 23931 45665 23977 45711
rect 24055 45665 24101 45711
rect 24179 45665 24225 45711
rect 24303 45665 24349 45711
rect 24427 45665 24473 45711
rect 24551 45665 24597 45711
rect 24675 45665 24721 45711
rect 24799 45665 24845 45711
rect 24923 45665 24969 45711
rect 25047 45665 25093 45711
rect 25171 45665 25217 45711
rect 25295 45665 25341 45711
rect 25419 45665 25465 45711
rect 25543 45665 25589 45711
rect 25667 45665 25713 45711
rect 25791 45665 25837 45711
rect 25915 45665 25961 45711
rect 26039 45665 26085 45711
rect 26163 45665 26209 45711
rect 26287 45665 26333 45711
rect 26411 45665 26457 45711
rect 26535 45665 26581 45711
rect 26659 45665 26705 45711
rect 26783 45665 26829 45711
rect 26907 45665 26953 45711
rect 27031 45665 27077 45711
rect 27155 45665 27201 45711
rect 27279 45665 27325 45711
rect 27403 45665 27449 45711
rect 27527 45665 27573 45711
rect 27651 45665 27697 45711
rect 27775 45665 27821 45711
rect 27899 45665 27945 45711
rect 28023 45665 28069 45711
rect 28147 45665 28193 45711
rect 28271 45665 28317 45711
rect 28395 45665 28441 45711
rect 28519 45665 28565 45711
rect 28643 45665 28689 45711
rect 28767 45665 28813 45711
rect 28891 45665 28937 45711
rect 29015 45665 29061 45711
rect 29139 45665 29185 45711
rect 29263 45665 29309 45711
rect 29387 45665 29433 45711
rect 29511 45665 29557 45711
rect 29635 45665 29681 45711
rect 29759 45665 29805 45711
rect 29883 45665 29929 45711
rect 30007 45665 30053 45711
rect 30131 45665 30177 45711
rect 30255 45665 30301 45711
rect 30379 45665 30425 45711
rect 30503 45665 30549 45711
rect 30627 45665 30673 45711
rect 30751 45665 30797 45711
rect 30875 45665 30921 45711
rect 30999 45665 31045 45711
rect 31123 45665 31169 45711
rect 31247 45665 31293 45711
rect 31371 45665 31417 45711
rect 31495 45665 31541 45711
rect 31619 45665 31665 45711
rect 31743 45665 31789 45711
rect 31867 45665 31913 45711
rect 31991 45665 32037 45711
rect 32115 45665 32161 45711
rect 32239 45665 32285 45711
rect 32363 45665 32409 45711
rect 32487 45665 32533 45711
rect 32611 45665 32657 45711
rect 32735 45665 32781 45711
rect 32859 45665 32905 45711
rect 32983 45665 33029 45711
rect 33107 45665 33153 45711
rect 33231 45665 33277 45711
rect 33355 45665 33401 45711
rect 33479 45665 33525 45711
rect 33603 45665 33649 45711
rect 33727 45665 33773 45711
rect 33851 45665 33897 45711
rect 33975 45665 34021 45711
rect 34099 45665 34145 45711
rect 34223 45665 34269 45711
rect 34347 45665 34393 45711
rect 34471 45665 34517 45711
rect 34595 45665 34641 45711
rect 34719 45665 34765 45711
rect 34843 45665 34889 45711
rect 34967 45665 35013 45711
rect 35091 45665 35137 45711
rect 35215 45665 35261 45711
rect 35339 45665 35385 45711
rect 35463 45665 35509 45711
rect 35587 45665 35633 45711
rect 35711 45665 35757 45711
rect 35835 45665 35881 45711
rect 35959 45665 36005 45711
rect 36083 45665 36129 45711
rect 36207 45665 36253 45711
rect 36331 45665 36377 45711
rect 36455 45665 36501 45711
rect 36579 45665 36625 45711
rect 36703 45665 36749 45711
rect 36827 45665 36873 45711
rect 36951 45665 36997 45711
rect 37075 45665 37121 45711
rect 37199 45665 37245 45711
rect 37323 45665 37369 45711
rect 37447 45665 37493 45711
rect 37571 45665 37617 45711
rect 37695 45665 37741 45711
rect 37819 45665 37865 45711
rect 37943 45665 37989 45711
rect 38067 45665 38113 45711
rect 38191 45665 38237 45711
rect 38315 45665 38361 45711
rect 38439 45665 38485 45711
rect 38563 45665 38609 45711
rect 38687 45665 38733 45711
rect 38811 45665 38857 45711
rect 38935 45665 38981 45711
rect 39059 45665 39105 45711
rect 39183 45665 39229 45711
rect 39307 45665 39353 45711
rect 39431 45665 39477 45711
rect 39555 45665 39601 45711
rect 39679 45665 39725 45711
rect 39803 45665 39849 45711
rect 39927 45665 39973 45711
rect 40051 45665 40097 45711
rect 40175 45665 40221 45711
rect 40299 45665 40345 45711
rect 40423 45665 40469 45711
rect 40547 45665 40593 45711
rect 40671 45665 40717 45711
rect 40795 45665 40841 45711
rect 40919 45665 40965 45711
rect 41043 45665 41089 45711
rect 41167 45665 41213 45711
rect 41291 45665 41337 45711
rect 41415 45665 41461 45711
rect 41539 45665 41585 45711
rect 41663 45665 41709 45711
rect 41787 45665 41833 45711
rect 41911 45665 41957 45711
rect 42035 45665 42081 45711
rect 42159 45665 42205 45711
rect 42283 45665 42329 45711
rect 42407 45665 42453 45711
rect 42531 45665 42577 45711
rect 42655 45665 42701 45711
rect 42779 45665 42825 45711
rect 42903 45665 42949 45711
rect 43027 45665 43073 45711
rect 43151 45665 43197 45711
rect 43275 45665 43321 45711
rect 43399 45665 43445 45711
rect 43523 45665 43569 45711
rect 43647 45665 43693 45711
rect 43771 45665 43817 45711
rect 43895 45665 43941 45711
rect 44019 45665 44065 45711
rect 44143 45665 44189 45711
rect 44267 45665 44313 45711
rect 44391 45665 44437 45711
rect 44515 45665 44561 45711
rect 44639 45665 44685 45711
rect 44763 45665 44809 45711
rect 44887 45665 44933 45711
rect 45011 45665 45057 45711
rect 45135 45665 45181 45711
rect 45259 45665 45305 45711
rect 45383 45665 45429 45711
rect 45507 45665 45553 45711
rect 45631 45665 45677 45711
rect 45755 45665 45801 45711
rect 45879 45665 45925 45711
rect 46003 45665 46049 45711
rect 46127 45665 46173 45711
rect 46251 45665 46297 45711
rect 46375 45665 46421 45711
rect 46499 45665 46545 45711
rect 46623 45665 46669 45711
rect 46747 45665 46793 45711
rect 46871 45665 46917 45711
rect 46995 45665 47041 45711
rect 47119 45665 47165 45711
rect 47243 45665 47289 45711
rect 47367 45665 47413 45711
rect 47491 45665 47537 45711
rect 47615 45665 47661 45711
rect 47739 45665 47785 45711
rect 47863 45665 47909 45711
rect 47987 45665 48033 45711
rect 48111 45665 48157 45711
rect 48235 45665 48281 45711
rect 48359 45665 48405 45711
rect 48483 45665 48529 45711
rect 48607 45665 48653 45711
rect 48731 45665 48777 45711
rect 48855 45665 48901 45711
rect 48979 45665 49025 45711
rect 49103 45665 49149 45711
rect 49227 45665 49273 45711
rect 49351 45665 49397 45711
rect 49475 45665 49521 45711
rect 49599 45665 49645 45711
rect 49723 45665 49769 45711
rect 49847 45665 49893 45711
rect 49971 45665 50017 45711
rect 50095 45665 50141 45711
rect 50219 45665 50265 45711
rect 50343 45665 50389 45711
rect 50467 45665 50513 45711
rect 50591 45665 50637 45711
rect 50715 45665 50761 45711
rect 50839 45665 50885 45711
rect 50963 45665 51009 45711
rect 51087 45665 51133 45711
rect 51211 45665 51257 45711
rect 51335 45665 51381 45711
rect 51459 45665 51505 45711
rect 51583 45665 51629 45711
rect 51707 45665 51753 45711
rect 51831 45665 51877 45711
rect 51955 45665 52001 45711
rect 52079 45665 52125 45711
rect 52203 45665 52249 45711
rect 52327 45665 52373 45711
rect 52451 45665 52497 45711
rect 52575 45665 52621 45711
rect 52699 45665 52745 45711
rect 52823 45665 52869 45711
rect 52947 45665 52993 45711
rect 53071 45665 53117 45711
rect 53195 45665 53241 45711
rect 53319 45665 53365 45711
rect 53443 45665 53489 45711
rect 53567 45665 53613 45711
rect 53691 45665 53737 45711
rect 53815 45665 53861 45711
rect 53939 45665 53985 45711
rect 54063 45665 54109 45711
rect 54187 45665 54233 45711
rect 54311 45665 54357 45711
rect 54435 45665 54481 45711
rect 54559 45665 54605 45711
rect 54683 45665 54729 45711
rect 54807 45665 54853 45711
rect 54931 45665 54977 45711
rect 55055 45665 55101 45711
rect 55179 45665 55225 45711
rect 55303 45665 55349 45711
rect 55427 45665 55473 45711
rect 55551 45665 55597 45711
rect 55675 45665 55721 45711
rect 55799 45665 55845 45711
rect 55923 45665 55969 45711
rect 56047 45665 56093 45711
rect 56171 45665 56217 45711
rect 56295 45665 56341 45711
rect 56419 45665 56465 45711
rect 56543 45665 56589 45711
rect 56667 45665 56713 45711
rect 56791 45665 56837 45711
rect 56915 45665 56961 45711
rect 57039 45665 57085 45711
rect 57163 45665 57209 45711
rect 57287 45665 57333 45711
rect 57411 45665 57457 45711
rect 57535 45665 57581 45711
rect 57659 45665 57705 45711
rect 57783 45665 57829 45711
rect 57907 45665 57953 45711
rect 58031 45665 58077 45711
rect 58155 45665 58201 45711
rect 58279 45665 58325 45711
rect 58403 45665 58449 45711
rect 58527 45665 58573 45711
rect 58651 45665 58697 45711
rect 58775 45665 58821 45711
rect 58899 45665 58945 45711
rect 59023 45665 59069 45711
rect 59147 45665 59193 45711
rect 59271 45665 59317 45711
rect 59395 45665 59441 45711
rect 59519 45665 59565 45711
rect 59643 45665 59689 45711
rect 59767 45665 59813 45711
rect 59891 45665 59937 45711
rect 60015 45665 60061 45711
rect 60139 45665 60185 45711
rect 60263 45665 60309 45711
rect 60387 45665 60433 45711
rect 60511 45665 60557 45711
rect 60635 45665 60681 45711
rect 60759 45665 60805 45711
rect 60883 45665 60929 45711
rect 61007 45665 61053 45711
rect 61131 45665 61177 45711
rect 61255 45665 61301 45711
rect 61379 45665 61425 45711
rect 61503 45665 61549 45711
rect 61627 45665 61673 45711
rect 61751 45665 61797 45711
rect 61875 45665 61921 45711
rect 61999 45665 62045 45711
rect 62123 45665 62169 45711
rect 62247 45665 62293 45711
rect 62371 45665 62417 45711
rect 62495 45665 62541 45711
rect 62619 45665 62665 45711
rect 62743 45665 62789 45711
rect 62867 45665 62913 45711
rect 62991 45665 63037 45711
rect 63115 45665 63161 45711
rect 63239 45665 63285 45711
rect 63363 45665 63409 45711
rect 63487 45665 63533 45711
rect 63611 45665 63657 45711
rect 63735 45665 63781 45711
rect 63859 45665 63905 45711
rect 63983 45665 64029 45711
rect 64107 45665 64153 45711
rect 64231 45665 64277 45711
rect 64355 45665 64401 45711
rect 64479 45665 64525 45711
rect 64603 45665 64649 45711
rect 64727 45665 64773 45711
rect 64851 45665 64897 45711
rect 64975 45665 65021 45711
rect 65099 45665 65145 45711
rect 65223 45665 65269 45711
rect 65347 45665 65393 45711
rect 65471 45665 65517 45711
rect 65595 45665 65641 45711
rect 65719 45665 65765 45711
rect 65843 45665 65889 45711
rect 65967 45665 66013 45711
rect 66091 45665 66137 45711
rect 66215 45665 66261 45711
rect 66339 45665 66385 45711
rect 66463 45665 66509 45711
rect 66587 45665 66633 45711
rect 66711 45665 66757 45711
rect 66835 45665 66881 45711
rect 66959 45665 67005 45711
rect 67083 45665 67129 45711
rect 67207 45665 67253 45711
rect 67331 45665 67377 45711
rect 67455 45665 67501 45711
rect 67579 45665 67625 45711
rect 67703 45665 67749 45711
rect 67827 45665 67873 45711
rect 67951 45665 67997 45711
rect 68075 45665 68121 45711
rect 68199 45665 68245 45711
rect 68323 45665 68369 45711
rect 68447 45665 68493 45711
rect 68571 45665 68617 45711
rect 68695 45665 68741 45711
rect 68819 45665 68865 45711
rect 68943 45665 68989 45711
rect 69067 45665 69113 45711
rect 69191 45665 69237 45711
rect 69315 45665 69361 45711
rect 69439 45665 69485 45711
rect 69563 45665 69609 45711
rect 69687 45665 69733 45711
rect 69811 45665 69857 45711
rect 69935 45665 69981 45711
rect 70059 45665 70105 45711
rect 70183 45665 70229 45711
rect 70307 45665 70353 45711
rect 70431 45665 70477 45711
rect 70555 45665 70601 45711
rect 70679 45665 70725 45711
rect 70803 45665 70849 45711
rect 70927 45665 70973 45711
rect 71051 45665 71097 45711
rect 71175 45665 71221 45711
rect 71299 45665 71345 45711
rect 71423 45665 71469 45711
rect 71547 45665 71593 45711
rect 71671 45665 71717 45711
rect 71795 45665 71841 45711
rect 71919 45665 71965 45711
rect 72043 45665 72089 45711
rect 72167 45665 72213 45711
rect 72291 45665 72337 45711
rect 72415 45665 72461 45711
rect 72539 45665 72585 45711
rect 72663 45665 72709 45711
rect 72787 45665 72833 45711
rect 72911 45665 72957 45711
rect 73035 45665 73081 45711
rect 73159 45665 73205 45711
rect 73283 45665 73329 45711
rect 73407 45665 73453 45711
rect 73531 45665 73577 45711
rect 73655 45665 73701 45711
rect 73779 45665 73825 45711
rect 73903 45665 73949 45711
rect 74027 45665 74073 45711
rect 74151 45665 74197 45711
rect 74275 45665 74321 45711
rect 74399 45665 74445 45711
rect 74523 45665 74569 45711
rect 74647 45665 74693 45711
rect 74771 45665 74817 45711
rect 74895 45665 74941 45711
rect 75019 45665 75065 45711
rect 75143 45665 75189 45711
rect 75267 45665 75313 45711
rect 75391 45665 75437 45711
rect 75515 45665 75561 45711
rect 75639 45665 75685 45711
rect 75763 45665 75809 45711
rect 75887 45665 75933 45711
rect 76011 45665 76057 45711
rect 76135 45665 76181 45711
rect 76259 45665 76305 45711
rect 76383 45665 76429 45711
rect 76507 45665 76553 45711
rect 76631 45665 76677 45711
rect 76755 45665 76801 45711
rect 76879 45665 76925 45711
rect 77003 45665 77049 45711
rect 77127 45665 77173 45711
rect 77251 45665 77297 45711
rect 77375 45665 77421 45711
rect 77499 45665 77545 45711
rect 77623 45665 77669 45711
rect 77747 45665 77793 45711
rect 77871 45665 77917 45711
rect 77995 45665 78041 45711
rect 78119 45665 78165 45711
rect 78243 45665 78289 45711
rect 78367 45665 78413 45711
rect 78491 45665 78537 45711
rect 78615 45665 78661 45711
rect 78739 45665 78785 45711
rect 78863 45665 78909 45711
rect 78987 45665 79033 45711
rect 79111 45665 79157 45711
rect 79235 45665 79281 45711
rect 79359 45665 79405 45711
rect 79483 45665 79529 45711
rect 79607 45665 79653 45711
rect 79731 45665 79777 45711
rect 79855 45665 79901 45711
rect 79979 45665 80025 45711
rect 80103 45665 80149 45711
rect 80227 45665 80273 45711
rect 80351 45665 80397 45711
rect 80475 45665 80521 45711
rect 80599 45665 80645 45711
rect 80723 45665 80769 45711
rect 80847 45665 80893 45711
rect 80971 45665 81017 45711
rect 81095 45665 81141 45711
rect 81219 45665 81265 45711
rect 81343 45665 81389 45711
rect 81467 45665 81513 45711
rect 81591 45665 81637 45711
rect 81715 45665 81761 45711
rect 81839 45665 81885 45711
rect 81963 45665 82009 45711
rect 82087 45665 82133 45711
rect 82211 45665 82257 45711
rect 82335 45665 82381 45711
rect 82459 45665 82505 45711
rect 82583 45665 82629 45711
rect 82707 45665 82753 45711
rect 82831 45665 82877 45711
rect 82955 45665 83001 45711
rect 83079 45665 83125 45711
rect 83203 45665 83249 45711
rect 83327 45665 83373 45711
rect 83451 45665 83497 45711
rect 83575 45665 83621 45711
rect 83699 45665 83745 45711
rect 83823 45665 83869 45711
rect 83947 45665 83993 45711
rect 84071 45665 84117 45711
rect 84195 45665 84241 45711
rect 84319 45665 84365 45711
rect 84443 45665 84489 45711
rect 84567 45665 84613 45711
rect 84691 45665 84737 45711
rect 84815 45665 84861 45711
rect 84939 45665 84985 45711
rect 85063 45665 85109 45711
rect 85187 45665 85233 45711
rect 85311 45665 85357 45711
rect 85435 45665 85481 45711
rect 85559 45665 85605 45711
rect 85683 45665 85729 45711
rect 85807 45665 85853 45711
rect 85931 45665 85977 45711
rect 371 1117 717 45563
rect 27498 1117 27744 45563
rect 27846 35996 28492 45442
rect 33044 44263 33090 44309
rect 33202 44263 33248 44309
rect 33360 44263 33406 44309
rect 33518 44263 33564 44309
rect 33677 44263 33723 44309
rect 33835 44263 33881 44309
rect 33993 44263 34039 44309
rect 34151 44263 34197 44309
rect 34309 44263 34355 44309
rect 34467 44263 34513 44309
rect 34625 44263 34671 44309
rect 34783 44263 34829 44309
rect 40117 44263 40163 44309
rect 40275 44263 40321 44309
rect 40433 44263 40479 44309
rect 40591 44263 40637 44309
rect 40750 44263 40796 44309
rect 40908 44263 40954 44309
rect 41066 44263 41112 44309
rect 41224 44263 41270 44309
rect 41382 44263 41428 44309
rect 41540 44263 41586 44309
rect 41698 44263 41744 44309
rect 41856 44263 41902 44309
rect 28810 44076 28856 44122
rect 28810 43912 28856 43958
rect 28810 43749 28856 43795
rect 28810 43586 28856 43632
rect 28810 43422 28856 43468
rect 44514 44263 44560 44309
rect 44672 44263 44718 44309
rect 44830 44263 44876 44309
rect 50129 44263 50175 44309
rect 50287 44263 50333 44309
rect 50445 44263 50491 44309
rect 50603 44263 50649 44309
rect 50762 44263 50808 44309
rect 50920 44263 50966 44309
rect 51078 44263 51124 44309
rect 51236 44263 51282 44309
rect 51394 44263 51440 44309
rect 51552 44263 51598 44309
rect 51710 44263 51756 44309
rect 51868 44263 51914 44309
rect 28810 43220 28856 43266
rect 28810 43057 28856 43103
rect 28810 42894 28856 42940
rect 28810 42731 28856 42777
rect 28810 42567 28856 42613
rect 37957 43304 38473 43350
rect 40836 43304 40882 43350
rect 40994 43304 41040 43350
rect 41152 43304 41198 43350
rect 41310 43304 41356 43350
rect 41469 43304 41515 43350
rect 41627 43304 41673 43350
rect 41785 43304 41831 43350
rect 41943 43304 41989 43350
rect 42101 43304 42147 43350
rect 42259 43304 42305 43350
rect 42418 43304 42464 43350
rect 42576 43304 42622 43350
rect 42734 43304 42780 43350
rect 42892 43304 42938 43350
rect 56267 44076 56313 44122
rect 56267 43912 56313 43958
rect 56267 43749 56313 43795
rect 56267 43586 56313 43632
rect 56267 43422 56313 43468
rect 28810 42404 28856 42450
rect 28810 42241 28856 42287
rect 28810 42077 28856 42123
rect 28810 41914 28856 41960
rect 28810 41751 28856 41797
rect 28810 41588 28856 41634
rect 34916 42404 34962 42450
rect 50160 42404 50206 42450
rect 56267 43220 56313 43266
rect 56267 43057 56313 43103
rect 56267 42894 56313 42940
rect 56267 42731 56313 42777
rect 56267 42567 56313 42613
rect 56267 42404 56313 42450
rect 28810 41420 28856 41466
rect 28810 41257 28856 41303
rect 28810 41094 28856 41140
rect 28810 40931 28856 40977
rect 28810 40767 28856 40813
rect 37957 41504 38473 41550
rect 40836 41504 40882 41550
rect 40994 41504 41040 41550
rect 41152 41504 41198 41550
rect 41310 41504 41356 41550
rect 41469 41504 41515 41550
rect 41627 41504 41673 41550
rect 41785 41504 41831 41550
rect 41943 41504 41989 41550
rect 42101 41504 42147 41550
rect 42259 41504 42305 41550
rect 42418 41504 42464 41550
rect 42576 41504 42622 41550
rect 42734 41504 42780 41550
rect 42892 41504 42938 41550
rect 56267 42241 56313 42287
rect 56267 42077 56313 42123
rect 56267 41914 56313 41960
rect 56267 41751 56313 41797
rect 56267 41588 56313 41634
rect 28810 40604 28856 40650
rect 28810 40441 28856 40487
rect 28810 40277 28856 40323
rect 28810 40114 28856 40160
rect 28810 39951 28856 39997
rect 28810 39788 28856 39834
rect 34916 40604 34962 40650
rect 50160 40604 50206 40650
rect 56267 41420 56313 41466
rect 56267 41257 56313 41303
rect 56267 41094 56313 41140
rect 56267 40931 56313 40977
rect 56267 40767 56313 40813
rect 56267 40604 56313 40650
rect 28810 39620 28856 39666
rect 28810 39457 28856 39503
rect 28810 39294 28856 39340
rect 28810 39131 28856 39177
rect 28810 38967 28856 39013
rect 37957 39704 38473 39750
rect 40836 39704 40882 39750
rect 40994 39704 41040 39750
rect 41152 39704 41198 39750
rect 41310 39704 41356 39750
rect 41469 39704 41515 39750
rect 41627 39704 41673 39750
rect 41785 39704 41831 39750
rect 41943 39704 41989 39750
rect 42101 39704 42147 39750
rect 42259 39704 42305 39750
rect 42418 39704 42464 39750
rect 42576 39704 42622 39750
rect 42734 39704 42780 39750
rect 42892 39704 42938 39750
rect 56267 40441 56313 40487
rect 56267 40277 56313 40323
rect 56267 40114 56313 40160
rect 56267 39951 56313 39997
rect 56267 39788 56313 39834
rect 28810 38804 28856 38850
rect 28810 38641 28856 38687
rect 28810 38477 28856 38523
rect 28810 38314 28856 38360
rect 28810 38151 28856 38197
rect 28810 37988 28856 38034
rect 34916 38804 34962 38850
rect 50160 38804 50206 38850
rect 56267 39620 56313 39666
rect 56267 39457 56313 39503
rect 56267 39294 56313 39340
rect 56267 39131 56313 39177
rect 56267 38967 56313 39013
rect 56267 38804 56313 38850
rect 28810 37820 28856 37866
rect 28810 37657 28856 37703
rect 28810 37494 28856 37540
rect 28810 37331 28856 37377
rect 28810 37167 28856 37213
rect 37957 37904 38473 37950
rect 40836 37904 40882 37950
rect 40994 37904 41040 37950
rect 41152 37904 41198 37950
rect 41310 37904 41356 37950
rect 41469 37904 41515 37950
rect 41627 37904 41673 37950
rect 41785 37904 41831 37950
rect 41943 37904 41989 37950
rect 42101 37904 42147 37950
rect 42259 37904 42305 37950
rect 42418 37904 42464 37950
rect 42576 37904 42622 37950
rect 42734 37904 42780 37950
rect 42892 37904 42938 37950
rect 56267 38641 56313 38687
rect 56267 38477 56313 38523
rect 56267 38314 56313 38360
rect 56267 38151 56313 38197
rect 56267 37988 56313 38034
rect 28810 37004 28856 37050
rect 28810 36841 28856 36887
rect 28810 36677 28856 36723
rect 28810 36514 28856 36560
rect 28810 36351 28856 36397
rect 28810 36188 28856 36234
rect 34916 37004 34962 37050
rect 50160 37004 50206 37050
rect 56267 37820 56313 37866
rect 56267 37657 56313 37703
rect 56267 37494 56313 37540
rect 56267 37331 56313 37377
rect 56267 37167 56313 37213
rect 56267 37004 56313 37050
rect 37957 36104 38473 36150
rect 40836 36104 40882 36150
rect 40994 36104 41040 36150
rect 41152 36104 41198 36150
rect 41310 36104 41356 36150
rect 41469 36104 41515 36150
rect 41627 36104 41673 36150
rect 41785 36104 41831 36150
rect 41943 36104 41989 36150
rect 42101 36104 42147 36150
rect 42259 36104 42305 36150
rect 42418 36104 42464 36150
rect 42576 36104 42622 36150
rect 42734 36104 42780 36150
rect 42892 36104 42938 36150
rect 56267 36841 56313 36887
rect 56267 36677 56313 36723
rect 56267 36514 56313 36560
rect 56267 36351 56313 36397
rect 56267 36188 56313 36234
rect 56632 35996 57278 45442
rect 27846 34256 57292 34602
rect 28639 3823 28685 3869
rect 28755 3823 28801 3869
rect 28871 3823 28917 3869
rect 28987 3823 29033 3869
rect 29103 3823 29149 3869
rect 29219 3823 29265 3869
rect 29335 3823 29381 3869
rect 29451 3823 29497 3869
rect 29567 3823 29613 3869
rect 29683 3823 29729 3869
rect 29799 3823 29845 3869
rect 29915 3823 29961 3869
rect 30031 3823 30077 3869
rect 30147 3823 30193 3869
rect 30263 3823 30309 3869
rect 30379 3823 30425 3869
rect 30495 3823 30541 3869
rect 30611 3823 30657 3869
rect 30727 3823 30773 3869
rect 30843 3823 30889 3869
rect 30959 3823 31005 3869
rect 31075 3823 31121 3869
rect 31191 3823 31237 3869
rect 31307 3823 31353 3869
rect 31423 3823 31469 3869
rect 31539 3823 31585 3869
rect 31655 3823 31701 3869
rect 31771 3823 31817 3869
rect 31887 3823 31933 3869
rect 32003 3823 32049 3869
rect 32119 3823 32165 3869
rect 32235 3823 32281 3869
rect 32351 3823 32397 3869
rect 32467 3823 32513 3869
rect 32583 3823 32629 3869
rect 32699 3823 32745 3869
rect 32815 3823 32861 3869
rect 32931 3823 32977 3869
rect 33047 3823 33093 3869
rect 33163 3823 33209 3869
rect 33279 3823 33325 3869
rect 33395 3823 33441 3869
rect 33511 3823 33557 3869
rect 33627 3823 33673 3869
rect 33743 3823 33789 3869
rect 33859 3823 33905 3869
rect 33975 3823 34021 3869
rect 34091 3823 34137 3869
rect 34207 3823 34253 3869
rect 34323 3823 34369 3869
rect 34439 3823 34485 3869
rect 34555 3823 34601 3869
rect 34671 3823 34717 3869
rect 34787 3823 34833 3869
rect 34903 3823 34949 3869
rect 35019 3823 35065 3869
rect 35135 3823 35181 3869
rect 35251 3823 35297 3869
rect 35367 3823 35413 3869
rect 35483 3823 35529 3869
rect 35599 3823 35645 3869
rect 35715 3823 35761 3869
rect 35831 3823 35877 3869
rect 35947 3823 35993 3869
rect 36063 3823 36109 3869
rect 36179 3823 36225 3869
rect 36295 3823 36341 3869
rect 36411 3823 36457 3869
rect 36527 3823 36573 3869
rect 36643 3823 36689 3869
rect 36759 3823 36805 3869
rect 36875 3823 36921 3869
rect 36991 3823 37037 3869
rect 37107 3823 37153 3869
rect 37223 3823 37269 3869
rect 37339 3823 37385 3869
rect 37455 3823 37501 3869
rect 37571 3823 37617 3869
rect 37687 3823 37733 3869
rect 37803 3823 37849 3869
rect 37919 3823 37965 3869
rect 38035 3823 38081 3869
rect 38151 3823 38197 3869
rect 38267 3823 38313 3869
rect 38383 3823 38429 3869
rect 38499 3823 38545 3869
rect 38615 3823 38661 3869
rect 38731 3823 38777 3869
rect 38847 3823 38893 3869
rect 38963 3823 39009 3869
rect 39079 3823 39125 3869
rect 39195 3823 39241 3869
rect 39311 3823 39357 3869
rect 39427 3823 39473 3869
rect 39543 3823 39589 3869
rect 39659 3823 39705 3869
rect 39775 3823 39821 3869
rect 39891 3823 39937 3869
rect 40007 3823 40053 3869
rect 40123 3823 40169 3869
rect 28639 3707 28685 3753
rect 28755 3707 28801 3753
rect 28871 3707 28917 3753
rect 28987 3707 29033 3753
rect 29103 3707 29149 3753
rect 29219 3707 29265 3753
rect 29335 3707 29381 3753
rect 29451 3707 29497 3753
rect 29567 3707 29613 3753
rect 29683 3707 29729 3753
rect 29799 3707 29845 3753
rect 29915 3707 29961 3753
rect 30031 3707 30077 3753
rect 30147 3707 30193 3753
rect 30263 3707 30309 3753
rect 30379 3707 30425 3753
rect 30495 3707 30541 3753
rect 30611 3707 30657 3753
rect 30727 3707 30773 3753
rect 30843 3707 30889 3753
rect 30959 3707 31005 3753
rect 31075 3707 31121 3753
rect 31191 3707 31237 3753
rect 31307 3707 31353 3753
rect 31423 3707 31469 3753
rect 31539 3707 31585 3753
rect 31655 3707 31701 3753
rect 31771 3707 31817 3753
rect 31887 3707 31933 3753
rect 32003 3707 32049 3753
rect 32119 3707 32165 3753
rect 32235 3707 32281 3753
rect 32351 3707 32397 3753
rect 32467 3707 32513 3753
rect 32583 3707 32629 3753
rect 32699 3707 32745 3753
rect 32815 3707 32861 3753
rect 32931 3707 32977 3753
rect 33047 3707 33093 3753
rect 33163 3707 33209 3753
rect 33279 3707 33325 3753
rect 33395 3707 33441 3753
rect 33511 3707 33557 3753
rect 33627 3707 33673 3753
rect 33743 3707 33789 3753
rect 33859 3707 33905 3753
rect 33975 3707 34021 3753
rect 34091 3707 34137 3753
rect 34207 3707 34253 3753
rect 34323 3707 34369 3753
rect 34439 3707 34485 3753
rect 34555 3707 34601 3753
rect 34671 3707 34717 3753
rect 34787 3707 34833 3753
rect 34903 3707 34949 3753
rect 35019 3707 35065 3753
rect 35135 3707 35181 3753
rect 35251 3707 35297 3753
rect 35367 3707 35413 3753
rect 35483 3707 35529 3753
rect 35599 3707 35645 3753
rect 35715 3707 35761 3753
rect 35831 3707 35877 3753
rect 35947 3707 35993 3753
rect 36063 3707 36109 3753
rect 36179 3707 36225 3753
rect 36295 3707 36341 3753
rect 36411 3707 36457 3753
rect 36527 3707 36573 3753
rect 36643 3707 36689 3753
rect 36759 3707 36805 3753
rect 36875 3707 36921 3753
rect 36991 3707 37037 3753
rect 37107 3707 37153 3753
rect 37223 3707 37269 3753
rect 37339 3707 37385 3753
rect 37455 3707 37501 3753
rect 37571 3707 37617 3753
rect 37687 3707 37733 3753
rect 37803 3707 37849 3753
rect 37919 3707 37965 3753
rect 38035 3707 38081 3753
rect 38151 3707 38197 3753
rect 38267 3707 38313 3753
rect 38383 3707 38429 3753
rect 38499 3707 38545 3753
rect 38615 3707 38661 3753
rect 38731 3707 38777 3753
rect 38847 3707 38893 3753
rect 38963 3707 39009 3753
rect 39079 3707 39125 3753
rect 39195 3707 39241 3753
rect 39311 3707 39357 3753
rect 39427 3707 39473 3753
rect 39543 3707 39589 3753
rect 39659 3707 39705 3753
rect 39775 3707 39821 3753
rect 39891 3707 39937 3753
rect 40007 3707 40053 3753
rect 40123 3707 40169 3753
rect 28639 3591 28685 3637
rect 28755 3591 28801 3637
rect 28871 3591 28917 3637
rect 28987 3591 29033 3637
rect 29103 3591 29149 3637
rect 29219 3591 29265 3637
rect 29335 3591 29381 3637
rect 29451 3591 29497 3637
rect 29567 3591 29613 3637
rect 29683 3591 29729 3637
rect 29799 3591 29845 3637
rect 29915 3591 29961 3637
rect 30031 3591 30077 3637
rect 30147 3591 30193 3637
rect 30263 3591 30309 3637
rect 30379 3591 30425 3637
rect 30495 3591 30541 3637
rect 30611 3591 30657 3637
rect 30727 3591 30773 3637
rect 30843 3591 30889 3637
rect 30959 3591 31005 3637
rect 31075 3591 31121 3637
rect 31191 3591 31237 3637
rect 31307 3591 31353 3637
rect 31423 3591 31469 3637
rect 31539 3591 31585 3637
rect 31655 3591 31701 3637
rect 31771 3591 31817 3637
rect 31887 3591 31933 3637
rect 32003 3591 32049 3637
rect 32119 3591 32165 3637
rect 32235 3591 32281 3637
rect 32351 3591 32397 3637
rect 32467 3591 32513 3637
rect 32583 3591 32629 3637
rect 32699 3591 32745 3637
rect 32815 3591 32861 3637
rect 32931 3591 32977 3637
rect 33047 3591 33093 3637
rect 33163 3591 33209 3637
rect 33279 3591 33325 3637
rect 33395 3591 33441 3637
rect 33511 3591 33557 3637
rect 33627 3591 33673 3637
rect 33743 3591 33789 3637
rect 33859 3591 33905 3637
rect 33975 3591 34021 3637
rect 34091 3591 34137 3637
rect 34207 3591 34253 3637
rect 34323 3591 34369 3637
rect 34439 3591 34485 3637
rect 34555 3591 34601 3637
rect 34671 3591 34717 3637
rect 34787 3591 34833 3637
rect 34903 3591 34949 3637
rect 35019 3591 35065 3637
rect 35135 3591 35181 3637
rect 35251 3591 35297 3637
rect 35367 3591 35413 3637
rect 35483 3591 35529 3637
rect 35599 3591 35645 3637
rect 35715 3591 35761 3637
rect 35831 3591 35877 3637
rect 35947 3591 35993 3637
rect 36063 3591 36109 3637
rect 36179 3591 36225 3637
rect 36295 3591 36341 3637
rect 36411 3591 36457 3637
rect 36527 3591 36573 3637
rect 36643 3591 36689 3637
rect 36759 3591 36805 3637
rect 36875 3591 36921 3637
rect 36991 3591 37037 3637
rect 37107 3591 37153 3637
rect 37223 3591 37269 3637
rect 37339 3591 37385 3637
rect 37455 3591 37501 3637
rect 37571 3591 37617 3637
rect 37687 3591 37733 3637
rect 37803 3591 37849 3637
rect 37919 3591 37965 3637
rect 38035 3591 38081 3637
rect 38151 3591 38197 3637
rect 38267 3591 38313 3637
rect 38383 3591 38429 3637
rect 38499 3591 38545 3637
rect 38615 3591 38661 3637
rect 38731 3591 38777 3637
rect 38847 3591 38893 3637
rect 38963 3591 39009 3637
rect 39079 3591 39125 3637
rect 39195 3591 39241 3637
rect 39311 3591 39357 3637
rect 39427 3591 39473 3637
rect 39543 3591 39589 3637
rect 39659 3591 39705 3637
rect 39775 3591 39821 3637
rect 39891 3591 39937 3637
rect 40007 3591 40053 3637
rect 40123 3591 40169 3637
rect 28639 3475 28685 3521
rect 28755 3475 28801 3521
rect 28871 3475 28917 3521
rect 28987 3475 29033 3521
rect 29103 3475 29149 3521
rect 29219 3475 29265 3521
rect 29335 3475 29381 3521
rect 29451 3475 29497 3521
rect 29567 3475 29613 3521
rect 29683 3475 29729 3521
rect 29799 3475 29845 3521
rect 29915 3475 29961 3521
rect 30031 3475 30077 3521
rect 30147 3475 30193 3521
rect 30263 3475 30309 3521
rect 30379 3475 30425 3521
rect 30495 3475 30541 3521
rect 30611 3475 30657 3521
rect 30727 3475 30773 3521
rect 30843 3475 30889 3521
rect 30959 3475 31005 3521
rect 31075 3475 31121 3521
rect 31191 3475 31237 3521
rect 31307 3475 31353 3521
rect 31423 3475 31469 3521
rect 31539 3475 31585 3521
rect 31655 3475 31701 3521
rect 31771 3475 31817 3521
rect 31887 3475 31933 3521
rect 32003 3475 32049 3521
rect 32119 3475 32165 3521
rect 32235 3475 32281 3521
rect 32351 3475 32397 3521
rect 32467 3475 32513 3521
rect 32583 3475 32629 3521
rect 32699 3475 32745 3521
rect 32815 3475 32861 3521
rect 32931 3475 32977 3521
rect 33047 3475 33093 3521
rect 33163 3475 33209 3521
rect 33279 3475 33325 3521
rect 33395 3475 33441 3521
rect 33511 3475 33557 3521
rect 33627 3475 33673 3521
rect 33743 3475 33789 3521
rect 33859 3475 33905 3521
rect 33975 3475 34021 3521
rect 34091 3475 34137 3521
rect 34207 3475 34253 3521
rect 34323 3475 34369 3521
rect 34439 3475 34485 3521
rect 34555 3475 34601 3521
rect 34671 3475 34717 3521
rect 34787 3475 34833 3521
rect 34903 3475 34949 3521
rect 35019 3475 35065 3521
rect 35135 3475 35181 3521
rect 35251 3475 35297 3521
rect 35367 3475 35413 3521
rect 35483 3475 35529 3521
rect 35599 3475 35645 3521
rect 35715 3475 35761 3521
rect 35831 3475 35877 3521
rect 35947 3475 35993 3521
rect 36063 3475 36109 3521
rect 36179 3475 36225 3521
rect 36295 3475 36341 3521
rect 36411 3475 36457 3521
rect 36527 3475 36573 3521
rect 36643 3475 36689 3521
rect 36759 3475 36805 3521
rect 36875 3475 36921 3521
rect 36991 3475 37037 3521
rect 37107 3475 37153 3521
rect 37223 3475 37269 3521
rect 37339 3475 37385 3521
rect 37455 3475 37501 3521
rect 37571 3475 37617 3521
rect 37687 3475 37733 3521
rect 37803 3475 37849 3521
rect 37919 3475 37965 3521
rect 38035 3475 38081 3521
rect 38151 3475 38197 3521
rect 38267 3475 38313 3521
rect 38383 3475 38429 3521
rect 38499 3475 38545 3521
rect 38615 3475 38661 3521
rect 38731 3475 38777 3521
rect 38847 3475 38893 3521
rect 38963 3475 39009 3521
rect 39079 3475 39125 3521
rect 39195 3475 39241 3521
rect 39311 3475 39357 3521
rect 39427 3475 39473 3521
rect 39543 3475 39589 3521
rect 39659 3475 39705 3521
rect 39775 3475 39821 3521
rect 39891 3475 39937 3521
rect 40007 3475 40053 3521
rect 40123 3475 40169 3521
rect 28639 3359 28685 3405
rect 28755 3359 28801 3405
rect 28871 3359 28917 3405
rect 28987 3359 29033 3405
rect 29103 3359 29149 3405
rect 29219 3359 29265 3405
rect 29335 3359 29381 3405
rect 29451 3359 29497 3405
rect 29567 3359 29613 3405
rect 29683 3359 29729 3405
rect 29799 3359 29845 3405
rect 29915 3359 29961 3405
rect 30031 3359 30077 3405
rect 30147 3359 30193 3405
rect 30263 3359 30309 3405
rect 30379 3359 30425 3405
rect 30495 3359 30541 3405
rect 30611 3359 30657 3405
rect 30727 3359 30773 3405
rect 30843 3359 30889 3405
rect 30959 3359 31005 3405
rect 31075 3359 31121 3405
rect 31191 3359 31237 3405
rect 31307 3359 31353 3405
rect 31423 3359 31469 3405
rect 31539 3359 31585 3405
rect 31655 3359 31701 3405
rect 31771 3359 31817 3405
rect 31887 3359 31933 3405
rect 32003 3359 32049 3405
rect 32119 3359 32165 3405
rect 32235 3359 32281 3405
rect 32351 3359 32397 3405
rect 32467 3359 32513 3405
rect 32583 3359 32629 3405
rect 32699 3359 32745 3405
rect 32815 3359 32861 3405
rect 32931 3359 32977 3405
rect 33047 3359 33093 3405
rect 33163 3359 33209 3405
rect 33279 3359 33325 3405
rect 33395 3359 33441 3405
rect 33511 3359 33557 3405
rect 33627 3359 33673 3405
rect 33743 3359 33789 3405
rect 33859 3359 33905 3405
rect 33975 3359 34021 3405
rect 34091 3359 34137 3405
rect 34207 3359 34253 3405
rect 34323 3359 34369 3405
rect 34439 3359 34485 3405
rect 34555 3359 34601 3405
rect 34671 3359 34717 3405
rect 34787 3359 34833 3405
rect 34903 3359 34949 3405
rect 35019 3359 35065 3405
rect 35135 3359 35181 3405
rect 35251 3359 35297 3405
rect 35367 3359 35413 3405
rect 35483 3359 35529 3405
rect 35599 3359 35645 3405
rect 35715 3359 35761 3405
rect 35831 3359 35877 3405
rect 35947 3359 35993 3405
rect 36063 3359 36109 3405
rect 36179 3359 36225 3405
rect 36295 3359 36341 3405
rect 36411 3359 36457 3405
rect 36527 3359 36573 3405
rect 36643 3359 36689 3405
rect 36759 3359 36805 3405
rect 36875 3359 36921 3405
rect 36991 3359 37037 3405
rect 37107 3359 37153 3405
rect 37223 3359 37269 3405
rect 37339 3359 37385 3405
rect 37455 3359 37501 3405
rect 37571 3359 37617 3405
rect 37687 3359 37733 3405
rect 37803 3359 37849 3405
rect 37919 3359 37965 3405
rect 38035 3359 38081 3405
rect 38151 3359 38197 3405
rect 38267 3359 38313 3405
rect 38383 3359 38429 3405
rect 38499 3359 38545 3405
rect 38615 3359 38661 3405
rect 38731 3359 38777 3405
rect 38847 3359 38893 3405
rect 38963 3359 39009 3405
rect 39079 3359 39125 3405
rect 39195 3359 39241 3405
rect 39311 3359 39357 3405
rect 39427 3359 39473 3405
rect 39543 3359 39589 3405
rect 39659 3359 39705 3405
rect 39775 3359 39821 3405
rect 39891 3359 39937 3405
rect 40007 3359 40053 3405
rect 40123 3359 40169 3405
rect 28639 3243 28685 3289
rect 28755 3243 28801 3289
rect 28871 3243 28917 3289
rect 28987 3243 29033 3289
rect 29103 3243 29149 3289
rect 29219 3243 29265 3289
rect 29335 3243 29381 3289
rect 29451 3243 29497 3289
rect 29567 3243 29613 3289
rect 29683 3243 29729 3289
rect 29799 3243 29845 3289
rect 29915 3243 29961 3289
rect 30031 3243 30077 3289
rect 30147 3243 30193 3289
rect 30263 3243 30309 3289
rect 30379 3243 30425 3289
rect 30495 3243 30541 3289
rect 30611 3243 30657 3289
rect 30727 3243 30773 3289
rect 30843 3243 30889 3289
rect 30959 3243 31005 3289
rect 31075 3243 31121 3289
rect 31191 3243 31237 3289
rect 31307 3243 31353 3289
rect 31423 3243 31469 3289
rect 31539 3243 31585 3289
rect 31655 3243 31701 3289
rect 31771 3243 31817 3289
rect 31887 3243 31933 3289
rect 32003 3243 32049 3289
rect 32119 3243 32165 3289
rect 32235 3243 32281 3289
rect 32351 3243 32397 3289
rect 32467 3243 32513 3289
rect 32583 3243 32629 3289
rect 32699 3243 32745 3289
rect 32815 3243 32861 3289
rect 32931 3243 32977 3289
rect 33047 3243 33093 3289
rect 33163 3243 33209 3289
rect 33279 3243 33325 3289
rect 33395 3243 33441 3289
rect 33511 3243 33557 3289
rect 33627 3243 33673 3289
rect 33743 3243 33789 3289
rect 33859 3243 33905 3289
rect 33975 3243 34021 3289
rect 34091 3243 34137 3289
rect 34207 3243 34253 3289
rect 34323 3243 34369 3289
rect 34439 3243 34485 3289
rect 34555 3243 34601 3289
rect 34671 3243 34717 3289
rect 34787 3243 34833 3289
rect 34903 3243 34949 3289
rect 35019 3243 35065 3289
rect 35135 3243 35181 3289
rect 35251 3243 35297 3289
rect 35367 3243 35413 3289
rect 35483 3243 35529 3289
rect 35599 3243 35645 3289
rect 35715 3243 35761 3289
rect 35831 3243 35877 3289
rect 35947 3243 35993 3289
rect 36063 3243 36109 3289
rect 36179 3243 36225 3289
rect 36295 3243 36341 3289
rect 36411 3243 36457 3289
rect 36527 3243 36573 3289
rect 36643 3243 36689 3289
rect 36759 3243 36805 3289
rect 36875 3243 36921 3289
rect 36991 3243 37037 3289
rect 37107 3243 37153 3289
rect 37223 3243 37269 3289
rect 37339 3243 37385 3289
rect 37455 3243 37501 3289
rect 37571 3243 37617 3289
rect 37687 3243 37733 3289
rect 37803 3243 37849 3289
rect 37919 3243 37965 3289
rect 38035 3243 38081 3289
rect 38151 3243 38197 3289
rect 38267 3243 38313 3289
rect 38383 3243 38429 3289
rect 38499 3243 38545 3289
rect 38615 3243 38661 3289
rect 38731 3243 38777 3289
rect 38847 3243 38893 3289
rect 38963 3243 39009 3289
rect 39079 3243 39125 3289
rect 39195 3243 39241 3289
rect 39311 3243 39357 3289
rect 39427 3243 39473 3289
rect 39543 3243 39589 3289
rect 39659 3243 39705 3289
rect 39775 3243 39821 3289
rect 39891 3243 39937 3289
rect 40007 3243 40053 3289
rect 40123 3243 40169 3289
rect 28639 3127 28685 3173
rect 28755 3127 28801 3173
rect 28871 3127 28917 3173
rect 28987 3127 29033 3173
rect 29103 3127 29149 3173
rect 29219 3127 29265 3173
rect 29335 3127 29381 3173
rect 29451 3127 29497 3173
rect 29567 3127 29613 3173
rect 29683 3127 29729 3173
rect 29799 3127 29845 3173
rect 29915 3127 29961 3173
rect 30031 3127 30077 3173
rect 30147 3127 30193 3173
rect 30263 3127 30309 3173
rect 30379 3127 30425 3173
rect 30495 3127 30541 3173
rect 30611 3127 30657 3173
rect 30727 3127 30773 3173
rect 30843 3127 30889 3173
rect 30959 3127 31005 3173
rect 31075 3127 31121 3173
rect 31191 3127 31237 3173
rect 31307 3127 31353 3173
rect 31423 3127 31469 3173
rect 31539 3127 31585 3173
rect 31655 3127 31701 3173
rect 31771 3127 31817 3173
rect 31887 3127 31933 3173
rect 32003 3127 32049 3173
rect 32119 3127 32165 3173
rect 32235 3127 32281 3173
rect 32351 3127 32397 3173
rect 32467 3127 32513 3173
rect 32583 3127 32629 3173
rect 32699 3127 32745 3173
rect 32815 3127 32861 3173
rect 32931 3127 32977 3173
rect 33047 3127 33093 3173
rect 33163 3127 33209 3173
rect 33279 3127 33325 3173
rect 33395 3127 33441 3173
rect 33511 3127 33557 3173
rect 33627 3127 33673 3173
rect 33743 3127 33789 3173
rect 33859 3127 33905 3173
rect 33975 3127 34021 3173
rect 34091 3127 34137 3173
rect 34207 3127 34253 3173
rect 34323 3127 34369 3173
rect 34439 3127 34485 3173
rect 34555 3127 34601 3173
rect 34671 3127 34717 3173
rect 34787 3127 34833 3173
rect 34903 3127 34949 3173
rect 35019 3127 35065 3173
rect 35135 3127 35181 3173
rect 35251 3127 35297 3173
rect 35367 3127 35413 3173
rect 35483 3127 35529 3173
rect 35599 3127 35645 3173
rect 35715 3127 35761 3173
rect 35831 3127 35877 3173
rect 35947 3127 35993 3173
rect 36063 3127 36109 3173
rect 36179 3127 36225 3173
rect 36295 3127 36341 3173
rect 36411 3127 36457 3173
rect 36527 3127 36573 3173
rect 36643 3127 36689 3173
rect 36759 3127 36805 3173
rect 36875 3127 36921 3173
rect 36991 3127 37037 3173
rect 37107 3127 37153 3173
rect 37223 3127 37269 3173
rect 37339 3127 37385 3173
rect 37455 3127 37501 3173
rect 37571 3127 37617 3173
rect 37687 3127 37733 3173
rect 37803 3127 37849 3173
rect 37919 3127 37965 3173
rect 38035 3127 38081 3173
rect 38151 3127 38197 3173
rect 38267 3127 38313 3173
rect 38383 3127 38429 3173
rect 38499 3127 38545 3173
rect 38615 3127 38661 3173
rect 38731 3127 38777 3173
rect 38847 3127 38893 3173
rect 38963 3127 39009 3173
rect 39079 3127 39125 3173
rect 39195 3127 39241 3173
rect 39311 3127 39357 3173
rect 39427 3127 39473 3173
rect 39543 3127 39589 3173
rect 39659 3127 39705 3173
rect 39775 3127 39821 3173
rect 39891 3127 39937 3173
rect 40007 3127 40053 3173
rect 40123 3127 40169 3173
rect 28639 3011 28685 3057
rect 28755 3011 28801 3057
rect 28871 3011 28917 3057
rect 28987 3011 29033 3057
rect 29103 3011 29149 3057
rect 29219 3011 29265 3057
rect 29335 3011 29381 3057
rect 29451 3011 29497 3057
rect 29567 3011 29613 3057
rect 29683 3011 29729 3057
rect 29799 3011 29845 3057
rect 29915 3011 29961 3057
rect 30031 3011 30077 3057
rect 30147 3011 30193 3057
rect 30263 3011 30309 3057
rect 30379 3011 30425 3057
rect 30495 3011 30541 3057
rect 30611 3011 30657 3057
rect 30727 3011 30773 3057
rect 30843 3011 30889 3057
rect 30959 3011 31005 3057
rect 31075 3011 31121 3057
rect 31191 3011 31237 3057
rect 31307 3011 31353 3057
rect 31423 3011 31469 3057
rect 31539 3011 31585 3057
rect 31655 3011 31701 3057
rect 31771 3011 31817 3057
rect 31887 3011 31933 3057
rect 32003 3011 32049 3057
rect 32119 3011 32165 3057
rect 32235 3011 32281 3057
rect 32351 3011 32397 3057
rect 32467 3011 32513 3057
rect 32583 3011 32629 3057
rect 32699 3011 32745 3057
rect 32815 3011 32861 3057
rect 32931 3011 32977 3057
rect 33047 3011 33093 3057
rect 33163 3011 33209 3057
rect 33279 3011 33325 3057
rect 33395 3011 33441 3057
rect 33511 3011 33557 3057
rect 33627 3011 33673 3057
rect 33743 3011 33789 3057
rect 33859 3011 33905 3057
rect 33975 3011 34021 3057
rect 34091 3011 34137 3057
rect 34207 3011 34253 3057
rect 34323 3011 34369 3057
rect 34439 3011 34485 3057
rect 34555 3011 34601 3057
rect 34671 3011 34717 3057
rect 34787 3011 34833 3057
rect 34903 3011 34949 3057
rect 35019 3011 35065 3057
rect 35135 3011 35181 3057
rect 35251 3011 35297 3057
rect 35367 3011 35413 3057
rect 35483 3011 35529 3057
rect 35599 3011 35645 3057
rect 35715 3011 35761 3057
rect 35831 3011 35877 3057
rect 35947 3011 35993 3057
rect 36063 3011 36109 3057
rect 36179 3011 36225 3057
rect 36295 3011 36341 3057
rect 36411 3011 36457 3057
rect 36527 3011 36573 3057
rect 36643 3011 36689 3057
rect 36759 3011 36805 3057
rect 36875 3011 36921 3057
rect 36991 3011 37037 3057
rect 37107 3011 37153 3057
rect 37223 3011 37269 3057
rect 37339 3011 37385 3057
rect 37455 3011 37501 3057
rect 37571 3011 37617 3057
rect 37687 3011 37733 3057
rect 37803 3011 37849 3057
rect 37919 3011 37965 3057
rect 38035 3011 38081 3057
rect 38151 3011 38197 3057
rect 38267 3011 38313 3057
rect 38383 3011 38429 3057
rect 38499 3011 38545 3057
rect 38615 3011 38661 3057
rect 38731 3011 38777 3057
rect 38847 3011 38893 3057
rect 38963 3011 39009 3057
rect 39079 3011 39125 3057
rect 39195 3011 39241 3057
rect 39311 3011 39357 3057
rect 39427 3011 39473 3057
rect 39543 3011 39589 3057
rect 39659 3011 39705 3057
rect 39775 3011 39821 3057
rect 39891 3011 39937 3057
rect 40007 3011 40053 3057
rect 40123 3011 40169 3057
rect 28639 2895 28685 2941
rect 28755 2895 28801 2941
rect 28871 2895 28917 2941
rect 28987 2895 29033 2941
rect 29103 2895 29149 2941
rect 29219 2895 29265 2941
rect 29335 2895 29381 2941
rect 29451 2895 29497 2941
rect 29567 2895 29613 2941
rect 29683 2895 29729 2941
rect 29799 2895 29845 2941
rect 29915 2895 29961 2941
rect 30031 2895 30077 2941
rect 30147 2895 30193 2941
rect 30263 2895 30309 2941
rect 30379 2895 30425 2941
rect 30495 2895 30541 2941
rect 30611 2895 30657 2941
rect 30727 2895 30773 2941
rect 30843 2895 30889 2941
rect 30959 2895 31005 2941
rect 31075 2895 31121 2941
rect 31191 2895 31237 2941
rect 31307 2895 31353 2941
rect 31423 2895 31469 2941
rect 31539 2895 31585 2941
rect 31655 2895 31701 2941
rect 31771 2895 31817 2941
rect 31887 2895 31933 2941
rect 32003 2895 32049 2941
rect 32119 2895 32165 2941
rect 32235 2895 32281 2941
rect 32351 2895 32397 2941
rect 32467 2895 32513 2941
rect 32583 2895 32629 2941
rect 32699 2895 32745 2941
rect 32815 2895 32861 2941
rect 32931 2895 32977 2941
rect 33047 2895 33093 2941
rect 33163 2895 33209 2941
rect 33279 2895 33325 2941
rect 33395 2895 33441 2941
rect 33511 2895 33557 2941
rect 33627 2895 33673 2941
rect 33743 2895 33789 2941
rect 33859 2895 33905 2941
rect 33975 2895 34021 2941
rect 34091 2895 34137 2941
rect 34207 2895 34253 2941
rect 34323 2895 34369 2941
rect 34439 2895 34485 2941
rect 34555 2895 34601 2941
rect 34671 2895 34717 2941
rect 34787 2895 34833 2941
rect 34903 2895 34949 2941
rect 35019 2895 35065 2941
rect 35135 2895 35181 2941
rect 35251 2895 35297 2941
rect 35367 2895 35413 2941
rect 35483 2895 35529 2941
rect 35599 2895 35645 2941
rect 35715 2895 35761 2941
rect 35831 2895 35877 2941
rect 35947 2895 35993 2941
rect 36063 2895 36109 2941
rect 36179 2895 36225 2941
rect 36295 2895 36341 2941
rect 36411 2895 36457 2941
rect 36527 2895 36573 2941
rect 36643 2895 36689 2941
rect 36759 2895 36805 2941
rect 36875 2895 36921 2941
rect 36991 2895 37037 2941
rect 37107 2895 37153 2941
rect 37223 2895 37269 2941
rect 37339 2895 37385 2941
rect 37455 2895 37501 2941
rect 37571 2895 37617 2941
rect 37687 2895 37733 2941
rect 37803 2895 37849 2941
rect 37919 2895 37965 2941
rect 38035 2895 38081 2941
rect 38151 2895 38197 2941
rect 38267 2895 38313 2941
rect 38383 2895 38429 2941
rect 38499 2895 38545 2941
rect 38615 2895 38661 2941
rect 38731 2895 38777 2941
rect 38847 2895 38893 2941
rect 38963 2895 39009 2941
rect 39079 2895 39125 2941
rect 39195 2895 39241 2941
rect 39311 2895 39357 2941
rect 39427 2895 39473 2941
rect 39543 2895 39589 2941
rect 39659 2895 39705 2941
rect 39775 2895 39821 2941
rect 39891 2895 39937 2941
rect 40007 2895 40053 2941
rect 40123 2895 40169 2941
rect 28639 2779 28685 2825
rect 28755 2779 28801 2825
rect 28871 2779 28917 2825
rect 28987 2779 29033 2825
rect 29103 2779 29149 2825
rect 29219 2779 29265 2825
rect 29335 2779 29381 2825
rect 29451 2779 29497 2825
rect 29567 2779 29613 2825
rect 29683 2779 29729 2825
rect 29799 2779 29845 2825
rect 29915 2779 29961 2825
rect 30031 2779 30077 2825
rect 30147 2779 30193 2825
rect 30263 2779 30309 2825
rect 30379 2779 30425 2825
rect 30495 2779 30541 2825
rect 30611 2779 30657 2825
rect 30727 2779 30773 2825
rect 30843 2779 30889 2825
rect 30959 2779 31005 2825
rect 31075 2779 31121 2825
rect 31191 2779 31237 2825
rect 31307 2779 31353 2825
rect 31423 2779 31469 2825
rect 31539 2779 31585 2825
rect 31655 2779 31701 2825
rect 31771 2779 31817 2825
rect 31887 2779 31933 2825
rect 32003 2779 32049 2825
rect 32119 2779 32165 2825
rect 32235 2779 32281 2825
rect 32351 2779 32397 2825
rect 32467 2779 32513 2825
rect 32583 2779 32629 2825
rect 32699 2779 32745 2825
rect 32815 2779 32861 2825
rect 32931 2779 32977 2825
rect 33047 2779 33093 2825
rect 33163 2779 33209 2825
rect 33279 2779 33325 2825
rect 33395 2779 33441 2825
rect 33511 2779 33557 2825
rect 33627 2779 33673 2825
rect 33743 2779 33789 2825
rect 33859 2779 33905 2825
rect 33975 2779 34021 2825
rect 34091 2779 34137 2825
rect 34207 2779 34253 2825
rect 34323 2779 34369 2825
rect 34439 2779 34485 2825
rect 34555 2779 34601 2825
rect 34671 2779 34717 2825
rect 34787 2779 34833 2825
rect 34903 2779 34949 2825
rect 35019 2779 35065 2825
rect 35135 2779 35181 2825
rect 35251 2779 35297 2825
rect 35367 2779 35413 2825
rect 35483 2779 35529 2825
rect 35599 2779 35645 2825
rect 35715 2779 35761 2825
rect 35831 2779 35877 2825
rect 35947 2779 35993 2825
rect 36063 2779 36109 2825
rect 36179 2779 36225 2825
rect 36295 2779 36341 2825
rect 36411 2779 36457 2825
rect 36527 2779 36573 2825
rect 36643 2779 36689 2825
rect 36759 2779 36805 2825
rect 36875 2779 36921 2825
rect 36991 2779 37037 2825
rect 37107 2779 37153 2825
rect 37223 2779 37269 2825
rect 37339 2779 37385 2825
rect 37455 2779 37501 2825
rect 37571 2779 37617 2825
rect 37687 2779 37733 2825
rect 37803 2779 37849 2825
rect 37919 2779 37965 2825
rect 38035 2779 38081 2825
rect 38151 2779 38197 2825
rect 38267 2779 38313 2825
rect 38383 2779 38429 2825
rect 38499 2779 38545 2825
rect 38615 2779 38661 2825
rect 38731 2779 38777 2825
rect 38847 2779 38893 2825
rect 38963 2779 39009 2825
rect 39079 2779 39125 2825
rect 39195 2779 39241 2825
rect 39311 2779 39357 2825
rect 39427 2779 39473 2825
rect 39543 2779 39589 2825
rect 39659 2779 39705 2825
rect 39775 2779 39821 2825
rect 39891 2779 39937 2825
rect 40007 2779 40053 2825
rect 40123 2779 40169 2825
rect 28639 2663 28685 2709
rect 28755 2663 28801 2709
rect 28871 2663 28917 2709
rect 28987 2663 29033 2709
rect 29103 2663 29149 2709
rect 29219 2663 29265 2709
rect 29335 2663 29381 2709
rect 29451 2663 29497 2709
rect 29567 2663 29613 2709
rect 29683 2663 29729 2709
rect 29799 2663 29845 2709
rect 29915 2663 29961 2709
rect 30031 2663 30077 2709
rect 30147 2663 30193 2709
rect 30263 2663 30309 2709
rect 30379 2663 30425 2709
rect 30495 2663 30541 2709
rect 30611 2663 30657 2709
rect 30727 2663 30773 2709
rect 30843 2663 30889 2709
rect 30959 2663 31005 2709
rect 31075 2663 31121 2709
rect 31191 2663 31237 2709
rect 31307 2663 31353 2709
rect 31423 2663 31469 2709
rect 31539 2663 31585 2709
rect 31655 2663 31701 2709
rect 31771 2663 31817 2709
rect 31887 2663 31933 2709
rect 32003 2663 32049 2709
rect 32119 2663 32165 2709
rect 32235 2663 32281 2709
rect 32351 2663 32397 2709
rect 32467 2663 32513 2709
rect 32583 2663 32629 2709
rect 32699 2663 32745 2709
rect 32815 2663 32861 2709
rect 32931 2663 32977 2709
rect 33047 2663 33093 2709
rect 33163 2663 33209 2709
rect 33279 2663 33325 2709
rect 33395 2663 33441 2709
rect 33511 2663 33557 2709
rect 33627 2663 33673 2709
rect 33743 2663 33789 2709
rect 33859 2663 33905 2709
rect 33975 2663 34021 2709
rect 34091 2663 34137 2709
rect 34207 2663 34253 2709
rect 34323 2663 34369 2709
rect 34439 2663 34485 2709
rect 34555 2663 34601 2709
rect 34671 2663 34717 2709
rect 34787 2663 34833 2709
rect 34903 2663 34949 2709
rect 35019 2663 35065 2709
rect 35135 2663 35181 2709
rect 35251 2663 35297 2709
rect 35367 2663 35413 2709
rect 35483 2663 35529 2709
rect 35599 2663 35645 2709
rect 35715 2663 35761 2709
rect 35831 2663 35877 2709
rect 35947 2663 35993 2709
rect 36063 2663 36109 2709
rect 36179 2663 36225 2709
rect 36295 2663 36341 2709
rect 36411 2663 36457 2709
rect 36527 2663 36573 2709
rect 36643 2663 36689 2709
rect 36759 2663 36805 2709
rect 36875 2663 36921 2709
rect 36991 2663 37037 2709
rect 37107 2663 37153 2709
rect 37223 2663 37269 2709
rect 37339 2663 37385 2709
rect 37455 2663 37501 2709
rect 37571 2663 37617 2709
rect 37687 2663 37733 2709
rect 37803 2663 37849 2709
rect 37919 2663 37965 2709
rect 38035 2663 38081 2709
rect 38151 2663 38197 2709
rect 38267 2663 38313 2709
rect 38383 2663 38429 2709
rect 38499 2663 38545 2709
rect 38615 2663 38661 2709
rect 38731 2663 38777 2709
rect 38847 2663 38893 2709
rect 38963 2663 39009 2709
rect 39079 2663 39125 2709
rect 39195 2663 39241 2709
rect 39311 2663 39357 2709
rect 39427 2663 39473 2709
rect 39543 2663 39589 2709
rect 39659 2663 39705 2709
rect 39775 2663 39821 2709
rect 39891 2663 39937 2709
rect 40007 2663 40053 2709
rect 40123 2663 40169 2709
rect 28639 2547 28685 2593
rect 28755 2547 28801 2593
rect 28871 2547 28917 2593
rect 28987 2547 29033 2593
rect 29103 2547 29149 2593
rect 29219 2547 29265 2593
rect 29335 2547 29381 2593
rect 29451 2547 29497 2593
rect 29567 2547 29613 2593
rect 29683 2547 29729 2593
rect 29799 2547 29845 2593
rect 29915 2547 29961 2593
rect 30031 2547 30077 2593
rect 30147 2547 30193 2593
rect 30263 2547 30309 2593
rect 30379 2547 30425 2593
rect 30495 2547 30541 2593
rect 30611 2547 30657 2593
rect 30727 2547 30773 2593
rect 30843 2547 30889 2593
rect 30959 2547 31005 2593
rect 31075 2547 31121 2593
rect 31191 2547 31237 2593
rect 31307 2547 31353 2593
rect 31423 2547 31469 2593
rect 31539 2547 31585 2593
rect 31655 2547 31701 2593
rect 31771 2547 31817 2593
rect 31887 2547 31933 2593
rect 32003 2547 32049 2593
rect 32119 2547 32165 2593
rect 32235 2547 32281 2593
rect 32351 2547 32397 2593
rect 32467 2547 32513 2593
rect 32583 2547 32629 2593
rect 32699 2547 32745 2593
rect 32815 2547 32861 2593
rect 32931 2547 32977 2593
rect 33047 2547 33093 2593
rect 33163 2547 33209 2593
rect 33279 2547 33325 2593
rect 33395 2547 33441 2593
rect 33511 2547 33557 2593
rect 33627 2547 33673 2593
rect 33743 2547 33789 2593
rect 33859 2547 33905 2593
rect 33975 2547 34021 2593
rect 34091 2547 34137 2593
rect 34207 2547 34253 2593
rect 34323 2547 34369 2593
rect 34439 2547 34485 2593
rect 34555 2547 34601 2593
rect 34671 2547 34717 2593
rect 34787 2547 34833 2593
rect 34903 2547 34949 2593
rect 35019 2547 35065 2593
rect 35135 2547 35181 2593
rect 35251 2547 35297 2593
rect 35367 2547 35413 2593
rect 35483 2547 35529 2593
rect 35599 2547 35645 2593
rect 35715 2547 35761 2593
rect 35831 2547 35877 2593
rect 35947 2547 35993 2593
rect 36063 2547 36109 2593
rect 36179 2547 36225 2593
rect 36295 2547 36341 2593
rect 36411 2547 36457 2593
rect 36527 2547 36573 2593
rect 36643 2547 36689 2593
rect 36759 2547 36805 2593
rect 36875 2547 36921 2593
rect 36991 2547 37037 2593
rect 37107 2547 37153 2593
rect 37223 2547 37269 2593
rect 37339 2547 37385 2593
rect 37455 2547 37501 2593
rect 37571 2547 37617 2593
rect 37687 2547 37733 2593
rect 37803 2547 37849 2593
rect 37919 2547 37965 2593
rect 38035 2547 38081 2593
rect 38151 2547 38197 2593
rect 38267 2547 38313 2593
rect 38383 2547 38429 2593
rect 38499 2547 38545 2593
rect 38615 2547 38661 2593
rect 38731 2547 38777 2593
rect 38847 2547 38893 2593
rect 38963 2547 39009 2593
rect 39079 2547 39125 2593
rect 39195 2547 39241 2593
rect 39311 2547 39357 2593
rect 39427 2547 39473 2593
rect 39543 2547 39589 2593
rect 39659 2547 39705 2593
rect 39775 2547 39821 2593
rect 39891 2547 39937 2593
rect 40007 2547 40053 2593
rect 40123 2547 40169 2593
rect 28639 2431 28685 2477
rect 28755 2431 28801 2477
rect 28871 2431 28917 2477
rect 28987 2431 29033 2477
rect 29103 2431 29149 2477
rect 29219 2431 29265 2477
rect 29335 2431 29381 2477
rect 29451 2431 29497 2477
rect 29567 2431 29613 2477
rect 29683 2431 29729 2477
rect 29799 2431 29845 2477
rect 29915 2431 29961 2477
rect 30031 2431 30077 2477
rect 30147 2431 30193 2477
rect 30263 2431 30309 2477
rect 30379 2431 30425 2477
rect 30495 2431 30541 2477
rect 30611 2431 30657 2477
rect 30727 2431 30773 2477
rect 30843 2431 30889 2477
rect 30959 2431 31005 2477
rect 31075 2431 31121 2477
rect 31191 2431 31237 2477
rect 31307 2431 31353 2477
rect 31423 2431 31469 2477
rect 31539 2431 31585 2477
rect 31655 2431 31701 2477
rect 31771 2431 31817 2477
rect 31887 2431 31933 2477
rect 32003 2431 32049 2477
rect 32119 2431 32165 2477
rect 32235 2431 32281 2477
rect 32351 2431 32397 2477
rect 32467 2431 32513 2477
rect 32583 2431 32629 2477
rect 32699 2431 32745 2477
rect 32815 2431 32861 2477
rect 32931 2431 32977 2477
rect 33047 2431 33093 2477
rect 33163 2431 33209 2477
rect 33279 2431 33325 2477
rect 33395 2431 33441 2477
rect 33511 2431 33557 2477
rect 33627 2431 33673 2477
rect 33743 2431 33789 2477
rect 33859 2431 33905 2477
rect 33975 2431 34021 2477
rect 34091 2431 34137 2477
rect 34207 2431 34253 2477
rect 34323 2431 34369 2477
rect 34439 2431 34485 2477
rect 34555 2431 34601 2477
rect 34671 2431 34717 2477
rect 34787 2431 34833 2477
rect 34903 2431 34949 2477
rect 35019 2431 35065 2477
rect 35135 2431 35181 2477
rect 35251 2431 35297 2477
rect 35367 2431 35413 2477
rect 35483 2431 35529 2477
rect 35599 2431 35645 2477
rect 35715 2431 35761 2477
rect 35831 2431 35877 2477
rect 35947 2431 35993 2477
rect 36063 2431 36109 2477
rect 36179 2431 36225 2477
rect 36295 2431 36341 2477
rect 36411 2431 36457 2477
rect 36527 2431 36573 2477
rect 36643 2431 36689 2477
rect 36759 2431 36805 2477
rect 36875 2431 36921 2477
rect 36991 2431 37037 2477
rect 37107 2431 37153 2477
rect 37223 2431 37269 2477
rect 37339 2431 37385 2477
rect 37455 2431 37501 2477
rect 37571 2431 37617 2477
rect 37687 2431 37733 2477
rect 37803 2431 37849 2477
rect 37919 2431 37965 2477
rect 38035 2431 38081 2477
rect 38151 2431 38197 2477
rect 38267 2431 38313 2477
rect 38383 2431 38429 2477
rect 38499 2431 38545 2477
rect 38615 2431 38661 2477
rect 38731 2431 38777 2477
rect 38847 2431 38893 2477
rect 38963 2431 39009 2477
rect 39079 2431 39125 2477
rect 39195 2431 39241 2477
rect 39311 2431 39357 2477
rect 39427 2431 39473 2477
rect 39543 2431 39589 2477
rect 39659 2431 39705 2477
rect 39775 2431 39821 2477
rect 39891 2431 39937 2477
rect 40007 2431 40053 2477
rect 40123 2431 40169 2477
rect 28639 2315 28685 2361
rect 28755 2315 28801 2361
rect 28871 2315 28917 2361
rect 28987 2315 29033 2361
rect 29103 2315 29149 2361
rect 29219 2315 29265 2361
rect 29335 2315 29381 2361
rect 29451 2315 29497 2361
rect 29567 2315 29613 2361
rect 29683 2315 29729 2361
rect 29799 2315 29845 2361
rect 29915 2315 29961 2361
rect 30031 2315 30077 2361
rect 30147 2315 30193 2361
rect 30263 2315 30309 2361
rect 30379 2315 30425 2361
rect 30495 2315 30541 2361
rect 30611 2315 30657 2361
rect 30727 2315 30773 2361
rect 30843 2315 30889 2361
rect 30959 2315 31005 2361
rect 31075 2315 31121 2361
rect 31191 2315 31237 2361
rect 31307 2315 31353 2361
rect 31423 2315 31469 2361
rect 31539 2315 31585 2361
rect 31655 2315 31701 2361
rect 31771 2315 31817 2361
rect 31887 2315 31933 2361
rect 32003 2315 32049 2361
rect 32119 2315 32165 2361
rect 32235 2315 32281 2361
rect 32351 2315 32397 2361
rect 32467 2315 32513 2361
rect 32583 2315 32629 2361
rect 32699 2315 32745 2361
rect 32815 2315 32861 2361
rect 32931 2315 32977 2361
rect 33047 2315 33093 2361
rect 33163 2315 33209 2361
rect 33279 2315 33325 2361
rect 33395 2315 33441 2361
rect 33511 2315 33557 2361
rect 33627 2315 33673 2361
rect 33743 2315 33789 2361
rect 33859 2315 33905 2361
rect 33975 2315 34021 2361
rect 34091 2315 34137 2361
rect 34207 2315 34253 2361
rect 34323 2315 34369 2361
rect 34439 2315 34485 2361
rect 34555 2315 34601 2361
rect 34671 2315 34717 2361
rect 34787 2315 34833 2361
rect 34903 2315 34949 2361
rect 35019 2315 35065 2361
rect 35135 2315 35181 2361
rect 35251 2315 35297 2361
rect 35367 2315 35413 2361
rect 35483 2315 35529 2361
rect 35599 2315 35645 2361
rect 35715 2315 35761 2361
rect 35831 2315 35877 2361
rect 35947 2315 35993 2361
rect 36063 2315 36109 2361
rect 36179 2315 36225 2361
rect 36295 2315 36341 2361
rect 36411 2315 36457 2361
rect 36527 2315 36573 2361
rect 36643 2315 36689 2361
rect 36759 2315 36805 2361
rect 36875 2315 36921 2361
rect 36991 2315 37037 2361
rect 37107 2315 37153 2361
rect 37223 2315 37269 2361
rect 37339 2315 37385 2361
rect 37455 2315 37501 2361
rect 37571 2315 37617 2361
rect 37687 2315 37733 2361
rect 37803 2315 37849 2361
rect 37919 2315 37965 2361
rect 38035 2315 38081 2361
rect 38151 2315 38197 2361
rect 38267 2315 38313 2361
rect 38383 2315 38429 2361
rect 38499 2315 38545 2361
rect 38615 2315 38661 2361
rect 38731 2315 38777 2361
rect 38847 2315 38893 2361
rect 38963 2315 39009 2361
rect 39079 2315 39125 2361
rect 39195 2315 39241 2361
rect 39311 2315 39357 2361
rect 39427 2315 39473 2361
rect 39543 2315 39589 2361
rect 39659 2315 39705 2361
rect 39775 2315 39821 2361
rect 39891 2315 39937 2361
rect 40007 2315 40053 2361
rect 40123 2315 40169 2361
rect 28639 2199 28685 2245
rect 28755 2199 28801 2245
rect 28871 2199 28917 2245
rect 28987 2199 29033 2245
rect 29103 2199 29149 2245
rect 29219 2199 29265 2245
rect 29335 2199 29381 2245
rect 29451 2199 29497 2245
rect 29567 2199 29613 2245
rect 29683 2199 29729 2245
rect 29799 2199 29845 2245
rect 29915 2199 29961 2245
rect 30031 2199 30077 2245
rect 30147 2199 30193 2245
rect 30263 2199 30309 2245
rect 30379 2199 30425 2245
rect 30495 2199 30541 2245
rect 30611 2199 30657 2245
rect 30727 2199 30773 2245
rect 30843 2199 30889 2245
rect 30959 2199 31005 2245
rect 31075 2199 31121 2245
rect 31191 2199 31237 2245
rect 31307 2199 31353 2245
rect 31423 2199 31469 2245
rect 31539 2199 31585 2245
rect 31655 2199 31701 2245
rect 31771 2199 31817 2245
rect 31887 2199 31933 2245
rect 32003 2199 32049 2245
rect 32119 2199 32165 2245
rect 32235 2199 32281 2245
rect 32351 2199 32397 2245
rect 32467 2199 32513 2245
rect 32583 2199 32629 2245
rect 32699 2199 32745 2245
rect 32815 2199 32861 2245
rect 32931 2199 32977 2245
rect 33047 2199 33093 2245
rect 33163 2199 33209 2245
rect 33279 2199 33325 2245
rect 33395 2199 33441 2245
rect 33511 2199 33557 2245
rect 33627 2199 33673 2245
rect 33743 2199 33789 2245
rect 33859 2199 33905 2245
rect 33975 2199 34021 2245
rect 34091 2199 34137 2245
rect 34207 2199 34253 2245
rect 34323 2199 34369 2245
rect 34439 2199 34485 2245
rect 34555 2199 34601 2245
rect 34671 2199 34717 2245
rect 34787 2199 34833 2245
rect 34903 2199 34949 2245
rect 35019 2199 35065 2245
rect 35135 2199 35181 2245
rect 35251 2199 35297 2245
rect 35367 2199 35413 2245
rect 35483 2199 35529 2245
rect 35599 2199 35645 2245
rect 35715 2199 35761 2245
rect 35831 2199 35877 2245
rect 35947 2199 35993 2245
rect 36063 2199 36109 2245
rect 36179 2199 36225 2245
rect 36295 2199 36341 2245
rect 36411 2199 36457 2245
rect 36527 2199 36573 2245
rect 36643 2199 36689 2245
rect 36759 2199 36805 2245
rect 36875 2199 36921 2245
rect 36991 2199 37037 2245
rect 37107 2199 37153 2245
rect 37223 2199 37269 2245
rect 37339 2199 37385 2245
rect 37455 2199 37501 2245
rect 37571 2199 37617 2245
rect 37687 2199 37733 2245
rect 37803 2199 37849 2245
rect 37919 2199 37965 2245
rect 38035 2199 38081 2245
rect 38151 2199 38197 2245
rect 38267 2199 38313 2245
rect 38383 2199 38429 2245
rect 38499 2199 38545 2245
rect 38615 2199 38661 2245
rect 38731 2199 38777 2245
rect 38847 2199 38893 2245
rect 38963 2199 39009 2245
rect 39079 2199 39125 2245
rect 39195 2199 39241 2245
rect 39311 2199 39357 2245
rect 39427 2199 39473 2245
rect 39543 2199 39589 2245
rect 39659 2199 39705 2245
rect 39775 2199 39821 2245
rect 39891 2199 39937 2245
rect 40007 2199 40053 2245
rect 40123 2199 40169 2245
rect 28639 2083 28685 2129
rect 28755 2083 28801 2129
rect 28871 2083 28917 2129
rect 28987 2083 29033 2129
rect 29103 2083 29149 2129
rect 29219 2083 29265 2129
rect 29335 2083 29381 2129
rect 29451 2083 29497 2129
rect 29567 2083 29613 2129
rect 29683 2083 29729 2129
rect 29799 2083 29845 2129
rect 29915 2083 29961 2129
rect 30031 2083 30077 2129
rect 30147 2083 30193 2129
rect 30263 2083 30309 2129
rect 30379 2083 30425 2129
rect 30495 2083 30541 2129
rect 30611 2083 30657 2129
rect 30727 2083 30773 2129
rect 30843 2083 30889 2129
rect 30959 2083 31005 2129
rect 31075 2083 31121 2129
rect 31191 2083 31237 2129
rect 31307 2083 31353 2129
rect 31423 2083 31469 2129
rect 31539 2083 31585 2129
rect 31655 2083 31701 2129
rect 31771 2083 31817 2129
rect 31887 2083 31933 2129
rect 32003 2083 32049 2129
rect 32119 2083 32165 2129
rect 32235 2083 32281 2129
rect 32351 2083 32397 2129
rect 32467 2083 32513 2129
rect 32583 2083 32629 2129
rect 32699 2083 32745 2129
rect 32815 2083 32861 2129
rect 32931 2083 32977 2129
rect 33047 2083 33093 2129
rect 33163 2083 33209 2129
rect 33279 2083 33325 2129
rect 33395 2083 33441 2129
rect 33511 2083 33557 2129
rect 33627 2083 33673 2129
rect 33743 2083 33789 2129
rect 33859 2083 33905 2129
rect 33975 2083 34021 2129
rect 34091 2083 34137 2129
rect 34207 2083 34253 2129
rect 34323 2083 34369 2129
rect 34439 2083 34485 2129
rect 34555 2083 34601 2129
rect 34671 2083 34717 2129
rect 34787 2083 34833 2129
rect 34903 2083 34949 2129
rect 35019 2083 35065 2129
rect 35135 2083 35181 2129
rect 35251 2083 35297 2129
rect 35367 2083 35413 2129
rect 35483 2083 35529 2129
rect 35599 2083 35645 2129
rect 35715 2083 35761 2129
rect 35831 2083 35877 2129
rect 35947 2083 35993 2129
rect 36063 2083 36109 2129
rect 36179 2083 36225 2129
rect 36295 2083 36341 2129
rect 36411 2083 36457 2129
rect 36527 2083 36573 2129
rect 36643 2083 36689 2129
rect 36759 2083 36805 2129
rect 36875 2083 36921 2129
rect 36991 2083 37037 2129
rect 37107 2083 37153 2129
rect 37223 2083 37269 2129
rect 37339 2083 37385 2129
rect 37455 2083 37501 2129
rect 37571 2083 37617 2129
rect 37687 2083 37733 2129
rect 37803 2083 37849 2129
rect 37919 2083 37965 2129
rect 38035 2083 38081 2129
rect 38151 2083 38197 2129
rect 38267 2083 38313 2129
rect 38383 2083 38429 2129
rect 38499 2083 38545 2129
rect 38615 2083 38661 2129
rect 38731 2083 38777 2129
rect 38847 2083 38893 2129
rect 38963 2083 39009 2129
rect 39079 2083 39125 2129
rect 39195 2083 39241 2129
rect 39311 2083 39357 2129
rect 39427 2083 39473 2129
rect 39543 2083 39589 2129
rect 39659 2083 39705 2129
rect 39775 2083 39821 2129
rect 39891 2083 39937 2129
rect 40007 2083 40053 2129
rect 40123 2083 40169 2129
rect 28639 1967 28685 2013
rect 28755 1967 28801 2013
rect 28871 1967 28917 2013
rect 28987 1967 29033 2013
rect 29103 1967 29149 2013
rect 29219 1967 29265 2013
rect 29335 1967 29381 2013
rect 29451 1967 29497 2013
rect 29567 1967 29613 2013
rect 29683 1967 29729 2013
rect 29799 1967 29845 2013
rect 29915 1967 29961 2013
rect 30031 1967 30077 2013
rect 30147 1967 30193 2013
rect 30263 1967 30309 2013
rect 30379 1967 30425 2013
rect 30495 1967 30541 2013
rect 30611 1967 30657 2013
rect 30727 1967 30773 2013
rect 30843 1967 30889 2013
rect 30959 1967 31005 2013
rect 31075 1967 31121 2013
rect 31191 1967 31237 2013
rect 31307 1967 31353 2013
rect 31423 1967 31469 2013
rect 31539 1967 31585 2013
rect 31655 1967 31701 2013
rect 31771 1967 31817 2013
rect 31887 1967 31933 2013
rect 32003 1967 32049 2013
rect 32119 1967 32165 2013
rect 32235 1967 32281 2013
rect 32351 1967 32397 2013
rect 32467 1967 32513 2013
rect 32583 1967 32629 2013
rect 32699 1967 32745 2013
rect 32815 1967 32861 2013
rect 32931 1967 32977 2013
rect 33047 1967 33093 2013
rect 33163 1967 33209 2013
rect 33279 1967 33325 2013
rect 33395 1967 33441 2013
rect 33511 1967 33557 2013
rect 33627 1967 33673 2013
rect 33743 1967 33789 2013
rect 33859 1967 33905 2013
rect 33975 1967 34021 2013
rect 34091 1967 34137 2013
rect 34207 1967 34253 2013
rect 34323 1967 34369 2013
rect 34439 1967 34485 2013
rect 34555 1967 34601 2013
rect 34671 1967 34717 2013
rect 34787 1967 34833 2013
rect 34903 1967 34949 2013
rect 35019 1967 35065 2013
rect 35135 1967 35181 2013
rect 35251 1967 35297 2013
rect 35367 1967 35413 2013
rect 35483 1967 35529 2013
rect 35599 1967 35645 2013
rect 35715 1967 35761 2013
rect 35831 1967 35877 2013
rect 35947 1967 35993 2013
rect 36063 1967 36109 2013
rect 36179 1967 36225 2013
rect 36295 1967 36341 2013
rect 36411 1967 36457 2013
rect 36527 1967 36573 2013
rect 36643 1967 36689 2013
rect 36759 1967 36805 2013
rect 36875 1967 36921 2013
rect 36991 1967 37037 2013
rect 37107 1967 37153 2013
rect 37223 1967 37269 2013
rect 37339 1967 37385 2013
rect 37455 1967 37501 2013
rect 37571 1967 37617 2013
rect 37687 1967 37733 2013
rect 37803 1967 37849 2013
rect 37919 1967 37965 2013
rect 38035 1967 38081 2013
rect 38151 1967 38197 2013
rect 38267 1967 38313 2013
rect 38383 1967 38429 2013
rect 38499 1967 38545 2013
rect 38615 1967 38661 2013
rect 38731 1967 38777 2013
rect 38847 1967 38893 2013
rect 38963 1967 39009 2013
rect 39079 1967 39125 2013
rect 39195 1967 39241 2013
rect 39311 1967 39357 2013
rect 39427 1967 39473 2013
rect 39543 1967 39589 2013
rect 39659 1967 39705 2013
rect 39775 1967 39821 2013
rect 39891 1967 39937 2013
rect 40007 1967 40053 2013
rect 40123 1967 40169 2013
rect 28639 1851 28685 1897
rect 28755 1851 28801 1897
rect 28871 1851 28917 1897
rect 28987 1851 29033 1897
rect 29103 1851 29149 1897
rect 29219 1851 29265 1897
rect 29335 1851 29381 1897
rect 29451 1851 29497 1897
rect 29567 1851 29613 1897
rect 29683 1851 29729 1897
rect 29799 1851 29845 1897
rect 29915 1851 29961 1897
rect 30031 1851 30077 1897
rect 30147 1851 30193 1897
rect 30263 1851 30309 1897
rect 30379 1851 30425 1897
rect 30495 1851 30541 1897
rect 30611 1851 30657 1897
rect 30727 1851 30773 1897
rect 30843 1851 30889 1897
rect 30959 1851 31005 1897
rect 31075 1851 31121 1897
rect 31191 1851 31237 1897
rect 31307 1851 31353 1897
rect 31423 1851 31469 1897
rect 31539 1851 31585 1897
rect 31655 1851 31701 1897
rect 31771 1851 31817 1897
rect 31887 1851 31933 1897
rect 32003 1851 32049 1897
rect 32119 1851 32165 1897
rect 32235 1851 32281 1897
rect 32351 1851 32397 1897
rect 32467 1851 32513 1897
rect 32583 1851 32629 1897
rect 32699 1851 32745 1897
rect 32815 1851 32861 1897
rect 32931 1851 32977 1897
rect 33047 1851 33093 1897
rect 33163 1851 33209 1897
rect 33279 1851 33325 1897
rect 33395 1851 33441 1897
rect 33511 1851 33557 1897
rect 33627 1851 33673 1897
rect 33743 1851 33789 1897
rect 33859 1851 33905 1897
rect 33975 1851 34021 1897
rect 34091 1851 34137 1897
rect 34207 1851 34253 1897
rect 34323 1851 34369 1897
rect 34439 1851 34485 1897
rect 34555 1851 34601 1897
rect 34671 1851 34717 1897
rect 34787 1851 34833 1897
rect 34903 1851 34949 1897
rect 35019 1851 35065 1897
rect 35135 1851 35181 1897
rect 35251 1851 35297 1897
rect 35367 1851 35413 1897
rect 35483 1851 35529 1897
rect 35599 1851 35645 1897
rect 35715 1851 35761 1897
rect 35831 1851 35877 1897
rect 35947 1851 35993 1897
rect 36063 1851 36109 1897
rect 36179 1851 36225 1897
rect 36295 1851 36341 1897
rect 36411 1851 36457 1897
rect 36527 1851 36573 1897
rect 36643 1851 36689 1897
rect 36759 1851 36805 1897
rect 36875 1851 36921 1897
rect 36991 1851 37037 1897
rect 37107 1851 37153 1897
rect 37223 1851 37269 1897
rect 37339 1851 37385 1897
rect 37455 1851 37501 1897
rect 37571 1851 37617 1897
rect 37687 1851 37733 1897
rect 37803 1851 37849 1897
rect 37919 1851 37965 1897
rect 38035 1851 38081 1897
rect 38151 1851 38197 1897
rect 38267 1851 38313 1897
rect 38383 1851 38429 1897
rect 38499 1851 38545 1897
rect 38615 1851 38661 1897
rect 38731 1851 38777 1897
rect 38847 1851 38893 1897
rect 38963 1851 39009 1897
rect 39079 1851 39125 1897
rect 39195 1851 39241 1897
rect 39311 1851 39357 1897
rect 39427 1851 39473 1897
rect 39543 1851 39589 1897
rect 39659 1851 39705 1897
rect 39775 1851 39821 1897
rect 39891 1851 39937 1897
rect 40007 1851 40053 1897
rect 40123 1851 40169 1897
rect 28639 1735 28685 1781
rect 28755 1735 28801 1781
rect 28871 1735 28917 1781
rect 28987 1735 29033 1781
rect 29103 1735 29149 1781
rect 29219 1735 29265 1781
rect 29335 1735 29381 1781
rect 29451 1735 29497 1781
rect 29567 1735 29613 1781
rect 29683 1735 29729 1781
rect 29799 1735 29845 1781
rect 29915 1735 29961 1781
rect 30031 1735 30077 1781
rect 30147 1735 30193 1781
rect 30263 1735 30309 1781
rect 30379 1735 30425 1781
rect 30495 1735 30541 1781
rect 30611 1735 30657 1781
rect 30727 1735 30773 1781
rect 30843 1735 30889 1781
rect 30959 1735 31005 1781
rect 31075 1735 31121 1781
rect 31191 1735 31237 1781
rect 31307 1735 31353 1781
rect 31423 1735 31469 1781
rect 31539 1735 31585 1781
rect 31655 1735 31701 1781
rect 31771 1735 31817 1781
rect 31887 1735 31933 1781
rect 32003 1735 32049 1781
rect 32119 1735 32165 1781
rect 32235 1735 32281 1781
rect 32351 1735 32397 1781
rect 32467 1735 32513 1781
rect 32583 1735 32629 1781
rect 32699 1735 32745 1781
rect 32815 1735 32861 1781
rect 32931 1735 32977 1781
rect 33047 1735 33093 1781
rect 33163 1735 33209 1781
rect 33279 1735 33325 1781
rect 33395 1735 33441 1781
rect 33511 1735 33557 1781
rect 33627 1735 33673 1781
rect 33743 1735 33789 1781
rect 33859 1735 33905 1781
rect 33975 1735 34021 1781
rect 34091 1735 34137 1781
rect 34207 1735 34253 1781
rect 34323 1735 34369 1781
rect 34439 1735 34485 1781
rect 34555 1735 34601 1781
rect 34671 1735 34717 1781
rect 34787 1735 34833 1781
rect 34903 1735 34949 1781
rect 35019 1735 35065 1781
rect 35135 1735 35181 1781
rect 35251 1735 35297 1781
rect 35367 1735 35413 1781
rect 35483 1735 35529 1781
rect 35599 1735 35645 1781
rect 35715 1735 35761 1781
rect 35831 1735 35877 1781
rect 35947 1735 35993 1781
rect 36063 1735 36109 1781
rect 36179 1735 36225 1781
rect 36295 1735 36341 1781
rect 36411 1735 36457 1781
rect 36527 1735 36573 1781
rect 36643 1735 36689 1781
rect 36759 1735 36805 1781
rect 36875 1735 36921 1781
rect 36991 1735 37037 1781
rect 37107 1735 37153 1781
rect 37223 1735 37269 1781
rect 37339 1735 37385 1781
rect 37455 1735 37501 1781
rect 37571 1735 37617 1781
rect 37687 1735 37733 1781
rect 37803 1735 37849 1781
rect 37919 1735 37965 1781
rect 38035 1735 38081 1781
rect 38151 1735 38197 1781
rect 38267 1735 38313 1781
rect 38383 1735 38429 1781
rect 38499 1735 38545 1781
rect 38615 1735 38661 1781
rect 38731 1735 38777 1781
rect 38847 1735 38893 1781
rect 38963 1735 39009 1781
rect 39079 1735 39125 1781
rect 39195 1735 39241 1781
rect 39311 1735 39357 1781
rect 39427 1735 39473 1781
rect 39543 1735 39589 1781
rect 39659 1735 39705 1781
rect 39775 1735 39821 1781
rect 39891 1735 39937 1781
rect 40007 1735 40053 1781
rect 40123 1735 40169 1781
rect 28639 1619 28685 1665
rect 28755 1619 28801 1665
rect 28871 1619 28917 1665
rect 28987 1619 29033 1665
rect 29103 1619 29149 1665
rect 29219 1619 29265 1665
rect 29335 1619 29381 1665
rect 29451 1619 29497 1665
rect 29567 1619 29613 1665
rect 29683 1619 29729 1665
rect 29799 1619 29845 1665
rect 29915 1619 29961 1665
rect 30031 1619 30077 1665
rect 30147 1619 30193 1665
rect 30263 1619 30309 1665
rect 30379 1619 30425 1665
rect 30495 1619 30541 1665
rect 30611 1619 30657 1665
rect 30727 1619 30773 1665
rect 30843 1619 30889 1665
rect 30959 1619 31005 1665
rect 31075 1619 31121 1665
rect 31191 1619 31237 1665
rect 31307 1619 31353 1665
rect 31423 1619 31469 1665
rect 31539 1619 31585 1665
rect 31655 1619 31701 1665
rect 31771 1619 31817 1665
rect 31887 1619 31933 1665
rect 32003 1619 32049 1665
rect 32119 1619 32165 1665
rect 32235 1619 32281 1665
rect 32351 1619 32397 1665
rect 32467 1619 32513 1665
rect 32583 1619 32629 1665
rect 32699 1619 32745 1665
rect 32815 1619 32861 1665
rect 32931 1619 32977 1665
rect 33047 1619 33093 1665
rect 33163 1619 33209 1665
rect 33279 1619 33325 1665
rect 33395 1619 33441 1665
rect 33511 1619 33557 1665
rect 33627 1619 33673 1665
rect 33743 1619 33789 1665
rect 33859 1619 33905 1665
rect 33975 1619 34021 1665
rect 34091 1619 34137 1665
rect 34207 1619 34253 1665
rect 34323 1619 34369 1665
rect 34439 1619 34485 1665
rect 34555 1619 34601 1665
rect 34671 1619 34717 1665
rect 34787 1619 34833 1665
rect 34903 1619 34949 1665
rect 35019 1619 35065 1665
rect 35135 1619 35181 1665
rect 35251 1619 35297 1665
rect 35367 1619 35413 1665
rect 35483 1619 35529 1665
rect 35599 1619 35645 1665
rect 35715 1619 35761 1665
rect 35831 1619 35877 1665
rect 35947 1619 35993 1665
rect 36063 1619 36109 1665
rect 36179 1619 36225 1665
rect 36295 1619 36341 1665
rect 36411 1619 36457 1665
rect 36527 1619 36573 1665
rect 36643 1619 36689 1665
rect 36759 1619 36805 1665
rect 36875 1619 36921 1665
rect 36991 1619 37037 1665
rect 37107 1619 37153 1665
rect 37223 1619 37269 1665
rect 37339 1619 37385 1665
rect 37455 1619 37501 1665
rect 37571 1619 37617 1665
rect 37687 1619 37733 1665
rect 37803 1619 37849 1665
rect 37919 1619 37965 1665
rect 38035 1619 38081 1665
rect 38151 1619 38197 1665
rect 38267 1619 38313 1665
rect 38383 1619 38429 1665
rect 38499 1619 38545 1665
rect 38615 1619 38661 1665
rect 38731 1619 38777 1665
rect 38847 1619 38893 1665
rect 38963 1619 39009 1665
rect 39079 1619 39125 1665
rect 39195 1619 39241 1665
rect 39311 1619 39357 1665
rect 39427 1619 39473 1665
rect 39543 1619 39589 1665
rect 39659 1619 39705 1665
rect 39775 1619 39821 1665
rect 39891 1619 39937 1665
rect 40007 1619 40053 1665
rect 40123 1619 40169 1665
rect 28639 1503 28685 1549
rect 28755 1503 28801 1549
rect 28871 1503 28917 1549
rect 28987 1503 29033 1549
rect 29103 1503 29149 1549
rect 29219 1503 29265 1549
rect 29335 1503 29381 1549
rect 29451 1503 29497 1549
rect 29567 1503 29613 1549
rect 29683 1503 29729 1549
rect 29799 1503 29845 1549
rect 29915 1503 29961 1549
rect 30031 1503 30077 1549
rect 30147 1503 30193 1549
rect 30263 1503 30309 1549
rect 30379 1503 30425 1549
rect 30495 1503 30541 1549
rect 30611 1503 30657 1549
rect 30727 1503 30773 1549
rect 30843 1503 30889 1549
rect 30959 1503 31005 1549
rect 31075 1503 31121 1549
rect 31191 1503 31237 1549
rect 31307 1503 31353 1549
rect 31423 1503 31469 1549
rect 31539 1503 31585 1549
rect 31655 1503 31701 1549
rect 31771 1503 31817 1549
rect 31887 1503 31933 1549
rect 32003 1503 32049 1549
rect 32119 1503 32165 1549
rect 32235 1503 32281 1549
rect 32351 1503 32397 1549
rect 32467 1503 32513 1549
rect 32583 1503 32629 1549
rect 32699 1503 32745 1549
rect 32815 1503 32861 1549
rect 32931 1503 32977 1549
rect 33047 1503 33093 1549
rect 33163 1503 33209 1549
rect 33279 1503 33325 1549
rect 33395 1503 33441 1549
rect 33511 1503 33557 1549
rect 33627 1503 33673 1549
rect 33743 1503 33789 1549
rect 33859 1503 33905 1549
rect 33975 1503 34021 1549
rect 34091 1503 34137 1549
rect 34207 1503 34253 1549
rect 34323 1503 34369 1549
rect 34439 1503 34485 1549
rect 34555 1503 34601 1549
rect 34671 1503 34717 1549
rect 34787 1503 34833 1549
rect 34903 1503 34949 1549
rect 35019 1503 35065 1549
rect 35135 1503 35181 1549
rect 35251 1503 35297 1549
rect 35367 1503 35413 1549
rect 35483 1503 35529 1549
rect 35599 1503 35645 1549
rect 35715 1503 35761 1549
rect 35831 1503 35877 1549
rect 35947 1503 35993 1549
rect 36063 1503 36109 1549
rect 36179 1503 36225 1549
rect 36295 1503 36341 1549
rect 36411 1503 36457 1549
rect 36527 1503 36573 1549
rect 36643 1503 36689 1549
rect 36759 1503 36805 1549
rect 36875 1503 36921 1549
rect 36991 1503 37037 1549
rect 37107 1503 37153 1549
rect 37223 1503 37269 1549
rect 37339 1503 37385 1549
rect 37455 1503 37501 1549
rect 37571 1503 37617 1549
rect 37687 1503 37733 1549
rect 37803 1503 37849 1549
rect 37919 1503 37965 1549
rect 38035 1503 38081 1549
rect 38151 1503 38197 1549
rect 38267 1503 38313 1549
rect 38383 1503 38429 1549
rect 38499 1503 38545 1549
rect 38615 1503 38661 1549
rect 38731 1503 38777 1549
rect 38847 1503 38893 1549
rect 38963 1503 39009 1549
rect 39079 1503 39125 1549
rect 39195 1503 39241 1549
rect 39311 1503 39357 1549
rect 39427 1503 39473 1549
rect 39543 1503 39589 1549
rect 39659 1503 39705 1549
rect 39775 1503 39821 1549
rect 39891 1503 39937 1549
rect 40007 1503 40053 1549
rect 40123 1503 40169 1549
rect 28639 1387 28685 1433
rect 28755 1387 28801 1433
rect 28871 1387 28917 1433
rect 28987 1387 29033 1433
rect 29103 1387 29149 1433
rect 29219 1387 29265 1433
rect 29335 1387 29381 1433
rect 29451 1387 29497 1433
rect 29567 1387 29613 1433
rect 29683 1387 29729 1433
rect 29799 1387 29845 1433
rect 29915 1387 29961 1433
rect 30031 1387 30077 1433
rect 30147 1387 30193 1433
rect 30263 1387 30309 1433
rect 30379 1387 30425 1433
rect 30495 1387 30541 1433
rect 30611 1387 30657 1433
rect 30727 1387 30773 1433
rect 30843 1387 30889 1433
rect 30959 1387 31005 1433
rect 31075 1387 31121 1433
rect 31191 1387 31237 1433
rect 31307 1387 31353 1433
rect 31423 1387 31469 1433
rect 31539 1387 31585 1433
rect 31655 1387 31701 1433
rect 31771 1387 31817 1433
rect 31887 1387 31933 1433
rect 32003 1387 32049 1433
rect 32119 1387 32165 1433
rect 32235 1387 32281 1433
rect 32351 1387 32397 1433
rect 32467 1387 32513 1433
rect 32583 1387 32629 1433
rect 32699 1387 32745 1433
rect 32815 1387 32861 1433
rect 32931 1387 32977 1433
rect 33047 1387 33093 1433
rect 33163 1387 33209 1433
rect 33279 1387 33325 1433
rect 33395 1387 33441 1433
rect 33511 1387 33557 1433
rect 33627 1387 33673 1433
rect 33743 1387 33789 1433
rect 33859 1387 33905 1433
rect 33975 1387 34021 1433
rect 34091 1387 34137 1433
rect 34207 1387 34253 1433
rect 34323 1387 34369 1433
rect 34439 1387 34485 1433
rect 34555 1387 34601 1433
rect 34671 1387 34717 1433
rect 34787 1387 34833 1433
rect 34903 1387 34949 1433
rect 35019 1387 35065 1433
rect 35135 1387 35181 1433
rect 35251 1387 35297 1433
rect 35367 1387 35413 1433
rect 35483 1387 35529 1433
rect 35599 1387 35645 1433
rect 35715 1387 35761 1433
rect 35831 1387 35877 1433
rect 35947 1387 35993 1433
rect 36063 1387 36109 1433
rect 36179 1387 36225 1433
rect 36295 1387 36341 1433
rect 36411 1387 36457 1433
rect 36527 1387 36573 1433
rect 36643 1387 36689 1433
rect 36759 1387 36805 1433
rect 36875 1387 36921 1433
rect 36991 1387 37037 1433
rect 37107 1387 37153 1433
rect 37223 1387 37269 1433
rect 37339 1387 37385 1433
rect 37455 1387 37501 1433
rect 37571 1387 37617 1433
rect 37687 1387 37733 1433
rect 37803 1387 37849 1433
rect 37919 1387 37965 1433
rect 38035 1387 38081 1433
rect 38151 1387 38197 1433
rect 38267 1387 38313 1433
rect 38383 1387 38429 1433
rect 38499 1387 38545 1433
rect 38615 1387 38661 1433
rect 38731 1387 38777 1433
rect 38847 1387 38893 1433
rect 38963 1387 39009 1433
rect 39079 1387 39125 1433
rect 39195 1387 39241 1433
rect 39311 1387 39357 1433
rect 39427 1387 39473 1433
rect 39543 1387 39589 1433
rect 39659 1387 39705 1433
rect 39775 1387 39821 1433
rect 39891 1387 39937 1433
rect 40007 1387 40053 1433
rect 40123 1387 40169 1433
rect 28639 1271 28685 1317
rect 28755 1271 28801 1317
rect 28871 1271 28917 1317
rect 28987 1271 29033 1317
rect 29103 1271 29149 1317
rect 29219 1271 29265 1317
rect 29335 1271 29381 1317
rect 29451 1271 29497 1317
rect 29567 1271 29613 1317
rect 29683 1271 29729 1317
rect 29799 1271 29845 1317
rect 29915 1271 29961 1317
rect 30031 1271 30077 1317
rect 30147 1271 30193 1317
rect 30263 1271 30309 1317
rect 30379 1271 30425 1317
rect 30495 1271 30541 1317
rect 30611 1271 30657 1317
rect 30727 1271 30773 1317
rect 30843 1271 30889 1317
rect 30959 1271 31005 1317
rect 31075 1271 31121 1317
rect 31191 1271 31237 1317
rect 31307 1271 31353 1317
rect 31423 1271 31469 1317
rect 31539 1271 31585 1317
rect 31655 1271 31701 1317
rect 31771 1271 31817 1317
rect 31887 1271 31933 1317
rect 32003 1271 32049 1317
rect 32119 1271 32165 1317
rect 32235 1271 32281 1317
rect 32351 1271 32397 1317
rect 32467 1271 32513 1317
rect 32583 1271 32629 1317
rect 32699 1271 32745 1317
rect 32815 1271 32861 1317
rect 32931 1271 32977 1317
rect 33047 1271 33093 1317
rect 33163 1271 33209 1317
rect 33279 1271 33325 1317
rect 33395 1271 33441 1317
rect 33511 1271 33557 1317
rect 33627 1271 33673 1317
rect 33743 1271 33789 1317
rect 33859 1271 33905 1317
rect 33975 1271 34021 1317
rect 34091 1271 34137 1317
rect 34207 1271 34253 1317
rect 34323 1271 34369 1317
rect 34439 1271 34485 1317
rect 34555 1271 34601 1317
rect 34671 1271 34717 1317
rect 34787 1271 34833 1317
rect 34903 1271 34949 1317
rect 35019 1271 35065 1317
rect 35135 1271 35181 1317
rect 35251 1271 35297 1317
rect 35367 1271 35413 1317
rect 35483 1271 35529 1317
rect 35599 1271 35645 1317
rect 35715 1271 35761 1317
rect 35831 1271 35877 1317
rect 35947 1271 35993 1317
rect 36063 1271 36109 1317
rect 36179 1271 36225 1317
rect 36295 1271 36341 1317
rect 36411 1271 36457 1317
rect 36527 1271 36573 1317
rect 36643 1271 36689 1317
rect 36759 1271 36805 1317
rect 36875 1271 36921 1317
rect 36991 1271 37037 1317
rect 37107 1271 37153 1317
rect 37223 1271 37269 1317
rect 37339 1271 37385 1317
rect 37455 1271 37501 1317
rect 37571 1271 37617 1317
rect 37687 1271 37733 1317
rect 37803 1271 37849 1317
rect 37919 1271 37965 1317
rect 38035 1271 38081 1317
rect 38151 1271 38197 1317
rect 38267 1271 38313 1317
rect 38383 1271 38429 1317
rect 38499 1271 38545 1317
rect 38615 1271 38661 1317
rect 38731 1271 38777 1317
rect 38847 1271 38893 1317
rect 38963 1271 39009 1317
rect 39079 1271 39125 1317
rect 39195 1271 39241 1317
rect 39311 1271 39357 1317
rect 39427 1271 39473 1317
rect 39543 1271 39589 1317
rect 39659 1271 39705 1317
rect 39775 1271 39821 1317
rect 39891 1271 39937 1317
rect 40007 1271 40053 1317
rect 40123 1271 40169 1317
rect 28639 1155 28685 1201
rect 28755 1155 28801 1201
rect 28871 1155 28917 1201
rect 28987 1155 29033 1201
rect 29103 1155 29149 1201
rect 29219 1155 29265 1201
rect 29335 1155 29381 1201
rect 29451 1155 29497 1201
rect 29567 1155 29613 1201
rect 29683 1155 29729 1201
rect 29799 1155 29845 1201
rect 29915 1155 29961 1201
rect 30031 1155 30077 1201
rect 30147 1155 30193 1201
rect 30263 1155 30309 1201
rect 30379 1155 30425 1201
rect 30495 1155 30541 1201
rect 30611 1155 30657 1201
rect 30727 1155 30773 1201
rect 30843 1155 30889 1201
rect 30959 1155 31005 1201
rect 31075 1155 31121 1201
rect 31191 1155 31237 1201
rect 31307 1155 31353 1201
rect 31423 1155 31469 1201
rect 31539 1155 31585 1201
rect 31655 1155 31701 1201
rect 31771 1155 31817 1201
rect 31887 1155 31933 1201
rect 32003 1155 32049 1201
rect 32119 1155 32165 1201
rect 32235 1155 32281 1201
rect 32351 1155 32397 1201
rect 32467 1155 32513 1201
rect 32583 1155 32629 1201
rect 32699 1155 32745 1201
rect 32815 1155 32861 1201
rect 32931 1155 32977 1201
rect 33047 1155 33093 1201
rect 33163 1155 33209 1201
rect 33279 1155 33325 1201
rect 33395 1155 33441 1201
rect 33511 1155 33557 1201
rect 33627 1155 33673 1201
rect 33743 1155 33789 1201
rect 33859 1155 33905 1201
rect 33975 1155 34021 1201
rect 34091 1155 34137 1201
rect 34207 1155 34253 1201
rect 34323 1155 34369 1201
rect 34439 1155 34485 1201
rect 34555 1155 34601 1201
rect 34671 1155 34717 1201
rect 34787 1155 34833 1201
rect 34903 1155 34949 1201
rect 35019 1155 35065 1201
rect 35135 1155 35181 1201
rect 35251 1155 35297 1201
rect 35367 1155 35413 1201
rect 35483 1155 35529 1201
rect 35599 1155 35645 1201
rect 35715 1155 35761 1201
rect 35831 1155 35877 1201
rect 35947 1155 35993 1201
rect 36063 1155 36109 1201
rect 36179 1155 36225 1201
rect 36295 1155 36341 1201
rect 36411 1155 36457 1201
rect 36527 1155 36573 1201
rect 36643 1155 36689 1201
rect 36759 1155 36805 1201
rect 36875 1155 36921 1201
rect 36991 1155 37037 1201
rect 37107 1155 37153 1201
rect 37223 1155 37269 1201
rect 37339 1155 37385 1201
rect 37455 1155 37501 1201
rect 37571 1155 37617 1201
rect 37687 1155 37733 1201
rect 37803 1155 37849 1201
rect 37919 1155 37965 1201
rect 38035 1155 38081 1201
rect 38151 1155 38197 1201
rect 38267 1155 38313 1201
rect 38383 1155 38429 1201
rect 38499 1155 38545 1201
rect 38615 1155 38661 1201
rect 38731 1155 38777 1201
rect 38847 1155 38893 1201
rect 38963 1155 39009 1201
rect 39079 1155 39125 1201
rect 39195 1155 39241 1201
rect 39311 1155 39357 1201
rect 39427 1155 39473 1201
rect 39543 1155 39589 1201
rect 39659 1155 39705 1201
rect 39775 1155 39821 1201
rect 39891 1155 39937 1201
rect 40007 1155 40053 1201
rect 40123 1155 40169 1201
rect 50845 3844 50891 3890
rect 50961 3844 51007 3890
rect 51077 3844 51123 3890
rect 51193 3844 51239 3890
rect 51309 3844 51355 3890
rect 51425 3844 51471 3890
rect 51541 3844 51587 3890
rect 51657 3844 51703 3890
rect 51773 3844 51819 3890
rect 51889 3844 51935 3890
rect 52005 3844 52051 3890
rect 52121 3844 52167 3890
rect 52237 3844 52283 3890
rect 52353 3844 52399 3890
rect 52469 3844 52515 3890
rect 52585 3844 52631 3890
rect 52701 3844 52747 3890
rect 52817 3844 52863 3890
rect 52933 3844 52979 3890
rect 53049 3844 53095 3890
rect 53165 3844 53211 3890
rect 53281 3844 53327 3890
rect 53397 3844 53443 3890
rect 53513 3844 53559 3890
rect 53629 3844 53675 3890
rect 53745 3844 53791 3890
rect 53861 3844 53907 3890
rect 53977 3844 54023 3890
rect 54093 3844 54139 3890
rect 54209 3844 54255 3890
rect 54325 3844 54371 3890
rect 54441 3844 54487 3890
rect 54557 3844 54603 3890
rect 54673 3844 54719 3890
rect 54789 3844 54835 3890
rect 54905 3844 54951 3890
rect 55021 3844 55067 3890
rect 55137 3844 55183 3890
rect 55253 3844 55299 3890
rect 55369 3844 55415 3890
rect 55485 3844 55531 3890
rect 55601 3844 55647 3890
rect 55717 3844 55763 3890
rect 55833 3844 55879 3890
rect 55949 3844 55995 3890
rect 56065 3844 56111 3890
rect 56181 3844 56227 3890
rect 56297 3844 56343 3890
rect 56413 3844 56459 3890
rect 56529 3844 56575 3890
rect 50845 3728 50891 3774
rect 50961 3728 51007 3774
rect 51077 3728 51123 3774
rect 51193 3728 51239 3774
rect 51309 3728 51355 3774
rect 51425 3728 51471 3774
rect 51541 3728 51587 3774
rect 51657 3728 51703 3774
rect 51773 3728 51819 3774
rect 51889 3728 51935 3774
rect 52005 3728 52051 3774
rect 52121 3728 52167 3774
rect 52237 3728 52283 3774
rect 52353 3728 52399 3774
rect 52469 3728 52515 3774
rect 52585 3728 52631 3774
rect 52701 3728 52747 3774
rect 52817 3728 52863 3774
rect 52933 3728 52979 3774
rect 53049 3728 53095 3774
rect 53165 3728 53211 3774
rect 53281 3728 53327 3774
rect 53397 3728 53443 3774
rect 53513 3728 53559 3774
rect 53629 3728 53675 3774
rect 53745 3728 53791 3774
rect 53861 3728 53907 3774
rect 53977 3728 54023 3774
rect 54093 3728 54139 3774
rect 54209 3728 54255 3774
rect 54325 3728 54371 3774
rect 54441 3728 54487 3774
rect 54557 3728 54603 3774
rect 54673 3728 54719 3774
rect 54789 3728 54835 3774
rect 54905 3728 54951 3774
rect 55021 3728 55067 3774
rect 55137 3728 55183 3774
rect 55253 3728 55299 3774
rect 55369 3728 55415 3774
rect 55485 3728 55531 3774
rect 55601 3728 55647 3774
rect 55717 3728 55763 3774
rect 55833 3728 55879 3774
rect 55949 3728 55995 3774
rect 56065 3728 56111 3774
rect 56181 3728 56227 3774
rect 56297 3728 56343 3774
rect 56413 3728 56459 3774
rect 56529 3728 56575 3774
rect 50845 3612 50891 3658
rect 50961 3612 51007 3658
rect 51077 3612 51123 3658
rect 51193 3612 51239 3658
rect 51309 3612 51355 3658
rect 51425 3612 51471 3658
rect 51541 3612 51587 3658
rect 51657 3612 51703 3658
rect 51773 3612 51819 3658
rect 51889 3612 51935 3658
rect 52005 3612 52051 3658
rect 52121 3612 52167 3658
rect 52237 3612 52283 3658
rect 52353 3612 52399 3658
rect 52469 3612 52515 3658
rect 52585 3612 52631 3658
rect 52701 3612 52747 3658
rect 52817 3612 52863 3658
rect 52933 3612 52979 3658
rect 53049 3612 53095 3658
rect 53165 3612 53211 3658
rect 53281 3612 53327 3658
rect 53397 3612 53443 3658
rect 53513 3612 53559 3658
rect 53629 3612 53675 3658
rect 53745 3612 53791 3658
rect 53861 3612 53907 3658
rect 53977 3612 54023 3658
rect 54093 3612 54139 3658
rect 54209 3612 54255 3658
rect 54325 3612 54371 3658
rect 54441 3612 54487 3658
rect 54557 3612 54603 3658
rect 54673 3612 54719 3658
rect 54789 3612 54835 3658
rect 54905 3612 54951 3658
rect 55021 3612 55067 3658
rect 55137 3612 55183 3658
rect 55253 3612 55299 3658
rect 55369 3612 55415 3658
rect 55485 3612 55531 3658
rect 55601 3612 55647 3658
rect 55717 3612 55763 3658
rect 55833 3612 55879 3658
rect 55949 3612 55995 3658
rect 56065 3612 56111 3658
rect 56181 3612 56227 3658
rect 56297 3612 56343 3658
rect 56413 3612 56459 3658
rect 56529 3612 56575 3658
rect 50845 3496 50891 3542
rect 50961 3496 51007 3542
rect 51077 3496 51123 3542
rect 51193 3496 51239 3542
rect 51309 3496 51355 3542
rect 51425 3496 51471 3542
rect 51541 3496 51587 3542
rect 51657 3496 51703 3542
rect 51773 3496 51819 3542
rect 51889 3496 51935 3542
rect 52005 3496 52051 3542
rect 52121 3496 52167 3542
rect 52237 3496 52283 3542
rect 52353 3496 52399 3542
rect 52469 3496 52515 3542
rect 52585 3496 52631 3542
rect 52701 3496 52747 3542
rect 52817 3496 52863 3542
rect 52933 3496 52979 3542
rect 53049 3496 53095 3542
rect 53165 3496 53211 3542
rect 53281 3496 53327 3542
rect 53397 3496 53443 3542
rect 53513 3496 53559 3542
rect 53629 3496 53675 3542
rect 53745 3496 53791 3542
rect 53861 3496 53907 3542
rect 53977 3496 54023 3542
rect 54093 3496 54139 3542
rect 54209 3496 54255 3542
rect 54325 3496 54371 3542
rect 54441 3496 54487 3542
rect 54557 3496 54603 3542
rect 54673 3496 54719 3542
rect 54789 3496 54835 3542
rect 54905 3496 54951 3542
rect 55021 3496 55067 3542
rect 55137 3496 55183 3542
rect 55253 3496 55299 3542
rect 55369 3496 55415 3542
rect 55485 3496 55531 3542
rect 55601 3496 55647 3542
rect 55717 3496 55763 3542
rect 55833 3496 55879 3542
rect 55949 3496 55995 3542
rect 56065 3496 56111 3542
rect 56181 3496 56227 3542
rect 56297 3496 56343 3542
rect 56413 3496 56459 3542
rect 56529 3496 56575 3542
rect 50845 3380 50891 3426
rect 50961 3380 51007 3426
rect 51077 3380 51123 3426
rect 51193 3380 51239 3426
rect 51309 3380 51355 3426
rect 51425 3380 51471 3426
rect 51541 3380 51587 3426
rect 51657 3380 51703 3426
rect 51773 3380 51819 3426
rect 51889 3380 51935 3426
rect 52005 3380 52051 3426
rect 52121 3380 52167 3426
rect 52237 3380 52283 3426
rect 52353 3380 52399 3426
rect 52469 3380 52515 3426
rect 52585 3380 52631 3426
rect 52701 3380 52747 3426
rect 52817 3380 52863 3426
rect 52933 3380 52979 3426
rect 53049 3380 53095 3426
rect 53165 3380 53211 3426
rect 53281 3380 53327 3426
rect 53397 3380 53443 3426
rect 53513 3380 53559 3426
rect 53629 3380 53675 3426
rect 53745 3380 53791 3426
rect 53861 3380 53907 3426
rect 53977 3380 54023 3426
rect 54093 3380 54139 3426
rect 54209 3380 54255 3426
rect 54325 3380 54371 3426
rect 54441 3380 54487 3426
rect 54557 3380 54603 3426
rect 54673 3380 54719 3426
rect 54789 3380 54835 3426
rect 54905 3380 54951 3426
rect 55021 3380 55067 3426
rect 55137 3380 55183 3426
rect 55253 3380 55299 3426
rect 55369 3380 55415 3426
rect 55485 3380 55531 3426
rect 55601 3380 55647 3426
rect 55717 3380 55763 3426
rect 55833 3380 55879 3426
rect 55949 3380 55995 3426
rect 56065 3380 56111 3426
rect 56181 3380 56227 3426
rect 56297 3380 56343 3426
rect 56413 3380 56459 3426
rect 56529 3380 56575 3426
rect 50845 3264 50891 3310
rect 50961 3264 51007 3310
rect 51077 3264 51123 3310
rect 51193 3264 51239 3310
rect 51309 3264 51355 3310
rect 51425 3264 51471 3310
rect 51541 3264 51587 3310
rect 51657 3264 51703 3310
rect 51773 3264 51819 3310
rect 51889 3264 51935 3310
rect 52005 3264 52051 3310
rect 52121 3264 52167 3310
rect 52237 3264 52283 3310
rect 52353 3264 52399 3310
rect 52469 3264 52515 3310
rect 52585 3264 52631 3310
rect 52701 3264 52747 3310
rect 52817 3264 52863 3310
rect 52933 3264 52979 3310
rect 53049 3264 53095 3310
rect 53165 3264 53211 3310
rect 53281 3264 53327 3310
rect 53397 3264 53443 3310
rect 53513 3264 53559 3310
rect 53629 3264 53675 3310
rect 53745 3264 53791 3310
rect 53861 3264 53907 3310
rect 53977 3264 54023 3310
rect 54093 3264 54139 3310
rect 54209 3264 54255 3310
rect 54325 3264 54371 3310
rect 54441 3264 54487 3310
rect 54557 3264 54603 3310
rect 54673 3264 54719 3310
rect 54789 3264 54835 3310
rect 54905 3264 54951 3310
rect 55021 3264 55067 3310
rect 55137 3264 55183 3310
rect 55253 3264 55299 3310
rect 55369 3264 55415 3310
rect 55485 3264 55531 3310
rect 55601 3264 55647 3310
rect 55717 3264 55763 3310
rect 55833 3264 55879 3310
rect 55949 3264 55995 3310
rect 56065 3264 56111 3310
rect 56181 3264 56227 3310
rect 56297 3264 56343 3310
rect 56413 3264 56459 3310
rect 56529 3264 56575 3310
rect 50845 3148 50891 3194
rect 50961 3148 51007 3194
rect 51077 3148 51123 3194
rect 51193 3148 51239 3194
rect 51309 3148 51355 3194
rect 51425 3148 51471 3194
rect 51541 3148 51587 3194
rect 51657 3148 51703 3194
rect 51773 3148 51819 3194
rect 51889 3148 51935 3194
rect 52005 3148 52051 3194
rect 52121 3148 52167 3194
rect 52237 3148 52283 3194
rect 52353 3148 52399 3194
rect 52469 3148 52515 3194
rect 52585 3148 52631 3194
rect 52701 3148 52747 3194
rect 52817 3148 52863 3194
rect 52933 3148 52979 3194
rect 53049 3148 53095 3194
rect 53165 3148 53211 3194
rect 53281 3148 53327 3194
rect 53397 3148 53443 3194
rect 53513 3148 53559 3194
rect 53629 3148 53675 3194
rect 53745 3148 53791 3194
rect 53861 3148 53907 3194
rect 53977 3148 54023 3194
rect 54093 3148 54139 3194
rect 54209 3148 54255 3194
rect 54325 3148 54371 3194
rect 54441 3148 54487 3194
rect 54557 3148 54603 3194
rect 54673 3148 54719 3194
rect 54789 3148 54835 3194
rect 54905 3148 54951 3194
rect 55021 3148 55067 3194
rect 55137 3148 55183 3194
rect 55253 3148 55299 3194
rect 55369 3148 55415 3194
rect 55485 3148 55531 3194
rect 55601 3148 55647 3194
rect 55717 3148 55763 3194
rect 55833 3148 55879 3194
rect 55949 3148 55995 3194
rect 56065 3148 56111 3194
rect 56181 3148 56227 3194
rect 56297 3148 56343 3194
rect 56413 3148 56459 3194
rect 56529 3148 56575 3194
rect 50845 3032 50891 3078
rect 50961 3032 51007 3078
rect 51077 3032 51123 3078
rect 51193 3032 51239 3078
rect 51309 3032 51355 3078
rect 51425 3032 51471 3078
rect 51541 3032 51587 3078
rect 51657 3032 51703 3078
rect 51773 3032 51819 3078
rect 51889 3032 51935 3078
rect 52005 3032 52051 3078
rect 52121 3032 52167 3078
rect 52237 3032 52283 3078
rect 52353 3032 52399 3078
rect 52469 3032 52515 3078
rect 52585 3032 52631 3078
rect 52701 3032 52747 3078
rect 52817 3032 52863 3078
rect 52933 3032 52979 3078
rect 53049 3032 53095 3078
rect 53165 3032 53211 3078
rect 53281 3032 53327 3078
rect 53397 3032 53443 3078
rect 53513 3032 53559 3078
rect 53629 3032 53675 3078
rect 53745 3032 53791 3078
rect 53861 3032 53907 3078
rect 53977 3032 54023 3078
rect 54093 3032 54139 3078
rect 54209 3032 54255 3078
rect 54325 3032 54371 3078
rect 54441 3032 54487 3078
rect 54557 3032 54603 3078
rect 54673 3032 54719 3078
rect 54789 3032 54835 3078
rect 54905 3032 54951 3078
rect 55021 3032 55067 3078
rect 55137 3032 55183 3078
rect 55253 3032 55299 3078
rect 55369 3032 55415 3078
rect 55485 3032 55531 3078
rect 55601 3032 55647 3078
rect 55717 3032 55763 3078
rect 55833 3032 55879 3078
rect 55949 3032 55995 3078
rect 56065 3032 56111 3078
rect 56181 3032 56227 3078
rect 56297 3032 56343 3078
rect 56413 3032 56459 3078
rect 56529 3032 56575 3078
rect 50845 2916 50891 2962
rect 50961 2916 51007 2962
rect 51077 2916 51123 2962
rect 51193 2916 51239 2962
rect 51309 2916 51355 2962
rect 51425 2916 51471 2962
rect 51541 2916 51587 2962
rect 51657 2916 51703 2962
rect 51773 2916 51819 2962
rect 51889 2916 51935 2962
rect 52005 2916 52051 2962
rect 52121 2916 52167 2962
rect 52237 2916 52283 2962
rect 52353 2916 52399 2962
rect 52469 2916 52515 2962
rect 52585 2916 52631 2962
rect 52701 2916 52747 2962
rect 52817 2916 52863 2962
rect 52933 2916 52979 2962
rect 53049 2916 53095 2962
rect 53165 2916 53211 2962
rect 53281 2916 53327 2962
rect 53397 2916 53443 2962
rect 53513 2916 53559 2962
rect 53629 2916 53675 2962
rect 53745 2916 53791 2962
rect 53861 2916 53907 2962
rect 53977 2916 54023 2962
rect 54093 2916 54139 2962
rect 54209 2916 54255 2962
rect 54325 2916 54371 2962
rect 54441 2916 54487 2962
rect 54557 2916 54603 2962
rect 54673 2916 54719 2962
rect 54789 2916 54835 2962
rect 54905 2916 54951 2962
rect 55021 2916 55067 2962
rect 55137 2916 55183 2962
rect 55253 2916 55299 2962
rect 55369 2916 55415 2962
rect 55485 2916 55531 2962
rect 55601 2916 55647 2962
rect 55717 2916 55763 2962
rect 55833 2916 55879 2962
rect 55949 2916 55995 2962
rect 56065 2916 56111 2962
rect 56181 2916 56227 2962
rect 56297 2916 56343 2962
rect 56413 2916 56459 2962
rect 56529 2916 56575 2962
rect 50845 2800 50891 2846
rect 50961 2800 51007 2846
rect 51077 2800 51123 2846
rect 51193 2800 51239 2846
rect 51309 2800 51355 2846
rect 51425 2800 51471 2846
rect 51541 2800 51587 2846
rect 51657 2800 51703 2846
rect 51773 2800 51819 2846
rect 51889 2800 51935 2846
rect 52005 2800 52051 2846
rect 52121 2800 52167 2846
rect 52237 2800 52283 2846
rect 52353 2800 52399 2846
rect 52469 2800 52515 2846
rect 52585 2800 52631 2846
rect 52701 2800 52747 2846
rect 52817 2800 52863 2846
rect 52933 2800 52979 2846
rect 53049 2800 53095 2846
rect 53165 2800 53211 2846
rect 53281 2800 53327 2846
rect 53397 2800 53443 2846
rect 53513 2800 53559 2846
rect 53629 2800 53675 2846
rect 53745 2800 53791 2846
rect 53861 2800 53907 2846
rect 53977 2800 54023 2846
rect 54093 2800 54139 2846
rect 54209 2800 54255 2846
rect 54325 2800 54371 2846
rect 54441 2800 54487 2846
rect 54557 2800 54603 2846
rect 54673 2800 54719 2846
rect 54789 2800 54835 2846
rect 54905 2800 54951 2846
rect 55021 2800 55067 2846
rect 55137 2800 55183 2846
rect 55253 2800 55299 2846
rect 55369 2800 55415 2846
rect 55485 2800 55531 2846
rect 55601 2800 55647 2846
rect 55717 2800 55763 2846
rect 55833 2800 55879 2846
rect 55949 2800 55995 2846
rect 56065 2800 56111 2846
rect 56181 2800 56227 2846
rect 56297 2800 56343 2846
rect 56413 2800 56459 2846
rect 56529 2800 56575 2846
rect 50845 2684 50891 2730
rect 50961 2684 51007 2730
rect 51077 2684 51123 2730
rect 51193 2684 51239 2730
rect 51309 2684 51355 2730
rect 51425 2684 51471 2730
rect 51541 2684 51587 2730
rect 51657 2684 51703 2730
rect 51773 2684 51819 2730
rect 51889 2684 51935 2730
rect 52005 2684 52051 2730
rect 52121 2684 52167 2730
rect 52237 2684 52283 2730
rect 52353 2684 52399 2730
rect 52469 2684 52515 2730
rect 52585 2684 52631 2730
rect 52701 2684 52747 2730
rect 52817 2684 52863 2730
rect 52933 2684 52979 2730
rect 53049 2684 53095 2730
rect 53165 2684 53211 2730
rect 53281 2684 53327 2730
rect 53397 2684 53443 2730
rect 53513 2684 53559 2730
rect 53629 2684 53675 2730
rect 53745 2684 53791 2730
rect 53861 2684 53907 2730
rect 53977 2684 54023 2730
rect 54093 2684 54139 2730
rect 54209 2684 54255 2730
rect 54325 2684 54371 2730
rect 54441 2684 54487 2730
rect 54557 2684 54603 2730
rect 54673 2684 54719 2730
rect 54789 2684 54835 2730
rect 54905 2684 54951 2730
rect 55021 2684 55067 2730
rect 55137 2684 55183 2730
rect 55253 2684 55299 2730
rect 55369 2684 55415 2730
rect 55485 2684 55531 2730
rect 55601 2684 55647 2730
rect 55717 2684 55763 2730
rect 55833 2684 55879 2730
rect 55949 2684 55995 2730
rect 56065 2684 56111 2730
rect 56181 2684 56227 2730
rect 56297 2684 56343 2730
rect 56413 2684 56459 2730
rect 56529 2684 56575 2730
rect 50845 2568 50891 2614
rect 50961 2568 51007 2614
rect 51077 2568 51123 2614
rect 51193 2568 51239 2614
rect 51309 2568 51355 2614
rect 51425 2568 51471 2614
rect 51541 2568 51587 2614
rect 51657 2568 51703 2614
rect 51773 2568 51819 2614
rect 51889 2568 51935 2614
rect 52005 2568 52051 2614
rect 52121 2568 52167 2614
rect 52237 2568 52283 2614
rect 52353 2568 52399 2614
rect 52469 2568 52515 2614
rect 52585 2568 52631 2614
rect 52701 2568 52747 2614
rect 52817 2568 52863 2614
rect 52933 2568 52979 2614
rect 53049 2568 53095 2614
rect 53165 2568 53211 2614
rect 53281 2568 53327 2614
rect 53397 2568 53443 2614
rect 53513 2568 53559 2614
rect 53629 2568 53675 2614
rect 53745 2568 53791 2614
rect 53861 2568 53907 2614
rect 53977 2568 54023 2614
rect 54093 2568 54139 2614
rect 54209 2568 54255 2614
rect 54325 2568 54371 2614
rect 54441 2568 54487 2614
rect 54557 2568 54603 2614
rect 54673 2568 54719 2614
rect 54789 2568 54835 2614
rect 54905 2568 54951 2614
rect 55021 2568 55067 2614
rect 55137 2568 55183 2614
rect 55253 2568 55299 2614
rect 55369 2568 55415 2614
rect 55485 2568 55531 2614
rect 55601 2568 55647 2614
rect 55717 2568 55763 2614
rect 55833 2568 55879 2614
rect 55949 2568 55995 2614
rect 56065 2568 56111 2614
rect 56181 2568 56227 2614
rect 56297 2568 56343 2614
rect 56413 2568 56459 2614
rect 56529 2568 56575 2614
rect 50845 2452 50891 2498
rect 50961 2452 51007 2498
rect 51077 2452 51123 2498
rect 51193 2452 51239 2498
rect 51309 2452 51355 2498
rect 51425 2452 51471 2498
rect 51541 2452 51587 2498
rect 51657 2452 51703 2498
rect 51773 2452 51819 2498
rect 51889 2452 51935 2498
rect 52005 2452 52051 2498
rect 52121 2452 52167 2498
rect 52237 2452 52283 2498
rect 52353 2452 52399 2498
rect 52469 2452 52515 2498
rect 52585 2452 52631 2498
rect 52701 2452 52747 2498
rect 52817 2452 52863 2498
rect 52933 2452 52979 2498
rect 53049 2452 53095 2498
rect 53165 2452 53211 2498
rect 53281 2452 53327 2498
rect 53397 2452 53443 2498
rect 53513 2452 53559 2498
rect 53629 2452 53675 2498
rect 53745 2452 53791 2498
rect 53861 2452 53907 2498
rect 53977 2452 54023 2498
rect 54093 2452 54139 2498
rect 54209 2452 54255 2498
rect 54325 2452 54371 2498
rect 54441 2452 54487 2498
rect 54557 2452 54603 2498
rect 54673 2452 54719 2498
rect 54789 2452 54835 2498
rect 54905 2452 54951 2498
rect 55021 2452 55067 2498
rect 55137 2452 55183 2498
rect 55253 2452 55299 2498
rect 55369 2452 55415 2498
rect 55485 2452 55531 2498
rect 55601 2452 55647 2498
rect 55717 2452 55763 2498
rect 55833 2452 55879 2498
rect 55949 2452 55995 2498
rect 56065 2452 56111 2498
rect 56181 2452 56227 2498
rect 56297 2452 56343 2498
rect 56413 2452 56459 2498
rect 56529 2452 56575 2498
rect 50845 2336 50891 2382
rect 50961 2336 51007 2382
rect 51077 2336 51123 2382
rect 51193 2336 51239 2382
rect 51309 2336 51355 2382
rect 51425 2336 51471 2382
rect 51541 2336 51587 2382
rect 51657 2336 51703 2382
rect 51773 2336 51819 2382
rect 51889 2336 51935 2382
rect 52005 2336 52051 2382
rect 52121 2336 52167 2382
rect 52237 2336 52283 2382
rect 52353 2336 52399 2382
rect 52469 2336 52515 2382
rect 52585 2336 52631 2382
rect 52701 2336 52747 2382
rect 52817 2336 52863 2382
rect 52933 2336 52979 2382
rect 53049 2336 53095 2382
rect 53165 2336 53211 2382
rect 53281 2336 53327 2382
rect 53397 2336 53443 2382
rect 53513 2336 53559 2382
rect 53629 2336 53675 2382
rect 53745 2336 53791 2382
rect 53861 2336 53907 2382
rect 53977 2336 54023 2382
rect 54093 2336 54139 2382
rect 54209 2336 54255 2382
rect 54325 2336 54371 2382
rect 54441 2336 54487 2382
rect 54557 2336 54603 2382
rect 54673 2336 54719 2382
rect 54789 2336 54835 2382
rect 54905 2336 54951 2382
rect 55021 2336 55067 2382
rect 55137 2336 55183 2382
rect 55253 2336 55299 2382
rect 55369 2336 55415 2382
rect 55485 2336 55531 2382
rect 55601 2336 55647 2382
rect 55717 2336 55763 2382
rect 55833 2336 55879 2382
rect 55949 2336 55995 2382
rect 56065 2336 56111 2382
rect 56181 2336 56227 2382
rect 56297 2336 56343 2382
rect 56413 2336 56459 2382
rect 56529 2336 56575 2382
rect 50845 2220 50891 2266
rect 50961 2220 51007 2266
rect 51077 2220 51123 2266
rect 51193 2220 51239 2266
rect 51309 2220 51355 2266
rect 51425 2220 51471 2266
rect 51541 2220 51587 2266
rect 51657 2220 51703 2266
rect 51773 2220 51819 2266
rect 51889 2220 51935 2266
rect 52005 2220 52051 2266
rect 52121 2220 52167 2266
rect 52237 2220 52283 2266
rect 52353 2220 52399 2266
rect 52469 2220 52515 2266
rect 52585 2220 52631 2266
rect 52701 2220 52747 2266
rect 52817 2220 52863 2266
rect 52933 2220 52979 2266
rect 53049 2220 53095 2266
rect 53165 2220 53211 2266
rect 53281 2220 53327 2266
rect 53397 2220 53443 2266
rect 53513 2220 53559 2266
rect 53629 2220 53675 2266
rect 53745 2220 53791 2266
rect 53861 2220 53907 2266
rect 53977 2220 54023 2266
rect 54093 2220 54139 2266
rect 54209 2220 54255 2266
rect 54325 2220 54371 2266
rect 54441 2220 54487 2266
rect 54557 2220 54603 2266
rect 54673 2220 54719 2266
rect 54789 2220 54835 2266
rect 54905 2220 54951 2266
rect 55021 2220 55067 2266
rect 55137 2220 55183 2266
rect 55253 2220 55299 2266
rect 55369 2220 55415 2266
rect 55485 2220 55531 2266
rect 55601 2220 55647 2266
rect 55717 2220 55763 2266
rect 55833 2220 55879 2266
rect 55949 2220 55995 2266
rect 56065 2220 56111 2266
rect 56181 2220 56227 2266
rect 56297 2220 56343 2266
rect 56413 2220 56459 2266
rect 56529 2220 56575 2266
rect 50845 2104 50891 2150
rect 50961 2104 51007 2150
rect 51077 2104 51123 2150
rect 51193 2104 51239 2150
rect 51309 2104 51355 2150
rect 51425 2104 51471 2150
rect 51541 2104 51587 2150
rect 51657 2104 51703 2150
rect 51773 2104 51819 2150
rect 51889 2104 51935 2150
rect 52005 2104 52051 2150
rect 52121 2104 52167 2150
rect 52237 2104 52283 2150
rect 52353 2104 52399 2150
rect 52469 2104 52515 2150
rect 52585 2104 52631 2150
rect 52701 2104 52747 2150
rect 52817 2104 52863 2150
rect 52933 2104 52979 2150
rect 53049 2104 53095 2150
rect 53165 2104 53211 2150
rect 53281 2104 53327 2150
rect 53397 2104 53443 2150
rect 53513 2104 53559 2150
rect 53629 2104 53675 2150
rect 53745 2104 53791 2150
rect 53861 2104 53907 2150
rect 53977 2104 54023 2150
rect 54093 2104 54139 2150
rect 54209 2104 54255 2150
rect 54325 2104 54371 2150
rect 54441 2104 54487 2150
rect 54557 2104 54603 2150
rect 54673 2104 54719 2150
rect 54789 2104 54835 2150
rect 54905 2104 54951 2150
rect 55021 2104 55067 2150
rect 55137 2104 55183 2150
rect 55253 2104 55299 2150
rect 55369 2104 55415 2150
rect 55485 2104 55531 2150
rect 55601 2104 55647 2150
rect 55717 2104 55763 2150
rect 55833 2104 55879 2150
rect 55949 2104 55995 2150
rect 56065 2104 56111 2150
rect 56181 2104 56227 2150
rect 56297 2104 56343 2150
rect 56413 2104 56459 2150
rect 56529 2104 56575 2150
rect 50845 1988 50891 2034
rect 50961 1988 51007 2034
rect 51077 1988 51123 2034
rect 51193 1988 51239 2034
rect 51309 1988 51355 2034
rect 51425 1988 51471 2034
rect 51541 1988 51587 2034
rect 51657 1988 51703 2034
rect 51773 1988 51819 2034
rect 51889 1988 51935 2034
rect 52005 1988 52051 2034
rect 52121 1988 52167 2034
rect 52237 1988 52283 2034
rect 52353 1988 52399 2034
rect 52469 1988 52515 2034
rect 52585 1988 52631 2034
rect 52701 1988 52747 2034
rect 52817 1988 52863 2034
rect 52933 1988 52979 2034
rect 53049 1988 53095 2034
rect 53165 1988 53211 2034
rect 53281 1988 53327 2034
rect 53397 1988 53443 2034
rect 53513 1988 53559 2034
rect 53629 1988 53675 2034
rect 53745 1988 53791 2034
rect 53861 1988 53907 2034
rect 53977 1988 54023 2034
rect 54093 1988 54139 2034
rect 54209 1988 54255 2034
rect 54325 1988 54371 2034
rect 54441 1988 54487 2034
rect 54557 1988 54603 2034
rect 54673 1988 54719 2034
rect 54789 1988 54835 2034
rect 54905 1988 54951 2034
rect 55021 1988 55067 2034
rect 55137 1988 55183 2034
rect 55253 1988 55299 2034
rect 55369 1988 55415 2034
rect 55485 1988 55531 2034
rect 55601 1988 55647 2034
rect 55717 1988 55763 2034
rect 55833 1988 55879 2034
rect 55949 1988 55995 2034
rect 56065 1988 56111 2034
rect 56181 1988 56227 2034
rect 56297 1988 56343 2034
rect 56413 1988 56459 2034
rect 56529 1988 56575 2034
rect 50845 1872 50891 1918
rect 50961 1872 51007 1918
rect 51077 1872 51123 1918
rect 51193 1872 51239 1918
rect 51309 1872 51355 1918
rect 51425 1872 51471 1918
rect 51541 1872 51587 1918
rect 51657 1872 51703 1918
rect 51773 1872 51819 1918
rect 51889 1872 51935 1918
rect 52005 1872 52051 1918
rect 52121 1872 52167 1918
rect 52237 1872 52283 1918
rect 52353 1872 52399 1918
rect 52469 1872 52515 1918
rect 52585 1872 52631 1918
rect 52701 1872 52747 1918
rect 52817 1872 52863 1918
rect 52933 1872 52979 1918
rect 53049 1872 53095 1918
rect 53165 1872 53211 1918
rect 53281 1872 53327 1918
rect 53397 1872 53443 1918
rect 53513 1872 53559 1918
rect 53629 1872 53675 1918
rect 53745 1872 53791 1918
rect 53861 1872 53907 1918
rect 53977 1872 54023 1918
rect 54093 1872 54139 1918
rect 54209 1872 54255 1918
rect 54325 1872 54371 1918
rect 54441 1872 54487 1918
rect 54557 1872 54603 1918
rect 54673 1872 54719 1918
rect 54789 1872 54835 1918
rect 54905 1872 54951 1918
rect 55021 1872 55067 1918
rect 55137 1872 55183 1918
rect 55253 1872 55299 1918
rect 55369 1872 55415 1918
rect 55485 1872 55531 1918
rect 55601 1872 55647 1918
rect 55717 1872 55763 1918
rect 55833 1872 55879 1918
rect 55949 1872 55995 1918
rect 56065 1872 56111 1918
rect 56181 1872 56227 1918
rect 56297 1872 56343 1918
rect 56413 1872 56459 1918
rect 56529 1872 56575 1918
rect 50845 1756 50891 1802
rect 50961 1756 51007 1802
rect 51077 1756 51123 1802
rect 51193 1756 51239 1802
rect 51309 1756 51355 1802
rect 51425 1756 51471 1802
rect 51541 1756 51587 1802
rect 51657 1756 51703 1802
rect 51773 1756 51819 1802
rect 51889 1756 51935 1802
rect 52005 1756 52051 1802
rect 52121 1756 52167 1802
rect 52237 1756 52283 1802
rect 52353 1756 52399 1802
rect 52469 1756 52515 1802
rect 52585 1756 52631 1802
rect 52701 1756 52747 1802
rect 52817 1756 52863 1802
rect 52933 1756 52979 1802
rect 53049 1756 53095 1802
rect 53165 1756 53211 1802
rect 53281 1756 53327 1802
rect 53397 1756 53443 1802
rect 53513 1756 53559 1802
rect 53629 1756 53675 1802
rect 53745 1756 53791 1802
rect 53861 1756 53907 1802
rect 53977 1756 54023 1802
rect 54093 1756 54139 1802
rect 54209 1756 54255 1802
rect 54325 1756 54371 1802
rect 54441 1756 54487 1802
rect 54557 1756 54603 1802
rect 54673 1756 54719 1802
rect 54789 1756 54835 1802
rect 54905 1756 54951 1802
rect 55021 1756 55067 1802
rect 55137 1756 55183 1802
rect 55253 1756 55299 1802
rect 55369 1756 55415 1802
rect 55485 1756 55531 1802
rect 55601 1756 55647 1802
rect 55717 1756 55763 1802
rect 55833 1756 55879 1802
rect 55949 1756 55995 1802
rect 56065 1756 56111 1802
rect 56181 1756 56227 1802
rect 56297 1756 56343 1802
rect 56413 1756 56459 1802
rect 56529 1756 56575 1802
rect 50845 1640 50891 1686
rect 50961 1640 51007 1686
rect 51077 1640 51123 1686
rect 51193 1640 51239 1686
rect 51309 1640 51355 1686
rect 51425 1640 51471 1686
rect 51541 1640 51587 1686
rect 51657 1640 51703 1686
rect 51773 1640 51819 1686
rect 51889 1640 51935 1686
rect 52005 1640 52051 1686
rect 52121 1640 52167 1686
rect 52237 1640 52283 1686
rect 52353 1640 52399 1686
rect 52469 1640 52515 1686
rect 52585 1640 52631 1686
rect 52701 1640 52747 1686
rect 52817 1640 52863 1686
rect 52933 1640 52979 1686
rect 53049 1640 53095 1686
rect 53165 1640 53211 1686
rect 53281 1640 53327 1686
rect 53397 1640 53443 1686
rect 53513 1640 53559 1686
rect 53629 1640 53675 1686
rect 53745 1640 53791 1686
rect 53861 1640 53907 1686
rect 53977 1640 54023 1686
rect 54093 1640 54139 1686
rect 54209 1640 54255 1686
rect 54325 1640 54371 1686
rect 54441 1640 54487 1686
rect 54557 1640 54603 1686
rect 54673 1640 54719 1686
rect 54789 1640 54835 1686
rect 54905 1640 54951 1686
rect 55021 1640 55067 1686
rect 55137 1640 55183 1686
rect 55253 1640 55299 1686
rect 55369 1640 55415 1686
rect 55485 1640 55531 1686
rect 55601 1640 55647 1686
rect 55717 1640 55763 1686
rect 55833 1640 55879 1686
rect 55949 1640 55995 1686
rect 56065 1640 56111 1686
rect 56181 1640 56227 1686
rect 56297 1640 56343 1686
rect 56413 1640 56459 1686
rect 56529 1640 56575 1686
rect 50845 1524 50891 1570
rect 50961 1524 51007 1570
rect 51077 1524 51123 1570
rect 51193 1524 51239 1570
rect 51309 1524 51355 1570
rect 51425 1524 51471 1570
rect 51541 1524 51587 1570
rect 51657 1524 51703 1570
rect 51773 1524 51819 1570
rect 51889 1524 51935 1570
rect 52005 1524 52051 1570
rect 52121 1524 52167 1570
rect 52237 1524 52283 1570
rect 52353 1524 52399 1570
rect 52469 1524 52515 1570
rect 52585 1524 52631 1570
rect 52701 1524 52747 1570
rect 52817 1524 52863 1570
rect 52933 1524 52979 1570
rect 53049 1524 53095 1570
rect 53165 1524 53211 1570
rect 53281 1524 53327 1570
rect 53397 1524 53443 1570
rect 53513 1524 53559 1570
rect 53629 1524 53675 1570
rect 53745 1524 53791 1570
rect 53861 1524 53907 1570
rect 53977 1524 54023 1570
rect 54093 1524 54139 1570
rect 54209 1524 54255 1570
rect 54325 1524 54371 1570
rect 54441 1524 54487 1570
rect 54557 1524 54603 1570
rect 54673 1524 54719 1570
rect 54789 1524 54835 1570
rect 54905 1524 54951 1570
rect 55021 1524 55067 1570
rect 55137 1524 55183 1570
rect 55253 1524 55299 1570
rect 55369 1524 55415 1570
rect 55485 1524 55531 1570
rect 55601 1524 55647 1570
rect 55717 1524 55763 1570
rect 55833 1524 55879 1570
rect 55949 1524 55995 1570
rect 56065 1524 56111 1570
rect 56181 1524 56227 1570
rect 56297 1524 56343 1570
rect 56413 1524 56459 1570
rect 56529 1524 56575 1570
rect 50845 1408 50891 1454
rect 50961 1408 51007 1454
rect 51077 1408 51123 1454
rect 51193 1408 51239 1454
rect 51309 1408 51355 1454
rect 51425 1408 51471 1454
rect 51541 1408 51587 1454
rect 51657 1408 51703 1454
rect 51773 1408 51819 1454
rect 51889 1408 51935 1454
rect 52005 1408 52051 1454
rect 52121 1408 52167 1454
rect 52237 1408 52283 1454
rect 52353 1408 52399 1454
rect 52469 1408 52515 1454
rect 52585 1408 52631 1454
rect 52701 1408 52747 1454
rect 52817 1408 52863 1454
rect 52933 1408 52979 1454
rect 53049 1408 53095 1454
rect 53165 1408 53211 1454
rect 53281 1408 53327 1454
rect 53397 1408 53443 1454
rect 53513 1408 53559 1454
rect 53629 1408 53675 1454
rect 53745 1408 53791 1454
rect 53861 1408 53907 1454
rect 53977 1408 54023 1454
rect 54093 1408 54139 1454
rect 54209 1408 54255 1454
rect 54325 1408 54371 1454
rect 54441 1408 54487 1454
rect 54557 1408 54603 1454
rect 54673 1408 54719 1454
rect 54789 1408 54835 1454
rect 54905 1408 54951 1454
rect 55021 1408 55067 1454
rect 55137 1408 55183 1454
rect 55253 1408 55299 1454
rect 55369 1408 55415 1454
rect 55485 1408 55531 1454
rect 55601 1408 55647 1454
rect 55717 1408 55763 1454
rect 55833 1408 55879 1454
rect 55949 1408 55995 1454
rect 56065 1408 56111 1454
rect 56181 1408 56227 1454
rect 56297 1408 56343 1454
rect 56413 1408 56459 1454
rect 56529 1408 56575 1454
rect 50845 1292 50891 1338
rect 50961 1292 51007 1338
rect 51077 1292 51123 1338
rect 51193 1292 51239 1338
rect 51309 1292 51355 1338
rect 51425 1292 51471 1338
rect 51541 1292 51587 1338
rect 51657 1292 51703 1338
rect 51773 1292 51819 1338
rect 51889 1292 51935 1338
rect 52005 1292 52051 1338
rect 52121 1292 52167 1338
rect 52237 1292 52283 1338
rect 52353 1292 52399 1338
rect 52469 1292 52515 1338
rect 52585 1292 52631 1338
rect 52701 1292 52747 1338
rect 52817 1292 52863 1338
rect 52933 1292 52979 1338
rect 53049 1292 53095 1338
rect 53165 1292 53211 1338
rect 53281 1292 53327 1338
rect 53397 1292 53443 1338
rect 53513 1292 53559 1338
rect 53629 1292 53675 1338
rect 53745 1292 53791 1338
rect 53861 1292 53907 1338
rect 53977 1292 54023 1338
rect 54093 1292 54139 1338
rect 54209 1292 54255 1338
rect 54325 1292 54371 1338
rect 54441 1292 54487 1338
rect 54557 1292 54603 1338
rect 54673 1292 54719 1338
rect 54789 1292 54835 1338
rect 54905 1292 54951 1338
rect 55021 1292 55067 1338
rect 55137 1292 55183 1338
rect 55253 1292 55299 1338
rect 55369 1292 55415 1338
rect 55485 1292 55531 1338
rect 55601 1292 55647 1338
rect 55717 1292 55763 1338
rect 55833 1292 55879 1338
rect 55949 1292 55995 1338
rect 56065 1292 56111 1338
rect 56181 1292 56227 1338
rect 56297 1292 56343 1338
rect 56413 1292 56459 1338
rect 56529 1292 56575 1338
rect 50845 1176 50891 1222
rect 50961 1176 51007 1222
rect 51077 1176 51123 1222
rect 51193 1176 51239 1222
rect 51309 1176 51355 1222
rect 51425 1176 51471 1222
rect 51541 1176 51587 1222
rect 51657 1176 51703 1222
rect 51773 1176 51819 1222
rect 51889 1176 51935 1222
rect 52005 1176 52051 1222
rect 52121 1176 52167 1222
rect 52237 1176 52283 1222
rect 52353 1176 52399 1222
rect 52469 1176 52515 1222
rect 52585 1176 52631 1222
rect 52701 1176 52747 1222
rect 52817 1176 52863 1222
rect 52933 1176 52979 1222
rect 53049 1176 53095 1222
rect 53165 1176 53211 1222
rect 53281 1176 53327 1222
rect 53397 1176 53443 1222
rect 53513 1176 53559 1222
rect 53629 1176 53675 1222
rect 53745 1176 53791 1222
rect 53861 1176 53907 1222
rect 53977 1176 54023 1222
rect 54093 1176 54139 1222
rect 54209 1176 54255 1222
rect 54325 1176 54371 1222
rect 54441 1176 54487 1222
rect 54557 1176 54603 1222
rect 54673 1176 54719 1222
rect 54789 1176 54835 1222
rect 54905 1176 54951 1222
rect 55021 1176 55067 1222
rect 55137 1176 55183 1222
rect 55253 1176 55299 1222
rect 55369 1176 55415 1222
rect 55485 1176 55531 1222
rect 55601 1176 55647 1222
rect 55717 1176 55763 1222
rect 55833 1176 55879 1222
rect 55949 1176 55995 1222
rect 56065 1176 56111 1222
rect 56181 1176 56227 1222
rect 56297 1176 56343 1222
rect 56413 1176 56459 1222
rect 56529 1176 56575 1222
rect 57380 1117 57626 45463
rect 85733 1117 86079 45563
rect 371 969 417 1015
rect 495 969 541 1015
rect 619 969 665 1015
rect 743 969 789 1015
rect 867 969 913 1015
rect 991 969 1037 1015
rect 1115 969 1161 1015
rect 1239 969 1285 1015
rect 1363 969 1409 1015
rect 1487 969 1533 1015
rect 1611 969 1657 1015
rect 1735 969 1781 1015
rect 1859 969 1905 1015
rect 1983 969 2029 1015
rect 2107 969 2153 1015
rect 2231 969 2277 1015
rect 2355 969 2401 1015
rect 2479 969 2525 1015
rect 2603 969 2649 1015
rect 2727 969 2773 1015
rect 2851 969 2897 1015
rect 2975 969 3021 1015
rect 3099 969 3145 1015
rect 3223 969 3269 1015
rect 3347 969 3393 1015
rect 3471 969 3517 1015
rect 3595 969 3641 1015
rect 3719 969 3765 1015
rect 3843 969 3889 1015
rect 3967 969 4013 1015
rect 4091 969 4137 1015
rect 4215 969 4261 1015
rect 4339 969 4385 1015
rect 4463 969 4509 1015
rect 4587 969 4633 1015
rect 4711 969 4757 1015
rect 4835 969 4881 1015
rect 4959 969 5005 1015
rect 5083 969 5129 1015
rect 5207 969 5253 1015
rect 5331 969 5377 1015
rect 5455 969 5501 1015
rect 5579 969 5625 1015
rect 5703 969 5749 1015
rect 5827 969 5873 1015
rect 5951 969 5997 1015
rect 6075 969 6121 1015
rect 6199 969 6245 1015
rect 6323 969 6369 1015
rect 6447 969 6493 1015
rect 6571 969 6617 1015
rect 6695 969 6741 1015
rect 6819 969 6865 1015
rect 6943 969 6989 1015
rect 7067 969 7113 1015
rect 7191 969 7237 1015
rect 7315 969 7361 1015
rect 7439 969 7485 1015
rect 7563 969 7609 1015
rect 7687 969 7733 1015
rect 7811 969 7857 1015
rect 7935 969 7981 1015
rect 8059 969 8105 1015
rect 8183 969 8229 1015
rect 8307 969 8353 1015
rect 8431 969 8477 1015
rect 8555 969 8601 1015
rect 8679 969 8725 1015
rect 8803 969 8849 1015
rect 8927 969 8973 1015
rect 9051 969 9097 1015
rect 9175 969 9221 1015
rect 9299 969 9345 1015
rect 9423 969 9469 1015
rect 9547 969 9593 1015
rect 9671 969 9717 1015
rect 9795 969 9841 1015
rect 9919 969 9965 1015
rect 10043 969 10089 1015
rect 10167 969 10213 1015
rect 10291 969 10337 1015
rect 10415 969 10461 1015
rect 10539 969 10585 1015
rect 10663 969 10709 1015
rect 10787 969 10833 1015
rect 10911 969 10957 1015
rect 11035 969 11081 1015
rect 11159 969 11205 1015
rect 11283 969 11329 1015
rect 11407 969 11453 1015
rect 11531 969 11577 1015
rect 11655 969 11701 1015
rect 11779 969 11825 1015
rect 11903 969 11949 1015
rect 12027 969 12073 1015
rect 12151 969 12197 1015
rect 12275 969 12321 1015
rect 12399 969 12445 1015
rect 12523 969 12569 1015
rect 12647 969 12693 1015
rect 12771 969 12817 1015
rect 12895 969 12941 1015
rect 13019 969 13065 1015
rect 13143 969 13189 1015
rect 13267 969 13313 1015
rect 13391 969 13437 1015
rect 13515 969 13561 1015
rect 13639 969 13685 1015
rect 13763 969 13809 1015
rect 13887 969 13933 1015
rect 14011 969 14057 1015
rect 14135 969 14181 1015
rect 14259 969 14305 1015
rect 14383 969 14429 1015
rect 14507 969 14553 1015
rect 14631 969 14677 1015
rect 14755 969 14801 1015
rect 14879 969 14925 1015
rect 15003 969 15049 1015
rect 15127 969 15173 1015
rect 15251 969 15297 1015
rect 15375 969 15421 1015
rect 15499 969 15545 1015
rect 15623 969 15669 1015
rect 15747 969 15793 1015
rect 15871 969 15917 1015
rect 15995 969 16041 1015
rect 16119 969 16165 1015
rect 16243 969 16289 1015
rect 16367 969 16413 1015
rect 16491 969 16537 1015
rect 16615 969 16661 1015
rect 16739 969 16785 1015
rect 16863 969 16909 1015
rect 16987 969 17033 1015
rect 17111 969 17157 1015
rect 17235 969 17281 1015
rect 17359 969 17405 1015
rect 17483 969 17529 1015
rect 17607 969 17653 1015
rect 17731 969 17777 1015
rect 17855 969 17901 1015
rect 17979 969 18025 1015
rect 18103 969 18149 1015
rect 18227 969 18273 1015
rect 18351 969 18397 1015
rect 18475 969 18521 1015
rect 18599 969 18645 1015
rect 18723 969 18769 1015
rect 18847 969 18893 1015
rect 18971 969 19017 1015
rect 19095 969 19141 1015
rect 19219 969 19265 1015
rect 19343 969 19389 1015
rect 19467 969 19513 1015
rect 19591 969 19637 1015
rect 19715 969 19761 1015
rect 19839 969 19885 1015
rect 19963 969 20009 1015
rect 20087 969 20133 1015
rect 20211 969 20257 1015
rect 20335 969 20381 1015
rect 20459 969 20505 1015
rect 20583 969 20629 1015
rect 20707 969 20753 1015
rect 20831 969 20877 1015
rect 20955 969 21001 1015
rect 21079 969 21125 1015
rect 21203 969 21249 1015
rect 21327 969 21373 1015
rect 21451 969 21497 1015
rect 21575 969 21621 1015
rect 21699 969 21745 1015
rect 21823 969 21869 1015
rect 21947 969 21993 1015
rect 22071 969 22117 1015
rect 22195 969 22241 1015
rect 22319 969 22365 1015
rect 22443 969 22489 1015
rect 22567 969 22613 1015
rect 22691 969 22737 1015
rect 22815 969 22861 1015
rect 22939 969 22985 1015
rect 23063 969 23109 1015
rect 23187 969 23233 1015
rect 23311 969 23357 1015
rect 23435 969 23481 1015
rect 23559 969 23605 1015
rect 23683 969 23729 1015
rect 23807 969 23853 1015
rect 23931 969 23977 1015
rect 24055 969 24101 1015
rect 24179 969 24225 1015
rect 24303 969 24349 1015
rect 24427 969 24473 1015
rect 24551 969 24597 1015
rect 24675 969 24721 1015
rect 24799 969 24845 1015
rect 24923 969 24969 1015
rect 25047 969 25093 1015
rect 25171 969 25217 1015
rect 25295 969 25341 1015
rect 25419 969 25465 1015
rect 25543 969 25589 1015
rect 25667 969 25713 1015
rect 25791 969 25837 1015
rect 25915 969 25961 1015
rect 26039 969 26085 1015
rect 26163 969 26209 1015
rect 26287 969 26333 1015
rect 26411 969 26457 1015
rect 26535 969 26581 1015
rect 26659 969 26705 1015
rect 26783 969 26829 1015
rect 26907 969 26953 1015
rect 27031 969 27077 1015
rect 27155 969 27201 1015
rect 27279 969 27325 1015
rect 27403 969 27449 1015
rect 27527 969 27573 1015
rect 27651 969 27697 1015
rect 27775 969 27821 1015
rect 27899 969 27945 1015
rect 28023 969 28069 1015
rect 28147 969 28193 1015
rect 28271 969 28317 1015
rect 28395 969 28441 1015
rect 28519 969 28565 1015
rect 28643 969 28689 1015
rect 28767 969 28813 1015
rect 28891 969 28937 1015
rect 29015 969 29061 1015
rect 29139 969 29185 1015
rect 29263 969 29309 1015
rect 29387 969 29433 1015
rect 29511 969 29557 1015
rect 29635 969 29681 1015
rect 29759 969 29805 1015
rect 29883 969 29929 1015
rect 30007 969 30053 1015
rect 30131 969 30177 1015
rect 30255 969 30301 1015
rect 30379 969 30425 1015
rect 30503 969 30549 1015
rect 30627 969 30673 1015
rect 30751 969 30797 1015
rect 30875 969 30921 1015
rect 30999 969 31045 1015
rect 31123 969 31169 1015
rect 31247 969 31293 1015
rect 31371 969 31417 1015
rect 31495 969 31541 1015
rect 31619 969 31665 1015
rect 31743 969 31789 1015
rect 31867 969 31913 1015
rect 31991 969 32037 1015
rect 32115 969 32161 1015
rect 32239 969 32285 1015
rect 32363 969 32409 1015
rect 32487 969 32533 1015
rect 32611 969 32657 1015
rect 32735 969 32781 1015
rect 32859 969 32905 1015
rect 32983 969 33029 1015
rect 33107 969 33153 1015
rect 33231 969 33277 1015
rect 33355 969 33401 1015
rect 33479 969 33525 1015
rect 33603 969 33649 1015
rect 33727 969 33773 1015
rect 33851 969 33897 1015
rect 33975 969 34021 1015
rect 34099 969 34145 1015
rect 34223 969 34269 1015
rect 34347 969 34393 1015
rect 34471 969 34517 1015
rect 34595 969 34641 1015
rect 34719 969 34765 1015
rect 34843 969 34889 1015
rect 34967 969 35013 1015
rect 35091 969 35137 1015
rect 35215 969 35261 1015
rect 35339 969 35385 1015
rect 35463 969 35509 1015
rect 35587 969 35633 1015
rect 35711 969 35757 1015
rect 35835 969 35881 1015
rect 35959 969 36005 1015
rect 36083 969 36129 1015
rect 36207 969 36253 1015
rect 36331 969 36377 1015
rect 36455 969 36501 1015
rect 36579 969 36625 1015
rect 36703 969 36749 1015
rect 36827 969 36873 1015
rect 36951 969 36997 1015
rect 37075 969 37121 1015
rect 37199 969 37245 1015
rect 37323 969 37369 1015
rect 37447 969 37493 1015
rect 37571 969 37617 1015
rect 37695 969 37741 1015
rect 37819 969 37865 1015
rect 37943 969 37989 1015
rect 38067 969 38113 1015
rect 38191 969 38237 1015
rect 38315 969 38361 1015
rect 38439 969 38485 1015
rect 38563 969 38609 1015
rect 38687 969 38733 1015
rect 38811 969 38857 1015
rect 38935 969 38981 1015
rect 39059 969 39105 1015
rect 39183 969 39229 1015
rect 39307 969 39353 1015
rect 39431 969 39477 1015
rect 39555 969 39601 1015
rect 39679 969 39725 1015
rect 39803 969 39849 1015
rect 39927 969 39973 1015
rect 40051 969 40097 1015
rect 40175 969 40221 1015
rect 40299 969 40345 1015
rect 40423 969 40469 1015
rect 40547 969 40593 1015
rect 40671 969 40717 1015
rect 40795 969 40841 1015
rect 40919 969 40965 1015
rect 41043 969 41089 1015
rect 41167 969 41213 1015
rect 41291 969 41337 1015
rect 41415 969 41461 1015
rect 41539 969 41585 1015
rect 41663 969 41709 1015
rect 41787 969 41833 1015
rect 41911 969 41957 1015
rect 42035 969 42081 1015
rect 42159 969 42205 1015
rect 42283 969 42329 1015
rect 42407 969 42453 1015
rect 42531 969 42577 1015
rect 42655 969 42701 1015
rect 42779 969 42825 1015
rect 42903 969 42949 1015
rect 43027 969 43073 1015
rect 43151 969 43197 1015
rect 43275 969 43321 1015
rect 43399 969 43445 1015
rect 43523 969 43569 1015
rect 43647 969 43693 1015
rect 43771 969 43817 1015
rect 43895 969 43941 1015
rect 44019 969 44065 1015
rect 44143 969 44189 1015
rect 44267 969 44313 1015
rect 44391 969 44437 1015
rect 44515 969 44561 1015
rect 44639 969 44685 1015
rect 44763 969 44809 1015
rect 44887 969 44933 1015
rect 45011 969 45057 1015
rect 45135 969 45181 1015
rect 45259 969 45305 1015
rect 45383 969 45429 1015
rect 45507 969 45553 1015
rect 45631 969 45677 1015
rect 45755 969 45801 1015
rect 45879 969 45925 1015
rect 46003 969 46049 1015
rect 46127 969 46173 1015
rect 46251 969 46297 1015
rect 46375 969 46421 1015
rect 46499 969 46545 1015
rect 46623 969 46669 1015
rect 46747 969 46793 1015
rect 46871 969 46917 1015
rect 46995 969 47041 1015
rect 47119 969 47165 1015
rect 47243 969 47289 1015
rect 47367 969 47413 1015
rect 47491 969 47537 1015
rect 47615 969 47661 1015
rect 47739 969 47785 1015
rect 47863 969 47909 1015
rect 47987 969 48033 1015
rect 48111 969 48157 1015
rect 48235 969 48281 1015
rect 48359 969 48405 1015
rect 48483 969 48529 1015
rect 48607 969 48653 1015
rect 48731 969 48777 1015
rect 48855 969 48901 1015
rect 48979 969 49025 1015
rect 49103 969 49149 1015
rect 49227 969 49273 1015
rect 49351 969 49397 1015
rect 49475 969 49521 1015
rect 49599 969 49645 1015
rect 49723 969 49769 1015
rect 49847 969 49893 1015
rect 49971 969 50017 1015
rect 50095 969 50141 1015
rect 50219 969 50265 1015
rect 50343 969 50389 1015
rect 50467 969 50513 1015
rect 50591 969 50637 1015
rect 50715 969 50761 1015
rect 50839 969 50885 1015
rect 50963 969 51009 1015
rect 51087 969 51133 1015
rect 51211 969 51257 1015
rect 51335 969 51381 1015
rect 51459 969 51505 1015
rect 51583 969 51629 1015
rect 51707 969 51753 1015
rect 51831 969 51877 1015
rect 51955 969 52001 1015
rect 52079 969 52125 1015
rect 52203 969 52249 1015
rect 52327 969 52373 1015
rect 52451 969 52497 1015
rect 52575 969 52621 1015
rect 52699 969 52745 1015
rect 52823 969 52869 1015
rect 52947 969 52993 1015
rect 53071 969 53117 1015
rect 53195 969 53241 1015
rect 53319 969 53365 1015
rect 53443 969 53489 1015
rect 53567 969 53613 1015
rect 53691 969 53737 1015
rect 53815 969 53861 1015
rect 53939 969 53985 1015
rect 54063 969 54109 1015
rect 54187 969 54233 1015
rect 54311 969 54357 1015
rect 54435 969 54481 1015
rect 54559 969 54605 1015
rect 54683 969 54729 1015
rect 54807 969 54853 1015
rect 54931 969 54977 1015
rect 55055 969 55101 1015
rect 55179 969 55225 1015
rect 55303 969 55349 1015
rect 55427 969 55473 1015
rect 55551 969 55597 1015
rect 55675 969 55721 1015
rect 55799 969 55845 1015
rect 55923 969 55969 1015
rect 56047 969 56093 1015
rect 56171 969 56217 1015
rect 56295 969 56341 1015
rect 56419 969 56465 1015
rect 56543 969 56589 1015
rect 56667 969 56713 1015
rect 56791 969 56837 1015
rect 56915 969 56961 1015
rect 57039 969 57085 1015
rect 57163 969 57209 1015
rect 57287 969 57333 1015
rect 57411 969 57457 1015
rect 57535 969 57581 1015
rect 57659 969 57705 1015
rect 57783 969 57829 1015
rect 57907 969 57953 1015
rect 58031 969 58077 1015
rect 58155 969 58201 1015
rect 58279 969 58325 1015
rect 58403 969 58449 1015
rect 58527 969 58573 1015
rect 58651 969 58697 1015
rect 58775 969 58821 1015
rect 58899 969 58945 1015
rect 59023 969 59069 1015
rect 59147 969 59193 1015
rect 59271 969 59317 1015
rect 59395 969 59441 1015
rect 59519 969 59565 1015
rect 59643 969 59689 1015
rect 59767 969 59813 1015
rect 59891 969 59937 1015
rect 60015 969 60061 1015
rect 60139 969 60185 1015
rect 60263 969 60309 1015
rect 60387 969 60433 1015
rect 60511 969 60557 1015
rect 60635 969 60681 1015
rect 60759 969 60805 1015
rect 60883 969 60929 1015
rect 61007 969 61053 1015
rect 61131 969 61177 1015
rect 61255 969 61301 1015
rect 61379 969 61425 1015
rect 61503 969 61549 1015
rect 61627 969 61673 1015
rect 61751 969 61797 1015
rect 61875 969 61921 1015
rect 61999 969 62045 1015
rect 62123 969 62169 1015
rect 62247 969 62293 1015
rect 62371 969 62417 1015
rect 62495 969 62541 1015
rect 62619 969 62665 1015
rect 62743 969 62789 1015
rect 62867 969 62913 1015
rect 62991 969 63037 1015
rect 63115 969 63161 1015
rect 63239 969 63285 1015
rect 63363 969 63409 1015
rect 63487 969 63533 1015
rect 63611 969 63657 1015
rect 63735 969 63781 1015
rect 63859 969 63905 1015
rect 63983 969 64029 1015
rect 64107 969 64153 1015
rect 64231 969 64277 1015
rect 64355 969 64401 1015
rect 64479 969 64525 1015
rect 64603 969 64649 1015
rect 64727 969 64773 1015
rect 64851 969 64897 1015
rect 64975 969 65021 1015
rect 65099 969 65145 1015
rect 65223 969 65269 1015
rect 65347 969 65393 1015
rect 65471 969 65517 1015
rect 65595 969 65641 1015
rect 65719 969 65765 1015
rect 65843 969 65889 1015
rect 65967 969 66013 1015
rect 66091 969 66137 1015
rect 66215 969 66261 1015
rect 66339 969 66385 1015
rect 66463 969 66509 1015
rect 66587 969 66633 1015
rect 66711 969 66757 1015
rect 66835 969 66881 1015
rect 66959 969 67005 1015
rect 67083 969 67129 1015
rect 67207 969 67253 1015
rect 67331 969 67377 1015
rect 67455 969 67501 1015
rect 67579 969 67625 1015
rect 67703 969 67749 1015
rect 67827 969 67873 1015
rect 67951 969 67997 1015
rect 68075 969 68121 1015
rect 68199 969 68245 1015
rect 68323 969 68369 1015
rect 68447 969 68493 1015
rect 68571 969 68617 1015
rect 68695 969 68741 1015
rect 68819 969 68865 1015
rect 68943 969 68989 1015
rect 69067 969 69113 1015
rect 69191 969 69237 1015
rect 69315 969 69361 1015
rect 69439 969 69485 1015
rect 69563 969 69609 1015
rect 69687 969 69733 1015
rect 69811 969 69857 1015
rect 69935 969 69981 1015
rect 70059 969 70105 1015
rect 70183 969 70229 1015
rect 70307 969 70353 1015
rect 70431 969 70477 1015
rect 70555 969 70601 1015
rect 70679 969 70725 1015
rect 70803 969 70849 1015
rect 70927 969 70973 1015
rect 71051 969 71097 1015
rect 71175 969 71221 1015
rect 71299 969 71345 1015
rect 71423 969 71469 1015
rect 71547 969 71593 1015
rect 71671 969 71717 1015
rect 71795 969 71841 1015
rect 71919 969 71965 1015
rect 72043 969 72089 1015
rect 72167 969 72213 1015
rect 72291 969 72337 1015
rect 72415 969 72461 1015
rect 72539 969 72585 1015
rect 72663 969 72709 1015
rect 72787 969 72833 1015
rect 72911 969 72957 1015
rect 73035 969 73081 1015
rect 73159 969 73205 1015
rect 73283 969 73329 1015
rect 73407 969 73453 1015
rect 73531 969 73577 1015
rect 73655 969 73701 1015
rect 73779 969 73825 1015
rect 73903 969 73949 1015
rect 74027 969 74073 1015
rect 74151 969 74197 1015
rect 74275 969 74321 1015
rect 74399 969 74445 1015
rect 74523 969 74569 1015
rect 74647 969 74693 1015
rect 74771 969 74817 1015
rect 74895 969 74941 1015
rect 75019 969 75065 1015
rect 75143 969 75189 1015
rect 75267 969 75313 1015
rect 75391 969 75437 1015
rect 75515 969 75561 1015
rect 75639 969 75685 1015
rect 75763 969 75809 1015
rect 75887 969 75933 1015
rect 76011 969 76057 1015
rect 76135 969 76181 1015
rect 76259 969 76305 1015
rect 76383 969 76429 1015
rect 76507 969 76553 1015
rect 76631 969 76677 1015
rect 76755 969 76801 1015
rect 76879 969 76925 1015
rect 77003 969 77049 1015
rect 77127 969 77173 1015
rect 77251 969 77297 1015
rect 77375 969 77421 1015
rect 77499 969 77545 1015
rect 77623 969 77669 1015
rect 77747 969 77793 1015
rect 77871 969 77917 1015
rect 77995 969 78041 1015
rect 78119 969 78165 1015
rect 78243 969 78289 1015
rect 78367 969 78413 1015
rect 78491 969 78537 1015
rect 78615 969 78661 1015
rect 78739 969 78785 1015
rect 78863 969 78909 1015
rect 78987 969 79033 1015
rect 79111 969 79157 1015
rect 79235 969 79281 1015
rect 79359 969 79405 1015
rect 79483 969 79529 1015
rect 79607 969 79653 1015
rect 79731 969 79777 1015
rect 79855 969 79901 1015
rect 79979 969 80025 1015
rect 80103 969 80149 1015
rect 80227 969 80273 1015
rect 80351 969 80397 1015
rect 80475 969 80521 1015
rect 80599 969 80645 1015
rect 80723 969 80769 1015
rect 80847 969 80893 1015
rect 80971 969 81017 1015
rect 81095 969 81141 1015
rect 81219 969 81265 1015
rect 81343 969 81389 1015
rect 81467 969 81513 1015
rect 81591 969 81637 1015
rect 81715 969 81761 1015
rect 81839 969 81885 1015
rect 81963 969 82009 1015
rect 82087 969 82133 1015
rect 82211 969 82257 1015
rect 82335 969 82381 1015
rect 82459 969 82505 1015
rect 82583 969 82629 1015
rect 82707 969 82753 1015
rect 82831 969 82877 1015
rect 82955 969 83001 1015
rect 83079 969 83125 1015
rect 83203 969 83249 1015
rect 83327 969 83373 1015
rect 83451 969 83497 1015
rect 83575 969 83621 1015
rect 83699 969 83745 1015
rect 83823 969 83869 1015
rect 83947 969 83993 1015
rect 84071 969 84117 1015
rect 84195 969 84241 1015
rect 84319 969 84365 1015
rect 84443 969 84489 1015
rect 84567 969 84613 1015
rect 84691 969 84737 1015
rect 84815 969 84861 1015
rect 84939 969 84985 1015
rect 85063 969 85109 1015
rect 85187 969 85233 1015
rect 85311 969 85357 1015
rect 85435 969 85481 1015
rect 85559 969 85605 1015
rect 85683 969 85729 1015
rect 85807 969 85853 1015
rect 85931 969 85977 1015
rect 371 845 417 891
rect 495 845 541 891
rect 619 845 665 891
rect 743 845 789 891
rect 867 845 913 891
rect 991 845 1037 891
rect 1115 845 1161 891
rect 1239 845 1285 891
rect 1363 845 1409 891
rect 1487 845 1533 891
rect 1611 845 1657 891
rect 1735 845 1781 891
rect 1859 845 1905 891
rect 1983 845 2029 891
rect 2107 845 2153 891
rect 2231 845 2277 891
rect 2355 845 2401 891
rect 2479 845 2525 891
rect 2603 845 2649 891
rect 2727 845 2773 891
rect 2851 845 2897 891
rect 2975 845 3021 891
rect 3099 845 3145 891
rect 3223 845 3269 891
rect 3347 845 3393 891
rect 3471 845 3517 891
rect 3595 845 3641 891
rect 3719 845 3765 891
rect 3843 845 3889 891
rect 3967 845 4013 891
rect 4091 845 4137 891
rect 4215 845 4261 891
rect 4339 845 4385 891
rect 4463 845 4509 891
rect 4587 845 4633 891
rect 4711 845 4757 891
rect 4835 845 4881 891
rect 4959 845 5005 891
rect 5083 845 5129 891
rect 5207 845 5253 891
rect 5331 845 5377 891
rect 5455 845 5501 891
rect 5579 845 5625 891
rect 5703 845 5749 891
rect 5827 845 5873 891
rect 5951 845 5997 891
rect 6075 845 6121 891
rect 6199 845 6245 891
rect 6323 845 6369 891
rect 6447 845 6493 891
rect 6571 845 6617 891
rect 6695 845 6741 891
rect 6819 845 6865 891
rect 6943 845 6989 891
rect 7067 845 7113 891
rect 7191 845 7237 891
rect 7315 845 7361 891
rect 7439 845 7485 891
rect 7563 845 7609 891
rect 7687 845 7733 891
rect 7811 845 7857 891
rect 7935 845 7981 891
rect 8059 845 8105 891
rect 8183 845 8229 891
rect 8307 845 8353 891
rect 8431 845 8477 891
rect 8555 845 8601 891
rect 8679 845 8725 891
rect 8803 845 8849 891
rect 8927 845 8973 891
rect 9051 845 9097 891
rect 9175 845 9221 891
rect 9299 845 9345 891
rect 9423 845 9469 891
rect 9547 845 9593 891
rect 9671 845 9717 891
rect 9795 845 9841 891
rect 9919 845 9965 891
rect 10043 845 10089 891
rect 10167 845 10213 891
rect 10291 845 10337 891
rect 10415 845 10461 891
rect 10539 845 10585 891
rect 10663 845 10709 891
rect 10787 845 10833 891
rect 10911 845 10957 891
rect 11035 845 11081 891
rect 11159 845 11205 891
rect 11283 845 11329 891
rect 11407 845 11453 891
rect 11531 845 11577 891
rect 11655 845 11701 891
rect 11779 845 11825 891
rect 11903 845 11949 891
rect 12027 845 12073 891
rect 12151 845 12197 891
rect 12275 845 12321 891
rect 12399 845 12445 891
rect 12523 845 12569 891
rect 12647 845 12693 891
rect 12771 845 12817 891
rect 12895 845 12941 891
rect 13019 845 13065 891
rect 13143 845 13189 891
rect 13267 845 13313 891
rect 13391 845 13437 891
rect 13515 845 13561 891
rect 13639 845 13685 891
rect 13763 845 13809 891
rect 13887 845 13933 891
rect 14011 845 14057 891
rect 14135 845 14181 891
rect 14259 845 14305 891
rect 14383 845 14429 891
rect 14507 845 14553 891
rect 14631 845 14677 891
rect 14755 845 14801 891
rect 14879 845 14925 891
rect 15003 845 15049 891
rect 15127 845 15173 891
rect 15251 845 15297 891
rect 15375 845 15421 891
rect 15499 845 15545 891
rect 15623 845 15669 891
rect 15747 845 15793 891
rect 15871 845 15917 891
rect 15995 845 16041 891
rect 16119 845 16165 891
rect 16243 845 16289 891
rect 16367 845 16413 891
rect 16491 845 16537 891
rect 16615 845 16661 891
rect 16739 845 16785 891
rect 16863 845 16909 891
rect 16987 845 17033 891
rect 17111 845 17157 891
rect 17235 845 17281 891
rect 17359 845 17405 891
rect 17483 845 17529 891
rect 17607 845 17653 891
rect 17731 845 17777 891
rect 17855 845 17901 891
rect 17979 845 18025 891
rect 18103 845 18149 891
rect 18227 845 18273 891
rect 18351 845 18397 891
rect 18475 845 18521 891
rect 18599 845 18645 891
rect 18723 845 18769 891
rect 18847 845 18893 891
rect 18971 845 19017 891
rect 19095 845 19141 891
rect 19219 845 19265 891
rect 19343 845 19389 891
rect 19467 845 19513 891
rect 19591 845 19637 891
rect 19715 845 19761 891
rect 19839 845 19885 891
rect 19963 845 20009 891
rect 20087 845 20133 891
rect 20211 845 20257 891
rect 20335 845 20381 891
rect 20459 845 20505 891
rect 20583 845 20629 891
rect 20707 845 20753 891
rect 20831 845 20877 891
rect 20955 845 21001 891
rect 21079 845 21125 891
rect 21203 845 21249 891
rect 21327 845 21373 891
rect 21451 845 21497 891
rect 21575 845 21621 891
rect 21699 845 21745 891
rect 21823 845 21869 891
rect 21947 845 21993 891
rect 22071 845 22117 891
rect 22195 845 22241 891
rect 22319 845 22365 891
rect 22443 845 22489 891
rect 22567 845 22613 891
rect 22691 845 22737 891
rect 22815 845 22861 891
rect 22939 845 22985 891
rect 23063 845 23109 891
rect 23187 845 23233 891
rect 23311 845 23357 891
rect 23435 845 23481 891
rect 23559 845 23605 891
rect 23683 845 23729 891
rect 23807 845 23853 891
rect 23931 845 23977 891
rect 24055 845 24101 891
rect 24179 845 24225 891
rect 24303 845 24349 891
rect 24427 845 24473 891
rect 24551 845 24597 891
rect 24675 845 24721 891
rect 24799 845 24845 891
rect 24923 845 24969 891
rect 25047 845 25093 891
rect 25171 845 25217 891
rect 25295 845 25341 891
rect 25419 845 25465 891
rect 25543 845 25589 891
rect 25667 845 25713 891
rect 25791 845 25837 891
rect 25915 845 25961 891
rect 26039 845 26085 891
rect 26163 845 26209 891
rect 26287 845 26333 891
rect 26411 845 26457 891
rect 26535 845 26581 891
rect 26659 845 26705 891
rect 26783 845 26829 891
rect 26907 845 26953 891
rect 27031 845 27077 891
rect 27155 845 27201 891
rect 27279 845 27325 891
rect 27403 845 27449 891
rect 27527 845 27573 891
rect 27651 845 27697 891
rect 27775 845 27821 891
rect 27899 845 27945 891
rect 28023 845 28069 891
rect 28147 845 28193 891
rect 28271 845 28317 891
rect 28395 845 28441 891
rect 28519 845 28565 891
rect 28643 845 28689 891
rect 28767 845 28813 891
rect 28891 845 28937 891
rect 29015 845 29061 891
rect 29139 845 29185 891
rect 29263 845 29309 891
rect 29387 845 29433 891
rect 29511 845 29557 891
rect 29635 845 29681 891
rect 29759 845 29805 891
rect 29883 845 29929 891
rect 30007 845 30053 891
rect 30131 845 30177 891
rect 30255 845 30301 891
rect 30379 845 30425 891
rect 30503 845 30549 891
rect 30627 845 30673 891
rect 30751 845 30797 891
rect 30875 845 30921 891
rect 30999 845 31045 891
rect 31123 845 31169 891
rect 31247 845 31293 891
rect 31371 845 31417 891
rect 31495 845 31541 891
rect 31619 845 31665 891
rect 31743 845 31789 891
rect 31867 845 31913 891
rect 31991 845 32037 891
rect 32115 845 32161 891
rect 32239 845 32285 891
rect 32363 845 32409 891
rect 32487 845 32533 891
rect 32611 845 32657 891
rect 32735 845 32781 891
rect 32859 845 32905 891
rect 32983 845 33029 891
rect 33107 845 33153 891
rect 33231 845 33277 891
rect 33355 845 33401 891
rect 33479 845 33525 891
rect 33603 845 33649 891
rect 33727 845 33773 891
rect 33851 845 33897 891
rect 33975 845 34021 891
rect 34099 845 34145 891
rect 34223 845 34269 891
rect 34347 845 34393 891
rect 34471 845 34517 891
rect 34595 845 34641 891
rect 34719 845 34765 891
rect 34843 845 34889 891
rect 34967 845 35013 891
rect 35091 845 35137 891
rect 35215 845 35261 891
rect 35339 845 35385 891
rect 35463 845 35509 891
rect 35587 845 35633 891
rect 35711 845 35757 891
rect 35835 845 35881 891
rect 35959 845 36005 891
rect 36083 845 36129 891
rect 36207 845 36253 891
rect 36331 845 36377 891
rect 36455 845 36501 891
rect 36579 845 36625 891
rect 36703 845 36749 891
rect 36827 845 36873 891
rect 36951 845 36997 891
rect 37075 845 37121 891
rect 37199 845 37245 891
rect 37323 845 37369 891
rect 37447 845 37493 891
rect 37571 845 37617 891
rect 37695 845 37741 891
rect 37819 845 37865 891
rect 37943 845 37989 891
rect 38067 845 38113 891
rect 38191 845 38237 891
rect 38315 845 38361 891
rect 38439 845 38485 891
rect 38563 845 38609 891
rect 38687 845 38733 891
rect 38811 845 38857 891
rect 38935 845 38981 891
rect 39059 845 39105 891
rect 39183 845 39229 891
rect 39307 845 39353 891
rect 39431 845 39477 891
rect 39555 845 39601 891
rect 39679 845 39725 891
rect 39803 845 39849 891
rect 39927 845 39973 891
rect 40051 845 40097 891
rect 40175 845 40221 891
rect 40299 845 40345 891
rect 40423 845 40469 891
rect 40547 845 40593 891
rect 40671 845 40717 891
rect 40795 845 40841 891
rect 40919 845 40965 891
rect 41043 845 41089 891
rect 41167 845 41213 891
rect 41291 845 41337 891
rect 41415 845 41461 891
rect 41539 845 41585 891
rect 41663 845 41709 891
rect 41787 845 41833 891
rect 41911 845 41957 891
rect 42035 845 42081 891
rect 42159 845 42205 891
rect 42283 845 42329 891
rect 42407 845 42453 891
rect 42531 845 42577 891
rect 42655 845 42701 891
rect 42779 845 42825 891
rect 42903 845 42949 891
rect 43027 845 43073 891
rect 43151 845 43197 891
rect 43275 845 43321 891
rect 43399 845 43445 891
rect 43523 845 43569 891
rect 43647 845 43693 891
rect 43771 845 43817 891
rect 43895 845 43941 891
rect 44019 845 44065 891
rect 44143 845 44189 891
rect 44267 845 44313 891
rect 44391 845 44437 891
rect 44515 845 44561 891
rect 44639 845 44685 891
rect 44763 845 44809 891
rect 44887 845 44933 891
rect 45011 845 45057 891
rect 45135 845 45181 891
rect 45259 845 45305 891
rect 45383 845 45429 891
rect 45507 845 45553 891
rect 45631 845 45677 891
rect 45755 845 45801 891
rect 45879 845 45925 891
rect 46003 845 46049 891
rect 46127 845 46173 891
rect 46251 845 46297 891
rect 46375 845 46421 891
rect 46499 845 46545 891
rect 46623 845 46669 891
rect 46747 845 46793 891
rect 46871 845 46917 891
rect 46995 845 47041 891
rect 47119 845 47165 891
rect 47243 845 47289 891
rect 47367 845 47413 891
rect 47491 845 47537 891
rect 47615 845 47661 891
rect 47739 845 47785 891
rect 47863 845 47909 891
rect 47987 845 48033 891
rect 48111 845 48157 891
rect 48235 845 48281 891
rect 48359 845 48405 891
rect 48483 845 48529 891
rect 48607 845 48653 891
rect 48731 845 48777 891
rect 48855 845 48901 891
rect 48979 845 49025 891
rect 49103 845 49149 891
rect 49227 845 49273 891
rect 49351 845 49397 891
rect 49475 845 49521 891
rect 49599 845 49645 891
rect 49723 845 49769 891
rect 49847 845 49893 891
rect 49971 845 50017 891
rect 50095 845 50141 891
rect 50219 845 50265 891
rect 50343 845 50389 891
rect 50467 845 50513 891
rect 50591 845 50637 891
rect 50715 845 50761 891
rect 50839 845 50885 891
rect 50963 845 51009 891
rect 51087 845 51133 891
rect 51211 845 51257 891
rect 51335 845 51381 891
rect 51459 845 51505 891
rect 51583 845 51629 891
rect 51707 845 51753 891
rect 51831 845 51877 891
rect 51955 845 52001 891
rect 52079 845 52125 891
rect 52203 845 52249 891
rect 52327 845 52373 891
rect 52451 845 52497 891
rect 52575 845 52621 891
rect 52699 845 52745 891
rect 52823 845 52869 891
rect 52947 845 52993 891
rect 53071 845 53117 891
rect 53195 845 53241 891
rect 53319 845 53365 891
rect 53443 845 53489 891
rect 53567 845 53613 891
rect 53691 845 53737 891
rect 53815 845 53861 891
rect 53939 845 53985 891
rect 54063 845 54109 891
rect 54187 845 54233 891
rect 54311 845 54357 891
rect 54435 845 54481 891
rect 54559 845 54605 891
rect 54683 845 54729 891
rect 54807 845 54853 891
rect 54931 845 54977 891
rect 55055 845 55101 891
rect 55179 845 55225 891
rect 55303 845 55349 891
rect 55427 845 55473 891
rect 55551 845 55597 891
rect 55675 845 55721 891
rect 55799 845 55845 891
rect 55923 845 55969 891
rect 56047 845 56093 891
rect 56171 845 56217 891
rect 56295 845 56341 891
rect 56419 845 56465 891
rect 56543 845 56589 891
rect 56667 845 56713 891
rect 56791 845 56837 891
rect 56915 845 56961 891
rect 57039 845 57085 891
rect 57163 845 57209 891
rect 57287 845 57333 891
rect 57411 845 57457 891
rect 57535 845 57581 891
rect 57659 845 57705 891
rect 57783 845 57829 891
rect 57907 845 57953 891
rect 58031 845 58077 891
rect 58155 845 58201 891
rect 58279 845 58325 891
rect 58403 845 58449 891
rect 58527 845 58573 891
rect 58651 845 58697 891
rect 58775 845 58821 891
rect 58899 845 58945 891
rect 59023 845 59069 891
rect 59147 845 59193 891
rect 59271 845 59317 891
rect 59395 845 59441 891
rect 59519 845 59565 891
rect 59643 845 59689 891
rect 59767 845 59813 891
rect 59891 845 59937 891
rect 60015 845 60061 891
rect 60139 845 60185 891
rect 60263 845 60309 891
rect 60387 845 60433 891
rect 60511 845 60557 891
rect 60635 845 60681 891
rect 60759 845 60805 891
rect 60883 845 60929 891
rect 61007 845 61053 891
rect 61131 845 61177 891
rect 61255 845 61301 891
rect 61379 845 61425 891
rect 61503 845 61549 891
rect 61627 845 61673 891
rect 61751 845 61797 891
rect 61875 845 61921 891
rect 61999 845 62045 891
rect 62123 845 62169 891
rect 62247 845 62293 891
rect 62371 845 62417 891
rect 62495 845 62541 891
rect 62619 845 62665 891
rect 62743 845 62789 891
rect 62867 845 62913 891
rect 62991 845 63037 891
rect 63115 845 63161 891
rect 63239 845 63285 891
rect 63363 845 63409 891
rect 63487 845 63533 891
rect 63611 845 63657 891
rect 63735 845 63781 891
rect 63859 845 63905 891
rect 63983 845 64029 891
rect 64107 845 64153 891
rect 64231 845 64277 891
rect 64355 845 64401 891
rect 64479 845 64525 891
rect 64603 845 64649 891
rect 64727 845 64773 891
rect 64851 845 64897 891
rect 64975 845 65021 891
rect 65099 845 65145 891
rect 65223 845 65269 891
rect 65347 845 65393 891
rect 65471 845 65517 891
rect 65595 845 65641 891
rect 65719 845 65765 891
rect 65843 845 65889 891
rect 65967 845 66013 891
rect 66091 845 66137 891
rect 66215 845 66261 891
rect 66339 845 66385 891
rect 66463 845 66509 891
rect 66587 845 66633 891
rect 66711 845 66757 891
rect 66835 845 66881 891
rect 66959 845 67005 891
rect 67083 845 67129 891
rect 67207 845 67253 891
rect 67331 845 67377 891
rect 67455 845 67501 891
rect 67579 845 67625 891
rect 67703 845 67749 891
rect 67827 845 67873 891
rect 67951 845 67997 891
rect 68075 845 68121 891
rect 68199 845 68245 891
rect 68323 845 68369 891
rect 68447 845 68493 891
rect 68571 845 68617 891
rect 68695 845 68741 891
rect 68819 845 68865 891
rect 68943 845 68989 891
rect 69067 845 69113 891
rect 69191 845 69237 891
rect 69315 845 69361 891
rect 69439 845 69485 891
rect 69563 845 69609 891
rect 69687 845 69733 891
rect 69811 845 69857 891
rect 69935 845 69981 891
rect 70059 845 70105 891
rect 70183 845 70229 891
rect 70307 845 70353 891
rect 70431 845 70477 891
rect 70555 845 70601 891
rect 70679 845 70725 891
rect 70803 845 70849 891
rect 70927 845 70973 891
rect 71051 845 71097 891
rect 71175 845 71221 891
rect 71299 845 71345 891
rect 71423 845 71469 891
rect 71547 845 71593 891
rect 71671 845 71717 891
rect 71795 845 71841 891
rect 71919 845 71965 891
rect 72043 845 72089 891
rect 72167 845 72213 891
rect 72291 845 72337 891
rect 72415 845 72461 891
rect 72539 845 72585 891
rect 72663 845 72709 891
rect 72787 845 72833 891
rect 72911 845 72957 891
rect 73035 845 73081 891
rect 73159 845 73205 891
rect 73283 845 73329 891
rect 73407 845 73453 891
rect 73531 845 73577 891
rect 73655 845 73701 891
rect 73779 845 73825 891
rect 73903 845 73949 891
rect 74027 845 74073 891
rect 74151 845 74197 891
rect 74275 845 74321 891
rect 74399 845 74445 891
rect 74523 845 74569 891
rect 74647 845 74693 891
rect 74771 845 74817 891
rect 74895 845 74941 891
rect 75019 845 75065 891
rect 75143 845 75189 891
rect 75267 845 75313 891
rect 75391 845 75437 891
rect 75515 845 75561 891
rect 75639 845 75685 891
rect 75763 845 75809 891
rect 75887 845 75933 891
rect 76011 845 76057 891
rect 76135 845 76181 891
rect 76259 845 76305 891
rect 76383 845 76429 891
rect 76507 845 76553 891
rect 76631 845 76677 891
rect 76755 845 76801 891
rect 76879 845 76925 891
rect 77003 845 77049 891
rect 77127 845 77173 891
rect 77251 845 77297 891
rect 77375 845 77421 891
rect 77499 845 77545 891
rect 77623 845 77669 891
rect 77747 845 77793 891
rect 77871 845 77917 891
rect 77995 845 78041 891
rect 78119 845 78165 891
rect 78243 845 78289 891
rect 78367 845 78413 891
rect 78491 845 78537 891
rect 78615 845 78661 891
rect 78739 845 78785 891
rect 78863 845 78909 891
rect 78987 845 79033 891
rect 79111 845 79157 891
rect 79235 845 79281 891
rect 79359 845 79405 891
rect 79483 845 79529 891
rect 79607 845 79653 891
rect 79731 845 79777 891
rect 79855 845 79901 891
rect 79979 845 80025 891
rect 80103 845 80149 891
rect 80227 845 80273 891
rect 80351 845 80397 891
rect 80475 845 80521 891
rect 80599 845 80645 891
rect 80723 845 80769 891
rect 80847 845 80893 891
rect 80971 845 81017 891
rect 81095 845 81141 891
rect 81219 845 81265 891
rect 81343 845 81389 891
rect 81467 845 81513 891
rect 81591 845 81637 891
rect 81715 845 81761 891
rect 81839 845 81885 891
rect 81963 845 82009 891
rect 82087 845 82133 891
rect 82211 845 82257 891
rect 82335 845 82381 891
rect 82459 845 82505 891
rect 82583 845 82629 891
rect 82707 845 82753 891
rect 82831 845 82877 891
rect 82955 845 83001 891
rect 83079 845 83125 891
rect 83203 845 83249 891
rect 83327 845 83373 891
rect 83451 845 83497 891
rect 83575 845 83621 891
rect 83699 845 83745 891
rect 83823 845 83869 891
rect 83947 845 83993 891
rect 84071 845 84117 891
rect 84195 845 84241 891
rect 84319 845 84365 891
rect 84443 845 84489 891
rect 84567 845 84613 891
rect 84691 845 84737 891
rect 84815 845 84861 891
rect 84939 845 84985 891
rect 85063 845 85109 891
rect 85187 845 85233 891
rect 85311 845 85357 891
rect 85435 845 85481 891
rect 85559 845 85605 891
rect 85683 845 85729 891
rect 85807 845 85853 891
rect 85931 845 85977 891
rect 371 721 417 767
rect 495 721 541 767
rect 619 721 665 767
rect 743 721 789 767
rect 867 721 913 767
rect 991 721 1037 767
rect 1115 721 1161 767
rect 1239 721 1285 767
rect 1363 721 1409 767
rect 1487 721 1533 767
rect 1611 721 1657 767
rect 1735 721 1781 767
rect 1859 721 1905 767
rect 1983 721 2029 767
rect 2107 721 2153 767
rect 2231 721 2277 767
rect 2355 721 2401 767
rect 2479 721 2525 767
rect 2603 721 2649 767
rect 2727 721 2773 767
rect 2851 721 2897 767
rect 2975 721 3021 767
rect 3099 721 3145 767
rect 3223 721 3269 767
rect 3347 721 3393 767
rect 3471 721 3517 767
rect 3595 721 3641 767
rect 3719 721 3765 767
rect 3843 721 3889 767
rect 3967 721 4013 767
rect 4091 721 4137 767
rect 4215 721 4261 767
rect 4339 721 4385 767
rect 4463 721 4509 767
rect 4587 721 4633 767
rect 4711 721 4757 767
rect 4835 721 4881 767
rect 4959 721 5005 767
rect 5083 721 5129 767
rect 5207 721 5253 767
rect 5331 721 5377 767
rect 5455 721 5501 767
rect 5579 721 5625 767
rect 5703 721 5749 767
rect 5827 721 5873 767
rect 5951 721 5997 767
rect 6075 721 6121 767
rect 6199 721 6245 767
rect 6323 721 6369 767
rect 6447 721 6493 767
rect 6571 721 6617 767
rect 6695 721 6741 767
rect 6819 721 6865 767
rect 6943 721 6989 767
rect 7067 721 7113 767
rect 7191 721 7237 767
rect 7315 721 7361 767
rect 7439 721 7485 767
rect 7563 721 7609 767
rect 7687 721 7733 767
rect 7811 721 7857 767
rect 7935 721 7981 767
rect 8059 721 8105 767
rect 8183 721 8229 767
rect 8307 721 8353 767
rect 8431 721 8477 767
rect 8555 721 8601 767
rect 8679 721 8725 767
rect 8803 721 8849 767
rect 8927 721 8973 767
rect 9051 721 9097 767
rect 9175 721 9221 767
rect 9299 721 9345 767
rect 9423 721 9469 767
rect 9547 721 9593 767
rect 9671 721 9717 767
rect 9795 721 9841 767
rect 9919 721 9965 767
rect 10043 721 10089 767
rect 10167 721 10213 767
rect 10291 721 10337 767
rect 10415 721 10461 767
rect 10539 721 10585 767
rect 10663 721 10709 767
rect 10787 721 10833 767
rect 10911 721 10957 767
rect 11035 721 11081 767
rect 11159 721 11205 767
rect 11283 721 11329 767
rect 11407 721 11453 767
rect 11531 721 11577 767
rect 11655 721 11701 767
rect 11779 721 11825 767
rect 11903 721 11949 767
rect 12027 721 12073 767
rect 12151 721 12197 767
rect 12275 721 12321 767
rect 12399 721 12445 767
rect 12523 721 12569 767
rect 12647 721 12693 767
rect 12771 721 12817 767
rect 12895 721 12941 767
rect 13019 721 13065 767
rect 13143 721 13189 767
rect 13267 721 13313 767
rect 13391 721 13437 767
rect 13515 721 13561 767
rect 13639 721 13685 767
rect 13763 721 13809 767
rect 13887 721 13933 767
rect 14011 721 14057 767
rect 14135 721 14181 767
rect 14259 721 14305 767
rect 14383 721 14429 767
rect 14507 721 14553 767
rect 14631 721 14677 767
rect 14755 721 14801 767
rect 14879 721 14925 767
rect 15003 721 15049 767
rect 15127 721 15173 767
rect 15251 721 15297 767
rect 15375 721 15421 767
rect 15499 721 15545 767
rect 15623 721 15669 767
rect 15747 721 15793 767
rect 15871 721 15917 767
rect 15995 721 16041 767
rect 16119 721 16165 767
rect 16243 721 16289 767
rect 16367 721 16413 767
rect 16491 721 16537 767
rect 16615 721 16661 767
rect 16739 721 16785 767
rect 16863 721 16909 767
rect 16987 721 17033 767
rect 17111 721 17157 767
rect 17235 721 17281 767
rect 17359 721 17405 767
rect 17483 721 17529 767
rect 17607 721 17653 767
rect 17731 721 17777 767
rect 17855 721 17901 767
rect 17979 721 18025 767
rect 18103 721 18149 767
rect 18227 721 18273 767
rect 18351 721 18397 767
rect 18475 721 18521 767
rect 18599 721 18645 767
rect 18723 721 18769 767
rect 18847 721 18893 767
rect 18971 721 19017 767
rect 19095 721 19141 767
rect 19219 721 19265 767
rect 19343 721 19389 767
rect 19467 721 19513 767
rect 19591 721 19637 767
rect 19715 721 19761 767
rect 19839 721 19885 767
rect 19963 721 20009 767
rect 20087 721 20133 767
rect 20211 721 20257 767
rect 20335 721 20381 767
rect 20459 721 20505 767
rect 20583 721 20629 767
rect 20707 721 20753 767
rect 20831 721 20877 767
rect 20955 721 21001 767
rect 21079 721 21125 767
rect 21203 721 21249 767
rect 21327 721 21373 767
rect 21451 721 21497 767
rect 21575 721 21621 767
rect 21699 721 21745 767
rect 21823 721 21869 767
rect 21947 721 21993 767
rect 22071 721 22117 767
rect 22195 721 22241 767
rect 22319 721 22365 767
rect 22443 721 22489 767
rect 22567 721 22613 767
rect 22691 721 22737 767
rect 22815 721 22861 767
rect 22939 721 22985 767
rect 23063 721 23109 767
rect 23187 721 23233 767
rect 23311 721 23357 767
rect 23435 721 23481 767
rect 23559 721 23605 767
rect 23683 721 23729 767
rect 23807 721 23853 767
rect 23931 721 23977 767
rect 24055 721 24101 767
rect 24179 721 24225 767
rect 24303 721 24349 767
rect 24427 721 24473 767
rect 24551 721 24597 767
rect 24675 721 24721 767
rect 24799 721 24845 767
rect 24923 721 24969 767
rect 25047 721 25093 767
rect 25171 721 25217 767
rect 25295 721 25341 767
rect 25419 721 25465 767
rect 25543 721 25589 767
rect 25667 721 25713 767
rect 25791 721 25837 767
rect 25915 721 25961 767
rect 26039 721 26085 767
rect 26163 721 26209 767
rect 26287 721 26333 767
rect 26411 721 26457 767
rect 26535 721 26581 767
rect 26659 721 26705 767
rect 26783 721 26829 767
rect 26907 721 26953 767
rect 27031 721 27077 767
rect 27155 721 27201 767
rect 27279 721 27325 767
rect 27403 721 27449 767
rect 27527 721 27573 767
rect 27651 721 27697 767
rect 27775 721 27821 767
rect 27899 721 27945 767
rect 28023 721 28069 767
rect 28147 721 28193 767
rect 28271 721 28317 767
rect 28395 721 28441 767
rect 28519 721 28565 767
rect 28643 721 28689 767
rect 28767 721 28813 767
rect 28891 721 28937 767
rect 29015 721 29061 767
rect 29139 721 29185 767
rect 29263 721 29309 767
rect 29387 721 29433 767
rect 29511 721 29557 767
rect 29635 721 29681 767
rect 29759 721 29805 767
rect 29883 721 29929 767
rect 30007 721 30053 767
rect 30131 721 30177 767
rect 30255 721 30301 767
rect 30379 721 30425 767
rect 30503 721 30549 767
rect 30627 721 30673 767
rect 30751 721 30797 767
rect 30875 721 30921 767
rect 30999 721 31045 767
rect 31123 721 31169 767
rect 31247 721 31293 767
rect 31371 721 31417 767
rect 31495 721 31541 767
rect 31619 721 31665 767
rect 31743 721 31789 767
rect 31867 721 31913 767
rect 31991 721 32037 767
rect 32115 721 32161 767
rect 32239 721 32285 767
rect 32363 721 32409 767
rect 32487 721 32533 767
rect 32611 721 32657 767
rect 32735 721 32781 767
rect 32859 721 32905 767
rect 32983 721 33029 767
rect 33107 721 33153 767
rect 33231 721 33277 767
rect 33355 721 33401 767
rect 33479 721 33525 767
rect 33603 721 33649 767
rect 33727 721 33773 767
rect 33851 721 33897 767
rect 33975 721 34021 767
rect 34099 721 34145 767
rect 34223 721 34269 767
rect 34347 721 34393 767
rect 34471 721 34517 767
rect 34595 721 34641 767
rect 34719 721 34765 767
rect 34843 721 34889 767
rect 34967 721 35013 767
rect 35091 721 35137 767
rect 35215 721 35261 767
rect 35339 721 35385 767
rect 35463 721 35509 767
rect 35587 721 35633 767
rect 35711 721 35757 767
rect 35835 721 35881 767
rect 35959 721 36005 767
rect 36083 721 36129 767
rect 36207 721 36253 767
rect 36331 721 36377 767
rect 36455 721 36501 767
rect 36579 721 36625 767
rect 36703 721 36749 767
rect 36827 721 36873 767
rect 36951 721 36997 767
rect 37075 721 37121 767
rect 37199 721 37245 767
rect 37323 721 37369 767
rect 37447 721 37493 767
rect 37571 721 37617 767
rect 37695 721 37741 767
rect 37819 721 37865 767
rect 37943 721 37989 767
rect 38067 721 38113 767
rect 38191 721 38237 767
rect 38315 721 38361 767
rect 38439 721 38485 767
rect 38563 721 38609 767
rect 38687 721 38733 767
rect 38811 721 38857 767
rect 38935 721 38981 767
rect 39059 721 39105 767
rect 39183 721 39229 767
rect 39307 721 39353 767
rect 39431 721 39477 767
rect 39555 721 39601 767
rect 39679 721 39725 767
rect 39803 721 39849 767
rect 39927 721 39973 767
rect 40051 721 40097 767
rect 40175 721 40221 767
rect 40299 721 40345 767
rect 40423 721 40469 767
rect 40547 721 40593 767
rect 40671 721 40717 767
rect 40795 721 40841 767
rect 40919 721 40965 767
rect 41043 721 41089 767
rect 41167 721 41213 767
rect 41291 721 41337 767
rect 41415 721 41461 767
rect 41539 721 41585 767
rect 41663 721 41709 767
rect 41787 721 41833 767
rect 41911 721 41957 767
rect 42035 721 42081 767
rect 42159 721 42205 767
rect 42283 721 42329 767
rect 42407 721 42453 767
rect 42531 721 42577 767
rect 42655 721 42701 767
rect 42779 721 42825 767
rect 42903 721 42949 767
rect 43027 721 43073 767
rect 43151 721 43197 767
rect 43275 721 43321 767
rect 43399 721 43445 767
rect 43523 721 43569 767
rect 43647 721 43693 767
rect 43771 721 43817 767
rect 43895 721 43941 767
rect 44019 721 44065 767
rect 44143 721 44189 767
rect 44267 721 44313 767
rect 44391 721 44437 767
rect 44515 721 44561 767
rect 44639 721 44685 767
rect 44763 721 44809 767
rect 44887 721 44933 767
rect 45011 721 45057 767
rect 45135 721 45181 767
rect 45259 721 45305 767
rect 45383 721 45429 767
rect 45507 721 45553 767
rect 45631 721 45677 767
rect 45755 721 45801 767
rect 45879 721 45925 767
rect 46003 721 46049 767
rect 46127 721 46173 767
rect 46251 721 46297 767
rect 46375 721 46421 767
rect 46499 721 46545 767
rect 46623 721 46669 767
rect 46747 721 46793 767
rect 46871 721 46917 767
rect 46995 721 47041 767
rect 47119 721 47165 767
rect 47243 721 47289 767
rect 47367 721 47413 767
rect 47491 721 47537 767
rect 47615 721 47661 767
rect 47739 721 47785 767
rect 47863 721 47909 767
rect 47987 721 48033 767
rect 48111 721 48157 767
rect 48235 721 48281 767
rect 48359 721 48405 767
rect 48483 721 48529 767
rect 48607 721 48653 767
rect 48731 721 48777 767
rect 48855 721 48901 767
rect 48979 721 49025 767
rect 49103 721 49149 767
rect 49227 721 49273 767
rect 49351 721 49397 767
rect 49475 721 49521 767
rect 49599 721 49645 767
rect 49723 721 49769 767
rect 49847 721 49893 767
rect 49971 721 50017 767
rect 50095 721 50141 767
rect 50219 721 50265 767
rect 50343 721 50389 767
rect 50467 721 50513 767
rect 50591 721 50637 767
rect 50715 721 50761 767
rect 50839 721 50885 767
rect 50963 721 51009 767
rect 51087 721 51133 767
rect 51211 721 51257 767
rect 51335 721 51381 767
rect 51459 721 51505 767
rect 51583 721 51629 767
rect 51707 721 51753 767
rect 51831 721 51877 767
rect 51955 721 52001 767
rect 52079 721 52125 767
rect 52203 721 52249 767
rect 52327 721 52373 767
rect 52451 721 52497 767
rect 52575 721 52621 767
rect 52699 721 52745 767
rect 52823 721 52869 767
rect 52947 721 52993 767
rect 53071 721 53117 767
rect 53195 721 53241 767
rect 53319 721 53365 767
rect 53443 721 53489 767
rect 53567 721 53613 767
rect 53691 721 53737 767
rect 53815 721 53861 767
rect 53939 721 53985 767
rect 54063 721 54109 767
rect 54187 721 54233 767
rect 54311 721 54357 767
rect 54435 721 54481 767
rect 54559 721 54605 767
rect 54683 721 54729 767
rect 54807 721 54853 767
rect 54931 721 54977 767
rect 55055 721 55101 767
rect 55179 721 55225 767
rect 55303 721 55349 767
rect 55427 721 55473 767
rect 55551 721 55597 767
rect 55675 721 55721 767
rect 55799 721 55845 767
rect 55923 721 55969 767
rect 56047 721 56093 767
rect 56171 721 56217 767
rect 56295 721 56341 767
rect 56419 721 56465 767
rect 56543 721 56589 767
rect 56667 721 56713 767
rect 56791 721 56837 767
rect 56915 721 56961 767
rect 57039 721 57085 767
rect 57163 721 57209 767
rect 57287 721 57333 767
rect 57411 721 57457 767
rect 57535 721 57581 767
rect 57659 721 57705 767
rect 57783 721 57829 767
rect 57907 721 57953 767
rect 58031 721 58077 767
rect 58155 721 58201 767
rect 58279 721 58325 767
rect 58403 721 58449 767
rect 58527 721 58573 767
rect 58651 721 58697 767
rect 58775 721 58821 767
rect 58899 721 58945 767
rect 59023 721 59069 767
rect 59147 721 59193 767
rect 59271 721 59317 767
rect 59395 721 59441 767
rect 59519 721 59565 767
rect 59643 721 59689 767
rect 59767 721 59813 767
rect 59891 721 59937 767
rect 60015 721 60061 767
rect 60139 721 60185 767
rect 60263 721 60309 767
rect 60387 721 60433 767
rect 60511 721 60557 767
rect 60635 721 60681 767
rect 60759 721 60805 767
rect 60883 721 60929 767
rect 61007 721 61053 767
rect 61131 721 61177 767
rect 61255 721 61301 767
rect 61379 721 61425 767
rect 61503 721 61549 767
rect 61627 721 61673 767
rect 61751 721 61797 767
rect 61875 721 61921 767
rect 61999 721 62045 767
rect 62123 721 62169 767
rect 62247 721 62293 767
rect 62371 721 62417 767
rect 62495 721 62541 767
rect 62619 721 62665 767
rect 62743 721 62789 767
rect 62867 721 62913 767
rect 62991 721 63037 767
rect 63115 721 63161 767
rect 63239 721 63285 767
rect 63363 721 63409 767
rect 63487 721 63533 767
rect 63611 721 63657 767
rect 63735 721 63781 767
rect 63859 721 63905 767
rect 63983 721 64029 767
rect 64107 721 64153 767
rect 64231 721 64277 767
rect 64355 721 64401 767
rect 64479 721 64525 767
rect 64603 721 64649 767
rect 64727 721 64773 767
rect 64851 721 64897 767
rect 64975 721 65021 767
rect 65099 721 65145 767
rect 65223 721 65269 767
rect 65347 721 65393 767
rect 65471 721 65517 767
rect 65595 721 65641 767
rect 65719 721 65765 767
rect 65843 721 65889 767
rect 65967 721 66013 767
rect 66091 721 66137 767
rect 66215 721 66261 767
rect 66339 721 66385 767
rect 66463 721 66509 767
rect 66587 721 66633 767
rect 66711 721 66757 767
rect 66835 721 66881 767
rect 66959 721 67005 767
rect 67083 721 67129 767
rect 67207 721 67253 767
rect 67331 721 67377 767
rect 67455 721 67501 767
rect 67579 721 67625 767
rect 67703 721 67749 767
rect 67827 721 67873 767
rect 67951 721 67997 767
rect 68075 721 68121 767
rect 68199 721 68245 767
rect 68323 721 68369 767
rect 68447 721 68493 767
rect 68571 721 68617 767
rect 68695 721 68741 767
rect 68819 721 68865 767
rect 68943 721 68989 767
rect 69067 721 69113 767
rect 69191 721 69237 767
rect 69315 721 69361 767
rect 69439 721 69485 767
rect 69563 721 69609 767
rect 69687 721 69733 767
rect 69811 721 69857 767
rect 69935 721 69981 767
rect 70059 721 70105 767
rect 70183 721 70229 767
rect 70307 721 70353 767
rect 70431 721 70477 767
rect 70555 721 70601 767
rect 70679 721 70725 767
rect 70803 721 70849 767
rect 70927 721 70973 767
rect 71051 721 71097 767
rect 71175 721 71221 767
rect 71299 721 71345 767
rect 71423 721 71469 767
rect 71547 721 71593 767
rect 71671 721 71717 767
rect 71795 721 71841 767
rect 71919 721 71965 767
rect 72043 721 72089 767
rect 72167 721 72213 767
rect 72291 721 72337 767
rect 72415 721 72461 767
rect 72539 721 72585 767
rect 72663 721 72709 767
rect 72787 721 72833 767
rect 72911 721 72957 767
rect 73035 721 73081 767
rect 73159 721 73205 767
rect 73283 721 73329 767
rect 73407 721 73453 767
rect 73531 721 73577 767
rect 73655 721 73701 767
rect 73779 721 73825 767
rect 73903 721 73949 767
rect 74027 721 74073 767
rect 74151 721 74197 767
rect 74275 721 74321 767
rect 74399 721 74445 767
rect 74523 721 74569 767
rect 74647 721 74693 767
rect 74771 721 74817 767
rect 74895 721 74941 767
rect 75019 721 75065 767
rect 75143 721 75189 767
rect 75267 721 75313 767
rect 75391 721 75437 767
rect 75515 721 75561 767
rect 75639 721 75685 767
rect 75763 721 75809 767
rect 75887 721 75933 767
rect 76011 721 76057 767
rect 76135 721 76181 767
rect 76259 721 76305 767
rect 76383 721 76429 767
rect 76507 721 76553 767
rect 76631 721 76677 767
rect 76755 721 76801 767
rect 76879 721 76925 767
rect 77003 721 77049 767
rect 77127 721 77173 767
rect 77251 721 77297 767
rect 77375 721 77421 767
rect 77499 721 77545 767
rect 77623 721 77669 767
rect 77747 721 77793 767
rect 77871 721 77917 767
rect 77995 721 78041 767
rect 78119 721 78165 767
rect 78243 721 78289 767
rect 78367 721 78413 767
rect 78491 721 78537 767
rect 78615 721 78661 767
rect 78739 721 78785 767
rect 78863 721 78909 767
rect 78987 721 79033 767
rect 79111 721 79157 767
rect 79235 721 79281 767
rect 79359 721 79405 767
rect 79483 721 79529 767
rect 79607 721 79653 767
rect 79731 721 79777 767
rect 79855 721 79901 767
rect 79979 721 80025 767
rect 80103 721 80149 767
rect 80227 721 80273 767
rect 80351 721 80397 767
rect 80475 721 80521 767
rect 80599 721 80645 767
rect 80723 721 80769 767
rect 80847 721 80893 767
rect 80971 721 81017 767
rect 81095 721 81141 767
rect 81219 721 81265 767
rect 81343 721 81389 767
rect 81467 721 81513 767
rect 81591 721 81637 767
rect 81715 721 81761 767
rect 81839 721 81885 767
rect 81963 721 82009 767
rect 82087 721 82133 767
rect 82211 721 82257 767
rect 82335 721 82381 767
rect 82459 721 82505 767
rect 82583 721 82629 767
rect 82707 721 82753 767
rect 82831 721 82877 767
rect 82955 721 83001 767
rect 83079 721 83125 767
rect 83203 721 83249 767
rect 83327 721 83373 767
rect 83451 721 83497 767
rect 83575 721 83621 767
rect 83699 721 83745 767
rect 83823 721 83869 767
rect 83947 721 83993 767
rect 84071 721 84117 767
rect 84195 721 84241 767
rect 84319 721 84365 767
rect 84443 721 84489 767
rect 84567 721 84613 767
rect 84691 721 84737 767
rect 84815 721 84861 767
rect 84939 721 84985 767
rect 85063 721 85109 767
rect 85187 721 85233 767
rect 85311 721 85357 767
rect 85435 721 85481 767
rect 85559 721 85605 767
rect 85683 721 85729 767
rect 85807 721 85853 767
rect 85931 721 85977 767
rect 371 597 417 643
rect 495 597 541 643
rect 619 597 665 643
rect 743 597 789 643
rect 867 597 913 643
rect 991 597 1037 643
rect 1115 597 1161 643
rect 1239 597 1285 643
rect 1363 597 1409 643
rect 1487 597 1533 643
rect 1611 597 1657 643
rect 1735 597 1781 643
rect 1859 597 1905 643
rect 1983 597 2029 643
rect 2107 597 2153 643
rect 2231 597 2277 643
rect 2355 597 2401 643
rect 2479 597 2525 643
rect 2603 597 2649 643
rect 2727 597 2773 643
rect 2851 597 2897 643
rect 2975 597 3021 643
rect 3099 597 3145 643
rect 3223 597 3269 643
rect 3347 597 3393 643
rect 3471 597 3517 643
rect 3595 597 3641 643
rect 3719 597 3765 643
rect 3843 597 3889 643
rect 3967 597 4013 643
rect 4091 597 4137 643
rect 4215 597 4261 643
rect 4339 597 4385 643
rect 4463 597 4509 643
rect 4587 597 4633 643
rect 4711 597 4757 643
rect 4835 597 4881 643
rect 4959 597 5005 643
rect 5083 597 5129 643
rect 5207 597 5253 643
rect 5331 597 5377 643
rect 5455 597 5501 643
rect 5579 597 5625 643
rect 5703 597 5749 643
rect 5827 597 5873 643
rect 5951 597 5997 643
rect 6075 597 6121 643
rect 6199 597 6245 643
rect 6323 597 6369 643
rect 6447 597 6493 643
rect 6571 597 6617 643
rect 6695 597 6741 643
rect 6819 597 6865 643
rect 6943 597 6989 643
rect 7067 597 7113 643
rect 7191 597 7237 643
rect 7315 597 7361 643
rect 7439 597 7485 643
rect 7563 597 7609 643
rect 7687 597 7733 643
rect 7811 597 7857 643
rect 7935 597 7981 643
rect 8059 597 8105 643
rect 8183 597 8229 643
rect 8307 597 8353 643
rect 8431 597 8477 643
rect 8555 597 8601 643
rect 8679 597 8725 643
rect 8803 597 8849 643
rect 8927 597 8973 643
rect 9051 597 9097 643
rect 9175 597 9221 643
rect 9299 597 9345 643
rect 9423 597 9469 643
rect 9547 597 9593 643
rect 9671 597 9717 643
rect 9795 597 9841 643
rect 9919 597 9965 643
rect 10043 597 10089 643
rect 10167 597 10213 643
rect 10291 597 10337 643
rect 10415 597 10461 643
rect 10539 597 10585 643
rect 10663 597 10709 643
rect 10787 597 10833 643
rect 10911 597 10957 643
rect 11035 597 11081 643
rect 11159 597 11205 643
rect 11283 597 11329 643
rect 11407 597 11453 643
rect 11531 597 11577 643
rect 11655 597 11701 643
rect 11779 597 11825 643
rect 11903 597 11949 643
rect 12027 597 12073 643
rect 12151 597 12197 643
rect 12275 597 12321 643
rect 12399 597 12445 643
rect 12523 597 12569 643
rect 12647 597 12693 643
rect 12771 597 12817 643
rect 12895 597 12941 643
rect 13019 597 13065 643
rect 13143 597 13189 643
rect 13267 597 13313 643
rect 13391 597 13437 643
rect 13515 597 13561 643
rect 13639 597 13685 643
rect 13763 597 13809 643
rect 13887 597 13933 643
rect 14011 597 14057 643
rect 14135 597 14181 643
rect 14259 597 14305 643
rect 14383 597 14429 643
rect 14507 597 14553 643
rect 14631 597 14677 643
rect 14755 597 14801 643
rect 14879 597 14925 643
rect 15003 597 15049 643
rect 15127 597 15173 643
rect 15251 597 15297 643
rect 15375 597 15421 643
rect 15499 597 15545 643
rect 15623 597 15669 643
rect 15747 597 15793 643
rect 15871 597 15917 643
rect 15995 597 16041 643
rect 16119 597 16165 643
rect 16243 597 16289 643
rect 16367 597 16413 643
rect 16491 597 16537 643
rect 16615 597 16661 643
rect 16739 597 16785 643
rect 16863 597 16909 643
rect 16987 597 17033 643
rect 17111 597 17157 643
rect 17235 597 17281 643
rect 17359 597 17405 643
rect 17483 597 17529 643
rect 17607 597 17653 643
rect 17731 597 17777 643
rect 17855 597 17901 643
rect 17979 597 18025 643
rect 18103 597 18149 643
rect 18227 597 18273 643
rect 18351 597 18397 643
rect 18475 597 18521 643
rect 18599 597 18645 643
rect 18723 597 18769 643
rect 18847 597 18893 643
rect 18971 597 19017 643
rect 19095 597 19141 643
rect 19219 597 19265 643
rect 19343 597 19389 643
rect 19467 597 19513 643
rect 19591 597 19637 643
rect 19715 597 19761 643
rect 19839 597 19885 643
rect 19963 597 20009 643
rect 20087 597 20133 643
rect 20211 597 20257 643
rect 20335 597 20381 643
rect 20459 597 20505 643
rect 20583 597 20629 643
rect 20707 597 20753 643
rect 20831 597 20877 643
rect 20955 597 21001 643
rect 21079 597 21125 643
rect 21203 597 21249 643
rect 21327 597 21373 643
rect 21451 597 21497 643
rect 21575 597 21621 643
rect 21699 597 21745 643
rect 21823 597 21869 643
rect 21947 597 21993 643
rect 22071 597 22117 643
rect 22195 597 22241 643
rect 22319 597 22365 643
rect 22443 597 22489 643
rect 22567 597 22613 643
rect 22691 597 22737 643
rect 22815 597 22861 643
rect 22939 597 22985 643
rect 23063 597 23109 643
rect 23187 597 23233 643
rect 23311 597 23357 643
rect 23435 597 23481 643
rect 23559 597 23605 643
rect 23683 597 23729 643
rect 23807 597 23853 643
rect 23931 597 23977 643
rect 24055 597 24101 643
rect 24179 597 24225 643
rect 24303 597 24349 643
rect 24427 597 24473 643
rect 24551 597 24597 643
rect 24675 597 24721 643
rect 24799 597 24845 643
rect 24923 597 24969 643
rect 25047 597 25093 643
rect 25171 597 25217 643
rect 25295 597 25341 643
rect 25419 597 25465 643
rect 25543 597 25589 643
rect 25667 597 25713 643
rect 25791 597 25837 643
rect 25915 597 25961 643
rect 26039 597 26085 643
rect 26163 597 26209 643
rect 26287 597 26333 643
rect 26411 597 26457 643
rect 26535 597 26581 643
rect 26659 597 26705 643
rect 26783 597 26829 643
rect 26907 597 26953 643
rect 27031 597 27077 643
rect 27155 597 27201 643
rect 27279 597 27325 643
rect 27403 597 27449 643
rect 27527 597 27573 643
rect 27651 597 27697 643
rect 27775 597 27821 643
rect 27899 597 27945 643
rect 28023 597 28069 643
rect 28147 597 28193 643
rect 28271 597 28317 643
rect 28395 597 28441 643
rect 28519 597 28565 643
rect 28643 597 28689 643
rect 28767 597 28813 643
rect 28891 597 28937 643
rect 29015 597 29061 643
rect 29139 597 29185 643
rect 29263 597 29309 643
rect 29387 597 29433 643
rect 29511 597 29557 643
rect 29635 597 29681 643
rect 29759 597 29805 643
rect 29883 597 29929 643
rect 30007 597 30053 643
rect 30131 597 30177 643
rect 30255 597 30301 643
rect 30379 597 30425 643
rect 30503 597 30549 643
rect 30627 597 30673 643
rect 30751 597 30797 643
rect 30875 597 30921 643
rect 30999 597 31045 643
rect 31123 597 31169 643
rect 31247 597 31293 643
rect 31371 597 31417 643
rect 31495 597 31541 643
rect 31619 597 31665 643
rect 31743 597 31789 643
rect 31867 597 31913 643
rect 31991 597 32037 643
rect 32115 597 32161 643
rect 32239 597 32285 643
rect 32363 597 32409 643
rect 32487 597 32533 643
rect 32611 597 32657 643
rect 32735 597 32781 643
rect 32859 597 32905 643
rect 32983 597 33029 643
rect 33107 597 33153 643
rect 33231 597 33277 643
rect 33355 597 33401 643
rect 33479 597 33525 643
rect 33603 597 33649 643
rect 33727 597 33773 643
rect 33851 597 33897 643
rect 33975 597 34021 643
rect 34099 597 34145 643
rect 34223 597 34269 643
rect 34347 597 34393 643
rect 34471 597 34517 643
rect 34595 597 34641 643
rect 34719 597 34765 643
rect 34843 597 34889 643
rect 34967 597 35013 643
rect 35091 597 35137 643
rect 35215 597 35261 643
rect 35339 597 35385 643
rect 35463 597 35509 643
rect 35587 597 35633 643
rect 35711 597 35757 643
rect 35835 597 35881 643
rect 35959 597 36005 643
rect 36083 597 36129 643
rect 36207 597 36253 643
rect 36331 597 36377 643
rect 36455 597 36501 643
rect 36579 597 36625 643
rect 36703 597 36749 643
rect 36827 597 36873 643
rect 36951 597 36997 643
rect 37075 597 37121 643
rect 37199 597 37245 643
rect 37323 597 37369 643
rect 37447 597 37493 643
rect 37571 597 37617 643
rect 37695 597 37741 643
rect 37819 597 37865 643
rect 37943 597 37989 643
rect 38067 597 38113 643
rect 38191 597 38237 643
rect 38315 597 38361 643
rect 38439 597 38485 643
rect 38563 597 38609 643
rect 38687 597 38733 643
rect 38811 597 38857 643
rect 38935 597 38981 643
rect 39059 597 39105 643
rect 39183 597 39229 643
rect 39307 597 39353 643
rect 39431 597 39477 643
rect 39555 597 39601 643
rect 39679 597 39725 643
rect 39803 597 39849 643
rect 39927 597 39973 643
rect 40051 597 40097 643
rect 40175 597 40221 643
rect 40299 597 40345 643
rect 40423 597 40469 643
rect 40547 597 40593 643
rect 40671 597 40717 643
rect 40795 597 40841 643
rect 40919 597 40965 643
rect 41043 597 41089 643
rect 41167 597 41213 643
rect 41291 597 41337 643
rect 41415 597 41461 643
rect 41539 597 41585 643
rect 41663 597 41709 643
rect 41787 597 41833 643
rect 41911 597 41957 643
rect 42035 597 42081 643
rect 42159 597 42205 643
rect 42283 597 42329 643
rect 42407 597 42453 643
rect 42531 597 42577 643
rect 42655 597 42701 643
rect 42779 597 42825 643
rect 42903 597 42949 643
rect 43027 597 43073 643
rect 43151 597 43197 643
rect 43275 597 43321 643
rect 43399 597 43445 643
rect 43523 597 43569 643
rect 43647 597 43693 643
rect 43771 597 43817 643
rect 43895 597 43941 643
rect 44019 597 44065 643
rect 44143 597 44189 643
rect 44267 597 44313 643
rect 44391 597 44437 643
rect 44515 597 44561 643
rect 44639 597 44685 643
rect 44763 597 44809 643
rect 44887 597 44933 643
rect 45011 597 45057 643
rect 45135 597 45181 643
rect 45259 597 45305 643
rect 45383 597 45429 643
rect 45507 597 45553 643
rect 45631 597 45677 643
rect 45755 597 45801 643
rect 45879 597 45925 643
rect 46003 597 46049 643
rect 46127 597 46173 643
rect 46251 597 46297 643
rect 46375 597 46421 643
rect 46499 597 46545 643
rect 46623 597 46669 643
rect 46747 597 46793 643
rect 46871 597 46917 643
rect 46995 597 47041 643
rect 47119 597 47165 643
rect 47243 597 47289 643
rect 47367 597 47413 643
rect 47491 597 47537 643
rect 47615 597 47661 643
rect 47739 597 47785 643
rect 47863 597 47909 643
rect 47987 597 48033 643
rect 48111 597 48157 643
rect 48235 597 48281 643
rect 48359 597 48405 643
rect 48483 597 48529 643
rect 48607 597 48653 643
rect 48731 597 48777 643
rect 48855 597 48901 643
rect 48979 597 49025 643
rect 49103 597 49149 643
rect 49227 597 49273 643
rect 49351 597 49397 643
rect 49475 597 49521 643
rect 49599 597 49645 643
rect 49723 597 49769 643
rect 49847 597 49893 643
rect 49971 597 50017 643
rect 50095 597 50141 643
rect 50219 597 50265 643
rect 50343 597 50389 643
rect 50467 597 50513 643
rect 50591 597 50637 643
rect 50715 597 50761 643
rect 50839 597 50885 643
rect 50963 597 51009 643
rect 51087 597 51133 643
rect 51211 597 51257 643
rect 51335 597 51381 643
rect 51459 597 51505 643
rect 51583 597 51629 643
rect 51707 597 51753 643
rect 51831 597 51877 643
rect 51955 597 52001 643
rect 52079 597 52125 643
rect 52203 597 52249 643
rect 52327 597 52373 643
rect 52451 597 52497 643
rect 52575 597 52621 643
rect 52699 597 52745 643
rect 52823 597 52869 643
rect 52947 597 52993 643
rect 53071 597 53117 643
rect 53195 597 53241 643
rect 53319 597 53365 643
rect 53443 597 53489 643
rect 53567 597 53613 643
rect 53691 597 53737 643
rect 53815 597 53861 643
rect 53939 597 53985 643
rect 54063 597 54109 643
rect 54187 597 54233 643
rect 54311 597 54357 643
rect 54435 597 54481 643
rect 54559 597 54605 643
rect 54683 597 54729 643
rect 54807 597 54853 643
rect 54931 597 54977 643
rect 55055 597 55101 643
rect 55179 597 55225 643
rect 55303 597 55349 643
rect 55427 597 55473 643
rect 55551 597 55597 643
rect 55675 597 55721 643
rect 55799 597 55845 643
rect 55923 597 55969 643
rect 56047 597 56093 643
rect 56171 597 56217 643
rect 56295 597 56341 643
rect 56419 597 56465 643
rect 56543 597 56589 643
rect 56667 597 56713 643
rect 56791 597 56837 643
rect 56915 597 56961 643
rect 57039 597 57085 643
rect 57163 597 57209 643
rect 57287 597 57333 643
rect 57411 597 57457 643
rect 57535 597 57581 643
rect 57659 597 57705 643
rect 57783 597 57829 643
rect 57907 597 57953 643
rect 58031 597 58077 643
rect 58155 597 58201 643
rect 58279 597 58325 643
rect 58403 597 58449 643
rect 58527 597 58573 643
rect 58651 597 58697 643
rect 58775 597 58821 643
rect 58899 597 58945 643
rect 59023 597 59069 643
rect 59147 597 59193 643
rect 59271 597 59317 643
rect 59395 597 59441 643
rect 59519 597 59565 643
rect 59643 597 59689 643
rect 59767 597 59813 643
rect 59891 597 59937 643
rect 60015 597 60061 643
rect 60139 597 60185 643
rect 60263 597 60309 643
rect 60387 597 60433 643
rect 60511 597 60557 643
rect 60635 597 60681 643
rect 60759 597 60805 643
rect 60883 597 60929 643
rect 61007 597 61053 643
rect 61131 597 61177 643
rect 61255 597 61301 643
rect 61379 597 61425 643
rect 61503 597 61549 643
rect 61627 597 61673 643
rect 61751 597 61797 643
rect 61875 597 61921 643
rect 61999 597 62045 643
rect 62123 597 62169 643
rect 62247 597 62293 643
rect 62371 597 62417 643
rect 62495 597 62541 643
rect 62619 597 62665 643
rect 62743 597 62789 643
rect 62867 597 62913 643
rect 62991 597 63037 643
rect 63115 597 63161 643
rect 63239 597 63285 643
rect 63363 597 63409 643
rect 63487 597 63533 643
rect 63611 597 63657 643
rect 63735 597 63781 643
rect 63859 597 63905 643
rect 63983 597 64029 643
rect 64107 597 64153 643
rect 64231 597 64277 643
rect 64355 597 64401 643
rect 64479 597 64525 643
rect 64603 597 64649 643
rect 64727 597 64773 643
rect 64851 597 64897 643
rect 64975 597 65021 643
rect 65099 597 65145 643
rect 65223 597 65269 643
rect 65347 597 65393 643
rect 65471 597 65517 643
rect 65595 597 65641 643
rect 65719 597 65765 643
rect 65843 597 65889 643
rect 65967 597 66013 643
rect 66091 597 66137 643
rect 66215 597 66261 643
rect 66339 597 66385 643
rect 66463 597 66509 643
rect 66587 597 66633 643
rect 66711 597 66757 643
rect 66835 597 66881 643
rect 66959 597 67005 643
rect 67083 597 67129 643
rect 67207 597 67253 643
rect 67331 597 67377 643
rect 67455 597 67501 643
rect 67579 597 67625 643
rect 67703 597 67749 643
rect 67827 597 67873 643
rect 67951 597 67997 643
rect 68075 597 68121 643
rect 68199 597 68245 643
rect 68323 597 68369 643
rect 68447 597 68493 643
rect 68571 597 68617 643
rect 68695 597 68741 643
rect 68819 597 68865 643
rect 68943 597 68989 643
rect 69067 597 69113 643
rect 69191 597 69237 643
rect 69315 597 69361 643
rect 69439 597 69485 643
rect 69563 597 69609 643
rect 69687 597 69733 643
rect 69811 597 69857 643
rect 69935 597 69981 643
rect 70059 597 70105 643
rect 70183 597 70229 643
rect 70307 597 70353 643
rect 70431 597 70477 643
rect 70555 597 70601 643
rect 70679 597 70725 643
rect 70803 597 70849 643
rect 70927 597 70973 643
rect 71051 597 71097 643
rect 71175 597 71221 643
rect 71299 597 71345 643
rect 71423 597 71469 643
rect 71547 597 71593 643
rect 71671 597 71717 643
rect 71795 597 71841 643
rect 71919 597 71965 643
rect 72043 597 72089 643
rect 72167 597 72213 643
rect 72291 597 72337 643
rect 72415 597 72461 643
rect 72539 597 72585 643
rect 72663 597 72709 643
rect 72787 597 72833 643
rect 72911 597 72957 643
rect 73035 597 73081 643
rect 73159 597 73205 643
rect 73283 597 73329 643
rect 73407 597 73453 643
rect 73531 597 73577 643
rect 73655 597 73701 643
rect 73779 597 73825 643
rect 73903 597 73949 643
rect 74027 597 74073 643
rect 74151 597 74197 643
rect 74275 597 74321 643
rect 74399 597 74445 643
rect 74523 597 74569 643
rect 74647 597 74693 643
rect 74771 597 74817 643
rect 74895 597 74941 643
rect 75019 597 75065 643
rect 75143 597 75189 643
rect 75267 597 75313 643
rect 75391 597 75437 643
rect 75515 597 75561 643
rect 75639 597 75685 643
rect 75763 597 75809 643
rect 75887 597 75933 643
rect 76011 597 76057 643
rect 76135 597 76181 643
rect 76259 597 76305 643
rect 76383 597 76429 643
rect 76507 597 76553 643
rect 76631 597 76677 643
rect 76755 597 76801 643
rect 76879 597 76925 643
rect 77003 597 77049 643
rect 77127 597 77173 643
rect 77251 597 77297 643
rect 77375 597 77421 643
rect 77499 597 77545 643
rect 77623 597 77669 643
rect 77747 597 77793 643
rect 77871 597 77917 643
rect 77995 597 78041 643
rect 78119 597 78165 643
rect 78243 597 78289 643
rect 78367 597 78413 643
rect 78491 597 78537 643
rect 78615 597 78661 643
rect 78739 597 78785 643
rect 78863 597 78909 643
rect 78987 597 79033 643
rect 79111 597 79157 643
rect 79235 597 79281 643
rect 79359 597 79405 643
rect 79483 597 79529 643
rect 79607 597 79653 643
rect 79731 597 79777 643
rect 79855 597 79901 643
rect 79979 597 80025 643
rect 80103 597 80149 643
rect 80227 597 80273 643
rect 80351 597 80397 643
rect 80475 597 80521 643
rect 80599 597 80645 643
rect 80723 597 80769 643
rect 80847 597 80893 643
rect 80971 597 81017 643
rect 81095 597 81141 643
rect 81219 597 81265 643
rect 81343 597 81389 643
rect 81467 597 81513 643
rect 81591 597 81637 643
rect 81715 597 81761 643
rect 81839 597 81885 643
rect 81963 597 82009 643
rect 82087 597 82133 643
rect 82211 597 82257 643
rect 82335 597 82381 643
rect 82459 597 82505 643
rect 82583 597 82629 643
rect 82707 597 82753 643
rect 82831 597 82877 643
rect 82955 597 83001 643
rect 83079 597 83125 643
rect 83203 597 83249 643
rect 83327 597 83373 643
rect 83451 597 83497 643
rect 83575 597 83621 643
rect 83699 597 83745 643
rect 83823 597 83869 643
rect 83947 597 83993 643
rect 84071 597 84117 643
rect 84195 597 84241 643
rect 84319 597 84365 643
rect 84443 597 84489 643
rect 84567 597 84613 643
rect 84691 597 84737 643
rect 84815 597 84861 643
rect 84939 597 84985 643
rect 85063 597 85109 643
rect 85187 597 85233 643
rect 85311 597 85357 643
rect 85435 597 85481 643
rect 85559 597 85605 643
rect 85683 597 85729 643
rect 85807 597 85853 643
rect 85931 597 85977 643
<< mvnsubdiffcont >>
rect 30854 44190 30900 44236
rect 31012 44190 31058 44236
rect 31170 44190 31216 44236
rect 31328 44190 31374 44236
rect 31487 44190 31533 44236
rect 31645 44190 31691 44236
rect 31803 44190 31849 44236
rect 31961 44190 32007 44236
rect 32119 44190 32165 44236
rect 32277 44190 32323 44236
rect 32435 44190 32481 44236
rect 32593 44190 32639 44236
rect 42717 44263 42763 44309
rect 42875 44263 42921 44309
rect 43033 44263 43079 44309
rect 43191 44263 43237 44309
rect 43350 44263 43396 44309
rect 43508 44263 43554 44309
rect 30637 44076 30683 44122
rect 30854 44027 30900 44073
rect 31012 44027 31058 44073
rect 31170 44027 31216 44073
rect 31328 44027 31374 44073
rect 31487 44027 31533 44073
rect 31645 44027 31691 44073
rect 31803 44027 31849 44073
rect 31961 44027 32007 44073
rect 32119 44027 32165 44073
rect 32277 44027 32323 44073
rect 32435 44027 32481 44073
rect 32593 44027 32639 44073
rect 30637 43912 30683 43958
rect 30854 43863 30900 43909
rect 31012 43863 31058 43909
rect 31170 43863 31216 43909
rect 31328 43863 31374 43909
rect 31487 43863 31533 43909
rect 31645 43863 31691 43909
rect 31803 43863 31849 43909
rect 31961 43863 32007 43909
rect 32119 43863 32165 43909
rect 32277 43863 32323 43909
rect 32435 43863 32481 43909
rect 32593 43863 32639 43909
rect 52483 44190 52529 44236
rect 52641 44190 52687 44236
rect 52799 44190 52845 44236
rect 52957 44190 53003 44236
rect 53115 44190 53161 44236
rect 53273 44190 53319 44236
rect 53431 44190 53477 44236
rect 53589 44190 53635 44236
rect 53748 44190 53794 44236
rect 53906 44190 53952 44236
rect 54064 44190 54110 44236
rect 54222 44190 54268 44236
rect 30637 43749 30683 43795
rect 30854 43700 30900 43746
rect 31012 43700 31058 43746
rect 31170 43700 31216 43746
rect 31328 43700 31374 43746
rect 31487 43700 31533 43746
rect 31645 43700 31691 43746
rect 31803 43700 31849 43746
rect 31961 43700 32007 43746
rect 32119 43700 32165 43746
rect 32277 43700 32323 43746
rect 32435 43700 32481 43746
rect 32593 43700 32639 43746
rect 54440 44076 54486 44122
rect 52483 44027 52529 44073
rect 52641 44027 52687 44073
rect 52799 44027 52845 44073
rect 52957 44027 53003 44073
rect 53115 44027 53161 44073
rect 53273 44027 53319 44073
rect 53431 44027 53477 44073
rect 53589 44027 53635 44073
rect 53748 44027 53794 44073
rect 53906 44027 53952 44073
rect 54064 44027 54110 44073
rect 54222 44027 54268 44073
rect 54440 43912 54486 43958
rect 52483 43863 52529 43909
rect 52641 43863 52687 43909
rect 52799 43863 52845 43909
rect 52957 43863 53003 43909
rect 53115 43863 53161 43909
rect 53273 43863 53319 43909
rect 53431 43863 53477 43909
rect 53589 43863 53635 43909
rect 53748 43863 53794 43909
rect 53906 43863 53952 43909
rect 54064 43863 54110 43909
rect 54222 43863 54268 43909
rect 54440 43749 54486 43795
rect 52483 43700 52529 43746
rect 52641 43700 52687 43746
rect 52799 43700 52845 43746
rect 52957 43700 53003 43746
rect 53115 43700 53161 43746
rect 53273 43700 53319 43746
rect 53431 43700 53477 43746
rect 53589 43700 53635 43746
rect 53748 43700 53794 43746
rect 53906 43700 53952 43746
rect 54064 43700 54110 43746
rect 54222 43700 54268 43746
rect 30637 43586 30683 43632
rect 30637 43422 30683 43468
rect 54440 43586 54486 43632
rect 54440 43422 54486 43468
rect 36489 43304 36723 43350
rect 30637 43220 30683 43266
rect 30855 43180 30901 43226
rect 30637 43057 30683 43103
rect 30855 43016 30901 43062
rect 30637 42894 30683 42940
rect 30855 42853 30901 42899
rect 30637 42731 30683 42777
rect 30855 42690 30901 42736
rect 39062 43304 39108 43350
rect 39220 43304 39266 43350
rect 45619 43304 45665 43350
rect 45777 43304 45823 43350
rect 45935 43304 45981 43350
rect 46093 43304 46139 43350
rect 46251 43304 46297 43350
rect 46409 43304 46455 43350
rect 46568 43304 46614 43350
rect 46726 43304 46772 43350
rect 46884 43304 46930 43350
rect 47042 43304 47088 43350
rect 47200 43304 47246 43350
rect 47358 43304 47404 43350
rect 47516 43304 47562 43350
rect 47675 43304 47721 43350
rect 47833 43304 47879 43350
rect 47991 43304 48037 43350
rect 48149 43304 48195 43350
rect 48307 43304 48353 43350
rect 48465 43304 48511 43350
rect 45619 43140 45665 43186
rect 45777 43140 45823 43186
rect 45935 43140 45981 43186
rect 46093 43140 46139 43186
rect 46251 43140 46297 43186
rect 46409 43140 46455 43186
rect 46568 43140 46614 43186
rect 46726 43140 46772 43186
rect 46884 43140 46930 43186
rect 47042 43140 47088 43186
rect 47200 43140 47246 43186
rect 47358 43140 47404 43186
rect 47516 43140 47562 43186
rect 47675 43140 47721 43186
rect 47833 43140 47879 43186
rect 47991 43140 48037 43186
rect 48149 43140 48195 43186
rect 48307 43140 48353 43186
rect 48465 43140 48511 43186
rect 54223 43180 54269 43226
rect 54440 43220 54486 43266
rect 30637 42567 30683 42613
rect 30855 42527 30901 42573
rect 54223 43016 54269 43062
rect 54440 43057 54486 43103
rect 54440 42894 54486 42940
rect 54440 42731 54486 42777
rect 54223 42527 54269 42573
rect 54440 42567 54486 42613
rect 30637 42404 30683 42450
rect 54440 42404 54486 42450
rect 30637 42241 30683 42287
rect 30855 42281 30901 42327
rect 30637 42077 30683 42123
rect 30855 42118 30901 42164
rect 30637 41914 30683 41960
rect 30855 41955 30901 42001
rect 30637 41751 30683 41797
rect 30855 41792 30901 41838
rect 30637 41588 30683 41634
rect 30855 41628 30901 41674
rect 54223 42281 54269 42327
rect 54440 42241 54486 42287
rect 36489 41504 36723 41550
rect 30637 41420 30683 41466
rect 30855 41380 30901 41426
rect 30637 41257 30683 41303
rect 30855 41216 30901 41262
rect 30637 41094 30683 41140
rect 30855 41053 30901 41099
rect 30637 40931 30683 40977
rect 30855 40890 30901 40936
rect 39062 41504 39108 41550
rect 39220 41504 39266 41550
rect 45619 41668 45665 41714
rect 45777 41668 45823 41714
rect 45935 41668 45981 41714
rect 46093 41668 46139 41714
rect 46251 41668 46297 41714
rect 46409 41668 46455 41714
rect 46568 41668 46614 41714
rect 46726 41668 46772 41714
rect 46884 41668 46930 41714
rect 47042 41668 47088 41714
rect 47200 41668 47246 41714
rect 47358 41668 47404 41714
rect 47516 41668 47562 41714
rect 47675 41668 47721 41714
rect 47833 41668 47879 41714
rect 47991 41668 48037 41714
rect 48149 41668 48195 41714
rect 48307 41668 48353 41714
rect 48465 41668 48511 41714
rect 54440 42077 54486 42123
rect 54440 41914 54486 41960
rect 54223 41792 54269 41838
rect 54440 41751 54486 41797
rect 54223 41628 54269 41674
rect 54440 41588 54486 41634
rect 45619 41504 45665 41550
rect 45777 41504 45823 41550
rect 45935 41504 45981 41550
rect 46093 41504 46139 41550
rect 46251 41504 46297 41550
rect 46409 41504 46455 41550
rect 46568 41504 46614 41550
rect 46726 41504 46772 41550
rect 46884 41504 46930 41550
rect 47042 41504 47088 41550
rect 47200 41504 47246 41550
rect 47358 41504 47404 41550
rect 47516 41504 47562 41550
rect 47675 41504 47721 41550
rect 47833 41504 47879 41550
rect 47991 41504 48037 41550
rect 48149 41504 48195 41550
rect 48307 41504 48353 41550
rect 48465 41504 48511 41550
rect 45619 41340 45665 41386
rect 45777 41340 45823 41386
rect 45935 41340 45981 41386
rect 46093 41340 46139 41386
rect 46251 41340 46297 41386
rect 46409 41340 46455 41386
rect 46568 41340 46614 41386
rect 46726 41340 46772 41386
rect 46884 41340 46930 41386
rect 47042 41340 47088 41386
rect 47200 41340 47246 41386
rect 47358 41340 47404 41386
rect 47516 41340 47562 41386
rect 47675 41340 47721 41386
rect 47833 41340 47879 41386
rect 47991 41340 48037 41386
rect 48149 41340 48195 41386
rect 48307 41340 48353 41386
rect 48465 41340 48511 41386
rect 54223 41380 54269 41426
rect 54440 41420 54486 41466
rect 30637 40767 30683 40813
rect 30855 40727 30901 40773
rect 54223 41216 54269 41262
rect 54440 41257 54486 41303
rect 54440 41094 54486 41140
rect 54440 40931 54486 40977
rect 54223 40727 54269 40773
rect 54440 40767 54486 40813
rect 30637 40604 30683 40650
rect 54440 40604 54486 40650
rect 30637 40441 30683 40487
rect 30855 40481 30901 40527
rect 30637 40277 30683 40323
rect 30855 40318 30901 40364
rect 30637 40114 30683 40160
rect 30855 40155 30901 40201
rect 30637 39951 30683 39997
rect 30855 39992 30901 40038
rect 30637 39788 30683 39834
rect 30855 39828 30901 39874
rect 54223 40481 54269 40527
rect 54440 40441 54486 40487
rect 36489 39704 36723 39750
rect 30637 39620 30683 39666
rect 30855 39580 30901 39626
rect 30637 39457 30683 39503
rect 30855 39416 30901 39462
rect 30637 39294 30683 39340
rect 30855 39253 30901 39299
rect 30637 39131 30683 39177
rect 30855 39090 30901 39136
rect 39062 39704 39108 39750
rect 39220 39704 39266 39750
rect 45619 39868 45665 39914
rect 45777 39868 45823 39914
rect 45935 39868 45981 39914
rect 46093 39868 46139 39914
rect 46251 39868 46297 39914
rect 46409 39868 46455 39914
rect 46568 39868 46614 39914
rect 46726 39868 46772 39914
rect 46884 39868 46930 39914
rect 47042 39868 47088 39914
rect 47200 39868 47246 39914
rect 47358 39868 47404 39914
rect 47516 39868 47562 39914
rect 47675 39868 47721 39914
rect 47833 39868 47879 39914
rect 47991 39868 48037 39914
rect 48149 39868 48195 39914
rect 48307 39868 48353 39914
rect 48465 39868 48511 39914
rect 54440 40277 54486 40323
rect 54440 40114 54486 40160
rect 54223 39992 54269 40038
rect 54440 39951 54486 39997
rect 54223 39828 54269 39874
rect 54440 39788 54486 39834
rect 45619 39704 45665 39750
rect 45777 39704 45823 39750
rect 45935 39704 45981 39750
rect 46093 39704 46139 39750
rect 46251 39704 46297 39750
rect 46409 39704 46455 39750
rect 46568 39704 46614 39750
rect 46726 39704 46772 39750
rect 46884 39704 46930 39750
rect 47042 39704 47088 39750
rect 47200 39704 47246 39750
rect 47358 39704 47404 39750
rect 47516 39704 47562 39750
rect 47675 39704 47721 39750
rect 47833 39704 47879 39750
rect 47991 39704 48037 39750
rect 48149 39704 48195 39750
rect 48307 39704 48353 39750
rect 48465 39704 48511 39750
rect 45619 39540 45665 39586
rect 45777 39540 45823 39586
rect 45935 39540 45981 39586
rect 46093 39540 46139 39586
rect 46251 39540 46297 39586
rect 46409 39540 46455 39586
rect 46568 39540 46614 39586
rect 46726 39540 46772 39586
rect 46884 39540 46930 39586
rect 47042 39540 47088 39586
rect 47200 39540 47246 39586
rect 47358 39540 47404 39586
rect 47516 39540 47562 39586
rect 47675 39540 47721 39586
rect 47833 39540 47879 39586
rect 47991 39540 48037 39586
rect 48149 39540 48195 39586
rect 48307 39540 48353 39586
rect 48465 39540 48511 39586
rect 54223 39580 54269 39626
rect 54440 39620 54486 39666
rect 30637 38967 30683 39013
rect 30855 38927 30901 38973
rect 54223 39416 54269 39462
rect 54440 39457 54486 39503
rect 54440 39294 54486 39340
rect 54440 39131 54486 39177
rect 54223 38927 54269 38973
rect 54440 38967 54486 39013
rect 30637 38804 30683 38850
rect 54440 38804 54486 38850
rect 30637 38641 30683 38687
rect 30855 38681 30901 38727
rect 30637 38477 30683 38523
rect 30855 38518 30901 38564
rect 30637 38314 30683 38360
rect 30855 38355 30901 38401
rect 30637 38151 30683 38197
rect 30855 38192 30901 38238
rect 30637 37988 30683 38034
rect 30855 38028 30901 38074
rect 54223 38681 54269 38727
rect 54440 38641 54486 38687
rect 36489 37904 36723 37950
rect 30637 37820 30683 37866
rect 30855 37780 30901 37826
rect 30637 37657 30683 37703
rect 30855 37616 30901 37662
rect 30637 37494 30683 37540
rect 30855 37453 30901 37499
rect 30637 37331 30683 37377
rect 30855 37290 30901 37336
rect 39062 37904 39108 37950
rect 39220 37904 39266 37950
rect 45619 38068 45665 38114
rect 45777 38068 45823 38114
rect 45935 38068 45981 38114
rect 46093 38068 46139 38114
rect 46251 38068 46297 38114
rect 46409 38068 46455 38114
rect 46568 38068 46614 38114
rect 46726 38068 46772 38114
rect 46884 38068 46930 38114
rect 47042 38068 47088 38114
rect 47200 38068 47246 38114
rect 47358 38068 47404 38114
rect 47516 38068 47562 38114
rect 47675 38068 47721 38114
rect 47833 38068 47879 38114
rect 47991 38068 48037 38114
rect 48149 38068 48195 38114
rect 48307 38068 48353 38114
rect 48465 38068 48511 38114
rect 54440 38477 54486 38523
rect 54440 38314 54486 38360
rect 54223 38192 54269 38238
rect 54440 38151 54486 38197
rect 54223 38028 54269 38074
rect 54440 37988 54486 38034
rect 45619 37904 45665 37950
rect 45777 37904 45823 37950
rect 45935 37904 45981 37950
rect 46093 37904 46139 37950
rect 46251 37904 46297 37950
rect 46409 37904 46455 37950
rect 46568 37904 46614 37950
rect 46726 37904 46772 37950
rect 46884 37904 46930 37950
rect 47042 37904 47088 37950
rect 47200 37904 47246 37950
rect 47358 37904 47404 37950
rect 47516 37904 47562 37950
rect 47675 37904 47721 37950
rect 47833 37904 47879 37950
rect 47991 37904 48037 37950
rect 48149 37904 48195 37950
rect 48307 37904 48353 37950
rect 48465 37904 48511 37950
rect 45619 37740 45665 37786
rect 45777 37740 45823 37786
rect 45935 37740 45981 37786
rect 46093 37740 46139 37786
rect 46251 37740 46297 37786
rect 46409 37740 46455 37786
rect 46568 37740 46614 37786
rect 46726 37740 46772 37786
rect 46884 37740 46930 37786
rect 47042 37740 47088 37786
rect 47200 37740 47246 37786
rect 47358 37740 47404 37786
rect 47516 37740 47562 37786
rect 47675 37740 47721 37786
rect 47833 37740 47879 37786
rect 47991 37740 48037 37786
rect 48149 37740 48195 37786
rect 48307 37740 48353 37786
rect 48465 37740 48511 37786
rect 54223 37780 54269 37826
rect 54440 37820 54486 37866
rect 30637 37167 30683 37213
rect 30855 37127 30901 37173
rect 54223 37616 54269 37662
rect 54440 37657 54486 37703
rect 54440 37494 54486 37540
rect 54440 37331 54486 37377
rect 54223 37127 54269 37173
rect 54440 37167 54486 37213
rect 30637 37004 30683 37050
rect 54440 37004 54486 37050
rect 30637 36841 30683 36887
rect 30855 36881 30901 36927
rect 30637 36677 30683 36723
rect 30855 36718 30901 36764
rect 30637 36514 30683 36560
rect 30855 36555 30901 36601
rect 30637 36351 30683 36397
rect 30855 36392 30901 36438
rect 30637 36188 30683 36234
rect 30855 36228 30901 36274
rect 54223 36881 54269 36927
rect 54440 36841 54486 36887
rect 36489 36104 36723 36150
rect 39062 36104 39108 36150
rect 39220 36104 39266 36150
rect 45619 36268 45665 36314
rect 45777 36268 45823 36314
rect 45935 36268 45981 36314
rect 46093 36268 46139 36314
rect 46251 36268 46297 36314
rect 46409 36268 46455 36314
rect 46568 36268 46614 36314
rect 46726 36268 46772 36314
rect 46884 36268 46930 36314
rect 47042 36268 47088 36314
rect 47200 36268 47246 36314
rect 47358 36268 47404 36314
rect 47516 36268 47562 36314
rect 47675 36268 47721 36314
rect 47833 36268 47879 36314
rect 47991 36268 48037 36314
rect 48149 36268 48195 36314
rect 48307 36268 48353 36314
rect 48465 36268 48511 36314
rect 54440 36677 54486 36723
rect 54440 36514 54486 36560
rect 54223 36392 54269 36438
rect 54440 36351 54486 36397
rect 54223 36228 54269 36274
rect 54440 36188 54486 36234
rect 45619 36104 45665 36150
rect 45777 36104 45823 36150
rect 45935 36104 45981 36150
rect 46093 36104 46139 36150
rect 46251 36104 46297 36150
rect 46409 36104 46455 36150
rect 46568 36104 46614 36150
rect 46726 36104 46772 36150
rect 46884 36104 46930 36150
rect 47042 36104 47088 36150
rect 47200 36104 47246 36150
rect 47358 36104 47404 36150
rect 47516 36104 47562 36150
rect 47675 36104 47721 36150
rect 47833 36104 47879 36150
rect 47991 36104 48037 36150
rect 48149 36104 48195 36150
rect 48307 36104 48353 36150
rect 48465 36104 48511 36150
<< polysilicon >>
rect 29072 44044 29274 44171
rect 29072 43998 29116 44044
rect 29162 43998 29274 44044
rect 29072 43881 29274 43998
rect 29072 43835 29116 43881
rect 29162 43835 29274 43881
rect 29072 43717 29274 43835
rect 29072 43671 29116 43717
rect 29162 43671 29274 43717
rect 29072 43554 29274 43671
rect 29072 43508 29116 43554
rect 29162 43508 29274 43554
rect 29072 43383 29274 43508
rect 30373 43383 30444 44171
rect 42300 44243 42478 44262
rect 42300 44197 42319 44243
rect 42459 44197 42478 44243
rect 44041 44291 44144 44310
rect 44041 44245 44067 44291
rect 44113 44245 44144 44291
rect 42300 44178 42478 44197
rect 37991 44143 38125 44150
rect 35233 44023 35396 44143
rect 37922 44045 38125 44143
rect 37922 44023 38035 44045
rect 35233 43919 35336 44023
rect 37991 43919 38035 44023
rect 32932 43799 33001 43919
rect 35023 43799 35396 43919
rect 37922 43905 38035 43919
rect 38081 43905 38125 44045
rect 40675 43958 40759 43977
rect 40675 43919 40694 43958
rect 37922 43800 38125 43905
rect 37922 43799 37993 43800
rect 38292 43799 38363 43919
rect 39681 43799 40062 43919
rect 40590 43818 40694 43919
rect 40740 43818 40759 43958
rect 42341 43920 42445 44178
rect 40590 43799 40759 43818
rect 40892 43800 40963 43920
rect 42281 43800 42445 43920
rect 44041 43919 44144 44245
rect 46948 44033 47101 44143
rect 42592 43799 42663 43919
rect 43981 43799 44144 43919
rect 44260 43998 44344 44017
rect 44260 43858 44279 43998
rect 44325 43919 44344 43998
rect 44325 43858 44432 43919
rect 44260 43799 44432 43858
rect 44960 43799 45333 43919
rect 46651 43799 46722 43919
rect 46948 43893 46967 44033
rect 47013 44023 47101 44033
rect 49627 44023 49790 44143
rect 47013 43919 47032 44023
rect 49687 43919 49790 44023
rect 47013 43893 47101 43919
rect 46948 43799 47101 43893
rect 49627 43799 50001 43919
rect 52023 43799 52094 43919
rect 29072 43144 29274 43271
rect 29072 43098 29116 43144
rect 29162 43098 29274 43144
rect 29072 42981 29274 43098
rect 29072 42935 29116 42981
rect 29162 42935 29274 42981
rect 29072 42817 29274 42935
rect 29072 42771 29116 42817
rect 29162 42771 29274 42817
rect 29072 42654 29274 42771
rect 29072 42608 29116 42654
rect 29162 42608 29274 42654
rect 29072 42483 29274 42608
rect 30373 42483 30444 43271
rect 31292 43155 31336 43275
rect 33336 43184 33671 43275
rect 33336 43155 33495 43184
rect 33476 43051 33495 43155
rect 31292 42931 31336 43051
rect 33336 42931 33495 43051
rect 33458 42827 33495 42931
rect 31292 42707 31336 42827
rect 33336 42762 33495 42827
rect 33541 43155 33671 43184
rect 34671 43155 34715 43275
rect 39657 43155 39727 43275
rect 40167 43155 40346 43275
rect 44451 43264 44799 43275
rect 33541 43051 33560 43155
rect 40262 43137 40346 43155
rect 43354 43209 43695 43264
rect 43354 43163 43373 43209
rect 43513 43163 43695 43209
rect 43354 43144 43695 43163
rect 44325 43155 44799 43264
rect 45323 43155 45393 43275
rect 44325 43144 44552 43155
rect 40262 43091 40281 43137
rect 40327 43091 40346 43137
rect 40262 43072 40346 43091
rect 33541 42931 33671 43051
rect 34671 42931 34715 43051
rect 50410 43155 50454 43275
rect 51454 43155 51789 43275
rect 53789 43155 53833 43275
rect 54679 43383 54750 44171
rect 55849 44044 56051 44171
rect 55849 43998 55961 44044
rect 56007 43998 56051 44044
rect 55849 43881 56051 43998
rect 55849 43835 55961 43881
rect 56007 43835 56051 43881
rect 55849 43717 56051 43835
rect 55849 43671 55961 43717
rect 56007 43671 56051 43717
rect 55849 43554 56051 43671
rect 55849 43508 55961 43554
rect 56007 43508 56051 43554
rect 55849 43383 56051 43508
rect 33541 42762 33560 42931
rect 35133 42844 35260 42964
rect 36360 42865 36540 42964
rect 36360 42844 36475 42865
rect 35133 42795 35192 42844
rect 33336 42707 33560 42762
rect 33620 42675 33671 42795
rect 34671 42740 35192 42795
rect 36431 42740 36475 42844
rect 34671 42675 35260 42740
rect 35133 42620 35260 42675
rect 36360 42725 36475 42740
rect 36521 42725 36540 42865
rect 36360 42620 36540 42725
rect 36678 42865 36841 42964
rect 36678 42725 36697 42865
rect 36743 42844 36841 42865
rect 37501 42844 37572 42964
rect 37826 42844 37896 42964
rect 38556 42867 38734 42964
rect 43625 42931 43695 43051
rect 44325 43014 44799 43051
rect 44325 42968 44358 43014
rect 44498 42968 44799 43014
rect 44325 42931 44799 42968
rect 45323 42931 45367 43051
rect 51556 43154 51665 43155
rect 51556 43051 51600 43154
rect 38556 42844 38669 42867
rect 36743 42740 36773 42844
rect 38627 42740 38669 42844
rect 36743 42725 36841 42740
rect 36678 42620 36841 42725
rect 37501 42620 37572 42740
rect 37826 42620 37896 42740
rect 38556 42727 38669 42740
rect 38715 42727 38734 42867
rect 48603 42892 48765 42964
rect 38556 42620 38734 42727
rect 38939 42620 39008 42740
rect 39326 42620 39598 42740
rect 39730 42706 39909 42740
rect 43625 42707 43695 42827
rect 44325 42707 44799 42827
rect 45323 42783 45623 42827
rect 45323 42737 45464 42783
rect 45604 42737 45623 42783
rect 45323 42707 45623 42737
rect 48603 42752 48622 42892
rect 48668 42844 48765 42892
rect 49865 42844 49991 42964
rect 50410 42931 50454 43051
rect 51454 42931 51600 43051
rect 48668 42752 48705 42844
rect 48603 42740 48705 42752
rect 49932 42795 49991 42844
rect 49932 42740 50454 42795
rect 39730 42660 39844 42706
rect 39890 42660 39909 42706
rect 39730 42620 39909 42660
rect 48603 42620 48765 42740
rect 49865 42675 50454 42740
rect 51454 42675 51498 42795
rect 51581 42732 51600 42931
rect 51646 43051 51665 43154
rect 51646 42931 51789 43051
rect 53789 42931 53833 43051
rect 51646 42827 51667 42931
rect 51646 42732 51789 42827
rect 51581 42707 51789 42732
rect 53789 42707 53833 42827
rect 49865 42620 49991 42675
rect 29072 42244 29274 42371
rect 29072 42198 29116 42244
rect 29162 42198 29274 42244
rect 29072 42081 29274 42198
rect 29072 42035 29116 42081
rect 29162 42035 29274 42081
rect 29072 41917 29274 42035
rect 29072 41871 29116 41917
rect 29162 41871 29274 41917
rect 29072 41754 29274 41871
rect 29072 41708 29116 41754
rect 29162 41708 29274 41754
rect 29072 41583 29274 41708
rect 30373 41583 30444 42371
rect 54679 42483 54750 43271
rect 55849 43144 56051 43271
rect 55849 43098 55961 43144
rect 56007 43098 56051 43144
rect 55849 42981 56051 43098
rect 55849 42935 55961 42981
rect 56007 42935 56051 42981
rect 55849 42817 56051 42935
rect 55849 42771 55961 42817
rect 56007 42771 56051 42817
rect 55849 42654 56051 42771
rect 55849 42608 55961 42654
rect 56007 42608 56051 42654
rect 55849 42483 56051 42608
rect 35133 42179 35260 42234
rect 31292 42027 31336 42147
rect 33336 42092 33560 42147
rect 33336 42027 33495 42092
rect 33458 41923 33495 42027
rect 31292 41803 31336 41923
rect 33336 41803 33495 41923
rect 33476 41699 33495 41803
rect 29072 41344 29274 41471
rect 29072 41298 29116 41344
rect 29162 41298 29274 41344
rect 29072 41181 29274 41298
rect 29072 41135 29116 41181
rect 29162 41135 29274 41181
rect 29072 41017 29274 41135
rect 29072 40971 29116 41017
rect 29162 40971 29274 41017
rect 29072 40854 29274 40971
rect 29072 40808 29116 40854
rect 29162 40808 29274 40854
rect 29072 40683 29274 40808
rect 30373 40683 30444 41471
rect 31292 41579 31336 41699
rect 33336 41670 33495 41699
rect 33541 41923 33560 42092
rect 33620 42059 33671 42179
rect 34671 42114 35260 42179
rect 36360 42129 36540 42234
rect 36360 42114 36475 42129
rect 34671 42059 35192 42114
rect 35133 42010 35192 42059
rect 36431 42010 36475 42114
rect 33541 41803 33671 41923
rect 34671 41803 34715 41923
rect 35133 41890 35260 42010
rect 36360 41989 36475 42010
rect 36521 41989 36540 42129
rect 36360 41890 36540 41989
rect 36678 42129 36841 42234
rect 36678 41989 36697 42129
rect 36743 42114 36841 42129
rect 37501 42114 37572 42234
rect 37826 42114 37896 42234
rect 38556 42127 38734 42234
rect 38556 42114 38669 42127
rect 36743 42010 36773 42114
rect 38627 42010 38669 42114
rect 36743 41989 36841 42010
rect 36678 41890 36841 41989
rect 37501 41890 37572 42010
rect 37826 41890 37896 42010
rect 38556 41987 38669 42010
rect 38715 41987 38734 42127
rect 38939 42114 39008 42234
rect 39326 42114 39598 42234
rect 39730 42194 39909 42234
rect 39730 42148 39844 42194
rect 39890 42148 39909 42194
rect 39730 42114 39909 42148
rect 43625 42027 43695 42147
rect 44325 42027 44799 42147
rect 45323 42117 45623 42147
rect 45323 42071 45464 42117
rect 45604 42071 45623 42117
rect 45323 42027 45623 42071
rect 48603 42114 48765 42234
rect 49865 42179 49991 42234
rect 49865 42114 50454 42179
rect 48603 42102 48705 42114
rect 38556 41890 38734 41987
rect 48603 41962 48622 42102
rect 48668 42010 48705 42102
rect 49932 42059 50454 42114
rect 51454 42059 51498 42179
rect 51581 42122 51789 42147
rect 49932 42010 49991 42059
rect 48668 41962 48765 42010
rect 33541 41699 33560 41803
rect 43625 41803 43695 41923
rect 44325 41886 44799 41923
rect 44325 41840 44358 41886
rect 44498 41840 44799 41886
rect 44325 41803 44799 41840
rect 45323 41803 45367 41923
rect 48603 41890 48765 41962
rect 49865 41890 49991 42010
rect 51581 41923 51600 42122
rect 40262 41763 40346 41782
rect 40262 41717 40281 41763
rect 40327 41717 40346 41763
rect 40262 41699 40346 41717
rect 50410 41803 50454 41923
rect 51454 41803 51600 41923
rect 33541 41670 33671 41699
rect 33336 41579 33671 41670
rect 34671 41579 34715 41699
rect 31292 41355 31336 41475
rect 33336 41384 33671 41475
rect 33336 41355 33495 41384
rect 33476 41251 33495 41355
rect 31292 41131 31336 41251
rect 33336 41131 33495 41251
rect 33458 41027 33495 41131
rect 31292 40907 31336 41027
rect 33336 40962 33495 41027
rect 33541 41355 33671 41384
rect 34671 41355 34715 41475
rect 39657 41579 39727 41699
rect 40167 41579 40346 41699
rect 43354 41691 43695 41710
rect 43354 41645 43373 41691
rect 43513 41645 43695 41691
rect 43354 41590 43695 41645
rect 44325 41699 44552 41710
rect 44325 41590 44799 41699
rect 39657 41355 39727 41475
rect 40167 41355 40346 41475
rect 44451 41579 44799 41590
rect 45323 41579 45393 41699
rect 51556 41700 51600 41803
rect 51646 42027 51789 42122
rect 53789 42027 53833 42147
rect 51646 41923 51667 42027
rect 51646 41803 51789 41923
rect 53789 41803 53833 41923
rect 51646 41700 51665 41803
rect 51556 41699 51665 41700
rect 50410 41579 50454 41699
rect 51454 41579 51789 41699
rect 53789 41579 53833 41699
rect 44451 41464 44799 41475
rect 33541 41251 33560 41355
rect 40262 41337 40346 41355
rect 43354 41409 43695 41464
rect 43354 41363 43373 41409
rect 43513 41363 43695 41409
rect 43354 41344 43695 41363
rect 44325 41355 44799 41464
rect 45323 41355 45393 41475
rect 44325 41344 44552 41355
rect 40262 41291 40281 41337
rect 40327 41291 40346 41337
rect 40262 41272 40346 41291
rect 33541 41131 33671 41251
rect 34671 41131 34715 41251
rect 50410 41355 50454 41475
rect 51454 41355 51789 41475
rect 53789 41355 53833 41475
rect 54679 41583 54750 42371
rect 55849 42244 56051 42371
rect 55849 42198 55961 42244
rect 56007 42198 56051 42244
rect 55849 42081 56051 42198
rect 55849 42035 55961 42081
rect 56007 42035 56051 42081
rect 55849 41917 56051 42035
rect 55849 41871 55961 41917
rect 56007 41871 56051 41917
rect 55849 41754 56051 41871
rect 55849 41708 55961 41754
rect 56007 41708 56051 41754
rect 55849 41583 56051 41708
rect 33541 40962 33560 41131
rect 35133 41044 35260 41164
rect 36360 41065 36540 41164
rect 36360 41044 36475 41065
rect 35133 40995 35192 41044
rect 33336 40907 33560 40962
rect 33620 40875 33671 40995
rect 34671 40940 35192 40995
rect 36431 40940 36475 41044
rect 34671 40875 35260 40940
rect 35133 40820 35260 40875
rect 36360 40925 36475 40940
rect 36521 40925 36540 41065
rect 36360 40820 36540 40925
rect 36678 41065 36841 41164
rect 36678 40925 36697 41065
rect 36743 41044 36841 41065
rect 37501 41044 37572 41164
rect 37826 41044 37896 41164
rect 38556 41067 38734 41164
rect 43625 41131 43695 41251
rect 44325 41214 44799 41251
rect 44325 41168 44358 41214
rect 44498 41168 44799 41214
rect 44325 41131 44799 41168
rect 45323 41131 45367 41251
rect 51556 41354 51665 41355
rect 51556 41251 51600 41354
rect 38556 41044 38669 41067
rect 36743 40940 36773 41044
rect 38627 40940 38669 41044
rect 36743 40925 36841 40940
rect 36678 40820 36841 40925
rect 37501 40820 37572 40940
rect 37826 40820 37896 40940
rect 38556 40927 38669 40940
rect 38715 40927 38734 41067
rect 48603 41092 48765 41164
rect 38556 40820 38734 40927
rect 38939 40820 39008 40940
rect 39326 40820 39598 40940
rect 39730 40906 39909 40940
rect 43625 40907 43695 41027
rect 44325 40907 44799 41027
rect 45323 40983 45623 41027
rect 45323 40937 45464 40983
rect 45604 40937 45623 40983
rect 45323 40907 45623 40937
rect 48603 40952 48622 41092
rect 48668 41044 48765 41092
rect 49865 41044 49991 41164
rect 50410 41131 50454 41251
rect 51454 41131 51600 41251
rect 48668 40952 48705 41044
rect 48603 40940 48705 40952
rect 49932 40995 49991 41044
rect 49932 40940 50454 40995
rect 39730 40860 39844 40906
rect 39890 40860 39909 40906
rect 39730 40820 39909 40860
rect 48603 40820 48765 40940
rect 49865 40875 50454 40940
rect 51454 40875 51498 40995
rect 51581 40932 51600 41131
rect 51646 41251 51665 41354
rect 51646 41131 51789 41251
rect 53789 41131 53833 41251
rect 51646 41027 51667 41131
rect 51646 40932 51789 41027
rect 51581 40907 51789 40932
rect 53789 40907 53833 41027
rect 49865 40820 49991 40875
rect 29072 40444 29274 40571
rect 29072 40398 29116 40444
rect 29162 40398 29274 40444
rect 29072 40281 29274 40398
rect 29072 40235 29116 40281
rect 29162 40235 29274 40281
rect 29072 40117 29274 40235
rect 29072 40071 29116 40117
rect 29162 40071 29274 40117
rect 29072 39954 29274 40071
rect 29072 39908 29116 39954
rect 29162 39908 29274 39954
rect 29072 39783 29274 39908
rect 30373 39783 30444 40571
rect 54679 40683 54750 41471
rect 55849 41344 56051 41471
rect 55849 41298 55961 41344
rect 56007 41298 56051 41344
rect 55849 41181 56051 41298
rect 55849 41135 55961 41181
rect 56007 41135 56051 41181
rect 55849 41017 56051 41135
rect 55849 40971 55961 41017
rect 56007 40971 56051 41017
rect 55849 40854 56051 40971
rect 55849 40808 55961 40854
rect 56007 40808 56051 40854
rect 55849 40683 56051 40808
rect 35133 40379 35260 40434
rect 31292 40227 31336 40347
rect 33336 40292 33560 40347
rect 33336 40227 33495 40292
rect 33458 40123 33495 40227
rect 31292 40003 31336 40123
rect 33336 40003 33495 40123
rect 33476 39899 33495 40003
rect 29072 39544 29274 39671
rect 29072 39498 29116 39544
rect 29162 39498 29274 39544
rect 29072 39381 29274 39498
rect 29072 39335 29116 39381
rect 29162 39335 29274 39381
rect 29072 39217 29274 39335
rect 29072 39171 29116 39217
rect 29162 39171 29274 39217
rect 29072 39054 29274 39171
rect 29072 39008 29116 39054
rect 29162 39008 29274 39054
rect 29072 38883 29274 39008
rect 30373 38883 30444 39671
rect 31292 39779 31336 39899
rect 33336 39870 33495 39899
rect 33541 40123 33560 40292
rect 33620 40259 33671 40379
rect 34671 40314 35260 40379
rect 36360 40329 36540 40434
rect 36360 40314 36475 40329
rect 34671 40259 35192 40314
rect 35133 40210 35192 40259
rect 36431 40210 36475 40314
rect 33541 40003 33671 40123
rect 34671 40003 34715 40123
rect 35133 40090 35260 40210
rect 36360 40189 36475 40210
rect 36521 40189 36540 40329
rect 36360 40090 36540 40189
rect 36678 40329 36841 40434
rect 36678 40189 36697 40329
rect 36743 40314 36841 40329
rect 37501 40314 37572 40434
rect 37826 40314 37896 40434
rect 38556 40327 38734 40434
rect 38556 40314 38669 40327
rect 36743 40210 36773 40314
rect 38627 40210 38669 40314
rect 36743 40189 36841 40210
rect 36678 40090 36841 40189
rect 37501 40090 37572 40210
rect 37826 40090 37896 40210
rect 38556 40187 38669 40210
rect 38715 40187 38734 40327
rect 38939 40314 39008 40434
rect 39326 40314 39598 40434
rect 39730 40394 39909 40434
rect 39730 40348 39844 40394
rect 39890 40348 39909 40394
rect 39730 40314 39909 40348
rect 43625 40227 43695 40347
rect 44325 40227 44799 40347
rect 45323 40317 45623 40347
rect 45323 40271 45464 40317
rect 45604 40271 45623 40317
rect 45323 40227 45623 40271
rect 48603 40314 48765 40434
rect 49865 40379 49991 40434
rect 49865 40314 50454 40379
rect 48603 40302 48705 40314
rect 38556 40090 38734 40187
rect 48603 40162 48622 40302
rect 48668 40210 48705 40302
rect 49932 40259 50454 40314
rect 51454 40259 51498 40379
rect 51581 40322 51789 40347
rect 49932 40210 49991 40259
rect 48668 40162 48765 40210
rect 33541 39899 33560 40003
rect 43625 40003 43695 40123
rect 44325 40086 44799 40123
rect 44325 40040 44358 40086
rect 44498 40040 44799 40086
rect 44325 40003 44799 40040
rect 45323 40003 45367 40123
rect 48603 40090 48765 40162
rect 49865 40090 49991 40210
rect 51581 40123 51600 40322
rect 40262 39963 40346 39982
rect 40262 39917 40281 39963
rect 40327 39917 40346 39963
rect 40262 39899 40346 39917
rect 50410 40003 50454 40123
rect 51454 40003 51600 40123
rect 33541 39870 33671 39899
rect 33336 39779 33671 39870
rect 34671 39779 34715 39899
rect 31292 39555 31336 39675
rect 33336 39584 33671 39675
rect 33336 39555 33495 39584
rect 33476 39451 33495 39555
rect 31292 39331 31336 39451
rect 33336 39331 33495 39451
rect 33458 39227 33495 39331
rect 31292 39107 31336 39227
rect 33336 39162 33495 39227
rect 33541 39555 33671 39584
rect 34671 39555 34715 39675
rect 39657 39779 39727 39899
rect 40167 39779 40346 39899
rect 43354 39891 43695 39910
rect 43354 39845 43373 39891
rect 43513 39845 43695 39891
rect 43354 39790 43695 39845
rect 44325 39899 44552 39910
rect 44325 39790 44799 39899
rect 39657 39555 39727 39675
rect 40167 39555 40346 39675
rect 44451 39779 44799 39790
rect 45323 39779 45393 39899
rect 51556 39900 51600 40003
rect 51646 40227 51789 40322
rect 53789 40227 53833 40347
rect 51646 40123 51667 40227
rect 51646 40003 51789 40123
rect 53789 40003 53833 40123
rect 51646 39900 51665 40003
rect 51556 39899 51665 39900
rect 50410 39779 50454 39899
rect 51454 39779 51789 39899
rect 53789 39779 53833 39899
rect 44451 39664 44799 39675
rect 33541 39451 33560 39555
rect 40262 39537 40346 39555
rect 43354 39609 43695 39664
rect 43354 39563 43373 39609
rect 43513 39563 43695 39609
rect 43354 39544 43695 39563
rect 44325 39555 44799 39664
rect 45323 39555 45393 39675
rect 44325 39544 44552 39555
rect 40262 39491 40281 39537
rect 40327 39491 40346 39537
rect 40262 39472 40346 39491
rect 33541 39331 33671 39451
rect 34671 39331 34715 39451
rect 50410 39555 50454 39675
rect 51454 39555 51789 39675
rect 53789 39555 53833 39675
rect 54679 39783 54750 40571
rect 55849 40444 56051 40571
rect 55849 40398 55961 40444
rect 56007 40398 56051 40444
rect 55849 40281 56051 40398
rect 55849 40235 55961 40281
rect 56007 40235 56051 40281
rect 55849 40117 56051 40235
rect 55849 40071 55961 40117
rect 56007 40071 56051 40117
rect 55849 39954 56051 40071
rect 55849 39908 55961 39954
rect 56007 39908 56051 39954
rect 55849 39783 56051 39908
rect 33541 39162 33560 39331
rect 35133 39244 35260 39364
rect 36360 39265 36540 39364
rect 36360 39244 36475 39265
rect 35133 39195 35192 39244
rect 33336 39107 33560 39162
rect 33620 39075 33671 39195
rect 34671 39140 35192 39195
rect 36431 39140 36475 39244
rect 34671 39075 35260 39140
rect 35133 39020 35260 39075
rect 36360 39125 36475 39140
rect 36521 39125 36540 39265
rect 36360 39020 36540 39125
rect 36678 39265 36841 39364
rect 36678 39125 36697 39265
rect 36743 39244 36841 39265
rect 37501 39244 37572 39364
rect 37826 39244 37896 39364
rect 38556 39267 38734 39364
rect 43625 39331 43695 39451
rect 44325 39414 44799 39451
rect 44325 39368 44358 39414
rect 44498 39368 44799 39414
rect 44325 39331 44799 39368
rect 45323 39331 45367 39451
rect 51556 39554 51665 39555
rect 51556 39451 51600 39554
rect 38556 39244 38669 39267
rect 36743 39140 36773 39244
rect 38627 39140 38669 39244
rect 36743 39125 36841 39140
rect 36678 39020 36841 39125
rect 37501 39020 37572 39140
rect 37826 39020 37896 39140
rect 38556 39127 38669 39140
rect 38715 39127 38734 39267
rect 48603 39292 48765 39364
rect 38556 39020 38734 39127
rect 38939 39020 39008 39140
rect 39326 39020 39598 39140
rect 39730 39106 39909 39140
rect 43625 39107 43695 39227
rect 44325 39107 44799 39227
rect 45323 39183 45623 39227
rect 45323 39137 45464 39183
rect 45604 39137 45623 39183
rect 45323 39107 45623 39137
rect 48603 39152 48622 39292
rect 48668 39244 48765 39292
rect 49865 39244 49991 39364
rect 50410 39331 50454 39451
rect 51454 39331 51600 39451
rect 48668 39152 48705 39244
rect 48603 39140 48705 39152
rect 49932 39195 49991 39244
rect 49932 39140 50454 39195
rect 39730 39060 39844 39106
rect 39890 39060 39909 39106
rect 39730 39020 39909 39060
rect 48603 39020 48765 39140
rect 49865 39075 50454 39140
rect 51454 39075 51498 39195
rect 51581 39132 51600 39331
rect 51646 39451 51665 39554
rect 51646 39331 51789 39451
rect 53789 39331 53833 39451
rect 51646 39227 51667 39331
rect 51646 39132 51789 39227
rect 51581 39107 51789 39132
rect 53789 39107 53833 39227
rect 49865 39020 49991 39075
rect 29072 38644 29274 38771
rect 29072 38598 29116 38644
rect 29162 38598 29274 38644
rect 29072 38481 29274 38598
rect 29072 38435 29116 38481
rect 29162 38435 29274 38481
rect 29072 38317 29274 38435
rect 29072 38271 29116 38317
rect 29162 38271 29274 38317
rect 29072 38154 29274 38271
rect 29072 38108 29116 38154
rect 29162 38108 29274 38154
rect 29072 37983 29274 38108
rect 30373 37983 30444 38771
rect 54679 38883 54750 39671
rect 55849 39544 56051 39671
rect 55849 39498 55961 39544
rect 56007 39498 56051 39544
rect 55849 39381 56051 39498
rect 55849 39335 55961 39381
rect 56007 39335 56051 39381
rect 55849 39217 56051 39335
rect 55849 39171 55961 39217
rect 56007 39171 56051 39217
rect 55849 39054 56051 39171
rect 55849 39008 55961 39054
rect 56007 39008 56051 39054
rect 55849 38883 56051 39008
rect 35133 38579 35260 38634
rect 31292 38427 31336 38547
rect 33336 38492 33560 38547
rect 33336 38427 33495 38492
rect 33458 38323 33495 38427
rect 31292 38203 31336 38323
rect 33336 38203 33495 38323
rect 33476 38099 33495 38203
rect 29072 37744 29274 37871
rect 29072 37698 29116 37744
rect 29162 37698 29274 37744
rect 29072 37581 29274 37698
rect 29072 37535 29116 37581
rect 29162 37535 29274 37581
rect 29072 37417 29274 37535
rect 29072 37371 29116 37417
rect 29162 37371 29274 37417
rect 29072 37254 29274 37371
rect 29072 37208 29116 37254
rect 29162 37208 29274 37254
rect 29072 37083 29274 37208
rect 30373 37083 30444 37871
rect 31292 37979 31336 38099
rect 33336 38070 33495 38099
rect 33541 38323 33560 38492
rect 33620 38459 33671 38579
rect 34671 38514 35260 38579
rect 36360 38529 36540 38634
rect 36360 38514 36475 38529
rect 34671 38459 35192 38514
rect 35133 38410 35192 38459
rect 36431 38410 36475 38514
rect 33541 38203 33671 38323
rect 34671 38203 34715 38323
rect 35133 38290 35260 38410
rect 36360 38389 36475 38410
rect 36521 38389 36540 38529
rect 36360 38290 36540 38389
rect 36678 38529 36841 38634
rect 36678 38389 36697 38529
rect 36743 38514 36841 38529
rect 37501 38514 37572 38634
rect 37826 38514 37896 38634
rect 38556 38527 38734 38634
rect 38556 38514 38669 38527
rect 36743 38410 36773 38514
rect 38627 38410 38669 38514
rect 36743 38389 36841 38410
rect 36678 38290 36841 38389
rect 37501 38290 37572 38410
rect 37826 38290 37896 38410
rect 38556 38387 38669 38410
rect 38715 38387 38734 38527
rect 38939 38514 39008 38634
rect 39326 38514 39598 38634
rect 39730 38594 39909 38634
rect 39730 38548 39844 38594
rect 39890 38548 39909 38594
rect 39730 38514 39909 38548
rect 43625 38427 43695 38547
rect 44325 38427 44799 38547
rect 45323 38517 45623 38547
rect 45323 38471 45464 38517
rect 45604 38471 45623 38517
rect 45323 38427 45623 38471
rect 48603 38514 48765 38634
rect 49865 38579 49991 38634
rect 49865 38514 50454 38579
rect 48603 38502 48705 38514
rect 38556 38290 38734 38387
rect 48603 38362 48622 38502
rect 48668 38410 48705 38502
rect 49932 38459 50454 38514
rect 51454 38459 51498 38579
rect 51581 38522 51789 38547
rect 49932 38410 49991 38459
rect 48668 38362 48765 38410
rect 33541 38099 33560 38203
rect 43625 38203 43695 38323
rect 44325 38286 44799 38323
rect 44325 38240 44358 38286
rect 44498 38240 44799 38286
rect 44325 38203 44799 38240
rect 45323 38203 45367 38323
rect 48603 38290 48765 38362
rect 49865 38290 49991 38410
rect 51581 38323 51600 38522
rect 40262 38163 40346 38182
rect 40262 38117 40281 38163
rect 40327 38117 40346 38163
rect 40262 38099 40346 38117
rect 50410 38203 50454 38323
rect 51454 38203 51600 38323
rect 33541 38070 33671 38099
rect 33336 37979 33671 38070
rect 34671 37979 34715 38099
rect 31292 37755 31336 37875
rect 33336 37784 33671 37875
rect 33336 37755 33495 37784
rect 33476 37651 33495 37755
rect 31292 37531 31336 37651
rect 33336 37531 33495 37651
rect 33458 37427 33495 37531
rect 31292 37307 31336 37427
rect 33336 37362 33495 37427
rect 33541 37755 33671 37784
rect 34671 37755 34715 37875
rect 39657 37979 39727 38099
rect 40167 37979 40346 38099
rect 43354 38091 43695 38110
rect 43354 38045 43373 38091
rect 43513 38045 43695 38091
rect 43354 37990 43695 38045
rect 44325 38099 44552 38110
rect 44325 37990 44799 38099
rect 39657 37755 39727 37875
rect 40167 37755 40346 37875
rect 44451 37979 44799 37990
rect 45323 37979 45393 38099
rect 51556 38100 51600 38203
rect 51646 38427 51789 38522
rect 53789 38427 53833 38547
rect 51646 38323 51667 38427
rect 51646 38203 51789 38323
rect 53789 38203 53833 38323
rect 51646 38100 51665 38203
rect 51556 38099 51665 38100
rect 50410 37979 50454 38099
rect 51454 37979 51789 38099
rect 53789 37979 53833 38099
rect 44451 37864 44799 37875
rect 33541 37651 33560 37755
rect 40262 37737 40346 37755
rect 43354 37809 43695 37864
rect 43354 37763 43373 37809
rect 43513 37763 43695 37809
rect 43354 37744 43695 37763
rect 44325 37755 44799 37864
rect 45323 37755 45393 37875
rect 44325 37744 44552 37755
rect 40262 37691 40281 37737
rect 40327 37691 40346 37737
rect 40262 37672 40346 37691
rect 33541 37531 33671 37651
rect 34671 37531 34715 37651
rect 50410 37755 50454 37875
rect 51454 37755 51789 37875
rect 53789 37755 53833 37875
rect 54679 37983 54750 38771
rect 55849 38644 56051 38771
rect 55849 38598 55961 38644
rect 56007 38598 56051 38644
rect 55849 38481 56051 38598
rect 55849 38435 55961 38481
rect 56007 38435 56051 38481
rect 55849 38317 56051 38435
rect 55849 38271 55961 38317
rect 56007 38271 56051 38317
rect 55849 38154 56051 38271
rect 55849 38108 55961 38154
rect 56007 38108 56051 38154
rect 55849 37983 56051 38108
rect 33541 37362 33560 37531
rect 35133 37444 35260 37564
rect 36360 37465 36540 37564
rect 36360 37444 36475 37465
rect 35133 37395 35192 37444
rect 33336 37307 33560 37362
rect 33620 37275 33671 37395
rect 34671 37340 35192 37395
rect 36431 37340 36475 37444
rect 34671 37275 35260 37340
rect 35133 37220 35260 37275
rect 36360 37325 36475 37340
rect 36521 37325 36540 37465
rect 36360 37220 36540 37325
rect 36678 37465 36841 37564
rect 36678 37325 36697 37465
rect 36743 37444 36841 37465
rect 37501 37444 37572 37564
rect 37826 37444 37896 37564
rect 38556 37467 38734 37564
rect 43625 37531 43695 37651
rect 44325 37614 44799 37651
rect 44325 37568 44358 37614
rect 44498 37568 44799 37614
rect 44325 37531 44799 37568
rect 45323 37531 45367 37651
rect 51556 37754 51665 37755
rect 51556 37651 51600 37754
rect 38556 37444 38669 37467
rect 36743 37340 36773 37444
rect 38627 37340 38669 37444
rect 36743 37325 36841 37340
rect 36678 37220 36841 37325
rect 37501 37220 37572 37340
rect 37826 37220 37896 37340
rect 38556 37327 38669 37340
rect 38715 37327 38734 37467
rect 48603 37492 48765 37564
rect 38556 37220 38734 37327
rect 38939 37220 39008 37340
rect 39326 37220 39598 37340
rect 39730 37306 39909 37340
rect 43625 37307 43695 37427
rect 44325 37307 44799 37427
rect 45323 37383 45623 37427
rect 45323 37337 45464 37383
rect 45604 37337 45623 37383
rect 45323 37307 45623 37337
rect 48603 37352 48622 37492
rect 48668 37444 48765 37492
rect 49865 37444 49991 37564
rect 50410 37531 50454 37651
rect 51454 37531 51600 37651
rect 48668 37352 48705 37444
rect 48603 37340 48705 37352
rect 49932 37395 49991 37444
rect 49932 37340 50454 37395
rect 39730 37260 39844 37306
rect 39890 37260 39909 37306
rect 39730 37220 39909 37260
rect 48603 37220 48765 37340
rect 49865 37275 50454 37340
rect 51454 37275 51498 37395
rect 51581 37332 51600 37531
rect 51646 37651 51665 37754
rect 51646 37531 51789 37651
rect 53789 37531 53833 37651
rect 51646 37427 51667 37531
rect 51646 37332 51789 37427
rect 51581 37307 51789 37332
rect 53789 37307 53833 37427
rect 49865 37220 49991 37275
rect 29072 36844 29274 36971
rect 29072 36798 29116 36844
rect 29162 36798 29274 36844
rect 29072 36681 29274 36798
rect 29072 36635 29116 36681
rect 29162 36635 29274 36681
rect 29072 36517 29274 36635
rect 29072 36471 29116 36517
rect 29162 36471 29274 36517
rect 29072 36354 29274 36471
rect 29072 36308 29116 36354
rect 29162 36308 29274 36354
rect 29072 36183 29274 36308
rect 30373 36183 30444 36971
rect 54679 37083 54750 37871
rect 55849 37744 56051 37871
rect 55849 37698 55961 37744
rect 56007 37698 56051 37744
rect 55849 37581 56051 37698
rect 55849 37535 55961 37581
rect 56007 37535 56051 37581
rect 55849 37417 56051 37535
rect 55849 37371 55961 37417
rect 56007 37371 56051 37417
rect 55849 37254 56051 37371
rect 55849 37208 55961 37254
rect 56007 37208 56051 37254
rect 55849 37083 56051 37208
rect 35133 36779 35260 36834
rect 31292 36627 31336 36747
rect 33336 36692 33560 36747
rect 33336 36627 33495 36692
rect 33458 36523 33495 36627
rect 31292 36403 31336 36523
rect 33336 36403 33495 36523
rect 33476 36299 33495 36403
rect 31292 36179 31336 36299
rect 33336 36270 33495 36299
rect 33541 36523 33560 36692
rect 33620 36659 33671 36779
rect 34671 36714 35260 36779
rect 36360 36729 36540 36834
rect 36360 36714 36475 36729
rect 34671 36659 35192 36714
rect 35133 36610 35192 36659
rect 36431 36610 36475 36714
rect 33541 36403 33671 36523
rect 34671 36403 34715 36523
rect 35133 36490 35260 36610
rect 36360 36589 36475 36610
rect 36521 36589 36540 36729
rect 36360 36490 36540 36589
rect 36678 36729 36841 36834
rect 36678 36589 36697 36729
rect 36743 36714 36841 36729
rect 37501 36714 37572 36834
rect 37826 36714 37896 36834
rect 38556 36727 38734 36834
rect 38556 36714 38669 36727
rect 36743 36610 36773 36714
rect 38627 36610 38669 36714
rect 36743 36589 36841 36610
rect 36678 36490 36841 36589
rect 37501 36490 37572 36610
rect 37826 36490 37896 36610
rect 38556 36587 38669 36610
rect 38715 36587 38734 36727
rect 38939 36714 39008 36834
rect 39326 36714 39598 36834
rect 39730 36794 39909 36834
rect 39730 36748 39844 36794
rect 39890 36748 39909 36794
rect 39730 36714 39909 36748
rect 43625 36627 43695 36747
rect 44325 36627 44799 36747
rect 45323 36717 45623 36747
rect 45323 36671 45464 36717
rect 45604 36671 45623 36717
rect 45323 36627 45623 36671
rect 48603 36714 48765 36834
rect 49865 36779 49991 36834
rect 49865 36714 50454 36779
rect 48603 36702 48705 36714
rect 38556 36490 38734 36587
rect 48603 36562 48622 36702
rect 48668 36610 48705 36702
rect 49932 36659 50454 36714
rect 51454 36659 51498 36779
rect 51581 36722 51789 36747
rect 49932 36610 49991 36659
rect 48668 36562 48765 36610
rect 33541 36299 33560 36403
rect 43625 36403 43695 36523
rect 44325 36486 44799 36523
rect 44325 36440 44358 36486
rect 44498 36440 44799 36486
rect 44325 36403 44799 36440
rect 45323 36403 45367 36523
rect 48603 36490 48765 36562
rect 49865 36490 49991 36610
rect 51581 36523 51600 36722
rect 40262 36363 40346 36382
rect 40262 36317 40281 36363
rect 40327 36317 40346 36363
rect 40262 36299 40346 36317
rect 50410 36403 50454 36523
rect 51454 36403 51600 36523
rect 33541 36270 33671 36299
rect 33336 36179 33671 36270
rect 34671 36179 34715 36299
rect 39657 36179 39727 36299
rect 40167 36179 40346 36299
rect 43354 36291 43695 36310
rect 43354 36245 43373 36291
rect 43513 36245 43695 36291
rect 43354 36190 43695 36245
rect 44325 36299 44552 36310
rect 44325 36190 44799 36299
rect 44451 36179 44799 36190
rect 45323 36179 45393 36299
rect 51556 36300 51600 36403
rect 51646 36627 51789 36722
rect 53789 36627 53833 36747
rect 51646 36523 51667 36627
rect 51646 36403 51789 36523
rect 53789 36403 53833 36523
rect 51646 36300 51665 36403
rect 51556 36299 51665 36300
rect 50410 36179 50454 36299
rect 51454 36179 51789 36299
rect 53789 36179 53833 36299
rect 54679 36183 54750 36971
rect 55849 36844 56051 36971
rect 55849 36798 55961 36844
rect 56007 36798 56051 36844
rect 55849 36681 56051 36798
rect 55849 36635 55961 36681
rect 56007 36635 56051 36681
rect 55849 36517 56051 36635
rect 55849 36471 55961 36517
rect 56007 36471 56051 36517
rect 55849 36354 56051 36471
rect 55849 36308 55961 36354
rect 56007 36308 56051 36354
rect 55849 36183 56051 36308
<< polycontact >>
rect 29116 43998 29162 44044
rect 29116 43835 29162 43881
rect 29116 43671 29162 43717
rect 29116 43508 29162 43554
rect 42319 44197 42459 44243
rect 44067 44245 44113 44291
rect 38035 43905 38081 44045
rect 40694 43818 40740 43958
rect 44279 43858 44325 43998
rect 46967 43893 47013 44033
rect 29116 43098 29162 43144
rect 29116 42935 29162 42981
rect 29116 42771 29162 42817
rect 29116 42608 29162 42654
rect 33495 42762 33541 43184
rect 43373 43163 43513 43209
rect 40281 43091 40327 43137
rect 55961 43998 56007 44044
rect 55961 43835 56007 43881
rect 55961 43671 56007 43717
rect 55961 43508 56007 43554
rect 36475 42725 36521 42865
rect 36697 42725 36743 42865
rect 44358 42968 44498 43014
rect 38669 42727 38715 42867
rect 45464 42737 45604 42783
rect 48622 42752 48668 42892
rect 39844 42660 39890 42706
rect 51600 42732 51646 43154
rect 29116 42198 29162 42244
rect 29116 42035 29162 42081
rect 29116 41871 29162 41917
rect 29116 41708 29162 41754
rect 55961 43098 56007 43144
rect 55961 42935 56007 42981
rect 55961 42771 56007 42817
rect 55961 42608 56007 42654
rect 29116 41298 29162 41344
rect 29116 41135 29162 41181
rect 29116 40971 29162 41017
rect 29116 40808 29162 40854
rect 33495 41670 33541 42092
rect 36475 41989 36521 42129
rect 36697 41989 36743 42129
rect 38669 41987 38715 42127
rect 39844 42148 39890 42194
rect 45464 42071 45604 42117
rect 48622 41962 48668 42102
rect 44358 41840 44498 41886
rect 40281 41717 40327 41763
rect 33495 40962 33541 41384
rect 43373 41645 43513 41691
rect 51600 41700 51646 42122
rect 43373 41363 43513 41409
rect 40281 41291 40327 41337
rect 55961 42198 56007 42244
rect 55961 42035 56007 42081
rect 55961 41871 56007 41917
rect 55961 41708 56007 41754
rect 36475 40925 36521 41065
rect 36697 40925 36743 41065
rect 44358 41168 44498 41214
rect 38669 40927 38715 41067
rect 45464 40937 45604 40983
rect 48622 40952 48668 41092
rect 39844 40860 39890 40906
rect 51600 40932 51646 41354
rect 29116 40398 29162 40444
rect 29116 40235 29162 40281
rect 29116 40071 29162 40117
rect 29116 39908 29162 39954
rect 55961 41298 56007 41344
rect 55961 41135 56007 41181
rect 55961 40971 56007 41017
rect 55961 40808 56007 40854
rect 29116 39498 29162 39544
rect 29116 39335 29162 39381
rect 29116 39171 29162 39217
rect 29116 39008 29162 39054
rect 33495 39870 33541 40292
rect 36475 40189 36521 40329
rect 36697 40189 36743 40329
rect 38669 40187 38715 40327
rect 39844 40348 39890 40394
rect 45464 40271 45604 40317
rect 48622 40162 48668 40302
rect 44358 40040 44498 40086
rect 40281 39917 40327 39963
rect 33495 39162 33541 39584
rect 43373 39845 43513 39891
rect 51600 39900 51646 40322
rect 43373 39563 43513 39609
rect 40281 39491 40327 39537
rect 55961 40398 56007 40444
rect 55961 40235 56007 40281
rect 55961 40071 56007 40117
rect 55961 39908 56007 39954
rect 36475 39125 36521 39265
rect 36697 39125 36743 39265
rect 44358 39368 44498 39414
rect 38669 39127 38715 39267
rect 45464 39137 45604 39183
rect 48622 39152 48668 39292
rect 39844 39060 39890 39106
rect 51600 39132 51646 39554
rect 29116 38598 29162 38644
rect 29116 38435 29162 38481
rect 29116 38271 29162 38317
rect 29116 38108 29162 38154
rect 55961 39498 56007 39544
rect 55961 39335 56007 39381
rect 55961 39171 56007 39217
rect 55961 39008 56007 39054
rect 29116 37698 29162 37744
rect 29116 37535 29162 37581
rect 29116 37371 29162 37417
rect 29116 37208 29162 37254
rect 33495 38070 33541 38492
rect 36475 38389 36521 38529
rect 36697 38389 36743 38529
rect 38669 38387 38715 38527
rect 39844 38548 39890 38594
rect 45464 38471 45604 38517
rect 48622 38362 48668 38502
rect 44358 38240 44498 38286
rect 40281 38117 40327 38163
rect 33495 37362 33541 37784
rect 43373 38045 43513 38091
rect 51600 38100 51646 38522
rect 43373 37763 43513 37809
rect 40281 37691 40327 37737
rect 55961 38598 56007 38644
rect 55961 38435 56007 38481
rect 55961 38271 56007 38317
rect 55961 38108 56007 38154
rect 36475 37325 36521 37465
rect 36697 37325 36743 37465
rect 44358 37568 44498 37614
rect 38669 37327 38715 37467
rect 45464 37337 45604 37383
rect 48622 37352 48668 37492
rect 39844 37260 39890 37306
rect 51600 37332 51646 37754
rect 29116 36798 29162 36844
rect 29116 36635 29162 36681
rect 29116 36471 29162 36517
rect 29116 36308 29162 36354
rect 55961 37698 56007 37744
rect 55961 37535 56007 37581
rect 55961 37371 56007 37417
rect 55961 37208 56007 37254
rect 33495 36270 33541 36692
rect 36475 36589 36521 36729
rect 36697 36589 36743 36729
rect 38669 36587 38715 36727
rect 39844 36748 39890 36794
rect 45464 36671 45604 36717
rect 48622 36562 48668 36702
rect 44358 36440 44498 36486
rect 40281 36317 40327 36363
rect 43373 36245 43513 36291
rect 51600 36300 51646 36722
rect 55961 36798 56007 36844
rect 55961 36635 56007 36681
rect 55961 36471 56007 36517
rect 55961 36308 56007 36354
<< metal1 >>
rect 282 46083 86090 46294
rect 282 46037 371 46083
rect 417 46037 495 46083
rect 541 46037 619 46083
rect 665 46037 743 46083
rect 789 46037 867 46083
rect 913 46037 991 46083
rect 1037 46037 1115 46083
rect 1161 46037 1239 46083
rect 1285 46037 1363 46083
rect 1409 46037 1487 46083
rect 1533 46037 1611 46083
rect 1657 46037 1735 46083
rect 1781 46037 1859 46083
rect 1905 46037 1983 46083
rect 2029 46037 2107 46083
rect 2153 46037 2231 46083
rect 2277 46037 2355 46083
rect 2401 46037 2479 46083
rect 2525 46037 2603 46083
rect 2649 46037 2727 46083
rect 2773 46037 2851 46083
rect 2897 46037 2975 46083
rect 3021 46037 3099 46083
rect 3145 46037 3223 46083
rect 3269 46037 3347 46083
rect 3393 46037 3471 46083
rect 3517 46037 3595 46083
rect 3641 46037 3719 46083
rect 3765 46037 3843 46083
rect 3889 46037 3967 46083
rect 4013 46037 4091 46083
rect 4137 46037 4215 46083
rect 4261 46037 4339 46083
rect 4385 46037 4463 46083
rect 4509 46037 4587 46083
rect 4633 46037 4711 46083
rect 4757 46037 4835 46083
rect 4881 46037 4959 46083
rect 5005 46037 5083 46083
rect 5129 46037 5207 46083
rect 5253 46037 5331 46083
rect 5377 46037 5455 46083
rect 5501 46037 5579 46083
rect 5625 46037 5703 46083
rect 5749 46037 5827 46083
rect 5873 46037 5951 46083
rect 5997 46037 6075 46083
rect 6121 46037 6199 46083
rect 6245 46037 6323 46083
rect 6369 46037 6447 46083
rect 6493 46037 6571 46083
rect 6617 46037 6695 46083
rect 6741 46037 6819 46083
rect 6865 46037 6943 46083
rect 6989 46037 7067 46083
rect 7113 46037 7191 46083
rect 7237 46037 7315 46083
rect 7361 46037 7439 46083
rect 7485 46037 7563 46083
rect 7609 46037 7687 46083
rect 7733 46037 7811 46083
rect 7857 46037 7935 46083
rect 7981 46037 8059 46083
rect 8105 46037 8183 46083
rect 8229 46037 8307 46083
rect 8353 46037 8431 46083
rect 8477 46037 8555 46083
rect 8601 46037 8679 46083
rect 8725 46037 8803 46083
rect 8849 46037 8927 46083
rect 8973 46037 9051 46083
rect 9097 46037 9175 46083
rect 9221 46037 9299 46083
rect 9345 46037 9423 46083
rect 9469 46037 9547 46083
rect 9593 46037 9671 46083
rect 9717 46037 9795 46083
rect 9841 46037 9919 46083
rect 9965 46037 10043 46083
rect 10089 46037 10167 46083
rect 10213 46037 10291 46083
rect 10337 46037 10415 46083
rect 10461 46037 10539 46083
rect 10585 46037 10663 46083
rect 10709 46037 10787 46083
rect 10833 46037 10911 46083
rect 10957 46037 11035 46083
rect 11081 46037 11159 46083
rect 11205 46037 11283 46083
rect 11329 46037 11407 46083
rect 11453 46037 11531 46083
rect 11577 46037 11655 46083
rect 11701 46037 11779 46083
rect 11825 46037 11903 46083
rect 11949 46037 12027 46083
rect 12073 46037 12151 46083
rect 12197 46037 12275 46083
rect 12321 46037 12399 46083
rect 12445 46037 12523 46083
rect 12569 46037 12647 46083
rect 12693 46037 12771 46083
rect 12817 46037 12895 46083
rect 12941 46037 13019 46083
rect 13065 46037 13143 46083
rect 13189 46037 13267 46083
rect 13313 46037 13391 46083
rect 13437 46037 13515 46083
rect 13561 46037 13639 46083
rect 13685 46037 13763 46083
rect 13809 46037 13887 46083
rect 13933 46037 14011 46083
rect 14057 46037 14135 46083
rect 14181 46037 14259 46083
rect 14305 46037 14383 46083
rect 14429 46037 14507 46083
rect 14553 46037 14631 46083
rect 14677 46037 14755 46083
rect 14801 46037 14879 46083
rect 14925 46037 15003 46083
rect 15049 46037 15127 46083
rect 15173 46037 15251 46083
rect 15297 46037 15375 46083
rect 15421 46037 15499 46083
rect 15545 46037 15623 46083
rect 15669 46037 15747 46083
rect 15793 46037 15871 46083
rect 15917 46037 15995 46083
rect 16041 46037 16119 46083
rect 16165 46037 16243 46083
rect 16289 46037 16367 46083
rect 16413 46037 16491 46083
rect 16537 46037 16615 46083
rect 16661 46037 16739 46083
rect 16785 46037 16863 46083
rect 16909 46037 16987 46083
rect 17033 46037 17111 46083
rect 17157 46037 17235 46083
rect 17281 46037 17359 46083
rect 17405 46037 17483 46083
rect 17529 46037 17607 46083
rect 17653 46037 17731 46083
rect 17777 46037 17855 46083
rect 17901 46037 17979 46083
rect 18025 46037 18103 46083
rect 18149 46037 18227 46083
rect 18273 46037 18351 46083
rect 18397 46037 18475 46083
rect 18521 46037 18599 46083
rect 18645 46037 18723 46083
rect 18769 46037 18847 46083
rect 18893 46037 18971 46083
rect 19017 46037 19095 46083
rect 19141 46037 19219 46083
rect 19265 46037 19343 46083
rect 19389 46037 19467 46083
rect 19513 46037 19591 46083
rect 19637 46037 19715 46083
rect 19761 46037 19839 46083
rect 19885 46037 19963 46083
rect 20009 46037 20087 46083
rect 20133 46037 20211 46083
rect 20257 46037 20335 46083
rect 20381 46037 20459 46083
rect 20505 46037 20583 46083
rect 20629 46037 20707 46083
rect 20753 46037 20831 46083
rect 20877 46037 20955 46083
rect 21001 46037 21079 46083
rect 21125 46037 21203 46083
rect 21249 46037 21327 46083
rect 21373 46037 21451 46083
rect 21497 46037 21575 46083
rect 21621 46037 21699 46083
rect 21745 46037 21823 46083
rect 21869 46037 21947 46083
rect 21993 46037 22071 46083
rect 22117 46037 22195 46083
rect 22241 46037 22319 46083
rect 22365 46037 22443 46083
rect 22489 46037 22567 46083
rect 22613 46037 22691 46083
rect 22737 46037 22815 46083
rect 22861 46037 22939 46083
rect 22985 46037 23063 46083
rect 23109 46037 23187 46083
rect 23233 46037 23311 46083
rect 23357 46037 23435 46083
rect 23481 46037 23559 46083
rect 23605 46037 23683 46083
rect 23729 46037 23807 46083
rect 23853 46037 23931 46083
rect 23977 46037 24055 46083
rect 24101 46037 24179 46083
rect 24225 46037 24303 46083
rect 24349 46037 24427 46083
rect 24473 46037 24551 46083
rect 24597 46037 24675 46083
rect 24721 46037 24799 46083
rect 24845 46037 24923 46083
rect 24969 46037 25047 46083
rect 25093 46037 25171 46083
rect 25217 46037 25295 46083
rect 25341 46037 25419 46083
rect 25465 46037 25543 46083
rect 25589 46037 25667 46083
rect 25713 46037 25791 46083
rect 25837 46037 25915 46083
rect 25961 46037 26039 46083
rect 26085 46037 26163 46083
rect 26209 46037 26287 46083
rect 26333 46037 26411 46083
rect 26457 46037 26535 46083
rect 26581 46037 26659 46083
rect 26705 46037 26783 46083
rect 26829 46037 26907 46083
rect 26953 46037 27031 46083
rect 27077 46037 27155 46083
rect 27201 46037 27279 46083
rect 27325 46037 27403 46083
rect 27449 46037 27527 46083
rect 27573 46037 27651 46083
rect 27697 46037 27775 46083
rect 27821 46037 27899 46083
rect 27945 46037 28023 46083
rect 28069 46037 28147 46083
rect 28193 46037 28271 46083
rect 28317 46037 28395 46083
rect 28441 46037 28519 46083
rect 28565 46037 28643 46083
rect 28689 46037 28767 46083
rect 28813 46037 28891 46083
rect 28937 46037 29015 46083
rect 29061 46037 29139 46083
rect 29185 46037 29263 46083
rect 29309 46037 29387 46083
rect 29433 46037 29511 46083
rect 29557 46037 29635 46083
rect 29681 46037 29759 46083
rect 29805 46037 29883 46083
rect 29929 46037 30007 46083
rect 30053 46037 30131 46083
rect 30177 46037 30255 46083
rect 30301 46037 30379 46083
rect 30425 46037 30503 46083
rect 30549 46037 30627 46083
rect 30673 46037 30751 46083
rect 30797 46037 30875 46083
rect 30921 46037 30999 46083
rect 31045 46037 31123 46083
rect 31169 46037 31247 46083
rect 31293 46037 31371 46083
rect 31417 46037 31495 46083
rect 31541 46037 31619 46083
rect 31665 46037 31743 46083
rect 31789 46037 31867 46083
rect 31913 46037 31991 46083
rect 32037 46037 32115 46083
rect 32161 46037 32239 46083
rect 32285 46037 32363 46083
rect 32409 46037 32487 46083
rect 32533 46037 32611 46083
rect 32657 46037 32735 46083
rect 32781 46037 32859 46083
rect 32905 46037 32983 46083
rect 33029 46037 33107 46083
rect 33153 46037 33231 46083
rect 33277 46037 33355 46083
rect 33401 46037 33479 46083
rect 33525 46037 33603 46083
rect 33649 46037 33727 46083
rect 33773 46037 33851 46083
rect 33897 46037 33975 46083
rect 34021 46037 34099 46083
rect 34145 46037 34223 46083
rect 34269 46037 34347 46083
rect 34393 46037 34471 46083
rect 34517 46037 34595 46083
rect 34641 46037 34719 46083
rect 34765 46037 34843 46083
rect 34889 46037 34967 46083
rect 35013 46037 35091 46083
rect 35137 46037 35215 46083
rect 35261 46037 35339 46083
rect 35385 46037 35463 46083
rect 35509 46037 35587 46083
rect 35633 46037 35711 46083
rect 35757 46037 35835 46083
rect 35881 46037 35959 46083
rect 36005 46037 36083 46083
rect 36129 46037 36207 46083
rect 36253 46037 36331 46083
rect 36377 46037 36455 46083
rect 36501 46037 36579 46083
rect 36625 46037 36703 46083
rect 36749 46037 36827 46083
rect 36873 46037 36951 46083
rect 36997 46037 37075 46083
rect 37121 46037 37199 46083
rect 37245 46037 37323 46083
rect 37369 46037 37447 46083
rect 37493 46037 37571 46083
rect 37617 46037 37695 46083
rect 37741 46037 37819 46083
rect 37865 46037 37943 46083
rect 37989 46037 38067 46083
rect 38113 46037 38191 46083
rect 38237 46037 38315 46083
rect 38361 46037 38439 46083
rect 38485 46037 38563 46083
rect 38609 46037 38687 46083
rect 38733 46037 38811 46083
rect 38857 46037 38935 46083
rect 38981 46037 39059 46083
rect 39105 46037 39183 46083
rect 39229 46037 39307 46083
rect 39353 46037 39431 46083
rect 39477 46037 39555 46083
rect 39601 46037 39679 46083
rect 39725 46037 39803 46083
rect 39849 46037 39927 46083
rect 39973 46037 40051 46083
rect 40097 46037 40175 46083
rect 40221 46037 40299 46083
rect 40345 46037 40423 46083
rect 40469 46037 40547 46083
rect 40593 46037 40671 46083
rect 40717 46037 40795 46083
rect 40841 46037 40919 46083
rect 40965 46037 41043 46083
rect 41089 46037 41167 46083
rect 41213 46037 41291 46083
rect 41337 46037 41415 46083
rect 41461 46037 41539 46083
rect 41585 46037 41663 46083
rect 41709 46037 41787 46083
rect 41833 46037 41911 46083
rect 41957 46037 42035 46083
rect 42081 46037 42159 46083
rect 42205 46037 42283 46083
rect 42329 46037 42407 46083
rect 42453 46037 42531 46083
rect 42577 46037 42655 46083
rect 42701 46037 42779 46083
rect 42825 46037 42903 46083
rect 42949 46037 43027 46083
rect 43073 46037 43151 46083
rect 43197 46037 43275 46083
rect 43321 46037 43399 46083
rect 43445 46037 43523 46083
rect 43569 46037 43647 46083
rect 43693 46037 43771 46083
rect 43817 46037 43895 46083
rect 43941 46037 44019 46083
rect 44065 46037 44143 46083
rect 44189 46037 44267 46083
rect 44313 46037 44391 46083
rect 44437 46037 44515 46083
rect 44561 46037 44639 46083
rect 44685 46037 44763 46083
rect 44809 46037 44887 46083
rect 44933 46037 45011 46083
rect 45057 46037 45135 46083
rect 45181 46037 45259 46083
rect 45305 46037 45383 46083
rect 45429 46037 45507 46083
rect 45553 46037 45631 46083
rect 45677 46037 45755 46083
rect 45801 46037 45879 46083
rect 45925 46037 46003 46083
rect 46049 46037 46127 46083
rect 46173 46037 46251 46083
rect 46297 46037 46375 46083
rect 46421 46037 46499 46083
rect 46545 46037 46623 46083
rect 46669 46037 46747 46083
rect 46793 46037 46871 46083
rect 46917 46037 46995 46083
rect 47041 46037 47119 46083
rect 47165 46037 47243 46083
rect 47289 46037 47367 46083
rect 47413 46037 47491 46083
rect 47537 46037 47615 46083
rect 47661 46037 47739 46083
rect 47785 46037 47863 46083
rect 47909 46037 47987 46083
rect 48033 46037 48111 46083
rect 48157 46037 48235 46083
rect 48281 46037 48359 46083
rect 48405 46037 48483 46083
rect 48529 46037 48607 46083
rect 48653 46037 48731 46083
rect 48777 46037 48855 46083
rect 48901 46037 48979 46083
rect 49025 46037 49103 46083
rect 49149 46037 49227 46083
rect 49273 46037 49351 46083
rect 49397 46037 49475 46083
rect 49521 46037 49599 46083
rect 49645 46037 49723 46083
rect 49769 46037 49847 46083
rect 49893 46037 49971 46083
rect 50017 46037 50095 46083
rect 50141 46037 50219 46083
rect 50265 46037 50343 46083
rect 50389 46037 50467 46083
rect 50513 46037 50591 46083
rect 50637 46037 50715 46083
rect 50761 46037 50839 46083
rect 50885 46037 50963 46083
rect 51009 46037 51087 46083
rect 51133 46037 51211 46083
rect 51257 46037 51335 46083
rect 51381 46037 51459 46083
rect 51505 46037 51583 46083
rect 51629 46037 51707 46083
rect 51753 46037 51831 46083
rect 51877 46037 51955 46083
rect 52001 46037 52079 46083
rect 52125 46037 52203 46083
rect 52249 46037 52327 46083
rect 52373 46037 52451 46083
rect 52497 46037 52575 46083
rect 52621 46037 52699 46083
rect 52745 46037 52823 46083
rect 52869 46037 52947 46083
rect 52993 46037 53071 46083
rect 53117 46037 53195 46083
rect 53241 46037 53319 46083
rect 53365 46037 53443 46083
rect 53489 46037 53567 46083
rect 53613 46037 53691 46083
rect 53737 46037 53815 46083
rect 53861 46037 53939 46083
rect 53985 46037 54063 46083
rect 54109 46037 54187 46083
rect 54233 46037 54311 46083
rect 54357 46037 54435 46083
rect 54481 46037 54559 46083
rect 54605 46037 54683 46083
rect 54729 46037 54807 46083
rect 54853 46037 54931 46083
rect 54977 46037 55055 46083
rect 55101 46037 55179 46083
rect 55225 46037 55303 46083
rect 55349 46037 55427 46083
rect 55473 46037 55551 46083
rect 55597 46037 55675 46083
rect 55721 46037 55799 46083
rect 55845 46037 55923 46083
rect 55969 46037 56047 46083
rect 56093 46037 56171 46083
rect 56217 46037 56295 46083
rect 56341 46037 56419 46083
rect 56465 46037 56543 46083
rect 56589 46037 56667 46083
rect 56713 46037 56791 46083
rect 56837 46037 56915 46083
rect 56961 46037 57039 46083
rect 57085 46037 57163 46083
rect 57209 46037 57287 46083
rect 57333 46037 57411 46083
rect 57457 46037 57535 46083
rect 57581 46037 57659 46083
rect 57705 46037 57783 46083
rect 57829 46037 57907 46083
rect 57953 46037 58031 46083
rect 58077 46037 58155 46083
rect 58201 46037 58279 46083
rect 58325 46037 58403 46083
rect 58449 46037 58527 46083
rect 58573 46037 58651 46083
rect 58697 46037 58775 46083
rect 58821 46037 58899 46083
rect 58945 46037 59023 46083
rect 59069 46037 59147 46083
rect 59193 46037 59271 46083
rect 59317 46037 59395 46083
rect 59441 46037 59519 46083
rect 59565 46037 59643 46083
rect 59689 46037 59767 46083
rect 59813 46037 59891 46083
rect 59937 46037 60015 46083
rect 60061 46037 60139 46083
rect 60185 46037 60263 46083
rect 60309 46037 60387 46083
rect 60433 46037 60511 46083
rect 60557 46037 60635 46083
rect 60681 46037 60759 46083
rect 60805 46037 60883 46083
rect 60929 46037 61007 46083
rect 61053 46037 61131 46083
rect 61177 46037 61255 46083
rect 61301 46037 61379 46083
rect 61425 46037 61503 46083
rect 61549 46037 61627 46083
rect 61673 46037 61751 46083
rect 61797 46037 61875 46083
rect 61921 46037 61999 46083
rect 62045 46037 62123 46083
rect 62169 46037 62247 46083
rect 62293 46037 62371 46083
rect 62417 46037 62495 46083
rect 62541 46037 62619 46083
rect 62665 46037 62743 46083
rect 62789 46037 62867 46083
rect 62913 46037 62991 46083
rect 63037 46037 63115 46083
rect 63161 46037 63239 46083
rect 63285 46037 63363 46083
rect 63409 46037 63487 46083
rect 63533 46037 63611 46083
rect 63657 46037 63735 46083
rect 63781 46037 63859 46083
rect 63905 46037 63983 46083
rect 64029 46037 64107 46083
rect 64153 46037 64231 46083
rect 64277 46037 64355 46083
rect 64401 46037 64479 46083
rect 64525 46037 64603 46083
rect 64649 46037 64727 46083
rect 64773 46037 64851 46083
rect 64897 46037 64975 46083
rect 65021 46037 65099 46083
rect 65145 46037 65223 46083
rect 65269 46037 65347 46083
rect 65393 46037 65471 46083
rect 65517 46037 65595 46083
rect 65641 46037 65719 46083
rect 65765 46037 65843 46083
rect 65889 46037 65967 46083
rect 66013 46037 66091 46083
rect 66137 46037 66215 46083
rect 66261 46037 66339 46083
rect 66385 46037 66463 46083
rect 66509 46037 66587 46083
rect 66633 46037 66711 46083
rect 66757 46037 66835 46083
rect 66881 46037 66959 46083
rect 67005 46037 67083 46083
rect 67129 46037 67207 46083
rect 67253 46037 67331 46083
rect 67377 46037 67455 46083
rect 67501 46037 67579 46083
rect 67625 46037 67703 46083
rect 67749 46037 67827 46083
rect 67873 46037 67951 46083
rect 67997 46037 68075 46083
rect 68121 46037 68199 46083
rect 68245 46037 68323 46083
rect 68369 46037 68447 46083
rect 68493 46037 68571 46083
rect 68617 46037 68695 46083
rect 68741 46037 68819 46083
rect 68865 46037 68943 46083
rect 68989 46037 69067 46083
rect 69113 46037 69191 46083
rect 69237 46037 69315 46083
rect 69361 46037 69439 46083
rect 69485 46037 69563 46083
rect 69609 46037 69687 46083
rect 69733 46037 69811 46083
rect 69857 46037 69935 46083
rect 69981 46037 70059 46083
rect 70105 46037 70183 46083
rect 70229 46037 70307 46083
rect 70353 46037 70431 46083
rect 70477 46037 70555 46083
rect 70601 46037 70679 46083
rect 70725 46037 70803 46083
rect 70849 46037 70927 46083
rect 70973 46037 71051 46083
rect 71097 46037 71175 46083
rect 71221 46037 71299 46083
rect 71345 46037 71423 46083
rect 71469 46037 71547 46083
rect 71593 46037 71671 46083
rect 71717 46037 71795 46083
rect 71841 46037 71919 46083
rect 71965 46037 72043 46083
rect 72089 46037 72167 46083
rect 72213 46037 72291 46083
rect 72337 46037 72415 46083
rect 72461 46037 72539 46083
rect 72585 46037 72663 46083
rect 72709 46037 72787 46083
rect 72833 46037 72911 46083
rect 72957 46037 73035 46083
rect 73081 46037 73159 46083
rect 73205 46037 73283 46083
rect 73329 46037 73407 46083
rect 73453 46037 73531 46083
rect 73577 46037 73655 46083
rect 73701 46037 73779 46083
rect 73825 46037 73903 46083
rect 73949 46037 74027 46083
rect 74073 46037 74151 46083
rect 74197 46037 74275 46083
rect 74321 46037 74399 46083
rect 74445 46037 74523 46083
rect 74569 46037 74647 46083
rect 74693 46037 74771 46083
rect 74817 46037 74895 46083
rect 74941 46037 75019 46083
rect 75065 46037 75143 46083
rect 75189 46037 75267 46083
rect 75313 46037 75391 46083
rect 75437 46037 75515 46083
rect 75561 46037 75639 46083
rect 75685 46037 75763 46083
rect 75809 46037 75887 46083
rect 75933 46037 76011 46083
rect 76057 46037 76135 46083
rect 76181 46037 76259 46083
rect 76305 46037 76383 46083
rect 76429 46037 76507 46083
rect 76553 46037 76631 46083
rect 76677 46037 76755 46083
rect 76801 46037 76879 46083
rect 76925 46037 77003 46083
rect 77049 46037 77127 46083
rect 77173 46037 77251 46083
rect 77297 46037 77375 46083
rect 77421 46037 77499 46083
rect 77545 46037 77623 46083
rect 77669 46037 77747 46083
rect 77793 46037 77871 46083
rect 77917 46037 77995 46083
rect 78041 46037 78119 46083
rect 78165 46037 78243 46083
rect 78289 46037 78367 46083
rect 78413 46037 78491 46083
rect 78537 46037 78615 46083
rect 78661 46037 78739 46083
rect 78785 46037 78863 46083
rect 78909 46037 78987 46083
rect 79033 46037 79111 46083
rect 79157 46037 79235 46083
rect 79281 46037 79359 46083
rect 79405 46037 79483 46083
rect 79529 46037 79607 46083
rect 79653 46037 79731 46083
rect 79777 46037 79855 46083
rect 79901 46037 79979 46083
rect 80025 46037 80103 46083
rect 80149 46037 80227 46083
rect 80273 46037 80351 46083
rect 80397 46037 80475 46083
rect 80521 46037 80599 46083
rect 80645 46037 80723 46083
rect 80769 46037 80847 46083
rect 80893 46037 80971 46083
rect 81017 46037 81095 46083
rect 81141 46037 81219 46083
rect 81265 46037 81343 46083
rect 81389 46037 81467 46083
rect 81513 46037 81591 46083
rect 81637 46037 81715 46083
rect 81761 46037 81839 46083
rect 81885 46037 81963 46083
rect 82009 46037 82087 46083
rect 82133 46037 82211 46083
rect 82257 46037 82335 46083
rect 82381 46037 82459 46083
rect 82505 46037 82583 46083
rect 82629 46037 82707 46083
rect 82753 46037 82831 46083
rect 82877 46037 82955 46083
rect 83001 46037 83079 46083
rect 83125 46037 83203 46083
rect 83249 46037 83327 46083
rect 83373 46037 83451 46083
rect 83497 46037 83575 46083
rect 83621 46037 83699 46083
rect 83745 46037 83823 46083
rect 83869 46037 83947 46083
rect 83993 46037 84071 46083
rect 84117 46037 84195 46083
rect 84241 46037 84319 46083
rect 84365 46037 84443 46083
rect 84489 46037 84567 46083
rect 84613 46037 84691 46083
rect 84737 46037 84815 46083
rect 84861 46037 84939 46083
rect 84985 46037 85063 46083
rect 85109 46037 85187 46083
rect 85233 46037 85311 46083
rect 85357 46037 85435 46083
rect 85481 46037 85559 46083
rect 85605 46037 85683 46083
rect 85729 46037 85807 46083
rect 85853 46037 85931 46083
rect 85977 46037 86090 46083
rect 282 45959 86090 46037
rect 282 45913 371 45959
rect 417 45913 495 45959
rect 541 45913 619 45959
rect 665 45913 743 45959
rect 789 45913 867 45959
rect 913 45913 991 45959
rect 1037 45913 1115 45959
rect 1161 45913 1239 45959
rect 1285 45913 1363 45959
rect 1409 45913 1487 45959
rect 1533 45913 1611 45959
rect 1657 45913 1735 45959
rect 1781 45913 1859 45959
rect 1905 45913 1983 45959
rect 2029 45913 2107 45959
rect 2153 45913 2231 45959
rect 2277 45913 2355 45959
rect 2401 45913 2479 45959
rect 2525 45913 2603 45959
rect 2649 45913 2727 45959
rect 2773 45913 2851 45959
rect 2897 45913 2975 45959
rect 3021 45913 3099 45959
rect 3145 45913 3223 45959
rect 3269 45913 3347 45959
rect 3393 45913 3471 45959
rect 3517 45913 3595 45959
rect 3641 45913 3719 45959
rect 3765 45913 3843 45959
rect 3889 45913 3967 45959
rect 4013 45913 4091 45959
rect 4137 45913 4215 45959
rect 4261 45913 4339 45959
rect 4385 45913 4463 45959
rect 4509 45913 4587 45959
rect 4633 45913 4711 45959
rect 4757 45913 4835 45959
rect 4881 45913 4959 45959
rect 5005 45913 5083 45959
rect 5129 45913 5207 45959
rect 5253 45913 5331 45959
rect 5377 45913 5455 45959
rect 5501 45913 5579 45959
rect 5625 45913 5703 45959
rect 5749 45913 5827 45959
rect 5873 45913 5951 45959
rect 5997 45913 6075 45959
rect 6121 45913 6199 45959
rect 6245 45913 6323 45959
rect 6369 45913 6447 45959
rect 6493 45913 6571 45959
rect 6617 45913 6695 45959
rect 6741 45913 6819 45959
rect 6865 45913 6943 45959
rect 6989 45913 7067 45959
rect 7113 45913 7191 45959
rect 7237 45913 7315 45959
rect 7361 45913 7439 45959
rect 7485 45913 7563 45959
rect 7609 45913 7687 45959
rect 7733 45913 7811 45959
rect 7857 45913 7935 45959
rect 7981 45913 8059 45959
rect 8105 45913 8183 45959
rect 8229 45913 8307 45959
rect 8353 45913 8431 45959
rect 8477 45913 8555 45959
rect 8601 45913 8679 45959
rect 8725 45913 8803 45959
rect 8849 45913 8927 45959
rect 8973 45913 9051 45959
rect 9097 45913 9175 45959
rect 9221 45913 9299 45959
rect 9345 45913 9423 45959
rect 9469 45913 9547 45959
rect 9593 45913 9671 45959
rect 9717 45913 9795 45959
rect 9841 45913 9919 45959
rect 9965 45913 10043 45959
rect 10089 45913 10167 45959
rect 10213 45913 10291 45959
rect 10337 45913 10415 45959
rect 10461 45913 10539 45959
rect 10585 45913 10663 45959
rect 10709 45913 10787 45959
rect 10833 45913 10911 45959
rect 10957 45913 11035 45959
rect 11081 45913 11159 45959
rect 11205 45913 11283 45959
rect 11329 45913 11407 45959
rect 11453 45913 11531 45959
rect 11577 45913 11655 45959
rect 11701 45913 11779 45959
rect 11825 45913 11903 45959
rect 11949 45913 12027 45959
rect 12073 45913 12151 45959
rect 12197 45913 12275 45959
rect 12321 45913 12399 45959
rect 12445 45913 12523 45959
rect 12569 45913 12647 45959
rect 12693 45913 12771 45959
rect 12817 45913 12895 45959
rect 12941 45913 13019 45959
rect 13065 45913 13143 45959
rect 13189 45913 13267 45959
rect 13313 45913 13391 45959
rect 13437 45913 13515 45959
rect 13561 45913 13639 45959
rect 13685 45913 13763 45959
rect 13809 45913 13887 45959
rect 13933 45913 14011 45959
rect 14057 45913 14135 45959
rect 14181 45913 14259 45959
rect 14305 45913 14383 45959
rect 14429 45913 14507 45959
rect 14553 45913 14631 45959
rect 14677 45913 14755 45959
rect 14801 45913 14879 45959
rect 14925 45913 15003 45959
rect 15049 45913 15127 45959
rect 15173 45913 15251 45959
rect 15297 45913 15375 45959
rect 15421 45913 15499 45959
rect 15545 45913 15623 45959
rect 15669 45913 15747 45959
rect 15793 45913 15871 45959
rect 15917 45913 15995 45959
rect 16041 45913 16119 45959
rect 16165 45913 16243 45959
rect 16289 45913 16367 45959
rect 16413 45913 16491 45959
rect 16537 45913 16615 45959
rect 16661 45913 16739 45959
rect 16785 45913 16863 45959
rect 16909 45913 16987 45959
rect 17033 45913 17111 45959
rect 17157 45913 17235 45959
rect 17281 45913 17359 45959
rect 17405 45913 17483 45959
rect 17529 45913 17607 45959
rect 17653 45913 17731 45959
rect 17777 45913 17855 45959
rect 17901 45913 17979 45959
rect 18025 45913 18103 45959
rect 18149 45913 18227 45959
rect 18273 45913 18351 45959
rect 18397 45913 18475 45959
rect 18521 45913 18599 45959
rect 18645 45913 18723 45959
rect 18769 45913 18847 45959
rect 18893 45913 18971 45959
rect 19017 45913 19095 45959
rect 19141 45913 19219 45959
rect 19265 45913 19343 45959
rect 19389 45913 19467 45959
rect 19513 45913 19591 45959
rect 19637 45913 19715 45959
rect 19761 45913 19839 45959
rect 19885 45913 19963 45959
rect 20009 45913 20087 45959
rect 20133 45913 20211 45959
rect 20257 45913 20335 45959
rect 20381 45913 20459 45959
rect 20505 45913 20583 45959
rect 20629 45913 20707 45959
rect 20753 45913 20831 45959
rect 20877 45913 20955 45959
rect 21001 45913 21079 45959
rect 21125 45913 21203 45959
rect 21249 45913 21327 45959
rect 21373 45913 21451 45959
rect 21497 45913 21575 45959
rect 21621 45913 21699 45959
rect 21745 45913 21823 45959
rect 21869 45913 21947 45959
rect 21993 45913 22071 45959
rect 22117 45913 22195 45959
rect 22241 45913 22319 45959
rect 22365 45913 22443 45959
rect 22489 45913 22567 45959
rect 22613 45913 22691 45959
rect 22737 45913 22815 45959
rect 22861 45913 22939 45959
rect 22985 45913 23063 45959
rect 23109 45913 23187 45959
rect 23233 45913 23311 45959
rect 23357 45913 23435 45959
rect 23481 45913 23559 45959
rect 23605 45913 23683 45959
rect 23729 45913 23807 45959
rect 23853 45913 23931 45959
rect 23977 45913 24055 45959
rect 24101 45913 24179 45959
rect 24225 45913 24303 45959
rect 24349 45913 24427 45959
rect 24473 45913 24551 45959
rect 24597 45913 24675 45959
rect 24721 45913 24799 45959
rect 24845 45913 24923 45959
rect 24969 45913 25047 45959
rect 25093 45913 25171 45959
rect 25217 45913 25295 45959
rect 25341 45913 25419 45959
rect 25465 45913 25543 45959
rect 25589 45913 25667 45959
rect 25713 45913 25791 45959
rect 25837 45913 25915 45959
rect 25961 45913 26039 45959
rect 26085 45913 26163 45959
rect 26209 45913 26287 45959
rect 26333 45913 26411 45959
rect 26457 45913 26535 45959
rect 26581 45913 26659 45959
rect 26705 45913 26783 45959
rect 26829 45913 26907 45959
rect 26953 45913 27031 45959
rect 27077 45913 27155 45959
rect 27201 45913 27279 45959
rect 27325 45913 27403 45959
rect 27449 45913 27527 45959
rect 27573 45913 27651 45959
rect 27697 45913 27775 45959
rect 27821 45913 27899 45959
rect 27945 45913 28023 45959
rect 28069 45913 28147 45959
rect 28193 45913 28271 45959
rect 28317 45913 28395 45959
rect 28441 45913 28519 45959
rect 28565 45913 28643 45959
rect 28689 45913 28767 45959
rect 28813 45913 28891 45959
rect 28937 45913 29015 45959
rect 29061 45913 29139 45959
rect 29185 45913 29263 45959
rect 29309 45913 29387 45959
rect 29433 45913 29511 45959
rect 29557 45913 29635 45959
rect 29681 45913 29759 45959
rect 29805 45913 29883 45959
rect 29929 45913 30007 45959
rect 30053 45913 30131 45959
rect 30177 45913 30255 45959
rect 30301 45913 30379 45959
rect 30425 45913 30503 45959
rect 30549 45913 30627 45959
rect 30673 45913 30751 45959
rect 30797 45913 30875 45959
rect 30921 45913 30999 45959
rect 31045 45913 31123 45959
rect 31169 45913 31247 45959
rect 31293 45913 31371 45959
rect 31417 45913 31495 45959
rect 31541 45913 31619 45959
rect 31665 45913 31743 45959
rect 31789 45913 31867 45959
rect 31913 45913 31991 45959
rect 32037 45913 32115 45959
rect 32161 45913 32239 45959
rect 32285 45913 32363 45959
rect 32409 45913 32487 45959
rect 32533 45913 32611 45959
rect 32657 45913 32735 45959
rect 32781 45913 32859 45959
rect 32905 45913 32983 45959
rect 33029 45913 33107 45959
rect 33153 45913 33231 45959
rect 33277 45913 33355 45959
rect 33401 45913 33479 45959
rect 33525 45913 33603 45959
rect 33649 45913 33727 45959
rect 33773 45913 33851 45959
rect 33897 45913 33975 45959
rect 34021 45913 34099 45959
rect 34145 45913 34223 45959
rect 34269 45913 34347 45959
rect 34393 45913 34471 45959
rect 34517 45913 34595 45959
rect 34641 45913 34719 45959
rect 34765 45913 34843 45959
rect 34889 45913 34967 45959
rect 35013 45913 35091 45959
rect 35137 45913 35215 45959
rect 35261 45913 35339 45959
rect 35385 45913 35463 45959
rect 35509 45913 35587 45959
rect 35633 45913 35711 45959
rect 35757 45913 35835 45959
rect 35881 45913 35959 45959
rect 36005 45913 36083 45959
rect 36129 45913 36207 45959
rect 36253 45913 36331 45959
rect 36377 45913 36455 45959
rect 36501 45913 36579 45959
rect 36625 45913 36703 45959
rect 36749 45913 36827 45959
rect 36873 45913 36951 45959
rect 36997 45913 37075 45959
rect 37121 45913 37199 45959
rect 37245 45913 37323 45959
rect 37369 45913 37447 45959
rect 37493 45913 37571 45959
rect 37617 45913 37695 45959
rect 37741 45913 37819 45959
rect 37865 45913 37943 45959
rect 37989 45913 38067 45959
rect 38113 45913 38191 45959
rect 38237 45913 38315 45959
rect 38361 45913 38439 45959
rect 38485 45913 38563 45959
rect 38609 45913 38687 45959
rect 38733 45913 38811 45959
rect 38857 45913 38935 45959
rect 38981 45913 39059 45959
rect 39105 45913 39183 45959
rect 39229 45913 39307 45959
rect 39353 45913 39431 45959
rect 39477 45913 39555 45959
rect 39601 45913 39679 45959
rect 39725 45913 39803 45959
rect 39849 45913 39927 45959
rect 39973 45913 40051 45959
rect 40097 45913 40175 45959
rect 40221 45913 40299 45959
rect 40345 45913 40423 45959
rect 40469 45913 40547 45959
rect 40593 45913 40671 45959
rect 40717 45913 40795 45959
rect 40841 45913 40919 45959
rect 40965 45913 41043 45959
rect 41089 45913 41167 45959
rect 41213 45913 41291 45959
rect 41337 45913 41415 45959
rect 41461 45913 41539 45959
rect 41585 45913 41663 45959
rect 41709 45913 41787 45959
rect 41833 45913 41911 45959
rect 41957 45913 42035 45959
rect 42081 45913 42159 45959
rect 42205 45913 42283 45959
rect 42329 45913 42407 45959
rect 42453 45913 42531 45959
rect 42577 45913 42655 45959
rect 42701 45913 42779 45959
rect 42825 45913 42903 45959
rect 42949 45913 43027 45959
rect 43073 45913 43151 45959
rect 43197 45913 43275 45959
rect 43321 45913 43399 45959
rect 43445 45913 43523 45959
rect 43569 45913 43647 45959
rect 43693 45913 43771 45959
rect 43817 45913 43895 45959
rect 43941 45913 44019 45959
rect 44065 45913 44143 45959
rect 44189 45913 44267 45959
rect 44313 45913 44391 45959
rect 44437 45913 44515 45959
rect 44561 45913 44639 45959
rect 44685 45913 44763 45959
rect 44809 45913 44887 45959
rect 44933 45913 45011 45959
rect 45057 45913 45135 45959
rect 45181 45913 45259 45959
rect 45305 45913 45383 45959
rect 45429 45913 45507 45959
rect 45553 45913 45631 45959
rect 45677 45913 45755 45959
rect 45801 45913 45879 45959
rect 45925 45913 46003 45959
rect 46049 45913 46127 45959
rect 46173 45913 46251 45959
rect 46297 45913 46375 45959
rect 46421 45913 46499 45959
rect 46545 45913 46623 45959
rect 46669 45913 46747 45959
rect 46793 45913 46871 45959
rect 46917 45913 46995 45959
rect 47041 45913 47119 45959
rect 47165 45913 47243 45959
rect 47289 45913 47367 45959
rect 47413 45913 47491 45959
rect 47537 45913 47615 45959
rect 47661 45913 47739 45959
rect 47785 45913 47863 45959
rect 47909 45913 47987 45959
rect 48033 45913 48111 45959
rect 48157 45913 48235 45959
rect 48281 45913 48359 45959
rect 48405 45913 48483 45959
rect 48529 45913 48607 45959
rect 48653 45913 48731 45959
rect 48777 45913 48855 45959
rect 48901 45913 48979 45959
rect 49025 45913 49103 45959
rect 49149 45913 49227 45959
rect 49273 45913 49351 45959
rect 49397 45913 49475 45959
rect 49521 45913 49599 45959
rect 49645 45913 49723 45959
rect 49769 45913 49847 45959
rect 49893 45913 49971 45959
rect 50017 45913 50095 45959
rect 50141 45913 50219 45959
rect 50265 45913 50343 45959
rect 50389 45913 50467 45959
rect 50513 45913 50591 45959
rect 50637 45913 50715 45959
rect 50761 45913 50839 45959
rect 50885 45913 50963 45959
rect 51009 45913 51087 45959
rect 51133 45913 51211 45959
rect 51257 45913 51335 45959
rect 51381 45913 51459 45959
rect 51505 45913 51583 45959
rect 51629 45913 51707 45959
rect 51753 45913 51831 45959
rect 51877 45913 51955 45959
rect 52001 45913 52079 45959
rect 52125 45913 52203 45959
rect 52249 45913 52327 45959
rect 52373 45913 52451 45959
rect 52497 45913 52575 45959
rect 52621 45913 52699 45959
rect 52745 45913 52823 45959
rect 52869 45913 52947 45959
rect 52993 45913 53071 45959
rect 53117 45913 53195 45959
rect 53241 45913 53319 45959
rect 53365 45913 53443 45959
rect 53489 45913 53567 45959
rect 53613 45913 53691 45959
rect 53737 45913 53815 45959
rect 53861 45913 53939 45959
rect 53985 45913 54063 45959
rect 54109 45913 54187 45959
rect 54233 45913 54311 45959
rect 54357 45913 54435 45959
rect 54481 45913 54559 45959
rect 54605 45913 54683 45959
rect 54729 45913 54807 45959
rect 54853 45913 54931 45959
rect 54977 45913 55055 45959
rect 55101 45913 55179 45959
rect 55225 45913 55303 45959
rect 55349 45913 55427 45959
rect 55473 45913 55551 45959
rect 55597 45913 55675 45959
rect 55721 45913 55799 45959
rect 55845 45913 55923 45959
rect 55969 45913 56047 45959
rect 56093 45913 56171 45959
rect 56217 45913 56295 45959
rect 56341 45913 56419 45959
rect 56465 45913 56543 45959
rect 56589 45913 56667 45959
rect 56713 45913 56791 45959
rect 56837 45913 56915 45959
rect 56961 45913 57039 45959
rect 57085 45913 57163 45959
rect 57209 45913 57287 45959
rect 57333 45913 57411 45959
rect 57457 45913 57535 45959
rect 57581 45913 57659 45959
rect 57705 45913 57783 45959
rect 57829 45913 57907 45959
rect 57953 45913 58031 45959
rect 58077 45913 58155 45959
rect 58201 45913 58279 45959
rect 58325 45913 58403 45959
rect 58449 45913 58527 45959
rect 58573 45913 58651 45959
rect 58697 45913 58775 45959
rect 58821 45913 58899 45959
rect 58945 45913 59023 45959
rect 59069 45913 59147 45959
rect 59193 45913 59271 45959
rect 59317 45913 59395 45959
rect 59441 45913 59519 45959
rect 59565 45913 59643 45959
rect 59689 45913 59767 45959
rect 59813 45913 59891 45959
rect 59937 45913 60015 45959
rect 60061 45913 60139 45959
rect 60185 45913 60263 45959
rect 60309 45913 60387 45959
rect 60433 45913 60511 45959
rect 60557 45913 60635 45959
rect 60681 45913 60759 45959
rect 60805 45913 60883 45959
rect 60929 45913 61007 45959
rect 61053 45913 61131 45959
rect 61177 45913 61255 45959
rect 61301 45913 61379 45959
rect 61425 45913 61503 45959
rect 61549 45913 61627 45959
rect 61673 45913 61751 45959
rect 61797 45913 61875 45959
rect 61921 45913 61999 45959
rect 62045 45913 62123 45959
rect 62169 45913 62247 45959
rect 62293 45913 62371 45959
rect 62417 45913 62495 45959
rect 62541 45913 62619 45959
rect 62665 45913 62743 45959
rect 62789 45913 62867 45959
rect 62913 45913 62991 45959
rect 63037 45913 63115 45959
rect 63161 45913 63239 45959
rect 63285 45913 63363 45959
rect 63409 45913 63487 45959
rect 63533 45913 63611 45959
rect 63657 45913 63735 45959
rect 63781 45913 63859 45959
rect 63905 45913 63983 45959
rect 64029 45913 64107 45959
rect 64153 45913 64231 45959
rect 64277 45913 64355 45959
rect 64401 45913 64479 45959
rect 64525 45913 64603 45959
rect 64649 45913 64727 45959
rect 64773 45913 64851 45959
rect 64897 45913 64975 45959
rect 65021 45913 65099 45959
rect 65145 45913 65223 45959
rect 65269 45913 65347 45959
rect 65393 45913 65471 45959
rect 65517 45913 65595 45959
rect 65641 45913 65719 45959
rect 65765 45913 65843 45959
rect 65889 45913 65967 45959
rect 66013 45913 66091 45959
rect 66137 45913 66215 45959
rect 66261 45913 66339 45959
rect 66385 45913 66463 45959
rect 66509 45913 66587 45959
rect 66633 45913 66711 45959
rect 66757 45913 66835 45959
rect 66881 45913 66959 45959
rect 67005 45913 67083 45959
rect 67129 45913 67207 45959
rect 67253 45913 67331 45959
rect 67377 45913 67455 45959
rect 67501 45913 67579 45959
rect 67625 45913 67703 45959
rect 67749 45913 67827 45959
rect 67873 45913 67951 45959
rect 67997 45913 68075 45959
rect 68121 45913 68199 45959
rect 68245 45913 68323 45959
rect 68369 45913 68447 45959
rect 68493 45913 68571 45959
rect 68617 45913 68695 45959
rect 68741 45913 68819 45959
rect 68865 45913 68943 45959
rect 68989 45913 69067 45959
rect 69113 45913 69191 45959
rect 69237 45913 69315 45959
rect 69361 45913 69439 45959
rect 69485 45913 69563 45959
rect 69609 45913 69687 45959
rect 69733 45913 69811 45959
rect 69857 45913 69935 45959
rect 69981 45913 70059 45959
rect 70105 45913 70183 45959
rect 70229 45913 70307 45959
rect 70353 45913 70431 45959
rect 70477 45913 70555 45959
rect 70601 45913 70679 45959
rect 70725 45913 70803 45959
rect 70849 45913 70927 45959
rect 70973 45913 71051 45959
rect 71097 45913 71175 45959
rect 71221 45913 71299 45959
rect 71345 45913 71423 45959
rect 71469 45913 71547 45959
rect 71593 45913 71671 45959
rect 71717 45913 71795 45959
rect 71841 45913 71919 45959
rect 71965 45913 72043 45959
rect 72089 45913 72167 45959
rect 72213 45913 72291 45959
rect 72337 45913 72415 45959
rect 72461 45913 72539 45959
rect 72585 45913 72663 45959
rect 72709 45913 72787 45959
rect 72833 45913 72911 45959
rect 72957 45913 73035 45959
rect 73081 45913 73159 45959
rect 73205 45913 73283 45959
rect 73329 45913 73407 45959
rect 73453 45913 73531 45959
rect 73577 45913 73655 45959
rect 73701 45913 73779 45959
rect 73825 45913 73903 45959
rect 73949 45913 74027 45959
rect 74073 45913 74151 45959
rect 74197 45913 74275 45959
rect 74321 45913 74399 45959
rect 74445 45913 74523 45959
rect 74569 45913 74647 45959
rect 74693 45913 74771 45959
rect 74817 45913 74895 45959
rect 74941 45913 75019 45959
rect 75065 45913 75143 45959
rect 75189 45913 75267 45959
rect 75313 45913 75391 45959
rect 75437 45913 75515 45959
rect 75561 45913 75639 45959
rect 75685 45913 75763 45959
rect 75809 45913 75887 45959
rect 75933 45913 76011 45959
rect 76057 45913 76135 45959
rect 76181 45913 76259 45959
rect 76305 45913 76383 45959
rect 76429 45913 76507 45959
rect 76553 45913 76631 45959
rect 76677 45913 76755 45959
rect 76801 45913 76879 45959
rect 76925 45913 77003 45959
rect 77049 45913 77127 45959
rect 77173 45913 77251 45959
rect 77297 45913 77375 45959
rect 77421 45913 77499 45959
rect 77545 45913 77623 45959
rect 77669 45913 77747 45959
rect 77793 45913 77871 45959
rect 77917 45913 77995 45959
rect 78041 45913 78119 45959
rect 78165 45913 78243 45959
rect 78289 45913 78367 45959
rect 78413 45913 78491 45959
rect 78537 45913 78615 45959
rect 78661 45913 78739 45959
rect 78785 45913 78863 45959
rect 78909 45913 78987 45959
rect 79033 45913 79111 45959
rect 79157 45913 79235 45959
rect 79281 45913 79359 45959
rect 79405 45913 79483 45959
rect 79529 45913 79607 45959
rect 79653 45913 79731 45959
rect 79777 45913 79855 45959
rect 79901 45913 79979 45959
rect 80025 45913 80103 45959
rect 80149 45913 80227 45959
rect 80273 45913 80351 45959
rect 80397 45913 80475 45959
rect 80521 45913 80599 45959
rect 80645 45913 80723 45959
rect 80769 45913 80847 45959
rect 80893 45913 80971 45959
rect 81017 45913 81095 45959
rect 81141 45913 81219 45959
rect 81265 45913 81343 45959
rect 81389 45913 81467 45959
rect 81513 45913 81591 45959
rect 81637 45913 81715 45959
rect 81761 45913 81839 45959
rect 81885 45913 81963 45959
rect 82009 45913 82087 45959
rect 82133 45913 82211 45959
rect 82257 45913 82335 45959
rect 82381 45913 82459 45959
rect 82505 45913 82583 45959
rect 82629 45913 82707 45959
rect 82753 45913 82831 45959
rect 82877 45913 82955 45959
rect 83001 45913 83079 45959
rect 83125 45913 83203 45959
rect 83249 45913 83327 45959
rect 83373 45913 83451 45959
rect 83497 45913 83575 45959
rect 83621 45913 83699 45959
rect 83745 45913 83823 45959
rect 83869 45913 83947 45959
rect 83993 45913 84071 45959
rect 84117 45913 84195 45959
rect 84241 45913 84319 45959
rect 84365 45913 84443 45959
rect 84489 45913 84567 45959
rect 84613 45913 84691 45959
rect 84737 45913 84815 45959
rect 84861 45913 84939 45959
rect 84985 45913 85063 45959
rect 85109 45913 85187 45959
rect 85233 45913 85311 45959
rect 85357 45913 85435 45959
rect 85481 45913 85559 45959
rect 85605 45913 85683 45959
rect 85729 45913 85807 45959
rect 85853 45913 85931 45959
rect 85977 45913 86090 45959
rect 282 45835 86090 45913
rect 282 45789 371 45835
rect 417 45789 495 45835
rect 541 45789 619 45835
rect 665 45789 743 45835
rect 789 45789 867 45835
rect 913 45789 991 45835
rect 1037 45789 1115 45835
rect 1161 45789 1239 45835
rect 1285 45789 1363 45835
rect 1409 45789 1487 45835
rect 1533 45789 1611 45835
rect 1657 45789 1735 45835
rect 1781 45789 1859 45835
rect 1905 45789 1983 45835
rect 2029 45789 2107 45835
rect 2153 45789 2231 45835
rect 2277 45789 2355 45835
rect 2401 45789 2479 45835
rect 2525 45789 2603 45835
rect 2649 45789 2727 45835
rect 2773 45789 2851 45835
rect 2897 45789 2975 45835
rect 3021 45789 3099 45835
rect 3145 45789 3223 45835
rect 3269 45789 3347 45835
rect 3393 45789 3471 45835
rect 3517 45789 3595 45835
rect 3641 45789 3719 45835
rect 3765 45789 3843 45835
rect 3889 45789 3967 45835
rect 4013 45789 4091 45835
rect 4137 45789 4215 45835
rect 4261 45789 4339 45835
rect 4385 45789 4463 45835
rect 4509 45789 4587 45835
rect 4633 45789 4711 45835
rect 4757 45789 4835 45835
rect 4881 45789 4959 45835
rect 5005 45789 5083 45835
rect 5129 45789 5207 45835
rect 5253 45789 5331 45835
rect 5377 45789 5455 45835
rect 5501 45789 5579 45835
rect 5625 45789 5703 45835
rect 5749 45789 5827 45835
rect 5873 45789 5951 45835
rect 5997 45789 6075 45835
rect 6121 45789 6199 45835
rect 6245 45789 6323 45835
rect 6369 45789 6447 45835
rect 6493 45789 6571 45835
rect 6617 45789 6695 45835
rect 6741 45789 6819 45835
rect 6865 45789 6943 45835
rect 6989 45789 7067 45835
rect 7113 45789 7191 45835
rect 7237 45789 7315 45835
rect 7361 45789 7439 45835
rect 7485 45789 7563 45835
rect 7609 45789 7687 45835
rect 7733 45789 7811 45835
rect 7857 45789 7935 45835
rect 7981 45789 8059 45835
rect 8105 45789 8183 45835
rect 8229 45789 8307 45835
rect 8353 45789 8431 45835
rect 8477 45789 8555 45835
rect 8601 45789 8679 45835
rect 8725 45789 8803 45835
rect 8849 45789 8927 45835
rect 8973 45789 9051 45835
rect 9097 45789 9175 45835
rect 9221 45789 9299 45835
rect 9345 45789 9423 45835
rect 9469 45789 9547 45835
rect 9593 45789 9671 45835
rect 9717 45789 9795 45835
rect 9841 45789 9919 45835
rect 9965 45789 10043 45835
rect 10089 45789 10167 45835
rect 10213 45789 10291 45835
rect 10337 45789 10415 45835
rect 10461 45789 10539 45835
rect 10585 45789 10663 45835
rect 10709 45789 10787 45835
rect 10833 45789 10911 45835
rect 10957 45789 11035 45835
rect 11081 45789 11159 45835
rect 11205 45789 11283 45835
rect 11329 45789 11407 45835
rect 11453 45789 11531 45835
rect 11577 45789 11655 45835
rect 11701 45789 11779 45835
rect 11825 45789 11903 45835
rect 11949 45789 12027 45835
rect 12073 45789 12151 45835
rect 12197 45789 12275 45835
rect 12321 45789 12399 45835
rect 12445 45789 12523 45835
rect 12569 45789 12647 45835
rect 12693 45789 12771 45835
rect 12817 45789 12895 45835
rect 12941 45789 13019 45835
rect 13065 45789 13143 45835
rect 13189 45789 13267 45835
rect 13313 45789 13391 45835
rect 13437 45789 13515 45835
rect 13561 45789 13639 45835
rect 13685 45789 13763 45835
rect 13809 45789 13887 45835
rect 13933 45789 14011 45835
rect 14057 45789 14135 45835
rect 14181 45789 14259 45835
rect 14305 45789 14383 45835
rect 14429 45789 14507 45835
rect 14553 45789 14631 45835
rect 14677 45789 14755 45835
rect 14801 45789 14879 45835
rect 14925 45789 15003 45835
rect 15049 45789 15127 45835
rect 15173 45789 15251 45835
rect 15297 45789 15375 45835
rect 15421 45789 15499 45835
rect 15545 45789 15623 45835
rect 15669 45789 15747 45835
rect 15793 45789 15871 45835
rect 15917 45789 15995 45835
rect 16041 45789 16119 45835
rect 16165 45789 16243 45835
rect 16289 45789 16367 45835
rect 16413 45789 16491 45835
rect 16537 45789 16615 45835
rect 16661 45789 16739 45835
rect 16785 45789 16863 45835
rect 16909 45789 16987 45835
rect 17033 45789 17111 45835
rect 17157 45789 17235 45835
rect 17281 45789 17359 45835
rect 17405 45789 17483 45835
rect 17529 45789 17607 45835
rect 17653 45789 17731 45835
rect 17777 45789 17855 45835
rect 17901 45789 17979 45835
rect 18025 45789 18103 45835
rect 18149 45789 18227 45835
rect 18273 45789 18351 45835
rect 18397 45789 18475 45835
rect 18521 45789 18599 45835
rect 18645 45789 18723 45835
rect 18769 45789 18847 45835
rect 18893 45789 18971 45835
rect 19017 45789 19095 45835
rect 19141 45789 19219 45835
rect 19265 45789 19343 45835
rect 19389 45789 19467 45835
rect 19513 45789 19591 45835
rect 19637 45789 19715 45835
rect 19761 45789 19839 45835
rect 19885 45789 19963 45835
rect 20009 45789 20087 45835
rect 20133 45789 20211 45835
rect 20257 45789 20335 45835
rect 20381 45789 20459 45835
rect 20505 45789 20583 45835
rect 20629 45789 20707 45835
rect 20753 45789 20831 45835
rect 20877 45789 20955 45835
rect 21001 45789 21079 45835
rect 21125 45789 21203 45835
rect 21249 45789 21327 45835
rect 21373 45789 21451 45835
rect 21497 45789 21575 45835
rect 21621 45789 21699 45835
rect 21745 45789 21823 45835
rect 21869 45789 21947 45835
rect 21993 45789 22071 45835
rect 22117 45789 22195 45835
rect 22241 45789 22319 45835
rect 22365 45789 22443 45835
rect 22489 45789 22567 45835
rect 22613 45789 22691 45835
rect 22737 45789 22815 45835
rect 22861 45789 22939 45835
rect 22985 45789 23063 45835
rect 23109 45789 23187 45835
rect 23233 45789 23311 45835
rect 23357 45789 23435 45835
rect 23481 45789 23559 45835
rect 23605 45789 23683 45835
rect 23729 45789 23807 45835
rect 23853 45789 23931 45835
rect 23977 45789 24055 45835
rect 24101 45789 24179 45835
rect 24225 45789 24303 45835
rect 24349 45789 24427 45835
rect 24473 45789 24551 45835
rect 24597 45789 24675 45835
rect 24721 45789 24799 45835
rect 24845 45789 24923 45835
rect 24969 45789 25047 45835
rect 25093 45789 25171 45835
rect 25217 45789 25295 45835
rect 25341 45789 25419 45835
rect 25465 45789 25543 45835
rect 25589 45789 25667 45835
rect 25713 45789 25791 45835
rect 25837 45789 25915 45835
rect 25961 45789 26039 45835
rect 26085 45789 26163 45835
rect 26209 45789 26287 45835
rect 26333 45789 26411 45835
rect 26457 45789 26535 45835
rect 26581 45789 26659 45835
rect 26705 45789 26783 45835
rect 26829 45789 26907 45835
rect 26953 45789 27031 45835
rect 27077 45789 27155 45835
rect 27201 45789 27279 45835
rect 27325 45789 27403 45835
rect 27449 45789 27527 45835
rect 27573 45789 27651 45835
rect 27697 45789 27775 45835
rect 27821 45789 27899 45835
rect 27945 45789 28023 45835
rect 28069 45789 28147 45835
rect 28193 45789 28271 45835
rect 28317 45789 28395 45835
rect 28441 45789 28519 45835
rect 28565 45789 28643 45835
rect 28689 45789 28767 45835
rect 28813 45789 28891 45835
rect 28937 45789 29015 45835
rect 29061 45789 29139 45835
rect 29185 45789 29263 45835
rect 29309 45789 29387 45835
rect 29433 45789 29511 45835
rect 29557 45789 29635 45835
rect 29681 45789 29759 45835
rect 29805 45789 29883 45835
rect 29929 45789 30007 45835
rect 30053 45789 30131 45835
rect 30177 45789 30255 45835
rect 30301 45789 30379 45835
rect 30425 45789 30503 45835
rect 30549 45789 30627 45835
rect 30673 45789 30751 45835
rect 30797 45789 30875 45835
rect 30921 45789 30999 45835
rect 31045 45789 31123 45835
rect 31169 45789 31247 45835
rect 31293 45789 31371 45835
rect 31417 45789 31495 45835
rect 31541 45789 31619 45835
rect 31665 45789 31743 45835
rect 31789 45789 31867 45835
rect 31913 45789 31991 45835
rect 32037 45789 32115 45835
rect 32161 45789 32239 45835
rect 32285 45789 32363 45835
rect 32409 45789 32487 45835
rect 32533 45789 32611 45835
rect 32657 45789 32735 45835
rect 32781 45789 32859 45835
rect 32905 45789 32983 45835
rect 33029 45789 33107 45835
rect 33153 45789 33231 45835
rect 33277 45789 33355 45835
rect 33401 45789 33479 45835
rect 33525 45789 33603 45835
rect 33649 45789 33727 45835
rect 33773 45789 33851 45835
rect 33897 45789 33975 45835
rect 34021 45789 34099 45835
rect 34145 45789 34223 45835
rect 34269 45789 34347 45835
rect 34393 45789 34471 45835
rect 34517 45789 34595 45835
rect 34641 45789 34719 45835
rect 34765 45789 34843 45835
rect 34889 45789 34967 45835
rect 35013 45789 35091 45835
rect 35137 45789 35215 45835
rect 35261 45789 35339 45835
rect 35385 45789 35463 45835
rect 35509 45789 35587 45835
rect 35633 45789 35711 45835
rect 35757 45789 35835 45835
rect 35881 45789 35959 45835
rect 36005 45789 36083 45835
rect 36129 45789 36207 45835
rect 36253 45789 36331 45835
rect 36377 45789 36455 45835
rect 36501 45789 36579 45835
rect 36625 45789 36703 45835
rect 36749 45789 36827 45835
rect 36873 45789 36951 45835
rect 36997 45789 37075 45835
rect 37121 45789 37199 45835
rect 37245 45789 37323 45835
rect 37369 45789 37447 45835
rect 37493 45789 37571 45835
rect 37617 45789 37695 45835
rect 37741 45789 37819 45835
rect 37865 45789 37943 45835
rect 37989 45789 38067 45835
rect 38113 45789 38191 45835
rect 38237 45789 38315 45835
rect 38361 45789 38439 45835
rect 38485 45789 38563 45835
rect 38609 45789 38687 45835
rect 38733 45789 38811 45835
rect 38857 45789 38935 45835
rect 38981 45789 39059 45835
rect 39105 45789 39183 45835
rect 39229 45789 39307 45835
rect 39353 45789 39431 45835
rect 39477 45789 39555 45835
rect 39601 45789 39679 45835
rect 39725 45789 39803 45835
rect 39849 45789 39927 45835
rect 39973 45789 40051 45835
rect 40097 45789 40175 45835
rect 40221 45789 40299 45835
rect 40345 45789 40423 45835
rect 40469 45789 40547 45835
rect 40593 45789 40671 45835
rect 40717 45789 40795 45835
rect 40841 45789 40919 45835
rect 40965 45789 41043 45835
rect 41089 45789 41167 45835
rect 41213 45789 41291 45835
rect 41337 45789 41415 45835
rect 41461 45789 41539 45835
rect 41585 45789 41663 45835
rect 41709 45789 41787 45835
rect 41833 45789 41911 45835
rect 41957 45789 42035 45835
rect 42081 45789 42159 45835
rect 42205 45789 42283 45835
rect 42329 45789 42407 45835
rect 42453 45789 42531 45835
rect 42577 45789 42655 45835
rect 42701 45789 42779 45835
rect 42825 45789 42903 45835
rect 42949 45789 43027 45835
rect 43073 45789 43151 45835
rect 43197 45789 43275 45835
rect 43321 45789 43399 45835
rect 43445 45789 43523 45835
rect 43569 45789 43647 45835
rect 43693 45789 43771 45835
rect 43817 45789 43895 45835
rect 43941 45789 44019 45835
rect 44065 45789 44143 45835
rect 44189 45789 44267 45835
rect 44313 45789 44391 45835
rect 44437 45789 44515 45835
rect 44561 45789 44639 45835
rect 44685 45789 44763 45835
rect 44809 45789 44887 45835
rect 44933 45789 45011 45835
rect 45057 45789 45135 45835
rect 45181 45789 45259 45835
rect 45305 45789 45383 45835
rect 45429 45789 45507 45835
rect 45553 45789 45631 45835
rect 45677 45789 45755 45835
rect 45801 45789 45879 45835
rect 45925 45789 46003 45835
rect 46049 45789 46127 45835
rect 46173 45789 46251 45835
rect 46297 45789 46375 45835
rect 46421 45789 46499 45835
rect 46545 45789 46623 45835
rect 46669 45789 46747 45835
rect 46793 45789 46871 45835
rect 46917 45789 46995 45835
rect 47041 45789 47119 45835
rect 47165 45789 47243 45835
rect 47289 45789 47367 45835
rect 47413 45789 47491 45835
rect 47537 45789 47615 45835
rect 47661 45789 47739 45835
rect 47785 45789 47863 45835
rect 47909 45789 47987 45835
rect 48033 45789 48111 45835
rect 48157 45789 48235 45835
rect 48281 45789 48359 45835
rect 48405 45789 48483 45835
rect 48529 45789 48607 45835
rect 48653 45789 48731 45835
rect 48777 45789 48855 45835
rect 48901 45789 48979 45835
rect 49025 45789 49103 45835
rect 49149 45789 49227 45835
rect 49273 45789 49351 45835
rect 49397 45789 49475 45835
rect 49521 45789 49599 45835
rect 49645 45789 49723 45835
rect 49769 45789 49847 45835
rect 49893 45789 49971 45835
rect 50017 45789 50095 45835
rect 50141 45789 50219 45835
rect 50265 45789 50343 45835
rect 50389 45789 50467 45835
rect 50513 45789 50591 45835
rect 50637 45789 50715 45835
rect 50761 45789 50839 45835
rect 50885 45789 50963 45835
rect 51009 45789 51087 45835
rect 51133 45789 51211 45835
rect 51257 45789 51335 45835
rect 51381 45789 51459 45835
rect 51505 45789 51583 45835
rect 51629 45789 51707 45835
rect 51753 45789 51831 45835
rect 51877 45789 51955 45835
rect 52001 45789 52079 45835
rect 52125 45789 52203 45835
rect 52249 45789 52327 45835
rect 52373 45789 52451 45835
rect 52497 45789 52575 45835
rect 52621 45789 52699 45835
rect 52745 45789 52823 45835
rect 52869 45789 52947 45835
rect 52993 45789 53071 45835
rect 53117 45789 53195 45835
rect 53241 45789 53319 45835
rect 53365 45789 53443 45835
rect 53489 45789 53567 45835
rect 53613 45789 53691 45835
rect 53737 45789 53815 45835
rect 53861 45789 53939 45835
rect 53985 45789 54063 45835
rect 54109 45789 54187 45835
rect 54233 45789 54311 45835
rect 54357 45789 54435 45835
rect 54481 45789 54559 45835
rect 54605 45789 54683 45835
rect 54729 45789 54807 45835
rect 54853 45789 54931 45835
rect 54977 45789 55055 45835
rect 55101 45789 55179 45835
rect 55225 45789 55303 45835
rect 55349 45789 55427 45835
rect 55473 45789 55551 45835
rect 55597 45789 55675 45835
rect 55721 45789 55799 45835
rect 55845 45789 55923 45835
rect 55969 45789 56047 45835
rect 56093 45789 56171 45835
rect 56217 45789 56295 45835
rect 56341 45789 56419 45835
rect 56465 45789 56543 45835
rect 56589 45789 56667 45835
rect 56713 45789 56791 45835
rect 56837 45789 56915 45835
rect 56961 45789 57039 45835
rect 57085 45789 57163 45835
rect 57209 45789 57287 45835
rect 57333 45789 57411 45835
rect 57457 45789 57535 45835
rect 57581 45789 57659 45835
rect 57705 45789 57783 45835
rect 57829 45789 57907 45835
rect 57953 45789 58031 45835
rect 58077 45789 58155 45835
rect 58201 45789 58279 45835
rect 58325 45789 58403 45835
rect 58449 45789 58527 45835
rect 58573 45789 58651 45835
rect 58697 45789 58775 45835
rect 58821 45789 58899 45835
rect 58945 45789 59023 45835
rect 59069 45789 59147 45835
rect 59193 45789 59271 45835
rect 59317 45789 59395 45835
rect 59441 45789 59519 45835
rect 59565 45789 59643 45835
rect 59689 45789 59767 45835
rect 59813 45789 59891 45835
rect 59937 45789 60015 45835
rect 60061 45789 60139 45835
rect 60185 45789 60263 45835
rect 60309 45789 60387 45835
rect 60433 45789 60511 45835
rect 60557 45789 60635 45835
rect 60681 45789 60759 45835
rect 60805 45789 60883 45835
rect 60929 45789 61007 45835
rect 61053 45789 61131 45835
rect 61177 45789 61255 45835
rect 61301 45789 61379 45835
rect 61425 45789 61503 45835
rect 61549 45789 61627 45835
rect 61673 45789 61751 45835
rect 61797 45789 61875 45835
rect 61921 45789 61999 45835
rect 62045 45789 62123 45835
rect 62169 45789 62247 45835
rect 62293 45789 62371 45835
rect 62417 45789 62495 45835
rect 62541 45789 62619 45835
rect 62665 45789 62743 45835
rect 62789 45789 62867 45835
rect 62913 45789 62991 45835
rect 63037 45789 63115 45835
rect 63161 45789 63239 45835
rect 63285 45789 63363 45835
rect 63409 45789 63487 45835
rect 63533 45789 63611 45835
rect 63657 45789 63735 45835
rect 63781 45789 63859 45835
rect 63905 45789 63983 45835
rect 64029 45789 64107 45835
rect 64153 45789 64231 45835
rect 64277 45789 64355 45835
rect 64401 45789 64479 45835
rect 64525 45789 64603 45835
rect 64649 45789 64727 45835
rect 64773 45789 64851 45835
rect 64897 45789 64975 45835
rect 65021 45789 65099 45835
rect 65145 45789 65223 45835
rect 65269 45789 65347 45835
rect 65393 45789 65471 45835
rect 65517 45789 65595 45835
rect 65641 45789 65719 45835
rect 65765 45789 65843 45835
rect 65889 45789 65967 45835
rect 66013 45789 66091 45835
rect 66137 45789 66215 45835
rect 66261 45789 66339 45835
rect 66385 45789 66463 45835
rect 66509 45789 66587 45835
rect 66633 45789 66711 45835
rect 66757 45789 66835 45835
rect 66881 45789 66959 45835
rect 67005 45789 67083 45835
rect 67129 45789 67207 45835
rect 67253 45789 67331 45835
rect 67377 45789 67455 45835
rect 67501 45789 67579 45835
rect 67625 45789 67703 45835
rect 67749 45789 67827 45835
rect 67873 45789 67951 45835
rect 67997 45789 68075 45835
rect 68121 45789 68199 45835
rect 68245 45789 68323 45835
rect 68369 45789 68447 45835
rect 68493 45789 68571 45835
rect 68617 45789 68695 45835
rect 68741 45789 68819 45835
rect 68865 45789 68943 45835
rect 68989 45789 69067 45835
rect 69113 45789 69191 45835
rect 69237 45789 69315 45835
rect 69361 45789 69439 45835
rect 69485 45789 69563 45835
rect 69609 45789 69687 45835
rect 69733 45789 69811 45835
rect 69857 45789 69935 45835
rect 69981 45789 70059 45835
rect 70105 45789 70183 45835
rect 70229 45789 70307 45835
rect 70353 45789 70431 45835
rect 70477 45789 70555 45835
rect 70601 45789 70679 45835
rect 70725 45789 70803 45835
rect 70849 45789 70927 45835
rect 70973 45789 71051 45835
rect 71097 45789 71175 45835
rect 71221 45789 71299 45835
rect 71345 45789 71423 45835
rect 71469 45789 71547 45835
rect 71593 45789 71671 45835
rect 71717 45789 71795 45835
rect 71841 45789 71919 45835
rect 71965 45789 72043 45835
rect 72089 45789 72167 45835
rect 72213 45789 72291 45835
rect 72337 45789 72415 45835
rect 72461 45789 72539 45835
rect 72585 45789 72663 45835
rect 72709 45789 72787 45835
rect 72833 45789 72911 45835
rect 72957 45789 73035 45835
rect 73081 45789 73159 45835
rect 73205 45789 73283 45835
rect 73329 45789 73407 45835
rect 73453 45789 73531 45835
rect 73577 45789 73655 45835
rect 73701 45789 73779 45835
rect 73825 45789 73903 45835
rect 73949 45789 74027 45835
rect 74073 45789 74151 45835
rect 74197 45789 74275 45835
rect 74321 45789 74399 45835
rect 74445 45789 74523 45835
rect 74569 45789 74647 45835
rect 74693 45789 74771 45835
rect 74817 45789 74895 45835
rect 74941 45789 75019 45835
rect 75065 45789 75143 45835
rect 75189 45789 75267 45835
rect 75313 45789 75391 45835
rect 75437 45789 75515 45835
rect 75561 45789 75639 45835
rect 75685 45789 75763 45835
rect 75809 45789 75887 45835
rect 75933 45789 76011 45835
rect 76057 45789 76135 45835
rect 76181 45789 76259 45835
rect 76305 45789 76383 45835
rect 76429 45789 76507 45835
rect 76553 45789 76631 45835
rect 76677 45789 76755 45835
rect 76801 45789 76879 45835
rect 76925 45789 77003 45835
rect 77049 45789 77127 45835
rect 77173 45789 77251 45835
rect 77297 45789 77375 45835
rect 77421 45789 77499 45835
rect 77545 45789 77623 45835
rect 77669 45789 77747 45835
rect 77793 45789 77871 45835
rect 77917 45789 77995 45835
rect 78041 45789 78119 45835
rect 78165 45789 78243 45835
rect 78289 45789 78367 45835
rect 78413 45789 78491 45835
rect 78537 45789 78615 45835
rect 78661 45789 78739 45835
rect 78785 45789 78863 45835
rect 78909 45789 78987 45835
rect 79033 45789 79111 45835
rect 79157 45789 79235 45835
rect 79281 45789 79359 45835
rect 79405 45789 79483 45835
rect 79529 45789 79607 45835
rect 79653 45789 79731 45835
rect 79777 45789 79855 45835
rect 79901 45789 79979 45835
rect 80025 45789 80103 45835
rect 80149 45789 80227 45835
rect 80273 45789 80351 45835
rect 80397 45789 80475 45835
rect 80521 45789 80599 45835
rect 80645 45789 80723 45835
rect 80769 45789 80847 45835
rect 80893 45789 80971 45835
rect 81017 45789 81095 45835
rect 81141 45789 81219 45835
rect 81265 45789 81343 45835
rect 81389 45789 81467 45835
rect 81513 45789 81591 45835
rect 81637 45789 81715 45835
rect 81761 45789 81839 45835
rect 81885 45789 81963 45835
rect 82009 45789 82087 45835
rect 82133 45789 82211 45835
rect 82257 45789 82335 45835
rect 82381 45789 82459 45835
rect 82505 45789 82583 45835
rect 82629 45789 82707 45835
rect 82753 45789 82831 45835
rect 82877 45789 82955 45835
rect 83001 45789 83079 45835
rect 83125 45789 83203 45835
rect 83249 45789 83327 45835
rect 83373 45789 83451 45835
rect 83497 45789 83575 45835
rect 83621 45789 83699 45835
rect 83745 45789 83823 45835
rect 83869 45789 83947 45835
rect 83993 45789 84071 45835
rect 84117 45789 84195 45835
rect 84241 45789 84319 45835
rect 84365 45789 84443 45835
rect 84489 45789 84567 45835
rect 84613 45789 84691 45835
rect 84737 45789 84815 45835
rect 84861 45789 84939 45835
rect 84985 45789 85063 45835
rect 85109 45789 85187 45835
rect 85233 45789 85311 45835
rect 85357 45789 85435 45835
rect 85481 45789 85559 45835
rect 85605 45789 85683 45835
rect 85729 45789 85807 45835
rect 85853 45789 85931 45835
rect 85977 45789 86090 45835
rect 282 45711 86090 45789
rect 282 45665 371 45711
rect 417 45665 495 45711
rect 541 45665 619 45711
rect 665 45665 743 45711
rect 789 45665 867 45711
rect 913 45665 991 45711
rect 1037 45665 1115 45711
rect 1161 45665 1239 45711
rect 1285 45665 1363 45711
rect 1409 45665 1487 45711
rect 1533 45665 1611 45711
rect 1657 45665 1735 45711
rect 1781 45665 1859 45711
rect 1905 45665 1983 45711
rect 2029 45665 2107 45711
rect 2153 45665 2231 45711
rect 2277 45665 2355 45711
rect 2401 45665 2479 45711
rect 2525 45665 2603 45711
rect 2649 45665 2727 45711
rect 2773 45665 2851 45711
rect 2897 45665 2975 45711
rect 3021 45665 3099 45711
rect 3145 45665 3223 45711
rect 3269 45665 3347 45711
rect 3393 45665 3471 45711
rect 3517 45665 3595 45711
rect 3641 45665 3719 45711
rect 3765 45665 3843 45711
rect 3889 45665 3967 45711
rect 4013 45665 4091 45711
rect 4137 45665 4215 45711
rect 4261 45665 4339 45711
rect 4385 45665 4463 45711
rect 4509 45665 4587 45711
rect 4633 45665 4711 45711
rect 4757 45665 4835 45711
rect 4881 45665 4959 45711
rect 5005 45665 5083 45711
rect 5129 45665 5207 45711
rect 5253 45665 5331 45711
rect 5377 45665 5455 45711
rect 5501 45665 5579 45711
rect 5625 45665 5703 45711
rect 5749 45665 5827 45711
rect 5873 45665 5951 45711
rect 5997 45665 6075 45711
rect 6121 45665 6199 45711
rect 6245 45665 6323 45711
rect 6369 45665 6447 45711
rect 6493 45665 6571 45711
rect 6617 45665 6695 45711
rect 6741 45665 6819 45711
rect 6865 45665 6943 45711
rect 6989 45665 7067 45711
rect 7113 45665 7191 45711
rect 7237 45665 7315 45711
rect 7361 45665 7439 45711
rect 7485 45665 7563 45711
rect 7609 45665 7687 45711
rect 7733 45665 7811 45711
rect 7857 45665 7935 45711
rect 7981 45665 8059 45711
rect 8105 45665 8183 45711
rect 8229 45665 8307 45711
rect 8353 45665 8431 45711
rect 8477 45665 8555 45711
rect 8601 45665 8679 45711
rect 8725 45665 8803 45711
rect 8849 45665 8927 45711
rect 8973 45665 9051 45711
rect 9097 45665 9175 45711
rect 9221 45665 9299 45711
rect 9345 45665 9423 45711
rect 9469 45665 9547 45711
rect 9593 45665 9671 45711
rect 9717 45665 9795 45711
rect 9841 45665 9919 45711
rect 9965 45665 10043 45711
rect 10089 45665 10167 45711
rect 10213 45665 10291 45711
rect 10337 45665 10415 45711
rect 10461 45665 10539 45711
rect 10585 45665 10663 45711
rect 10709 45665 10787 45711
rect 10833 45665 10911 45711
rect 10957 45665 11035 45711
rect 11081 45665 11159 45711
rect 11205 45665 11283 45711
rect 11329 45665 11407 45711
rect 11453 45665 11531 45711
rect 11577 45665 11655 45711
rect 11701 45665 11779 45711
rect 11825 45665 11903 45711
rect 11949 45665 12027 45711
rect 12073 45665 12151 45711
rect 12197 45665 12275 45711
rect 12321 45665 12399 45711
rect 12445 45665 12523 45711
rect 12569 45665 12647 45711
rect 12693 45665 12771 45711
rect 12817 45665 12895 45711
rect 12941 45665 13019 45711
rect 13065 45665 13143 45711
rect 13189 45665 13267 45711
rect 13313 45665 13391 45711
rect 13437 45665 13515 45711
rect 13561 45665 13639 45711
rect 13685 45665 13763 45711
rect 13809 45665 13887 45711
rect 13933 45665 14011 45711
rect 14057 45665 14135 45711
rect 14181 45665 14259 45711
rect 14305 45665 14383 45711
rect 14429 45665 14507 45711
rect 14553 45665 14631 45711
rect 14677 45665 14755 45711
rect 14801 45665 14879 45711
rect 14925 45665 15003 45711
rect 15049 45665 15127 45711
rect 15173 45665 15251 45711
rect 15297 45665 15375 45711
rect 15421 45665 15499 45711
rect 15545 45665 15623 45711
rect 15669 45665 15747 45711
rect 15793 45665 15871 45711
rect 15917 45665 15995 45711
rect 16041 45665 16119 45711
rect 16165 45665 16243 45711
rect 16289 45665 16367 45711
rect 16413 45665 16491 45711
rect 16537 45665 16615 45711
rect 16661 45665 16739 45711
rect 16785 45665 16863 45711
rect 16909 45665 16987 45711
rect 17033 45665 17111 45711
rect 17157 45665 17235 45711
rect 17281 45665 17359 45711
rect 17405 45665 17483 45711
rect 17529 45665 17607 45711
rect 17653 45665 17731 45711
rect 17777 45665 17855 45711
rect 17901 45665 17979 45711
rect 18025 45665 18103 45711
rect 18149 45665 18227 45711
rect 18273 45665 18351 45711
rect 18397 45665 18475 45711
rect 18521 45665 18599 45711
rect 18645 45665 18723 45711
rect 18769 45665 18847 45711
rect 18893 45665 18971 45711
rect 19017 45665 19095 45711
rect 19141 45665 19219 45711
rect 19265 45665 19343 45711
rect 19389 45665 19467 45711
rect 19513 45665 19591 45711
rect 19637 45665 19715 45711
rect 19761 45665 19839 45711
rect 19885 45665 19963 45711
rect 20009 45665 20087 45711
rect 20133 45665 20211 45711
rect 20257 45665 20335 45711
rect 20381 45665 20459 45711
rect 20505 45665 20583 45711
rect 20629 45665 20707 45711
rect 20753 45665 20831 45711
rect 20877 45665 20955 45711
rect 21001 45665 21079 45711
rect 21125 45665 21203 45711
rect 21249 45665 21327 45711
rect 21373 45665 21451 45711
rect 21497 45665 21575 45711
rect 21621 45665 21699 45711
rect 21745 45665 21823 45711
rect 21869 45665 21947 45711
rect 21993 45665 22071 45711
rect 22117 45665 22195 45711
rect 22241 45665 22319 45711
rect 22365 45665 22443 45711
rect 22489 45665 22567 45711
rect 22613 45665 22691 45711
rect 22737 45665 22815 45711
rect 22861 45665 22939 45711
rect 22985 45665 23063 45711
rect 23109 45665 23187 45711
rect 23233 45665 23311 45711
rect 23357 45665 23435 45711
rect 23481 45665 23559 45711
rect 23605 45665 23683 45711
rect 23729 45665 23807 45711
rect 23853 45665 23931 45711
rect 23977 45665 24055 45711
rect 24101 45665 24179 45711
rect 24225 45665 24303 45711
rect 24349 45665 24427 45711
rect 24473 45665 24551 45711
rect 24597 45665 24675 45711
rect 24721 45665 24799 45711
rect 24845 45665 24923 45711
rect 24969 45665 25047 45711
rect 25093 45665 25171 45711
rect 25217 45665 25295 45711
rect 25341 45665 25419 45711
rect 25465 45665 25543 45711
rect 25589 45665 25667 45711
rect 25713 45665 25791 45711
rect 25837 45665 25915 45711
rect 25961 45665 26039 45711
rect 26085 45665 26163 45711
rect 26209 45665 26287 45711
rect 26333 45665 26411 45711
rect 26457 45665 26535 45711
rect 26581 45665 26659 45711
rect 26705 45665 26783 45711
rect 26829 45665 26907 45711
rect 26953 45665 27031 45711
rect 27077 45665 27155 45711
rect 27201 45665 27279 45711
rect 27325 45665 27403 45711
rect 27449 45665 27527 45711
rect 27573 45665 27651 45711
rect 27697 45665 27775 45711
rect 27821 45665 27899 45711
rect 27945 45665 28023 45711
rect 28069 45665 28147 45711
rect 28193 45665 28271 45711
rect 28317 45665 28395 45711
rect 28441 45665 28519 45711
rect 28565 45665 28643 45711
rect 28689 45665 28767 45711
rect 28813 45665 28891 45711
rect 28937 45665 29015 45711
rect 29061 45665 29139 45711
rect 29185 45665 29263 45711
rect 29309 45665 29387 45711
rect 29433 45665 29511 45711
rect 29557 45665 29635 45711
rect 29681 45665 29759 45711
rect 29805 45665 29883 45711
rect 29929 45665 30007 45711
rect 30053 45665 30131 45711
rect 30177 45665 30255 45711
rect 30301 45665 30379 45711
rect 30425 45665 30503 45711
rect 30549 45665 30627 45711
rect 30673 45665 30751 45711
rect 30797 45665 30875 45711
rect 30921 45665 30999 45711
rect 31045 45665 31123 45711
rect 31169 45665 31247 45711
rect 31293 45665 31371 45711
rect 31417 45665 31495 45711
rect 31541 45665 31619 45711
rect 31665 45665 31743 45711
rect 31789 45665 31867 45711
rect 31913 45665 31991 45711
rect 32037 45665 32115 45711
rect 32161 45665 32239 45711
rect 32285 45665 32363 45711
rect 32409 45665 32487 45711
rect 32533 45665 32611 45711
rect 32657 45665 32735 45711
rect 32781 45665 32859 45711
rect 32905 45665 32983 45711
rect 33029 45665 33107 45711
rect 33153 45665 33231 45711
rect 33277 45665 33355 45711
rect 33401 45665 33479 45711
rect 33525 45665 33603 45711
rect 33649 45665 33727 45711
rect 33773 45665 33851 45711
rect 33897 45665 33975 45711
rect 34021 45665 34099 45711
rect 34145 45665 34223 45711
rect 34269 45665 34347 45711
rect 34393 45665 34471 45711
rect 34517 45665 34595 45711
rect 34641 45665 34719 45711
rect 34765 45665 34843 45711
rect 34889 45665 34967 45711
rect 35013 45665 35091 45711
rect 35137 45665 35215 45711
rect 35261 45665 35339 45711
rect 35385 45665 35463 45711
rect 35509 45665 35587 45711
rect 35633 45665 35711 45711
rect 35757 45665 35835 45711
rect 35881 45665 35959 45711
rect 36005 45665 36083 45711
rect 36129 45665 36207 45711
rect 36253 45665 36331 45711
rect 36377 45665 36455 45711
rect 36501 45665 36579 45711
rect 36625 45665 36703 45711
rect 36749 45665 36827 45711
rect 36873 45665 36951 45711
rect 36997 45665 37075 45711
rect 37121 45665 37199 45711
rect 37245 45665 37323 45711
rect 37369 45665 37447 45711
rect 37493 45665 37571 45711
rect 37617 45665 37695 45711
rect 37741 45665 37819 45711
rect 37865 45665 37943 45711
rect 37989 45665 38067 45711
rect 38113 45665 38191 45711
rect 38237 45665 38315 45711
rect 38361 45665 38439 45711
rect 38485 45665 38563 45711
rect 38609 45665 38687 45711
rect 38733 45665 38811 45711
rect 38857 45665 38935 45711
rect 38981 45665 39059 45711
rect 39105 45665 39183 45711
rect 39229 45665 39307 45711
rect 39353 45665 39431 45711
rect 39477 45665 39555 45711
rect 39601 45665 39679 45711
rect 39725 45665 39803 45711
rect 39849 45665 39927 45711
rect 39973 45665 40051 45711
rect 40097 45665 40175 45711
rect 40221 45665 40299 45711
rect 40345 45665 40423 45711
rect 40469 45665 40547 45711
rect 40593 45665 40671 45711
rect 40717 45665 40795 45711
rect 40841 45665 40919 45711
rect 40965 45665 41043 45711
rect 41089 45665 41167 45711
rect 41213 45665 41291 45711
rect 41337 45665 41415 45711
rect 41461 45665 41539 45711
rect 41585 45665 41663 45711
rect 41709 45665 41787 45711
rect 41833 45665 41911 45711
rect 41957 45665 42035 45711
rect 42081 45665 42159 45711
rect 42205 45665 42283 45711
rect 42329 45665 42407 45711
rect 42453 45665 42531 45711
rect 42577 45665 42655 45711
rect 42701 45665 42779 45711
rect 42825 45665 42903 45711
rect 42949 45665 43027 45711
rect 43073 45665 43151 45711
rect 43197 45665 43275 45711
rect 43321 45665 43399 45711
rect 43445 45665 43523 45711
rect 43569 45665 43647 45711
rect 43693 45665 43771 45711
rect 43817 45665 43895 45711
rect 43941 45665 44019 45711
rect 44065 45665 44143 45711
rect 44189 45665 44267 45711
rect 44313 45665 44391 45711
rect 44437 45665 44515 45711
rect 44561 45665 44639 45711
rect 44685 45665 44763 45711
rect 44809 45665 44887 45711
rect 44933 45665 45011 45711
rect 45057 45665 45135 45711
rect 45181 45665 45259 45711
rect 45305 45665 45383 45711
rect 45429 45665 45507 45711
rect 45553 45665 45631 45711
rect 45677 45665 45755 45711
rect 45801 45665 45879 45711
rect 45925 45665 46003 45711
rect 46049 45665 46127 45711
rect 46173 45665 46251 45711
rect 46297 45665 46375 45711
rect 46421 45665 46499 45711
rect 46545 45665 46623 45711
rect 46669 45665 46747 45711
rect 46793 45665 46871 45711
rect 46917 45665 46995 45711
rect 47041 45665 47119 45711
rect 47165 45665 47243 45711
rect 47289 45665 47367 45711
rect 47413 45665 47491 45711
rect 47537 45665 47615 45711
rect 47661 45665 47739 45711
rect 47785 45665 47863 45711
rect 47909 45665 47987 45711
rect 48033 45665 48111 45711
rect 48157 45665 48235 45711
rect 48281 45665 48359 45711
rect 48405 45665 48483 45711
rect 48529 45665 48607 45711
rect 48653 45665 48731 45711
rect 48777 45665 48855 45711
rect 48901 45665 48979 45711
rect 49025 45665 49103 45711
rect 49149 45665 49227 45711
rect 49273 45665 49351 45711
rect 49397 45665 49475 45711
rect 49521 45665 49599 45711
rect 49645 45665 49723 45711
rect 49769 45665 49847 45711
rect 49893 45665 49971 45711
rect 50017 45665 50095 45711
rect 50141 45665 50219 45711
rect 50265 45665 50343 45711
rect 50389 45665 50467 45711
rect 50513 45665 50591 45711
rect 50637 45665 50715 45711
rect 50761 45665 50839 45711
rect 50885 45665 50963 45711
rect 51009 45665 51087 45711
rect 51133 45665 51211 45711
rect 51257 45665 51335 45711
rect 51381 45665 51459 45711
rect 51505 45665 51583 45711
rect 51629 45665 51707 45711
rect 51753 45665 51831 45711
rect 51877 45665 51955 45711
rect 52001 45665 52079 45711
rect 52125 45665 52203 45711
rect 52249 45665 52327 45711
rect 52373 45665 52451 45711
rect 52497 45665 52575 45711
rect 52621 45665 52699 45711
rect 52745 45665 52823 45711
rect 52869 45665 52947 45711
rect 52993 45665 53071 45711
rect 53117 45665 53195 45711
rect 53241 45665 53319 45711
rect 53365 45665 53443 45711
rect 53489 45665 53567 45711
rect 53613 45665 53691 45711
rect 53737 45665 53815 45711
rect 53861 45665 53939 45711
rect 53985 45665 54063 45711
rect 54109 45665 54187 45711
rect 54233 45665 54311 45711
rect 54357 45665 54435 45711
rect 54481 45665 54559 45711
rect 54605 45665 54683 45711
rect 54729 45665 54807 45711
rect 54853 45665 54931 45711
rect 54977 45665 55055 45711
rect 55101 45665 55179 45711
rect 55225 45665 55303 45711
rect 55349 45665 55427 45711
rect 55473 45665 55551 45711
rect 55597 45665 55675 45711
rect 55721 45665 55799 45711
rect 55845 45665 55923 45711
rect 55969 45665 56047 45711
rect 56093 45665 56171 45711
rect 56217 45665 56295 45711
rect 56341 45665 56419 45711
rect 56465 45665 56543 45711
rect 56589 45665 56667 45711
rect 56713 45665 56791 45711
rect 56837 45665 56915 45711
rect 56961 45665 57039 45711
rect 57085 45665 57163 45711
rect 57209 45665 57287 45711
rect 57333 45665 57411 45711
rect 57457 45665 57535 45711
rect 57581 45665 57659 45711
rect 57705 45665 57783 45711
rect 57829 45665 57907 45711
rect 57953 45665 58031 45711
rect 58077 45665 58155 45711
rect 58201 45665 58279 45711
rect 58325 45665 58403 45711
rect 58449 45665 58527 45711
rect 58573 45665 58651 45711
rect 58697 45665 58775 45711
rect 58821 45665 58899 45711
rect 58945 45665 59023 45711
rect 59069 45665 59147 45711
rect 59193 45665 59271 45711
rect 59317 45665 59395 45711
rect 59441 45665 59519 45711
rect 59565 45665 59643 45711
rect 59689 45665 59767 45711
rect 59813 45665 59891 45711
rect 59937 45665 60015 45711
rect 60061 45665 60139 45711
rect 60185 45665 60263 45711
rect 60309 45665 60387 45711
rect 60433 45665 60511 45711
rect 60557 45665 60635 45711
rect 60681 45665 60759 45711
rect 60805 45665 60883 45711
rect 60929 45665 61007 45711
rect 61053 45665 61131 45711
rect 61177 45665 61255 45711
rect 61301 45665 61379 45711
rect 61425 45665 61503 45711
rect 61549 45665 61627 45711
rect 61673 45665 61751 45711
rect 61797 45665 61875 45711
rect 61921 45665 61999 45711
rect 62045 45665 62123 45711
rect 62169 45665 62247 45711
rect 62293 45665 62371 45711
rect 62417 45665 62495 45711
rect 62541 45665 62619 45711
rect 62665 45665 62743 45711
rect 62789 45665 62867 45711
rect 62913 45665 62991 45711
rect 63037 45665 63115 45711
rect 63161 45665 63239 45711
rect 63285 45665 63363 45711
rect 63409 45665 63487 45711
rect 63533 45665 63611 45711
rect 63657 45665 63735 45711
rect 63781 45665 63859 45711
rect 63905 45665 63983 45711
rect 64029 45665 64107 45711
rect 64153 45665 64231 45711
rect 64277 45665 64355 45711
rect 64401 45665 64479 45711
rect 64525 45665 64603 45711
rect 64649 45665 64727 45711
rect 64773 45665 64851 45711
rect 64897 45665 64975 45711
rect 65021 45665 65099 45711
rect 65145 45665 65223 45711
rect 65269 45665 65347 45711
rect 65393 45665 65471 45711
rect 65517 45665 65595 45711
rect 65641 45665 65719 45711
rect 65765 45665 65843 45711
rect 65889 45665 65967 45711
rect 66013 45665 66091 45711
rect 66137 45665 66215 45711
rect 66261 45665 66339 45711
rect 66385 45665 66463 45711
rect 66509 45665 66587 45711
rect 66633 45665 66711 45711
rect 66757 45665 66835 45711
rect 66881 45665 66959 45711
rect 67005 45665 67083 45711
rect 67129 45665 67207 45711
rect 67253 45665 67331 45711
rect 67377 45665 67455 45711
rect 67501 45665 67579 45711
rect 67625 45665 67703 45711
rect 67749 45665 67827 45711
rect 67873 45665 67951 45711
rect 67997 45665 68075 45711
rect 68121 45665 68199 45711
rect 68245 45665 68323 45711
rect 68369 45665 68447 45711
rect 68493 45665 68571 45711
rect 68617 45665 68695 45711
rect 68741 45665 68819 45711
rect 68865 45665 68943 45711
rect 68989 45665 69067 45711
rect 69113 45665 69191 45711
rect 69237 45665 69315 45711
rect 69361 45665 69439 45711
rect 69485 45665 69563 45711
rect 69609 45665 69687 45711
rect 69733 45665 69811 45711
rect 69857 45665 69935 45711
rect 69981 45665 70059 45711
rect 70105 45665 70183 45711
rect 70229 45665 70307 45711
rect 70353 45665 70431 45711
rect 70477 45665 70555 45711
rect 70601 45665 70679 45711
rect 70725 45665 70803 45711
rect 70849 45665 70927 45711
rect 70973 45665 71051 45711
rect 71097 45665 71175 45711
rect 71221 45665 71299 45711
rect 71345 45665 71423 45711
rect 71469 45665 71547 45711
rect 71593 45665 71671 45711
rect 71717 45665 71795 45711
rect 71841 45665 71919 45711
rect 71965 45665 72043 45711
rect 72089 45665 72167 45711
rect 72213 45665 72291 45711
rect 72337 45665 72415 45711
rect 72461 45665 72539 45711
rect 72585 45665 72663 45711
rect 72709 45665 72787 45711
rect 72833 45665 72911 45711
rect 72957 45665 73035 45711
rect 73081 45665 73159 45711
rect 73205 45665 73283 45711
rect 73329 45665 73407 45711
rect 73453 45665 73531 45711
rect 73577 45665 73655 45711
rect 73701 45665 73779 45711
rect 73825 45665 73903 45711
rect 73949 45665 74027 45711
rect 74073 45665 74151 45711
rect 74197 45665 74275 45711
rect 74321 45665 74399 45711
rect 74445 45665 74523 45711
rect 74569 45665 74647 45711
rect 74693 45665 74771 45711
rect 74817 45665 74895 45711
rect 74941 45665 75019 45711
rect 75065 45665 75143 45711
rect 75189 45665 75267 45711
rect 75313 45665 75391 45711
rect 75437 45665 75515 45711
rect 75561 45665 75639 45711
rect 75685 45665 75763 45711
rect 75809 45665 75887 45711
rect 75933 45665 76011 45711
rect 76057 45665 76135 45711
rect 76181 45665 76259 45711
rect 76305 45665 76383 45711
rect 76429 45665 76507 45711
rect 76553 45665 76631 45711
rect 76677 45665 76755 45711
rect 76801 45665 76879 45711
rect 76925 45665 77003 45711
rect 77049 45665 77127 45711
rect 77173 45665 77251 45711
rect 77297 45665 77375 45711
rect 77421 45665 77499 45711
rect 77545 45665 77623 45711
rect 77669 45665 77747 45711
rect 77793 45665 77871 45711
rect 77917 45665 77995 45711
rect 78041 45665 78119 45711
rect 78165 45665 78243 45711
rect 78289 45665 78367 45711
rect 78413 45665 78491 45711
rect 78537 45665 78615 45711
rect 78661 45665 78739 45711
rect 78785 45665 78863 45711
rect 78909 45665 78987 45711
rect 79033 45665 79111 45711
rect 79157 45665 79235 45711
rect 79281 45665 79359 45711
rect 79405 45665 79483 45711
rect 79529 45665 79607 45711
rect 79653 45665 79731 45711
rect 79777 45665 79855 45711
rect 79901 45665 79979 45711
rect 80025 45665 80103 45711
rect 80149 45665 80227 45711
rect 80273 45665 80351 45711
rect 80397 45665 80475 45711
rect 80521 45665 80599 45711
rect 80645 45665 80723 45711
rect 80769 45665 80847 45711
rect 80893 45665 80971 45711
rect 81017 45665 81095 45711
rect 81141 45665 81219 45711
rect 81265 45665 81343 45711
rect 81389 45665 81467 45711
rect 81513 45665 81591 45711
rect 81637 45665 81715 45711
rect 81761 45665 81839 45711
rect 81885 45665 81963 45711
rect 82009 45665 82087 45711
rect 82133 45665 82211 45711
rect 82257 45665 82335 45711
rect 82381 45665 82459 45711
rect 82505 45665 82583 45711
rect 82629 45665 82707 45711
rect 82753 45665 82831 45711
rect 82877 45665 82955 45711
rect 83001 45665 83079 45711
rect 83125 45665 83203 45711
rect 83249 45665 83327 45711
rect 83373 45665 83451 45711
rect 83497 45665 83575 45711
rect 83621 45665 83699 45711
rect 83745 45665 83823 45711
rect 83869 45665 83947 45711
rect 83993 45665 84071 45711
rect 84117 45665 84195 45711
rect 84241 45665 84319 45711
rect 84365 45665 84443 45711
rect 84489 45665 84567 45711
rect 84613 45665 84691 45711
rect 84737 45665 84815 45711
rect 84861 45665 84939 45711
rect 84985 45665 85063 45711
rect 85109 45665 85187 45711
rect 85233 45665 85311 45711
rect 85357 45665 85435 45711
rect 85481 45665 85559 45711
rect 85605 45665 85683 45711
rect 85729 45665 85807 45711
rect 85853 45665 85931 45711
rect 85977 45665 86090 45711
rect 282 45563 86090 45665
rect 282 1117 371 45563
rect 717 45294 27498 45563
rect 717 1282 1282 45294
rect 25313 44338 26040 45294
rect 25313 44286 25337 44338
rect 25389 44286 25461 44338
rect 25513 44286 25585 44338
rect 25637 44286 25709 44338
rect 25761 44286 25833 44338
rect 25885 44286 25957 44338
rect 26009 44286 26040 44338
rect 25313 44214 26040 44286
rect 25313 44162 25337 44214
rect 25389 44162 25461 44214
rect 25513 44162 25585 44214
rect 25637 44162 25709 44214
rect 25761 44162 25833 44214
rect 25885 44162 25957 44214
rect 26009 44162 26040 44214
rect 25313 44076 26040 44162
rect 25388 34972 25960 34984
rect 25388 34920 25400 34972
rect 25452 34920 25524 34972
rect 25576 34920 25648 34972
rect 25700 34920 25772 34972
rect 25824 34920 25896 34972
rect 25948 34920 25960 34972
rect 25388 34909 25960 34920
rect 27387 34938 27498 45294
rect 27744 45463 85733 45563
rect 27744 45442 57380 45463
rect 27744 44253 27846 45442
rect 28492 45294 56632 45442
rect 28492 44253 29196 45294
rect 34227 44366 35024 45294
rect 33001 44309 35024 44366
rect 27744 44201 27790 44253
rect 27842 44201 27846 44253
rect 28492 44201 28634 44253
rect 28686 44201 28845 44253
rect 28897 44201 29056 44253
rect 29108 44201 29196 44253
rect 27744 42453 27846 44201
rect 28492 44122 29196 44201
rect 29283 44253 30365 44294
rect 29283 44250 29582 44253
rect 29283 44204 29317 44250
rect 29363 44204 29478 44250
rect 29524 44204 29582 44250
rect 29283 44201 29582 44204
rect 29634 44250 29793 44253
rect 29845 44250 30005 44253
rect 29634 44204 29638 44250
rect 29684 44204 29793 44250
rect 29845 44204 29959 44250
rect 29634 44201 29793 44204
rect 29845 44201 30005 44204
rect 30057 44250 30216 44253
rect 30057 44204 30121 44250
rect 30167 44204 30216 44250
rect 30057 44201 30216 44204
rect 30268 44250 30365 44253
rect 30268 44204 30284 44250
rect 30330 44204 30365 44250
rect 30268 44201 30365 44204
rect 29283 44161 30365 44201
rect 30583 44253 32694 44294
rect 30583 44201 30807 44253
rect 30859 44236 31018 44253
rect 31070 44236 31229 44253
rect 30583 44190 30854 44201
rect 30900 44190 31012 44236
rect 31070 44201 31170 44236
rect 31058 44190 31170 44201
rect 31216 44201 31229 44236
rect 31281 44236 31440 44253
rect 31492 44236 31651 44253
rect 31703 44236 31861 44253
rect 31281 44201 31328 44236
rect 31216 44190 31328 44201
rect 31374 44201 31440 44236
rect 31374 44190 31487 44201
rect 31533 44190 31645 44236
rect 31703 44201 31803 44236
rect 31691 44190 31803 44201
rect 31849 44201 31861 44236
rect 31913 44236 32072 44253
rect 32124 44236 32283 44253
rect 32335 44236 32494 44253
rect 31913 44201 31961 44236
rect 31849 44190 31961 44201
rect 32007 44201 32072 44236
rect 32007 44190 32119 44201
rect 32165 44190 32277 44236
rect 32335 44201 32435 44236
rect 32323 44190 32435 44201
rect 32481 44201 32494 44236
rect 32546 44236 32694 44253
rect 32546 44201 32593 44236
rect 32481 44190 32593 44201
rect 32639 44190 32694 44236
rect 29544 44160 30306 44161
rect 28492 44076 28810 44122
rect 28856 44076 29196 44122
rect 28492 44044 29196 44076
rect 28492 43998 29116 44044
rect 29162 43998 29196 44044
rect 28492 43958 29196 43998
rect 28492 43912 28810 43958
rect 28856 43912 29196 43958
rect 28492 43881 29196 43912
rect 28492 43835 29116 43881
rect 29162 43835 29196 43881
rect 28492 43795 29196 43835
rect 28492 43749 28810 43795
rect 28856 43749 29196 43795
rect 28492 43717 29196 43749
rect 28492 43671 29116 43717
rect 29162 43671 29196 43717
rect 28492 43632 29196 43671
rect 28492 43586 28810 43632
rect 28856 43586 29196 43632
rect 28492 43554 29196 43586
rect 28492 43508 29116 43554
rect 29162 43508 29196 43554
rect 28492 43468 29196 43508
rect 28492 43422 28810 43468
rect 28856 43422 29196 43468
rect 28492 43266 29196 43422
rect 30583 44122 32694 44190
rect 30583 44076 30637 44122
rect 30683 44076 32694 44122
rect 30583 44073 32694 44076
rect 30583 44035 30854 44073
rect 30583 43983 30807 44035
rect 30900 44027 31012 44073
rect 31058 44035 31170 44073
rect 31070 44027 31170 44035
rect 31216 44035 31328 44073
rect 31216 44027 31229 44035
rect 30859 43983 31018 44027
rect 31070 43983 31229 44027
rect 31281 44027 31328 44035
rect 31374 44035 31487 44073
rect 31374 44027 31440 44035
rect 31533 44027 31645 44073
rect 31691 44035 31803 44073
rect 31703 44027 31803 44035
rect 31849 44035 31961 44073
rect 31849 44027 31861 44035
rect 31281 43983 31440 44027
rect 31492 43983 31651 44027
rect 31703 43983 31861 44027
rect 31913 44027 31961 44035
rect 32007 44035 32119 44073
rect 32007 44027 32072 44035
rect 32165 44027 32277 44073
rect 32323 44035 32435 44073
rect 32335 44027 32435 44035
rect 32481 44035 32593 44073
rect 32481 44027 32494 44035
rect 31913 43983 32072 44027
rect 32124 43983 32283 44027
rect 32335 43983 32494 44027
rect 32546 44027 32593 44035
rect 32639 44027 32694 44073
rect 32546 43983 32694 44027
rect 30583 43958 32694 43983
rect 30583 43912 30637 43958
rect 30683 43912 32694 43958
rect 33001 44263 33044 44309
rect 33090 44263 33202 44309
rect 33248 44263 33360 44309
rect 33406 44263 33518 44309
rect 33564 44263 33677 44309
rect 33723 44263 33835 44309
rect 33881 44263 33993 44309
rect 34039 44263 34151 44309
rect 34197 44263 34309 44309
rect 34355 44263 34467 44309
rect 34513 44263 34625 44309
rect 34671 44263 34783 44309
rect 34829 44271 35024 44309
rect 40062 44346 40590 45294
rect 43738 44346 44599 45294
rect 50558 44346 51373 45294
rect 40062 44309 41937 44346
rect 34829 44263 35013 44271
rect 33001 44253 35013 44263
rect 33001 44201 34290 44253
rect 34342 44201 34501 44253
rect 34553 44201 34712 44253
rect 34764 44201 34923 44253
rect 34975 44201 35013 44253
rect 35405 44233 36377 44273
rect 35405 44218 35443 44233
rect 35495 44218 35654 44233
rect 35706 44218 35865 44233
rect 35917 44218 36076 44233
rect 36128 44218 36287 44233
rect 36339 44218 36377 44233
rect 40062 44263 40117 44309
rect 40163 44263 40275 44309
rect 40321 44263 40433 44309
rect 40479 44263 40591 44309
rect 40637 44263 40750 44309
rect 40796 44263 40908 44309
rect 40954 44263 41066 44309
rect 41112 44263 41224 44309
rect 41270 44263 41382 44309
rect 41428 44263 41540 44309
rect 41586 44263 41698 44309
rect 41744 44263 41856 44309
rect 41902 44263 41937 44309
rect 40062 44258 41937 44263
rect 33001 44035 35013 44201
rect 35396 44172 35409 44218
rect 37291 44172 37348 44218
rect 37394 44172 37451 44218
rect 37497 44172 37554 44218
rect 37600 44172 37657 44218
rect 37703 44172 37760 44218
rect 37806 44172 37863 44218
rect 37909 44172 37922 44218
rect 40062 44206 40252 44258
rect 40304 44206 40432 44258
rect 40484 44226 41937 44258
rect 42208 44309 43589 44346
rect 42208 44305 42717 44309
rect 42208 44253 42710 44305
rect 42763 44263 42875 44309
rect 42921 44305 43033 44309
rect 42762 44253 42921 44263
rect 42973 44263 43033 44305
rect 43079 44305 43191 44309
rect 43079 44263 43132 44305
rect 42973 44253 43132 44263
rect 43184 44263 43191 44305
rect 43237 44263 43350 44309
rect 43396 44263 43508 44309
rect 43554 44263 43589 44309
rect 43184 44253 43589 44263
rect 42208 44244 43589 44253
rect 40484 44206 40590 44226
rect 35405 44141 36377 44172
rect 38000 44045 38116 44112
rect 33001 43994 34290 44035
rect 33001 43948 33014 43994
rect 33774 43948 33831 43994
rect 33877 43948 33934 43994
rect 33980 43948 34037 43994
rect 34083 43948 34140 43994
rect 34186 43948 34243 43994
rect 34289 43983 34290 43994
rect 34342 43994 34501 44035
rect 34553 43994 34712 44035
rect 34764 43994 34923 44035
rect 34975 43994 35013 44035
rect 35159 43994 35444 44035
rect 34342 43983 34346 43994
rect 34289 43948 34346 43983
rect 34392 43948 34449 43994
rect 34495 43983 34501 43994
rect 34495 43948 34552 43983
rect 34598 43948 34655 43994
rect 34701 43983 34712 43994
rect 34701 43948 34758 43983
rect 34804 43948 34861 43994
rect 34907 43983 34923 43994
rect 34907 43948 34964 43983
rect 35010 43948 35023 43994
rect 35159 43948 35409 43994
rect 37291 43948 37348 43994
rect 37394 43948 37451 43994
rect 37497 43948 37554 43994
rect 37600 43948 37657 43994
rect 37703 43948 37760 43994
rect 37806 43948 37863 43994
rect 37909 43948 37922 43994
rect 34251 43943 35013 43948
rect 30583 43909 32694 43912
rect 30583 43863 30854 43909
rect 30900 43863 31012 43909
rect 31058 43863 31170 43909
rect 31216 43863 31328 43909
rect 31374 43863 31487 43909
rect 31533 43863 31645 43909
rect 31691 43863 31803 43909
rect 31849 43863 31961 43909
rect 32007 43863 32119 43909
rect 32165 43863 32277 43909
rect 32323 43863 32435 43909
rect 32481 43863 32593 43909
rect 32639 43863 32694 43909
rect 30583 43818 32694 43863
rect 30583 43795 30807 43818
rect 30583 43749 30637 43795
rect 30683 43766 30807 43795
rect 30859 43766 31018 43818
rect 31070 43766 31229 43818
rect 31281 43766 31440 43818
rect 31492 43766 31651 43818
rect 31703 43766 31861 43818
rect 31913 43766 32072 43818
rect 32124 43766 32283 43818
rect 32335 43766 32494 43818
rect 32546 43766 32694 43818
rect 35159 43915 35444 43948
rect 33012 43772 33984 43812
rect 35159 43804 35275 43915
rect 38000 43905 38035 44045
rect 38081 43905 38116 44045
rect 39015 44035 39565 44042
rect 39014 44001 39565 44035
rect 39014 43994 39053 44001
rect 39105 43994 39264 44001
rect 39316 43994 39475 44001
rect 39527 43994 39565 44001
rect 40062 44040 40590 44206
rect 42208 44192 42246 44244
rect 42298 44243 42458 44244
rect 42298 44197 42319 44243
rect 42510 44226 43589 44244
rect 43738 44309 44960 44346
rect 43738 44305 44514 44309
rect 43738 44253 43777 44305
rect 43829 44253 43988 44305
rect 44040 44291 44199 44305
rect 44040 44253 44067 44291
rect 43738 44245 44067 44253
rect 44113 44253 44199 44291
rect 44251 44253 44410 44305
rect 44462 44263 44514 44305
rect 44560 44263 44672 44309
rect 44718 44263 44830 44309
rect 44876 44263 44960 44309
rect 50001 44309 52023 44346
rect 56212 44328 56632 45294
rect 48789 44267 49551 44273
rect 44462 44253 44960 44263
rect 44113 44245 44960 44253
rect 42510 44213 43222 44226
rect 42510 44212 42717 44213
rect 43738 44212 44960 44245
rect 42298 44192 42458 44197
rect 42510 44192 42548 44212
rect 42208 44151 42548 44192
rect 40062 43994 40252 44040
rect 40304 43994 40432 44040
rect 40484 43994 40590 44040
rect 44268 43998 44336 44009
rect 38363 43948 38376 43994
rect 38422 43948 38479 43994
rect 38525 43948 38582 43994
rect 38628 43948 38686 43994
rect 38732 43948 38790 43994
rect 38836 43948 38894 43994
rect 38940 43948 38998 43994
rect 39044 43949 39053 43994
rect 39044 43948 39102 43949
rect 39148 43948 39206 43994
rect 39252 43949 39264 43994
rect 39252 43948 39310 43949
rect 39356 43948 39414 43994
rect 39460 43949 39475 43994
rect 39460 43948 39518 43949
rect 39564 43948 39622 43994
rect 39668 43948 39681 43994
rect 40062 43948 40075 43994
rect 40121 43948 40189 43994
rect 40235 43988 40252 43994
rect 40235 43948 40303 43988
rect 40349 43948 40417 43994
rect 40484 43988 40531 43994
rect 40463 43948 40531 43988
rect 40577 43948 40590 43994
rect 40683 43958 40976 43995
rect 39014 43915 39565 43948
rect 39015 43909 39565 43915
rect 33012 43770 33050 43772
rect 33102 43770 33261 43772
rect 33313 43770 33472 43772
rect 33524 43770 33683 43772
rect 33735 43770 33894 43772
rect 33946 43770 33984 43772
rect 34917 43770 35275 43804
rect 35405 43770 36377 43810
rect 38000 43804 38116 43905
rect 40683 43818 40694 43958
rect 40740 43949 40976 43958
rect 41022 43949 41079 43995
rect 41125 43949 41182 43995
rect 41228 43949 41286 43995
rect 41332 43949 41390 43995
rect 41436 43949 41494 43995
rect 41540 43949 41598 43995
rect 41644 43949 41702 43995
rect 41748 43949 41806 43995
rect 41852 43949 41910 43995
rect 41956 43949 42014 43995
rect 42060 43949 42118 43995
rect 42164 43949 42222 43995
rect 42268 43994 42851 43995
rect 44268 43994 44279 43998
rect 42268 43949 42676 43994
rect 40740 43818 40751 43949
rect 42663 43948 42676 43949
rect 42722 43948 42779 43994
rect 42825 43948 42882 43994
rect 42928 43948 42986 43994
rect 43032 43948 43090 43994
rect 43136 43948 43194 43994
rect 43240 43948 43298 43994
rect 43344 43948 43402 43994
rect 43448 43948 43506 43994
rect 43552 43948 43610 43994
rect 43656 43948 43714 43994
rect 43760 43948 43818 43994
rect 43864 43948 43922 43994
rect 43968 43948 44279 43994
rect 44268 43858 44279 43948
rect 44325 43858 44336 43998
rect 44432 43994 44960 44212
rect 44432 43948 44445 43994
rect 44491 43948 44559 43994
rect 44605 43948 44673 43994
rect 44719 43948 44787 43994
rect 44833 43948 44901 43994
rect 44947 43948 44960 43994
rect 45333 44233 49619 44267
rect 45333 44218 48828 44233
rect 48880 44218 49039 44233
rect 49091 44218 49250 44233
rect 49302 44218 49461 44233
rect 49513 44218 49619 44233
rect 50001 44263 50129 44309
rect 50175 44263 50287 44309
rect 50333 44263 50445 44309
rect 50491 44263 50603 44309
rect 50649 44263 50762 44309
rect 50808 44263 50920 44309
rect 50966 44263 51078 44309
rect 51124 44263 51236 44309
rect 51282 44263 51394 44309
rect 51440 44263 51552 44309
rect 51598 44263 51710 44309
rect 51756 44263 51868 44309
rect 51914 44263 52023 44309
rect 50001 44253 52023 44263
rect 45333 44172 47114 44218
rect 48996 44181 49039 44218
rect 48996 44172 49053 44181
rect 49099 44172 49156 44218
rect 49202 44181 49250 44218
rect 49202 44172 49259 44181
rect 49305 44172 49362 44218
rect 49408 44181 49461 44218
rect 49513 44181 49568 44218
rect 49408 44172 49465 44181
rect 49511 44172 49568 44181
rect 49614 44172 49627 44218
rect 50001 44201 50137 44253
rect 50189 44201 50348 44253
rect 50400 44201 50559 44253
rect 50611 44201 50770 44253
rect 50822 44201 52023 44253
rect 45333 44147 49619 44172
rect 45333 43994 46651 44147
rect 48789 44140 49551 44147
rect 45333 43948 45346 43994
rect 45392 43948 45449 43994
rect 45495 43948 45552 43994
rect 45598 43948 45656 43994
rect 45702 43948 45760 43994
rect 45806 43948 45864 43994
rect 45910 43948 45968 43994
rect 46014 43948 46072 43994
rect 46118 43948 46176 43994
rect 46222 43948 46280 43994
rect 46326 43948 46384 43994
rect 46430 43948 46488 43994
rect 46534 43948 46592 43994
rect 46638 43948 46651 43994
rect 46956 44033 47024 44044
rect 44432 43915 44960 43948
rect 44268 43847 44336 43858
rect 46956 43893 46967 44033
rect 47013 43893 47024 44033
rect 50001 44035 52023 44201
rect 50001 43994 50137 44035
rect 50189 43994 50348 44035
rect 50400 43994 50559 44035
rect 50611 43994 50770 44035
rect 50822 43994 52023 44035
rect 47101 43948 47114 43994
rect 48996 43948 49053 43994
rect 49099 43948 49156 43994
rect 49202 43948 49259 43994
rect 49305 43948 49362 43994
rect 49408 43948 49465 43994
rect 49511 43948 49568 43994
rect 49614 43948 49861 43994
rect 46956 43882 47024 43893
rect 40683 43807 40751 43818
rect 38000 43770 40590 43804
rect 40971 43771 42155 43811
rect 46956 43804 47023 43882
rect 30683 43749 32694 43766
rect 30583 43746 32694 43749
rect 30583 43700 30854 43746
rect 30900 43700 31012 43746
rect 31058 43700 31170 43746
rect 31216 43700 31328 43746
rect 31374 43700 31487 43746
rect 31533 43700 31645 43746
rect 31691 43700 31803 43746
rect 31849 43700 31961 43746
rect 32007 43700 32119 43746
rect 32165 43700 32277 43746
rect 32323 43700 32435 43746
rect 32481 43700 32593 43746
rect 32639 43700 32694 43746
rect 33001 43724 33014 43770
rect 33774 43724 33831 43770
rect 33877 43724 33894 43770
rect 33980 43724 34037 43770
rect 34083 43724 34140 43770
rect 34186 43724 34243 43770
rect 34289 43724 34346 43770
rect 34392 43724 34449 43770
rect 34495 43724 34552 43770
rect 34598 43724 34655 43770
rect 34701 43724 34758 43770
rect 34804 43724 34861 43770
rect 34907 43724 34964 43770
rect 35010 43724 35275 43770
rect 35396 43724 35409 43770
rect 37291 43724 37348 43770
rect 37394 43724 37451 43770
rect 37497 43724 37554 43770
rect 37600 43724 37657 43770
rect 37703 43724 37760 43770
rect 37806 43724 37863 43770
rect 37909 43724 37922 43770
rect 38000 43724 38376 43770
rect 38422 43724 38479 43770
rect 38525 43724 38582 43770
rect 38628 43724 38686 43770
rect 38732 43724 38790 43770
rect 38836 43724 38894 43770
rect 38940 43724 38998 43770
rect 39044 43724 39102 43770
rect 39148 43724 39206 43770
rect 39252 43724 39310 43770
rect 39356 43724 39414 43770
rect 39460 43724 39518 43770
rect 39564 43724 39622 43770
rect 39668 43724 40075 43770
rect 40121 43724 40189 43770
rect 40235 43724 40303 43770
rect 40349 43724 40417 43770
rect 40463 43724 40531 43770
rect 40577 43724 40590 43770
rect 40963 43725 40976 43771
rect 41022 43770 41079 43771
rect 41062 43725 41079 43770
rect 41125 43725 41182 43771
rect 41228 43770 41286 43771
rect 41273 43725 41286 43770
rect 41332 43725 41390 43771
rect 41436 43770 41494 43771
rect 41484 43725 41494 43770
rect 41540 43725 41598 43771
rect 41644 43770 41702 43771
rect 41695 43725 41702 43770
rect 41748 43725 41806 43771
rect 41852 43770 41910 43771
rect 41852 43725 41854 43770
rect 30583 43643 32694 43700
rect 33012 43720 33050 43724
rect 33102 43720 33261 43724
rect 33313 43720 33472 43724
rect 33524 43720 33683 43724
rect 33735 43720 33894 43724
rect 33946 43720 33984 43724
rect 33012 43680 33984 43720
rect 34917 43684 35275 43724
rect 35405 43718 35443 43724
rect 35495 43718 35654 43724
rect 35706 43718 35865 43724
rect 35917 43718 36076 43724
rect 36128 43718 36287 43724
rect 36339 43718 36377 43724
rect 35405 43678 36377 43718
rect 38000 43684 40590 43724
rect 40971 43718 41010 43725
rect 41062 43718 41221 43725
rect 41273 43718 41432 43725
rect 41484 43718 41643 43725
rect 41695 43718 41854 43725
rect 41906 43725 41910 43770
rect 41956 43725 42014 43771
rect 42060 43770 42118 43771
rect 42060 43725 42064 43770
rect 41906 43718 42064 43725
rect 42116 43725 42118 43770
rect 42164 43725 42222 43771
rect 42268 43770 42851 43771
rect 44432 43770 47023 43804
rect 48789 43770 49551 43810
rect 49744 43770 49861 43948
rect 50001 43948 50014 43994
rect 50822 43983 50831 43994
rect 50774 43948 50831 43983
rect 50877 43948 50934 43994
rect 50980 43948 51037 43994
rect 51083 43948 51140 43994
rect 51186 43948 51243 43994
rect 51289 43948 51346 43994
rect 51392 43948 51449 43994
rect 51495 43948 51552 43994
rect 51598 43948 51655 43994
rect 51701 43948 51758 43994
rect 51804 43948 51861 43994
rect 51907 43948 51964 43994
rect 52010 43948 52023 43994
rect 50001 43929 52023 43948
rect 52428 44253 54540 44294
rect 52428 44236 52576 44253
rect 52428 44190 52483 44236
rect 52529 44201 52576 44236
rect 52628 44236 52787 44253
rect 52839 44236 52998 44253
rect 53050 44236 53209 44253
rect 52628 44201 52641 44236
rect 52529 44190 52641 44201
rect 52687 44201 52787 44236
rect 52687 44190 52799 44201
rect 52845 44190 52957 44236
rect 53050 44201 53115 44236
rect 53003 44190 53115 44201
rect 53161 44201 53209 44236
rect 53261 44236 53419 44253
rect 53471 44236 53630 44253
rect 53682 44236 53841 44253
rect 53261 44201 53273 44236
rect 53161 44190 53273 44201
rect 53319 44201 53419 44236
rect 53319 44190 53431 44201
rect 53477 44190 53589 44236
rect 53682 44201 53748 44236
rect 53635 44190 53748 44201
rect 53794 44201 53841 44236
rect 53893 44236 54052 44253
rect 54104 44236 54263 44253
rect 53893 44201 53906 44236
rect 53794 44190 53906 44201
rect 53952 44201 54052 44236
rect 53952 44190 54064 44201
rect 54110 44190 54222 44236
rect 54315 44201 54540 44253
rect 54268 44190 54540 44201
rect 52428 44122 54540 44190
rect 54758 44253 55840 44294
rect 54758 44250 54855 44253
rect 54758 44204 54793 44250
rect 54839 44204 54855 44250
rect 54758 44201 54855 44204
rect 54907 44250 55066 44253
rect 54907 44204 54956 44250
rect 55002 44204 55066 44250
rect 54907 44201 55066 44204
rect 55118 44250 55278 44253
rect 55330 44250 55489 44253
rect 55164 44204 55278 44250
rect 55330 44204 55439 44250
rect 55485 44204 55489 44250
rect 55118 44201 55278 44204
rect 55330 44201 55489 44204
rect 55541 44250 55840 44253
rect 55541 44204 55599 44250
rect 55645 44204 55760 44250
rect 55806 44204 55840 44250
rect 55541 44201 55840 44204
rect 54758 44161 55840 44201
rect 55927 44253 56632 44328
rect 57278 44253 57380 45442
rect 55927 44201 56015 44253
rect 56067 44201 56226 44253
rect 56278 44201 56437 44253
rect 56489 44201 56632 44253
rect 57278 44201 57281 44253
rect 57333 44201 57380 44253
rect 54817 44160 55579 44161
rect 52428 44076 54440 44122
rect 54486 44076 54540 44122
rect 52428 44073 54540 44076
rect 52428 44027 52483 44073
rect 52529 44035 52641 44073
rect 52529 44027 52576 44035
rect 52428 43983 52576 44027
rect 52628 44027 52641 44035
rect 52687 44035 52799 44073
rect 52687 44027 52787 44035
rect 52845 44027 52957 44073
rect 53003 44035 53115 44073
rect 53050 44027 53115 44035
rect 53161 44035 53273 44073
rect 53161 44027 53209 44035
rect 52628 43983 52787 44027
rect 52839 43983 52998 44027
rect 53050 43983 53209 44027
rect 53261 44027 53273 44035
rect 53319 44035 53431 44073
rect 53319 44027 53419 44035
rect 53477 44027 53589 44073
rect 53635 44035 53748 44073
rect 53682 44027 53748 44035
rect 53794 44035 53906 44073
rect 53794 44027 53841 44035
rect 53261 43983 53419 44027
rect 53471 43983 53630 44027
rect 53682 43983 53841 44027
rect 53893 44027 53906 44035
rect 53952 44035 54064 44073
rect 53952 44027 54052 44035
rect 54110 44027 54222 44073
rect 54268 44035 54540 44073
rect 53893 43983 54052 44027
rect 54104 43983 54263 44027
rect 54315 43983 54540 44035
rect 52428 43958 54540 43983
rect 52428 43912 54440 43958
rect 54486 43912 54540 43958
rect 52428 43909 54540 43912
rect 52428 43863 52483 43909
rect 52529 43863 52641 43909
rect 52687 43863 52799 43909
rect 52845 43863 52957 43909
rect 53003 43863 53115 43909
rect 53161 43863 53273 43909
rect 53319 43863 53431 43909
rect 53477 43863 53589 43909
rect 53635 43863 53748 43909
rect 53794 43863 53906 43909
rect 53952 43863 54064 43909
rect 54110 43863 54222 43909
rect 54268 43863 54540 43909
rect 52428 43818 54540 43863
rect 51043 43770 52015 43810
rect 42268 43725 42676 43770
rect 42116 43718 42155 43725
rect 42663 43724 42676 43725
rect 42722 43724 42779 43770
rect 42825 43724 42882 43770
rect 42928 43724 42986 43770
rect 43032 43724 43090 43770
rect 43136 43724 43194 43770
rect 43240 43724 43298 43770
rect 43344 43724 43402 43770
rect 43448 43724 43506 43770
rect 43552 43724 43610 43770
rect 43656 43724 43714 43770
rect 43760 43724 43818 43770
rect 43864 43724 43922 43770
rect 43968 43724 43981 43770
rect 44432 43724 44445 43770
rect 44491 43724 44559 43770
rect 44605 43724 44673 43770
rect 44719 43724 44787 43770
rect 44833 43724 44901 43770
rect 44947 43724 45346 43770
rect 45392 43724 45449 43770
rect 45495 43724 45552 43770
rect 45598 43724 45656 43770
rect 45702 43724 45760 43770
rect 45806 43724 45864 43770
rect 45910 43724 45968 43770
rect 46014 43724 46072 43770
rect 46118 43724 46176 43770
rect 46222 43724 46280 43770
rect 46326 43724 46384 43770
rect 46430 43724 46488 43770
rect 46534 43724 46592 43770
rect 46638 43724 47023 43770
rect 47101 43724 47114 43770
rect 48996 43724 49039 43770
rect 49099 43724 49156 43770
rect 49202 43724 49250 43770
rect 49305 43724 49362 43770
rect 49408 43724 49461 43770
rect 49513 43724 49568 43770
rect 49614 43724 49627 43770
rect 49744 43724 50014 43770
rect 50774 43724 50831 43770
rect 50877 43724 50934 43770
rect 50980 43724 51037 43770
rect 51133 43724 51140 43770
rect 51186 43724 51243 43770
rect 51289 43724 51292 43770
rect 40971 43677 42155 43718
rect 44432 43684 47023 43724
rect 48789 43718 48828 43724
rect 48880 43718 49039 43724
rect 49091 43718 49250 43724
rect 49302 43718 49461 43724
rect 49513 43718 49551 43724
rect 48789 43677 49551 43718
rect 51043 43718 51081 43724
rect 51133 43718 51292 43724
rect 51344 43724 51346 43770
rect 51392 43724 51449 43770
rect 51495 43724 51503 43770
rect 51598 43724 51655 43770
rect 51701 43724 51714 43770
rect 51804 43724 51861 43770
rect 51907 43724 51925 43770
rect 52010 43724 52023 43770
rect 52428 43766 52576 43818
rect 52628 43766 52787 43818
rect 52839 43766 52998 43818
rect 53050 43766 53209 43818
rect 53261 43766 53419 43818
rect 53471 43766 53630 43818
rect 53682 43766 53841 43818
rect 53893 43766 54052 43818
rect 54104 43766 54263 43818
rect 54315 43795 54540 43818
rect 54315 43766 54440 43795
rect 52428 43749 54440 43766
rect 54486 43749 54540 43795
rect 52428 43746 54540 43749
rect 51344 43718 51503 43724
rect 51555 43718 51714 43724
rect 51766 43718 51925 43724
rect 51977 43718 52015 43724
rect 51043 43678 52015 43718
rect 52428 43700 52483 43746
rect 52529 43700 52641 43746
rect 52687 43700 52799 43746
rect 52845 43700 52957 43746
rect 53003 43700 53115 43746
rect 53161 43700 53273 43746
rect 53319 43700 53431 43746
rect 53477 43700 53589 43746
rect 53635 43700 53748 43746
rect 53794 43700 53906 43746
rect 53952 43700 54064 43746
rect 54110 43700 54222 43746
rect 54268 43700 54540 43746
rect 52428 43643 54540 43700
rect 30583 43632 30955 43643
rect 30583 43586 30637 43632
rect 30683 43586 30955 43632
rect 30583 43468 30955 43586
rect 30583 43422 30637 43468
rect 30683 43422 30955 43468
rect 30583 43394 30955 43422
rect 54167 43632 54540 43643
rect 54167 43586 54440 43632
rect 54486 43586 54540 43632
rect 54167 43468 54540 43586
rect 54167 43422 54440 43468
rect 54486 43422 54540 43468
rect 28492 43220 28810 43266
rect 28856 43220 29196 43266
rect 29283 43353 30365 43394
rect 29283 43350 29582 43353
rect 29283 43304 29317 43350
rect 29363 43304 29478 43350
rect 29524 43304 29582 43350
rect 29283 43301 29582 43304
rect 29634 43350 29793 43353
rect 29845 43350 30005 43353
rect 29634 43304 29638 43350
rect 29684 43304 29793 43350
rect 29845 43304 29959 43350
rect 29634 43301 29793 43304
rect 29845 43301 30005 43304
rect 30057 43350 30216 43353
rect 30057 43304 30121 43350
rect 30167 43304 30216 43350
rect 30057 43301 30216 43304
rect 30268 43350 30365 43353
rect 30268 43304 30284 43350
rect 30330 43304 30365 43350
rect 30268 43301 30365 43304
rect 29283 43261 30365 43301
rect 30583 43353 32842 43394
rect 34247 43387 35008 43393
rect 30583 43301 30854 43353
rect 30906 43301 31065 43353
rect 31117 43301 31276 43353
rect 31328 43350 31486 43353
rect 31538 43350 31697 43353
rect 31749 43350 31909 43353
rect 31961 43350 32120 43353
rect 32172 43350 32330 43353
rect 32382 43350 32541 43353
rect 32593 43350 32752 43353
rect 32804 43350 32842 43353
rect 34246 43353 35008 43387
rect 34246 43350 34284 43353
rect 34336 43350 34495 43353
rect 34547 43350 34707 43353
rect 31328 43304 31349 43350
rect 33323 43304 33336 43350
rect 33671 43304 33684 43350
rect 33730 43304 33787 43350
rect 33833 43304 33890 43350
rect 33936 43304 33993 43350
rect 34039 43304 34096 43350
rect 34142 43304 34199 43350
rect 34245 43304 34284 43350
rect 34348 43304 34405 43350
rect 34451 43304 34495 43350
rect 34554 43304 34612 43350
rect 34658 43304 34707 43350
rect 31328 43301 31486 43304
rect 31538 43301 31697 43304
rect 31749 43301 31909 43304
rect 31961 43301 32120 43304
rect 32172 43301 32330 43304
rect 32382 43301 32541 43304
rect 32593 43301 32752 43304
rect 32804 43301 32842 43304
rect 30583 43266 32842 43301
rect 34246 43301 34284 43304
rect 34336 43301 34495 43304
rect 34547 43301 34707 43304
rect 34759 43301 34918 43353
rect 34970 43301 35008 43353
rect 34246 43267 35008 43301
rect 29544 43260 30306 43261
rect 28492 43144 29196 43220
rect 28492 43103 29116 43144
rect 28492 43057 28810 43103
rect 28856 43098 29116 43103
rect 29162 43098 29196 43144
rect 28856 43057 29196 43098
rect 28492 42981 29196 43057
rect 28492 42940 29116 42981
rect 28492 42894 28810 42940
rect 28856 42935 29116 42940
rect 29162 42935 29196 42981
rect 28856 42894 29196 42935
rect 28492 42817 29196 42894
rect 28492 42777 29116 42817
rect 28492 42731 28810 42777
rect 28856 42771 29116 42777
rect 29162 42771 29196 42817
rect 28856 42731 29196 42771
rect 28492 42654 29196 42731
rect 28492 42613 29116 42654
rect 28492 42567 28810 42613
rect 28856 42608 29116 42613
rect 29162 42608 29196 42654
rect 28856 42567 29196 42608
rect 28492 42453 29196 42567
rect 30583 43220 30637 43266
rect 30683 43260 32842 43266
rect 34247 43260 35008 43267
rect 35182 43387 36364 43394
rect 37946 43393 38324 43394
rect 35182 43353 36958 43387
rect 35182 43301 35220 43353
rect 35272 43301 35430 43353
rect 35482 43301 35641 43353
rect 35693 43301 35853 43353
rect 35905 43301 36064 43353
rect 36116 43301 36274 43353
rect 36326 43350 36958 43353
rect 36326 43304 36489 43350
rect 36723 43304 36958 43350
rect 36326 43301 36958 43304
rect 35182 43267 36958 43301
rect 37946 43353 38842 43393
rect 37946 43350 38330 43353
rect 38382 43350 38541 43353
rect 37946 43304 37957 43350
rect 38473 43304 38541 43350
rect 37946 43301 38330 43304
rect 38382 43301 38541 43304
rect 38593 43301 38752 43353
rect 38804 43301 38842 43353
rect 35182 43260 36364 43267
rect 37946 43260 38842 43301
rect 39014 43387 39322 43394
rect 40215 43387 40523 43394
rect 40788 43387 42986 43401
rect 54167 43394 54540 43422
rect 55927 44122 56632 44201
rect 55927 44076 56267 44122
rect 56313 44076 56632 44122
rect 55927 44044 56632 44076
rect 55927 43998 55961 44044
rect 56007 43998 56632 44044
rect 55927 43958 56632 43998
rect 55927 43912 56267 43958
rect 56313 43912 56632 43958
rect 55927 43881 56632 43912
rect 55927 43835 55961 43881
rect 56007 43835 56632 43881
rect 55927 43795 56632 43835
rect 55927 43749 56267 43795
rect 56313 43749 56632 43795
rect 55927 43717 56632 43749
rect 55927 43671 55961 43717
rect 56007 43671 56632 43717
rect 55927 43632 56632 43671
rect 55927 43586 56267 43632
rect 56313 43586 56632 43632
rect 55927 43554 56632 43586
rect 55927 43508 55961 43554
rect 56007 43508 56632 43554
rect 55927 43468 56632 43508
rect 55927 43422 56267 43468
rect 56313 43422 56632 43468
rect 43753 43387 44514 43393
rect 39014 43353 39323 43387
rect 39014 43301 39052 43353
rect 39104 43350 39232 43353
rect 39108 43304 39220 43350
rect 39104 43301 39232 43304
rect 39284 43301 39323 43353
rect 30683 43226 31040 43260
rect 30683 43220 30855 43226
rect 30583 43180 30855 43220
rect 30901 43180 31040 43226
rect 30583 43103 31040 43180
rect 33484 43184 33552 43195
rect 33019 43129 33327 43170
rect 33019 43126 33057 43129
rect 33109 43126 33237 43129
rect 33289 43126 33327 43129
rect 30583 43057 30637 43103
rect 30683 43062 31040 43103
rect 31336 43080 31349 43126
rect 33323 43080 33336 43126
rect 30683 43057 30855 43062
rect 30583 43016 30855 43057
rect 30901 43016 31040 43062
rect 33019 43077 33057 43080
rect 33109 43077 33237 43080
rect 33289 43077 33327 43080
rect 33019 43037 33327 43077
rect 30583 42940 31040 43016
rect 30583 42894 30637 42940
rect 30683 42924 31040 42940
rect 30683 42902 31493 42924
rect 30683 42899 31349 42902
rect 30683 42894 30855 42899
rect 30583 42853 30855 42894
rect 30901 42856 31349 42899
rect 33323 42856 33336 42902
rect 30901 42853 31493 42856
rect 30583 42805 31493 42853
rect 30583 42777 31040 42805
rect 30583 42731 30637 42777
rect 30683 42736 31040 42777
rect 30683 42731 30855 42736
rect 30583 42690 30855 42731
rect 30901 42690 31040 42736
rect 33484 42762 33495 43184
rect 33541 42762 33552 43184
rect 33781 43137 34089 43178
rect 33781 43126 33819 43137
rect 33871 43126 33999 43137
rect 34051 43126 34089 43137
rect 33671 43080 33684 43126
rect 33730 43080 33787 43126
rect 33871 43085 33890 43126
rect 33833 43080 33890 43085
rect 33936 43080 33993 43126
rect 34051 43085 34096 43126
rect 34039 43080 34096 43085
rect 34142 43080 34199 43126
rect 34245 43080 34302 43126
rect 34348 43080 34405 43126
rect 34451 43080 34508 43126
rect 34554 43080 34612 43126
rect 34658 43080 34671 43126
rect 33781 43045 34089 43080
rect 35294 43051 36266 43091
rect 37853 43088 38161 43104
rect 35294 43039 35332 43051
rect 35384 43039 35543 43051
rect 35595 43039 35754 43051
rect 35806 43039 35965 43051
rect 36017 43039 36176 43051
rect 36228 43039 36266 43051
rect 36438 43039 36953 43088
rect 37439 43063 38161 43088
rect 37439 43039 37891 43063
rect 37943 43039 38071 43063
rect 38123 43039 38161 43063
rect 35260 42993 35273 43039
rect 35523 42999 35543 43039
rect 35523 42993 35580 42999
rect 35626 42993 35683 43039
rect 35729 42999 35754 43039
rect 35729 42993 35786 42999
rect 35832 42993 35889 43039
rect 35935 42999 35965 43039
rect 35935 42993 35992 42999
rect 36038 42993 36095 43039
rect 36141 42999 36176 43039
rect 36141 42993 36198 42999
rect 36244 42993 36301 43039
rect 36347 42993 36360 43039
rect 36438 42993 36854 43039
rect 36900 42993 36971 43039
rect 37017 42993 37088 43039
rect 37134 42993 37206 43039
rect 37252 42993 37324 43039
rect 37370 42993 37442 43039
rect 37488 43011 37891 43039
rect 37488 42993 37909 43011
rect 37955 42993 38026 43039
rect 38123 43011 38143 43039
rect 38072 42993 38143 43011
rect 38189 42993 38261 43039
rect 38307 42993 38379 43039
rect 38425 42993 38497 43039
rect 38543 42993 38556 43039
rect 35294 42959 36266 42993
rect 36438 42968 36953 42993
rect 37439 42971 38161 42993
rect 37439 42968 37931 42971
rect 34228 42902 34718 42931
rect 33671 42856 33684 42902
rect 33730 42856 33787 42902
rect 33833 42856 33890 42902
rect 33936 42856 33993 42902
rect 34039 42856 34096 42902
rect 34142 42856 34199 42902
rect 34245 42891 34302 42902
rect 34245 42856 34267 42891
rect 34348 42856 34405 42902
rect 34451 42891 34508 42902
rect 34499 42856 34508 42891
rect 34554 42856 34612 42902
rect 34658 42891 34718 42902
rect 34228 42839 34267 42856
rect 34319 42839 34447 42856
rect 34499 42839 34627 42856
rect 34679 42839 34718 42891
rect 36438 42865 36554 42968
rect 34228 42798 34718 42839
rect 34964 42815 36360 42859
rect 30583 42613 31040 42690
rect 33019 42681 33327 42722
rect 33019 42678 33057 42681
rect 33109 42678 33237 42681
rect 33289 42678 33327 42681
rect 33484 42680 33552 42762
rect 34964 42769 35273 42815
rect 35523 42769 35580 42815
rect 35626 42769 35683 42815
rect 35729 42769 35786 42815
rect 35832 42769 35889 42815
rect 35935 42769 35992 42815
rect 36038 42769 36095 42815
rect 36141 42769 36198 42815
rect 36244 42769 36301 42815
rect 36347 42769 36360 42815
rect 34964 42737 36360 42769
rect 34964 42680 35082 42737
rect 31336 42632 31349 42678
rect 33323 42632 33336 42678
rect 33484 42643 35082 42680
rect 30583 42567 30637 42613
rect 30683 42573 31040 42613
rect 33019 42629 33057 42632
rect 33109 42629 33237 42632
rect 33289 42629 33327 42632
rect 33019 42589 33327 42629
rect 33484 42597 33816 42643
rect 33862 42597 34002 42643
rect 34048 42597 34189 42643
rect 34235 42597 34376 42643
rect 34422 42597 34562 42643
rect 34608 42597 35082 42643
rect 36438 42725 36475 42865
rect 36521 42725 36554 42865
rect 33484 42589 35082 42597
rect 35294 42591 36266 42631
rect 36438 42625 36554 42725
rect 36640 42865 36773 42888
rect 36640 42816 36697 42865
rect 36640 42764 36678 42816
rect 36640 42725 36697 42764
rect 36743 42725 36773 42865
rect 38658 42867 38726 42878
rect 36924 42857 37685 42863
rect 36923 42856 37685 42857
rect 36923 42823 37931 42856
rect 36923 42815 36961 42823
rect 37013 42815 37172 42823
rect 37224 42815 37384 42823
rect 36841 42769 36854 42815
rect 36900 42771 36961 42815
rect 36900 42769 36971 42771
rect 37017 42769 37088 42815
rect 37134 42771 37172 42815
rect 37134 42769 37206 42771
rect 37252 42769 37324 42815
rect 37370 42771 37384 42815
rect 37436 42815 37595 42823
rect 37436 42771 37442 42815
rect 37370 42769 37442 42771
rect 37488 42771 37595 42815
rect 37647 42815 37931 42823
rect 37647 42771 37909 42815
rect 37488 42769 37909 42771
rect 37955 42769 38026 42815
rect 38072 42769 38143 42815
rect 38189 42769 38261 42815
rect 38307 42769 38379 42815
rect 38425 42769 38497 42815
rect 38543 42769 38556 42815
rect 36923 42737 37931 42769
rect 36924 42730 37685 42737
rect 36640 42705 36773 42725
rect 38658 42727 38669 42867
rect 38715 42727 38726 42867
rect 39014 42815 39323 43301
rect 39492 43364 42986 43387
rect 43704 43364 44514 43387
rect 39492 43353 44514 43364
rect 39492 43350 40253 43353
rect 39492 43304 39740 43350
rect 39786 43304 39862 43350
rect 39908 43304 39985 43350
rect 40031 43304 40108 43350
rect 40154 43304 40253 43350
rect 39492 43301 40253 43304
rect 40305 43301 40433 43353
rect 40485 43350 43790 43353
rect 40485 43304 40836 43350
rect 40882 43304 40994 43350
rect 41040 43304 41152 43350
rect 41198 43304 41310 43350
rect 41356 43304 41469 43350
rect 41515 43304 41627 43350
rect 41673 43304 41785 43350
rect 41831 43304 41943 43350
rect 41989 43304 42101 43350
rect 42147 43304 42259 43350
rect 42305 43304 42418 43350
rect 42464 43304 42576 43350
rect 42622 43304 42734 43350
rect 42780 43304 42892 43350
rect 42938 43304 43739 43350
rect 43785 43304 43790 43350
rect 40485 43301 43790 43304
rect 43842 43350 44001 43353
rect 43842 43304 43906 43350
rect 43952 43304 44001 43350
rect 43842 43301 44001 43304
rect 44053 43350 44213 43353
rect 44265 43350 44424 43353
rect 44053 43304 44071 43350
rect 44117 43304 44213 43350
rect 44282 43304 44424 43350
rect 44053 43301 44213 43304
rect 44265 43301 44424 43304
rect 44476 43301 44514 43353
rect 39492 43290 44514 43301
rect 39492 43267 42986 43290
rect 43704 43267 44514 43290
rect 39492 42815 39608 43267
rect 40215 43261 40523 43267
rect 40788 43253 42986 43267
rect 43753 43260 44514 43267
rect 44796 43387 45346 43393
rect 48800 43387 49982 43394
rect 50308 43387 50859 43394
rect 44796 43353 49982 43387
rect 44796 43350 44834 43353
rect 44886 43350 45045 43353
rect 45097 43350 45256 43353
rect 45308 43350 48838 43353
rect 44796 43304 44812 43350
rect 44886 43304 44925 43350
rect 44971 43304 45038 43350
rect 45097 43304 45151 43350
rect 45197 43304 45256 43350
rect 45310 43304 45619 43350
rect 45665 43304 45777 43350
rect 45823 43304 45935 43350
rect 45981 43304 46093 43350
rect 46139 43304 46251 43350
rect 46297 43304 46409 43350
rect 46455 43304 46568 43350
rect 46614 43304 46726 43350
rect 46772 43304 46884 43350
rect 46930 43304 47042 43350
rect 47088 43304 47200 43350
rect 47246 43304 47358 43350
rect 47404 43304 47516 43350
rect 47562 43304 47675 43350
rect 47721 43304 47833 43350
rect 47879 43304 47991 43350
rect 48037 43304 48149 43350
rect 48195 43304 48307 43350
rect 48353 43304 48465 43350
rect 48511 43304 48838 43350
rect 44796 43301 44834 43304
rect 44886 43301 45045 43304
rect 45097 43301 45256 43304
rect 45308 43301 48838 43304
rect 48890 43301 49048 43353
rect 49100 43301 49259 43353
rect 49311 43301 49471 43353
rect 49523 43301 49682 43353
rect 49734 43301 49892 43353
rect 49944 43301 49982 43353
rect 44796 43267 49982 43301
rect 50307 43353 50859 43387
rect 50307 43301 50346 43353
rect 50398 43350 50557 43353
rect 50609 43350 50768 43353
rect 50820 43350 50859 43353
rect 52278 43353 54540 43394
rect 52278 43350 52316 43353
rect 52368 43350 52527 43353
rect 52579 43350 52738 43353
rect 52790 43350 52948 43353
rect 53000 43350 53159 43353
rect 53211 43350 53371 43353
rect 53423 43350 53582 43353
rect 53634 43350 53792 43353
rect 50398 43304 50467 43350
rect 50513 43304 50557 43350
rect 50617 43304 50674 43350
rect 50720 43304 50768 43350
rect 50823 43304 50880 43350
rect 50926 43304 50983 43350
rect 51029 43304 51086 43350
rect 51132 43304 51189 43350
rect 51235 43304 51292 43350
rect 51338 43304 51395 43350
rect 51441 43304 51454 43350
rect 51789 43304 51802 43350
rect 53776 43304 53792 43350
rect 50398 43301 50557 43304
rect 50609 43301 50768 43304
rect 50820 43301 50859 43304
rect 50307 43267 50859 43301
rect 44796 43260 45346 43267
rect 43362 43209 43524 43220
rect 39737 43126 39866 43155
rect 40246 43137 40362 43174
rect 43362 43163 43373 43209
rect 43513 43163 43524 43209
rect 43362 43156 43524 43163
rect 39727 43080 39740 43126
rect 39786 43115 39862 43126
rect 39827 43080 39862 43115
rect 39908 43080 39985 43126
rect 40031 43080 40108 43126
rect 40154 43080 40167 43126
rect 40246 43091 40281 43137
rect 40327 43091 40362 43137
rect 39737 43063 39775 43080
rect 39827 43063 39866 43080
rect 39737 43036 39866 43063
rect 39737 43023 39865 43036
rect 39923 42900 40085 42940
rect 39923 42848 39994 42900
rect 40046 42848 40085 42900
rect 39008 42769 39021 42815
rect 39067 42769 39144 42815
rect 39190 42769 39267 42815
rect 39313 42769 39326 42815
rect 39492 42769 39641 42815
rect 39687 42769 39730 42815
rect 39014 42737 39323 42769
rect 39492 42737 39608 42769
rect 37853 42625 38161 42630
rect 36438 42591 36953 42625
rect 37439 42591 38161 42625
rect 38658 42605 38726 42727
rect 39923 42717 40085 42848
rect 39809 42714 40085 42717
rect 39809 42706 39994 42714
rect 39809 42660 39844 42706
rect 39890 42662 39994 42706
rect 40046 42693 40085 42714
rect 40246 42693 40362 43091
rect 40718 43115 43524 43156
rect 45584 43186 48546 43267
rect 48800 43260 49982 43267
rect 50308 43260 50859 43267
rect 52278 43301 52316 43304
rect 52368 43301 52527 43304
rect 52579 43301 52738 43304
rect 52790 43301 52948 43304
rect 53000 43301 53159 43304
rect 53211 43301 53371 43304
rect 53423 43301 53582 43304
rect 53634 43301 53792 43304
rect 53844 43301 54003 43353
rect 54055 43301 54214 43353
rect 54266 43301 54540 43353
rect 52278 43266 54540 43301
rect 52278 43260 54440 43266
rect 45584 43140 45619 43186
rect 45665 43140 45777 43186
rect 45823 43140 45935 43186
rect 45981 43140 46093 43186
rect 46139 43140 46251 43186
rect 46297 43140 46409 43186
rect 46455 43140 46568 43186
rect 46614 43140 46726 43186
rect 46772 43140 46884 43186
rect 46930 43140 47042 43186
rect 47088 43140 47200 43186
rect 47246 43140 47358 43186
rect 47404 43140 47516 43186
rect 47562 43140 47675 43186
rect 47721 43140 47833 43186
rect 47879 43140 47991 43186
rect 48037 43140 48149 43186
rect 48195 43140 48307 43186
rect 48353 43140 48465 43186
rect 48511 43140 48546 43186
rect 54085 43226 54440 43260
rect 54085 43180 54223 43226
rect 54269 43220 54440 43226
rect 54486 43220 54540 43266
rect 54758 43353 55840 43394
rect 54758 43350 54855 43353
rect 54758 43304 54793 43350
rect 54839 43304 54855 43350
rect 54758 43301 54855 43304
rect 54907 43350 55066 43353
rect 54907 43304 54956 43350
rect 55002 43304 55066 43350
rect 54907 43301 55066 43304
rect 55118 43350 55278 43353
rect 55330 43350 55489 43353
rect 55164 43304 55278 43350
rect 55330 43304 55439 43350
rect 55485 43304 55489 43350
rect 55118 43301 55278 43304
rect 55330 43301 55489 43304
rect 55541 43350 55840 43353
rect 55541 43304 55599 43350
rect 55645 43304 55760 43350
rect 55806 43304 55840 43350
rect 55541 43301 55840 43304
rect 54758 43261 55840 43301
rect 55927 43266 56632 43422
rect 54817 43260 55579 43261
rect 54269 43180 54540 43220
rect 40718 43063 41935 43115
rect 41987 43063 43524 43115
rect 40718 43022 43524 43063
rect 44605 43080 44812 43126
rect 44858 43080 44925 43126
rect 44971 43080 45038 43126
rect 45084 43080 45151 43126
rect 45197 43080 45264 43126
rect 45310 43080 45323 43126
rect 45584 43104 48546 43140
rect 51035 43129 51343 43170
rect 51035 43126 51073 43129
rect 51125 43126 51253 43129
rect 51305 43126 51343 43129
rect 51589 43154 51657 43165
rect 44341 43014 44509 43025
rect 44341 42968 44358 43014
rect 44498 42968 44509 43014
rect 44341 42924 44509 42968
rect 42229 42884 44509 42924
rect 42229 42832 43445 42884
rect 43497 42832 44509 42884
rect 42229 42791 44509 42832
rect 44605 42693 44721 43080
rect 48905 43054 49877 43094
rect 50454 43080 50467 43126
rect 50513 43080 50571 43126
rect 50617 43080 50674 43126
rect 50720 43080 50777 43126
rect 50823 43080 50880 43126
rect 50926 43080 50983 43126
rect 51029 43080 51073 43126
rect 51132 43080 51189 43126
rect 51235 43080 51253 43126
rect 51338 43080 51395 43126
rect 51441 43080 51454 43126
rect 48905 43039 48943 43054
rect 48995 43039 49154 43054
rect 49206 43039 49365 43054
rect 49417 43039 49576 43054
rect 49628 43039 49787 43054
rect 49839 43039 49877 43054
rect 48765 42993 48778 43039
rect 48824 42993 48881 43039
rect 48927 43002 48943 43039
rect 48927 42993 48984 43002
rect 49030 42993 49087 43039
rect 49133 43002 49154 43039
rect 49133 42993 49190 43002
rect 49236 42993 49293 43039
rect 49339 43002 49365 43039
rect 49339 42993 49396 43002
rect 49442 42993 49499 43039
rect 49545 43002 49576 43039
rect 49545 42993 49602 43002
rect 49852 42993 49877 43039
rect 51035 43077 51073 43080
rect 51125 43077 51253 43080
rect 51305 43077 51343 43080
rect 51035 43037 51343 43077
rect 48557 42947 48687 42988
rect 48905 42962 49877 42993
rect 44901 42902 45241 42931
rect 44799 42856 44812 42902
rect 44858 42856 44925 42902
rect 44971 42891 45038 42902
rect 44991 42856 45038 42891
rect 45084 42856 45151 42902
rect 45197 42891 45264 42902
rect 45203 42856 45264 42891
rect 45310 42856 45323 42902
rect 48557 42895 48596 42947
rect 48648 42895 48687 42947
rect 48557 42892 48687 42895
rect 44901 42839 44939 42856
rect 44991 42839 45151 42856
rect 45203 42839 45241 42856
rect 44901 42798 45241 42839
rect 45400 42783 48379 42816
rect 45400 42737 45464 42783
rect 45604 42775 48379 42783
rect 45400 42723 45597 42737
rect 45649 42723 48379 42775
rect 40046 42678 44918 42693
rect 45400 42682 48379 42723
rect 48557 42752 48622 42892
rect 48668 42752 48687 42892
rect 50262 42902 50812 42931
rect 50262 42891 50467 42902
rect 50513 42891 50571 42902
rect 49820 42815 50160 42856
rect 48765 42769 48778 42815
rect 48824 42769 48881 42815
rect 48927 42769 48984 42815
rect 49030 42769 49087 42815
rect 49133 42769 49190 42815
rect 49236 42769 49293 42815
rect 49339 42769 49396 42815
rect 49442 42769 49499 42815
rect 49545 42769 49602 42815
rect 49852 42769 50160 42815
rect 50262 42839 50300 42891
rect 50352 42856 50467 42891
rect 50563 42856 50571 42891
rect 50617 42856 50674 42902
rect 50720 42891 50777 42902
rect 50720 42856 50722 42891
rect 50352 42839 50511 42856
rect 50563 42839 50722 42856
rect 50774 42856 50777 42891
rect 50823 42856 50880 42902
rect 50926 42856 50983 42902
rect 51029 42856 51086 42902
rect 51132 42856 51189 42902
rect 51235 42856 51292 42902
rect 51338 42856 51395 42902
rect 51441 42856 51454 42902
rect 50774 42839 50812 42856
rect 50262 42798 50812 42839
rect 48557 42729 48687 42752
rect 49820 42737 50160 42769
rect 40046 42662 44812 42678
rect 39890 42660 44812 42662
rect 39809 42657 44812 42660
rect 39809 42611 43739 42657
rect 43785 42611 43906 42657
rect 43952 42611 44071 42657
rect 44117 42611 44236 42657
rect 44282 42632 44812 42657
rect 44858 42632 44925 42678
rect 44971 42632 45038 42678
rect 45084 42632 45151 42678
rect 45197 42632 45264 42678
rect 45310 42632 45323 42678
rect 48557 42677 48596 42729
rect 48648 42677 48687 42729
rect 48557 42637 48687 42677
rect 50044 42680 50160 42737
rect 51589 42732 51600 43154
rect 51646 42732 51657 43154
rect 51797 43126 52105 43163
rect 51789 43080 51802 43126
rect 53776 43080 53789 43126
rect 54085 43103 54540 43180
rect 51797 43070 51835 43080
rect 51887 43070 52015 43080
rect 52067 43070 52105 43080
rect 51797 43030 52105 43070
rect 54085 43062 54440 43103
rect 54085 43016 54223 43062
rect 54269 43057 54440 43062
rect 54486 43057 54540 43103
rect 54269 43016 54540 43057
rect 54085 42940 54540 43016
rect 54085 42924 54440 42940
rect 53585 42902 54440 42924
rect 51789 42856 51802 42902
rect 53776 42894 54440 42902
rect 54486 42894 54540 42940
rect 53776 42856 54540 42894
rect 53585 42805 54540 42856
rect 51589 42680 51657 42732
rect 54085 42777 54540 42805
rect 54085 42731 54440 42777
rect 54486 42731 54540 42777
rect 50044 42643 51657 42680
rect 51797 42678 52105 42700
rect 44282 42611 44918 42632
rect 38658 42591 39723 42605
rect 30683 42567 30855 42573
rect 30583 42527 30855 42567
rect 30901 42527 31040 42573
rect 33484 42560 34643 42589
rect 35260 42545 35273 42591
rect 35523 42545 35543 42591
rect 35626 42545 35683 42591
rect 35729 42545 35754 42591
rect 35832 42545 35889 42591
rect 35935 42545 35965 42591
rect 36038 42545 36095 42591
rect 36141 42545 36176 42591
rect 36244 42545 36301 42591
rect 36347 42545 36360 42591
rect 36438 42545 36854 42591
rect 36900 42545 36971 42591
rect 37017 42545 37088 42591
rect 37134 42545 37206 42591
rect 37252 42545 37324 42591
rect 37370 42545 37442 42591
rect 37488 42589 37909 42591
rect 37488 42545 37891 42589
rect 37955 42545 38026 42591
rect 38072 42589 38143 42591
rect 38123 42545 38143 42589
rect 38189 42545 38261 42591
rect 38307 42545 38379 42591
rect 38425 42545 38497 42591
rect 38543 42545 38556 42591
rect 38658 42545 39021 42591
rect 39067 42545 39144 42591
rect 39190 42545 39267 42591
rect 39313 42545 39641 42591
rect 39687 42545 39730 42591
rect 39809 42573 44918 42611
rect 48905 42591 49877 42631
rect 48765 42545 48778 42591
rect 48824 42545 48881 42591
rect 48927 42545 48943 42591
rect 49030 42545 49087 42591
rect 49133 42545 49154 42591
rect 49236 42545 49293 42591
rect 49339 42545 49365 42591
rect 49442 42545 49499 42591
rect 49545 42545 49576 42591
rect 49852 42545 49877 42591
rect 50044 42597 50516 42643
rect 50562 42597 50703 42643
rect 50749 42597 50890 42643
rect 50936 42597 51076 42643
rect 51122 42597 51263 42643
rect 51309 42597 51657 42643
rect 51789 42632 51802 42678
rect 53776 42632 53789 42678
rect 50044 42587 51657 42597
rect 50481 42560 51657 42587
rect 51797 42607 51835 42632
rect 51887 42607 52015 42632
rect 52067 42607 52105 42632
rect 51797 42567 52105 42607
rect 54085 42613 54540 42731
rect 54085 42573 54440 42613
rect 30583 42494 31040 42527
rect 35294 42539 35332 42545
rect 35384 42539 35543 42545
rect 35595 42539 35754 42545
rect 35806 42539 35965 42545
rect 36017 42539 36176 42545
rect 36228 42539 36266 42545
rect 34870 42494 35025 42501
rect 35294 42499 36266 42539
rect 36438 42505 36953 42545
rect 37439 42537 37891 42545
rect 37943 42537 38071 42545
rect 38123 42537 38161 42545
rect 37439 42505 38161 42537
rect 37853 42497 38161 42505
rect 27744 42401 27790 42453
rect 27842 42401 27846 42453
rect 28492 42401 28634 42453
rect 28686 42450 28845 42453
rect 28686 42404 28810 42450
rect 28686 42401 28845 42404
rect 28897 42401 29056 42453
rect 29108 42401 29196 42453
rect 27744 40653 27846 42401
rect 28492 42287 29196 42401
rect 29283 42453 30365 42494
rect 29283 42450 29582 42453
rect 29283 42404 29317 42450
rect 29363 42404 29478 42450
rect 29524 42404 29582 42450
rect 29283 42401 29582 42404
rect 29634 42450 29793 42453
rect 29845 42450 30005 42453
rect 29634 42404 29638 42450
rect 29684 42404 29793 42450
rect 29845 42404 29959 42450
rect 29634 42401 29793 42404
rect 29845 42401 30005 42404
rect 30057 42450 30216 42453
rect 30057 42404 30121 42450
rect 30167 42404 30216 42450
rect 30057 42401 30216 42404
rect 30268 42450 30365 42453
rect 30268 42404 30284 42450
rect 30330 42404 30365 42450
rect 30268 42401 30365 42404
rect 29283 42361 30365 42401
rect 30583 42453 32842 42494
rect 30583 42450 30854 42453
rect 30583 42404 30637 42450
rect 30683 42404 30854 42450
rect 30583 42401 30854 42404
rect 30906 42401 31065 42453
rect 31117 42401 31276 42453
rect 31328 42401 31486 42453
rect 31538 42401 31697 42453
rect 31749 42401 31909 42453
rect 31961 42401 32120 42453
rect 32172 42401 32330 42453
rect 32382 42401 32541 42453
rect 32593 42401 32752 42453
rect 32804 42401 32842 42453
rect 29544 42360 30306 42361
rect 30583 42360 32842 42401
rect 34717 42453 35025 42494
rect 38658 42485 39723 42545
rect 48905 42539 48943 42545
rect 48995 42539 49154 42545
rect 49206 42539 49365 42545
rect 49417 42539 49576 42545
rect 49628 42539 49787 42545
rect 49839 42539 49877 42545
rect 48905 42499 49877 42539
rect 54085 42527 54223 42573
rect 54269 42567 54440 42573
rect 54486 42567 54540 42613
rect 54269 42527 54540 42567
rect 50099 42494 50255 42501
rect 54085 42494 54540 42527
rect 55927 43220 56267 43266
rect 56313 43220 56632 43266
rect 55927 43144 56632 43220
rect 55927 43098 55961 43144
rect 56007 43103 56632 43144
rect 56007 43098 56267 43103
rect 55927 43057 56267 43098
rect 56313 43057 56632 43103
rect 55927 42981 56632 43057
rect 55927 42935 55961 42981
rect 56007 42940 56632 42981
rect 56007 42935 56267 42940
rect 55927 42894 56267 42935
rect 56313 42894 56632 42940
rect 55927 42817 56632 42894
rect 55927 42771 55961 42817
rect 56007 42777 56632 42817
rect 56007 42771 56267 42777
rect 55927 42731 56267 42771
rect 56313 42731 56632 42777
rect 55927 42654 56632 42731
rect 55927 42608 55961 42654
rect 56007 42613 56632 42654
rect 56007 42608 56267 42613
rect 55927 42567 56267 42608
rect 56313 42567 56632 42613
rect 34717 42401 34755 42453
rect 34807 42450 34935 42453
rect 34807 42404 34916 42450
rect 34807 42401 34935 42404
rect 34987 42401 35025 42453
rect 34717 42360 35025 42401
rect 50099 42453 50408 42494
rect 50099 42401 50138 42453
rect 50190 42450 50318 42453
rect 50206 42404 50318 42450
rect 50190 42401 50318 42404
rect 50370 42401 50408 42453
rect 28492 42241 28810 42287
rect 28856 42244 29196 42287
rect 28856 42241 29116 42244
rect 28492 42198 29116 42241
rect 29162 42198 29196 42244
rect 28492 42123 29196 42198
rect 28492 42077 28810 42123
rect 28856 42081 29196 42123
rect 28856 42077 29116 42081
rect 28492 42035 29116 42077
rect 29162 42035 29196 42081
rect 28492 41960 29196 42035
rect 28492 41914 28810 41960
rect 28856 41917 29196 41960
rect 28856 41914 29116 41917
rect 28492 41871 29116 41914
rect 29162 41871 29196 41917
rect 28492 41797 29196 41871
rect 28492 41751 28810 41797
rect 28856 41754 29196 41797
rect 28856 41751 29116 41754
rect 28492 41708 29116 41751
rect 29162 41708 29196 41754
rect 28492 41634 29196 41708
rect 28492 41588 28810 41634
rect 28856 41588 29196 41634
rect 30583 42327 31040 42360
rect 34870 42353 35025 42360
rect 30583 42287 30855 42327
rect 30583 42241 30637 42287
rect 30683 42281 30855 42287
rect 30901 42281 31040 42327
rect 35294 42315 36266 42355
rect 37853 42349 38161 42357
rect 35294 42309 35332 42315
rect 35384 42309 35543 42315
rect 35595 42309 35754 42315
rect 35806 42309 35965 42315
rect 36017 42309 36176 42315
rect 36228 42309 36266 42315
rect 36438 42309 36953 42349
rect 37439 42317 38161 42349
rect 37439 42309 37891 42317
rect 37943 42309 38071 42317
rect 38123 42309 38161 42317
rect 38658 42309 39723 42369
rect 50099 42360 50408 42401
rect 52278 42453 54540 42494
rect 52278 42401 52316 42453
rect 52368 42401 52527 42453
rect 52579 42401 52738 42453
rect 52790 42401 52948 42453
rect 53000 42401 53159 42453
rect 53211 42401 53371 42453
rect 53423 42401 53582 42453
rect 53634 42401 53792 42453
rect 53844 42401 54003 42453
rect 54055 42401 54214 42453
rect 54266 42450 54540 42453
rect 54266 42404 54440 42450
rect 54486 42404 54540 42450
rect 54266 42401 54540 42404
rect 52278 42360 54540 42401
rect 54758 42453 55840 42494
rect 54758 42450 54855 42453
rect 54758 42404 54793 42450
rect 54839 42404 54855 42450
rect 54758 42401 54855 42404
rect 54907 42450 55066 42453
rect 54907 42404 54956 42450
rect 55002 42404 55066 42450
rect 54907 42401 55066 42404
rect 55118 42450 55278 42453
rect 55330 42450 55489 42453
rect 55164 42404 55278 42450
rect 55330 42404 55439 42450
rect 55485 42404 55489 42450
rect 55118 42401 55278 42404
rect 55330 42401 55489 42404
rect 55541 42450 55840 42453
rect 55541 42404 55599 42450
rect 55645 42404 55760 42450
rect 55806 42404 55840 42450
rect 55541 42401 55840 42404
rect 54758 42361 55840 42401
rect 55927 42453 56632 42567
rect 57278 42453 57380 44201
rect 55927 42401 56015 42453
rect 56067 42401 56226 42453
rect 56278 42450 56437 42453
rect 56313 42404 56437 42450
rect 56278 42401 56437 42404
rect 56489 42401 56632 42453
rect 57278 42401 57281 42453
rect 57333 42401 57380 42453
rect 54817 42360 55579 42361
rect 48905 42315 49877 42355
rect 50099 42353 50255 42360
rect 48905 42309 48943 42315
rect 48995 42309 49154 42315
rect 49206 42309 49365 42315
rect 49417 42309 49576 42315
rect 49628 42309 49787 42315
rect 49839 42309 49877 42315
rect 30683 42241 31040 42281
rect 33484 42265 34643 42294
rect 30583 42164 31040 42241
rect 33019 42225 33327 42265
rect 33019 42222 33057 42225
rect 33109 42222 33237 42225
rect 33289 42222 33327 42225
rect 33484 42257 35082 42265
rect 35260 42263 35273 42309
rect 35523 42263 35543 42309
rect 35626 42263 35683 42309
rect 35729 42263 35754 42309
rect 35832 42263 35889 42309
rect 35935 42263 35965 42309
rect 36038 42263 36095 42309
rect 36141 42263 36176 42309
rect 36244 42263 36301 42309
rect 36347 42263 36360 42309
rect 36438 42263 36854 42309
rect 36900 42263 36971 42309
rect 37017 42263 37088 42309
rect 37134 42263 37206 42309
rect 37252 42263 37324 42309
rect 37370 42263 37442 42309
rect 37488 42265 37891 42309
rect 37488 42263 37909 42265
rect 37955 42263 38026 42309
rect 38123 42265 38143 42309
rect 38072 42263 38143 42265
rect 38189 42263 38261 42309
rect 38307 42263 38379 42309
rect 38425 42263 38497 42309
rect 38543 42263 38556 42309
rect 38658 42263 39021 42309
rect 39067 42263 39144 42309
rect 39190 42263 39267 42309
rect 39313 42263 39641 42309
rect 39687 42263 39730 42309
rect 31336 42176 31349 42222
rect 33323 42176 33336 42222
rect 33484 42211 33816 42257
rect 33862 42211 34002 42257
rect 34048 42211 34189 42257
rect 34235 42211 34376 42257
rect 34422 42211 34562 42257
rect 34608 42211 35082 42257
rect 35294 42223 36266 42263
rect 36438 42229 36953 42263
rect 37439 42229 38161 42263
rect 30583 42123 30855 42164
rect 30583 42077 30637 42123
rect 30683 42118 30855 42123
rect 30901 42118 31040 42164
rect 33019 42173 33057 42176
rect 33109 42173 33237 42176
rect 33289 42173 33327 42176
rect 33019 42132 33327 42173
rect 33484 42174 35082 42211
rect 30683 42077 31040 42118
rect 30583 42049 31040 42077
rect 33484 42092 33552 42174
rect 30583 42001 31493 42049
rect 30583 41960 30855 42001
rect 30583 41914 30637 41960
rect 30683 41955 30855 41960
rect 30901 41998 31493 42001
rect 30901 41955 31349 41998
rect 30683 41952 31349 41955
rect 33323 41952 33336 41998
rect 30683 41930 31493 41952
rect 30683 41914 31040 41930
rect 30583 41838 31040 41914
rect 30583 41797 30855 41838
rect 30583 41751 30637 41797
rect 30683 41792 30855 41797
rect 30901 41792 31040 41838
rect 30683 41751 31040 41792
rect 33019 41777 33327 41817
rect 33019 41774 33057 41777
rect 33109 41774 33237 41777
rect 33289 41774 33327 41777
rect 30583 41674 31040 41751
rect 31336 41728 31349 41774
rect 33323 41728 33336 41774
rect 33019 41725 33057 41728
rect 33109 41725 33237 41728
rect 33289 41725 33327 41728
rect 33019 41684 33327 41725
rect 30583 41634 30855 41674
rect 28492 41466 29196 41588
rect 28492 41420 28810 41466
rect 28856 41420 29196 41466
rect 29283 41553 30365 41594
rect 29283 41550 29582 41553
rect 29283 41504 29317 41550
rect 29363 41504 29478 41550
rect 29524 41504 29582 41550
rect 29283 41501 29582 41504
rect 29634 41550 29793 41553
rect 29845 41550 30005 41553
rect 29634 41504 29638 41550
rect 29684 41504 29793 41550
rect 29845 41504 29959 41550
rect 29634 41501 29793 41504
rect 29845 41501 30005 41504
rect 30057 41550 30216 41553
rect 30057 41504 30121 41550
rect 30167 41504 30216 41550
rect 30057 41501 30216 41504
rect 30268 41550 30365 41553
rect 30268 41504 30284 41550
rect 30330 41504 30365 41550
rect 30268 41501 30365 41504
rect 29283 41461 30365 41501
rect 30583 41588 30637 41634
rect 30683 41628 30855 41634
rect 30901 41628 31040 41674
rect 33484 41670 33495 42092
rect 33541 41670 33552 42092
rect 34964 42117 35082 42174
rect 36438 42129 36554 42229
rect 37853 42224 38161 42229
rect 38658 42249 39723 42263
rect 34964 42085 36360 42117
rect 34228 42015 34718 42056
rect 34228 41998 34267 42015
rect 34319 41998 34447 42015
rect 34499 41998 34627 42015
rect 33671 41952 33684 41998
rect 33730 41952 33787 41998
rect 33833 41952 33890 41998
rect 33936 41952 33993 41998
rect 34039 41952 34096 41998
rect 34142 41952 34199 41998
rect 34245 41963 34267 41998
rect 34245 41952 34302 41963
rect 34348 41952 34405 41998
rect 34499 41963 34508 41998
rect 34451 41952 34508 41963
rect 34554 41952 34612 41998
rect 34679 41963 34718 42015
rect 34964 42039 35273 42085
rect 35523 42039 35580 42085
rect 35626 42039 35683 42085
rect 35729 42039 35786 42085
rect 35832 42039 35889 42085
rect 35935 42039 35992 42085
rect 36038 42039 36095 42085
rect 36141 42039 36198 42085
rect 36244 42039 36301 42085
rect 36347 42039 36360 42085
rect 34964 41995 36360 42039
rect 34658 41952 34718 41963
rect 34228 41923 34718 41952
rect 36438 41989 36475 42129
rect 36521 41989 36554 42129
rect 35294 41861 36266 41895
rect 36438 41886 36554 41989
rect 36640 42129 36773 42149
rect 36640 42090 36697 42129
rect 36640 42038 36678 42090
rect 36640 41989 36697 42038
rect 36743 41989 36773 42129
rect 38658 42127 38726 42249
rect 39809 42243 44918 42281
rect 48765 42263 48778 42309
rect 48824 42263 48881 42309
rect 48927 42263 48943 42309
rect 49030 42263 49087 42309
rect 49133 42263 49154 42309
rect 49236 42263 49293 42309
rect 49339 42263 49365 42309
rect 49442 42263 49499 42309
rect 49545 42263 49576 42309
rect 49852 42263 49877 42309
rect 54085 42327 54540 42360
rect 50481 42267 51657 42294
rect 39809 42197 43739 42243
rect 43785 42197 43906 42243
rect 43952 42197 44071 42243
rect 44117 42197 44236 42243
rect 44282 42222 44918 42243
rect 48905 42223 49877 42263
rect 50044 42257 51657 42267
rect 44282 42197 44812 42222
rect 39809 42194 44812 42197
rect 39809 42148 39844 42194
rect 39890 42192 44812 42194
rect 39890 42148 39994 42192
rect 39809 42140 39994 42148
rect 40046 42176 44812 42192
rect 44858 42176 44925 42222
rect 44971 42176 45038 42222
rect 45084 42176 45151 42222
rect 45197 42176 45264 42222
rect 45310 42176 45323 42222
rect 48557 42177 48687 42217
rect 40046 42161 44918 42176
rect 40046 42140 40085 42161
rect 39809 42137 40085 42140
rect 36924 42117 37685 42124
rect 36923 42085 37931 42117
rect 36841 42039 36854 42085
rect 36900 42083 36971 42085
rect 36900 42039 36961 42083
rect 37017 42039 37088 42085
rect 37134 42083 37206 42085
rect 37134 42039 37172 42083
rect 37252 42039 37324 42085
rect 37370 42083 37442 42085
rect 37370 42039 37384 42083
rect 36923 42031 36961 42039
rect 37013 42031 37172 42039
rect 37224 42031 37384 42039
rect 37436 42039 37442 42083
rect 37488 42083 37909 42085
rect 37488 42039 37595 42083
rect 37436 42031 37595 42039
rect 37647 42039 37909 42083
rect 37955 42039 38026 42085
rect 38072 42039 38143 42085
rect 38189 42039 38261 42085
rect 38307 42039 38379 42085
rect 38425 42039 38497 42085
rect 38543 42039 38556 42085
rect 37647 42031 37931 42039
rect 36923 41998 37931 42031
rect 36923 41997 37685 41998
rect 36924 41991 37685 41997
rect 36640 41966 36773 41989
rect 38658 41987 38669 42127
rect 38715 41987 38726 42127
rect 39014 42085 39323 42117
rect 39492 42085 39608 42117
rect 39008 42039 39021 42085
rect 39067 42039 39144 42085
rect 39190 42039 39267 42085
rect 39313 42039 39326 42085
rect 39492 42039 39641 42085
rect 39687 42039 39730 42085
rect 38658 41976 38726 41987
rect 36438 41861 36953 41886
rect 37439 41883 37931 41886
rect 37439 41861 38161 41883
rect 35260 41815 35273 41861
rect 35523 41855 35580 41861
rect 35523 41815 35543 41855
rect 35626 41815 35683 41861
rect 35729 41855 35786 41861
rect 35729 41815 35754 41855
rect 35832 41815 35889 41861
rect 35935 41855 35992 41861
rect 35935 41815 35965 41855
rect 36038 41815 36095 41861
rect 36141 41855 36198 41861
rect 36141 41815 36176 41855
rect 36244 41815 36301 41861
rect 36347 41815 36360 41861
rect 36438 41815 36854 41861
rect 36900 41815 36971 41861
rect 37017 41815 37088 41861
rect 37134 41815 37206 41861
rect 37252 41815 37324 41861
rect 37370 41815 37442 41861
rect 37488 41843 37909 41861
rect 37488 41815 37891 41843
rect 37955 41815 38026 41861
rect 38072 41843 38143 41861
rect 38123 41815 38143 41843
rect 38189 41815 38261 41861
rect 38307 41815 38379 41861
rect 38425 41815 38497 41861
rect 38543 41815 38556 41861
rect 33781 41774 34089 41809
rect 35294 41803 35332 41815
rect 35384 41803 35543 41815
rect 35595 41803 35754 41815
rect 35806 41803 35965 41815
rect 36017 41803 36176 41815
rect 36228 41803 36266 41815
rect 33671 41728 33684 41774
rect 33730 41728 33787 41774
rect 33833 41769 33890 41774
rect 33871 41728 33890 41769
rect 33936 41728 33993 41774
rect 34039 41769 34096 41774
rect 34051 41728 34096 41769
rect 34142 41728 34199 41774
rect 34245 41728 34302 41774
rect 34348 41728 34405 41774
rect 34451 41728 34508 41774
rect 34554 41728 34612 41774
rect 34658 41728 34671 41774
rect 35294 41763 36266 41803
rect 36438 41766 36953 41815
rect 37439 41791 37891 41815
rect 37943 41791 38071 41815
rect 38123 41791 38161 41815
rect 37439 41766 38161 41791
rect 37853 41750 38161 41766
rect 33781 41717 33819 41728
rect 33871 41717 33999 41728
rect 34051 41717 34089 41728
rect 33781 41676 34089 41717
rect 33484 41659 33552 41670
rect 30683 41594 31040 41628
rect 30683 41588 32842 41594
rect 30583 41553 32842 41588
rect 34247 41587 35008 41594
rect 30583 41501 30854 41553
rect 30906 41501 31065 41553
rect 31117 41501 31276 41553
rect 31328 41550 31486 41553
rect 31538 41550 31697 41553
rect 31749 41550 31909 41553
rect 31961 41550 32120 41553
rect 32172 41550 32330 41553
rect 32382 41550 32541 41553
rect 32593 41550 32752 41553
rect 32804 41550 32842 41553
rect 34246 41553 35008 41587
rect 34246 41550 34284 41553
rect 34336 41550 34495 41553
rect 34547 41550 34707 41553
rect 31328 41504 31349 41550
rect 33323 41504 33336 41550
rect 33671 41504 33684 41550
rect 33730 41504 33787 41550
rect 33833 41504 33890 41550
rect 33936 41504 33993 41550
rect 34039 41504 34096 41550
rect 34142 41504 34199 41550
rect 34245 41504 34284 41550
rect 34348 41504 34405 41550
rect 34451 41504 34495 41550
rect 34554 41504 34612 41550
rect 34658 41504 34707 41550
rect 31328 41501 31486 41504
rect 31538 41501 31697 41504
rect 31749 41501 31909 41504
rect 31961 41501 32120 41504
rect 32172 41501 32330 41504
rect 32382 41501 32541 41504
rect 32593 41501 32752 41504
rect 32804 41501 32842 41504
rect 30583 41466 32842 41501
rect 34246 41501 34284 41504
rect 34336 41501 34495 41504
rect 34547 41501 34707 41504
rect 34759 41501 34918 41553
rect 34970 41501 35008 41553
rect 34246 41467 35008 41501
rect 29544 41460 30306 41461
rect 28492 41344 29196 41420
rect 28492 41303 29116 41344
rect 28492 41257 28810 41303
rect 28856 41298 29116 41303
rect 29162 41298 29196 41344
rect 28856 41257 29196 41298
rect 28492 41181 29196 41257
rect 28492 41140 29116 41181
rect 28492 41094 28810 41140
rect 28856 41135 29116 41140
rect 29162 41135 29196 41181
rect 28856 41094 29196 41135
rect 28492 41017 29196 41094
rect 28492 40977 29116 41017
rect 28492 40931 28810 40977
rect 28856 40971 29116 40977
rect 29162 40971 29196 41017
rect 28856 40931 29196 40971
rect 28492 40854 29196 40931
rect 28492 40813 29116 40854
rect 28492 40767 28810 40813
rect 28856 40808 29116 40813
rect 29162 40808 29196 40854
rect 28856 40767 29196 40808
rect 28492 40653 29196 40767
rect 30583 41420 30637 41466
rect 30683 41460 32842 41466
rect 34247 41460 35008 41467
rect 35182 41587 36364 41594
rect 35182 41553 36958 41587
rect 35182 41501 35220 41553
rect 35272 41501 35430 41553
rect 35482 41501 35641 41553
rect 35693 41501 35853 41553
rect 35905 41501 36064 41553
rect 36116 41501 36274 41553
rect 36326 41550 36958 41553
rect 36326 41504 36489 41550
rect 36723 41504 36958 41550
rect 36326 41501 36958 41504
rect 35182 41467 36958 41501
rect 37946 41553 38842 41594
rect 37946 41550 38330 41553
rect 38382 41550 38541 41553
rect 37946 41504 37957 41550
rect 38473 41504 38541 41550
rect 37946 41501 38330 41504
rect 38382 41501 38541 41504
rect 38593 41501 38752 41553
rect 38804 41501 38842 41553
rect 35182 41460 36364 41467
rect 37946 41460 38842 41501
rect 39014 41553 39323 42039
rect 39014 41501 39052 41553
rect 39104 41550 39232 41553
rect 39108 41504 39220 41550
rect 39104 41501 39232 41504
rect 39284 41501 39323 41553
rect 30683 41426 31040 41460
rect 30683 41420 30855 41426
rect 30583 41380 30855 41420
rect 30901 41380 31040 41426
rect 30583 41303 31040 41380
rect 33484 41384 33552 41395
rect 33019 41329 33327 41370
rect 33019 41326 33057 41329
rect 33109 41326 33237 41329
rect 33289 41326 33327 41329
rect 30583 41257 30637 41303
rect 30683 41262 31040 41303
rect 31336 41280 31349 41326
rect 33323 41280 33336 41326
rect 30683 41257 30855 41262
rect 30583 41216 30855 41257
rect 30901 41216 31040 41262
rect 33019 41277 33057 41280
rect 33109 41277 33237 41280
rect 33289 41277 33327 41280
rect 33019 41237 33327 41277
rect 30583 41140 31040 41216
rect 30583 41094 30637 41140
rect 30683 41124 31040 41140
rect 30683 41102 31493 41124
rect 30683 41099 31349 41102
rect 30683 41094 30855 41099
rect 30583 41053 30855 41094
rect 30901 41056 31349 41099
rect 33323 41056 33336 41102
rect 30901 41053 31493 41056
rect 30583 41005 31493 41053
rect 30583 40977 31040 41005
rect 30583 40931 30637 40977
rect 30683 40936 31040 40977
rect 30683 40931 30855 40936
rect 30583 40890 30855 40931
rect 30901 40890 31040 40936
rect 33484 40962 33495 41384
rect 33541 40962 33552 41384
rect 33781 41337 34089 41378
rect 33781 41326 33819 41337
rect 33871 41326 33999 41337
rect 34051 41326 34089 41337
rect 33671 41280 33684 41326
rect 33730 41280 33787 41326
rect 33871 41285 33890 41326
rect 33833 41280 33890 41285
rect 33936 41280 33993 41326
rect 34051 41285 34096 41326
rect 34039 41280 34096 41285
rect 34142 41280 34199 41326
rect 34245 41280 34302 41326
rect 34348 41280 34405 41326
rect 34451 41280 34508 41326
rect 34554 41280 34612 41326
rect 34658 41280 34671 41326
rect 33781 41245 34089 41280
rect 35294 41251 36266 41291
rect 37853 41288 38161 41304
rect 35294 41239 35332 41251
rect 35384 41239 35543 41251
rect 35595 41239 35754 41251
rect 35806 41239 35965 41251
rect 36017 41239 36176 41251
rect 36228 41239 36266 41251
rect 36438 41239 36953 41288
rect 37439 41263 38161 41288
rect 37439 41239 37891 41263
rect 37943 41239 38071 41263
rect 38123 41239 38161 41263
rect 35260 41193 35273 41239
rect 35523 41199 35543 41239
rect 35523 41193 35580 41199
rect 35626 41193 35683 41239
rect 35729 41199 35754 41239
rect 35729 41193 35786 41199
rect 35832 41193 35889 41239
rect 35935 41199 35965 41239
rect 35935 41193 35992 41199
rect 36038 41193 36095 41239
rect 36141 41199 36176 41239
rect 36141 41193 36198 41199
rect 36244 41193 36301 41239
rect 36347 41193 36360 41239
rect 36438 41193 36854 41239
rect 36900 41193 36971 41239
rect 37017 41193 37088 41239
rect 37134 41193 37206 41239
rect 37252 41193 37324 41239
rect 37370 41193 37442 41239
rect 37488 41211 37891 41239
rect 37488 41193 37909 41211
rect 37955 41193 38026 41239
rect 38123 41211 38143 41239
rect 38072 41193 38143 41211
rect 38189 41193 38261 41239
rect 38307 41193 38379 41239
rect 38425 41193 38497 41239
rect 38543 41193 38556 41239
rect 35294 41159 36266 41193
rect 36438 41168 36953 41193
rect 37439 41171 38161 41193
rect 37439 41168 37931 41171
rect 34228 41102 34718 41131
rect 33671 41056 33684 41102
rect 33730 41056 33787 41102
rect 33833 41056 33890 41102
rect 33936 41056 33993 41102
rect 34039 41056 34096 41102
rect 34142 41056 34199 41102
rect 34245 41091 34302 41102
rect 34245 41056 34267 41091
rect 34348 41056 34405 41102
rect 34451 41091 34508 41102
rect 34499 41056 34508 41091
rect 34554 41056 34612 41102
rect 34658 41091 34718 41102
rect 34228 41039 34267 41056
rect 34319 41039 34447 41056
rect 34499 41039 34627 41056
rect 34679 41039 34718 41091
rect 36438 41065 36554 41168
rect 34228 40998 34718 41039
rect 34964 41015 36360 41059
rect 30583 40813 31040 40890
rect 33019 40881 33327 40922
rect 33019 40878 33057 40881
rect 33109 40878 33237 40881
rect 33289 40878 33327 40881
rect 33484 40880 33552 40962
rect 34964 40969 35273 41015
rect 35523 40969 35580 41015
rect 35626 40969 35683 41015
rect 35729 40969 35786 41015
rect 35832 40969 35889 41015
rect 35935 40969 35992 41015
rect 36038 40969 36095 41015
rect 36141 40969 36198 41015
rect 36244 40969 36301 41015
rect 36347 40969 36360 41015
rect 34964 40937 36360 40969
rect 34964 40880 35082 40937
rect 31336 40832 31349 40878
rect 33323 40832 33336 40878
rect 33484 40843 35082 40880
rect 30583 40767 30637 40813
rect 30683 40773 31040 40813
rect 33019 40829 33057 40832
rect 33109 40829 33237 40832
rect 33289 40829 33327 40832
rect 33019 40789 33327 40829
rect 33484 40797 33816 40843
rect 33862 40797 34002 40843
rect 34048 40797 34189 40843
rect 34235 40797 34376 40843
rect 34422 40797 34562 40843
rect 34608 40797 35082 40843
rect 36438 40925 36475 41065
rect 36521 40925 36554 41065
rect 33484 40789 35082 40797
rect 35294 40791 36266 40831
rect 36438 40825 36554 40925
rect 36640 41065 36773 41088
rect 36640 41016 36697 41065
rect 36640 40964 36678 41016
rect 36640 40925 36697 40964
rect 36743 40925 36773 41065
rect 38658 41067 38726 41078
rect 36924 41057 37685 41063
rect 36923 41056 37685 41057
rect 36923 41023 37931 41056
rect 36923 41015 36961 41023
rect 37013 41015 37172 41023
rect 37224 41015 37384 41023
rect 36841 40969 36854 41015
rect 36900 40971 36961 41015
rect 36900 40969 36971 40971
rect 37017 40969 37088 41015
rect 37134 40971 37172 41015
rect 37134 40969 37206 40971
rect 37252 40969 37324 41015
rect 37370 40971 37384 41015
rect 37436 41015 37595 41023
rect 37436 40971 37442 41015
rect 37370 40969 37442 40971
rect 37488 40971 37595 41015
rect 37647 41015 37931 41023
rect 37647 40971 37909 41015
rect 37488 40969 37909 40971
rect 37955 40969 38026 41015
rect 38072 40969 38143 41015
rect 38189 40969 38261 41015
rect 38307 40969 38379 41015
rect 38425 40969 38497 41015
rect 38543 40969 38556 41015
rect 36923 40937 37931 40969
rect 36924 40930 37685 40937
rect 36640 40905 36773 40925
rect 38658 40927 38669 41067
rect 38715 40927 38726 41067
rect 39014 41015 39323 41501
rect 39492 41587 39608 42039
rect 39923 42006 40085 42137
rect 39923 41954 39994 42006
rect 40046 41954 40085 42006
rect 39923 41914 40085 41954
rect 39737 41818 39865 41831
rect 39737 41791 39866 41818
rect 39737 41774 39775 41791
rect 39827 41774 39866 41791
rect 39727 41728 39740 41774
rect 39827 41739 39862 41774
rect 39786 41728 39862 41739
rect 39908 41728 39985 41774
rect 40031 41728 40108 41774
rect 40154 41728 40167 41774
rect 40246 41763 40362 42161
rect 42229 42022 44509 42063
rect 42229 41970 43445 42022
rect 43497 41970 44509 42022
rect 42229 41930 44509 41970
rect 44341 41886 44509 41930
rect 44341 41840 44358 41886
rect 44498 41840 44509 41886
rect 39737 41699 39866 41728
rect 40246 41717 40281 41763
rect 40327 41717 40362 41763
rect 40246 41680 40362 41717
rect 40718 41791 43524 41832
rect 44341 41829 44509 41840
rect 40718 41739 41935 41791
rect 41987 41739 43524 41791
rect 40718 41698 43524 41739
rect 44605 41774 44721 42161
rect 45400 42131 48379 42172
rect 45400 42117 45975 42131
rect 45400 42071 45464 42117
rect 45604 42079 45975 42117
rect 46027 42079 48379 42131
rect 45604 42071 48379 42079
rect 44901 42015 45241 42056
rect 45400 42038 48379 42071
rect 48557 42125 48596 42177
rect 48648 42125 48687 42177
rect 48557 42102 48687 42125
rect 50044 42211 50516 42257
rect 50562 42211 50703 42257
rect 50749 42211 50890 42257
rect 50936 42211 51076 42257
rect 51122 42211 51263 42257
rect 51309 42211 51657 42257
rect 51797 42247 52105 42287
rect 51797 42222 51835 42247
rect 51887 42222 52015 42247
rect 52067 42222 52105 42247
rect 54085 42281 54223 42327
rect 54269 42287 54540 42327
rect 54269 42281 54440 42287
rect 54085 42241 54440 42281
rect 54486 42241 54540 42287
rect 50044 42174 51657 42211
rect 51789 42176 51802 42222
rect 53776 42176 53789 42222
rect 50044 42117 50160 42174
rect 44901 41998 44939 42015
rect 44991 41998 45151 42015
rect 45203 41998 45241 42015
rect 44799 41952 44812 41998
rect 44858 41952 44925 41998
rect 44991 41963 45038 41998
rect 44971 41952 45038 41963
rect 45084 41952 45151 41998
rect 45203 41963 45264 41998
rect 45197 41952 45264 41963
rect 45310 41952 45323 41998
rect 48557 41962 48622 42102
rect 48668 41962 48687 42102
rect 49820 42085 50160 42117
rect 48765 42039 48778 42085
rect 48824 42039 48881 42085
rect 48927 42039 48984 42085
rect 49030 42039 49087 42085
rect 49133 42039 49190 42085
rect 49236 42039 49293 42085
rect 49339 42039 49396 42085
rect 49442 42039 49499 42085
rect 49545 42039 49602 42085
rect 49852 42039 50160 42085
rect 51589 42122 51657 42174
rect 51797 42154 52105 42176
rect 49820 41998 50160 42039
rect 50262 42015 50812 42056
rect 48557 41959 48687 41962
rect 44901 41923 45241 41952
rect 48557 41907 48596 41959
rect 48648 41907 48687 41959
rect 50262 41963 50300 42015
rect 50352 41998 50511 42015
rect 50563 41998 50722 42015
rect 50352 41963 50467 41998
rect 50563 41963 50571 41998
rect 50262 41952 50467 41963
rect 50513 41952 50571 41963
rect 50617 41952 50674 41998
rect 50720 41963 50722 41998
rect 50774 41998 50812 42015
rect 50774 41963 50777 41998
rect 50720 41952 50777 41963
rect 50823 41952 50880 41998
rect 50926 41952 50983 41998
rect 51029 41952 51086 41998
rect 51132 41952 51189 41998
rect 51235 41952 51292 41998
rect 51338 41952 51395 41998
rect 51441 41952 51454 41998
rect 50262 41923 50812 41952
rect 48557 41866 48687 41907
rect 48905 41861 49877 41892
rect 48765 41815 48778 41861
rect 48824 41815 48881 41861
rect 48927 41852 48984 41861
rect 48927 41815 48943 41852
rect 49030 41815 49087 41861
rect 49133 41852 49190 41861
rect 49133 41815 49154 41852
rect 49236 41815 49293 41861
rect 49339 41852 49396 41861
rect 49339 41815 49365 41852
rect 49442 41815 49499 41861
rect 49545 41852 49602 41861
rect 49545 41815 49576 41852
rect 49852 41815 49877 41861
rect 48905 41800 48943 41815
rect 48995 41800 49154 41815
rect 49206 41800 49365 41815
rect 49417 41800 49576 41815
rect 49628 41800 49787 41815
rect 49839 41800 49877 41815
rect 44605 41728 44812 41774
rect 44858 41728 44925 41774
rect 44971 41728 45038 41774
rect 45084 41728 45151 41774
rect 45197 41728 45264 41774
rect 45310 41728 45323 41774
rect 48905 41760 49877 41800
rect 51035 41777 51343 41817
rect 51035 41774 51073 41777
rect 51125 41774 51253 41777
rect 51305 41774 51343 41777
rect 43362 41691 43524 41698
rect 43362 41645 43373 41691
rect 43513 41645 43524 41691
rect 43362 41634 43524 41645
rect 45584 41714 48546 41750
rect 50454 41728 50467 41774
rect 50513 41728 50571 41774
rect 50617 41728 50674 41774
rect 50720 41728 50777 41774
rect 50823 41728 50880 41774
rect 50926 41728 50983 41774
rect 51029 41728 51073 41774
rect 51132 41728 51189 41774
rect 51235 41728 51253 41774
rect 51338 41728 51395 41774
rect 51441 41728 51454 41774
rect 45584 41668 45619 41714
rect 45665 41668 45777 41714
rect 45823 41668 45935 41714
rect 45981 41668 46093 41714
rect 46139 41668 46251 41714
rect 46297 41668 46409 41714
rect 46455 41668 46568 41714
rect 46614 41668 46726 41714
rect 46772 41668 46884 41714
rect 46930 41668 47042 41714
rect 47088 41668 47200 41714
rect 47246 41668 47358 41714
rect 47404 41668 47516 41714
rect 47562 41668 47675 41714
rect 47721 41668 47833 41714
rect 47879 41668 47991 41714
rect 48037 41668 48149 41714
rect 48195 41668 48307 41714
rect 48353 41668 48465 41714
rect 48511 41668 48546 41714
rect 51035 41725 51073 41728
rect 51125 41725 51253 41728
rect 51305 41725 51343 41728
rect 51035 41684 51343 41725
rect 51589 41700 51600 42122
rect 51646 41700 51657 42122
rect 54085 42123 54540 42241
rect 54085 42077 54440 42123
rect 54486 42077 54540 42123
rect 54085 42049 54540 42077
rect 53585 41998 54540 42049
rect 51789 41952 51802 41998
rect 53776 41960 54540 41998
rect 53776 41952 54440 41960
rect 53585 41930 54440 41952
rect 54085 41914 54440 41930
rect 54486 41914 54540 41960
rect 54085 41838 54540 41914
rect 51797 41784 52105 41824
rect 51797 41774 51835 41784
rect 51887 41774 52015 41784
rect 52067 41774 52105 41784
rect 54085 41792 54223 41838
rect 54269 41797 54540 41838
rect 54269 41792 54440 41797
rect 51789 41728 51802 41774
rect 53776 41728 53789 41774
rect 54085 41751 54440 41792
rect 54486 41751 54540 41797
rect 51589 41689 51657 41700
rect 51797 41691 52105 41728
rect 40215 41587 40523 41594
rect 40788 41587 42986 41601
rect 43753 41587 44514 41594
rect 39492 41564 42986 41587
rect 43704 41564 44514 41587
rect 39492 41553 44514 41564
rect 39492 41550 40253 41553
rect 39492 41504 39740 41550
rect 39786 41504 39862 41550
rect 39908 41504 39985 41550
rect 40031 41504 40108 41550
rect 40154 41504 40253 41550
rect 39492 41501 40253 41504
rect 40305 41501 40433 41553
rect 40485 41550 43790 41553
rect 40485 41504 40836 41550
rect 40882 41504 40994 41550
rect 41040 41504 41152 41550
rect 41198 41504 41310 41550
rect 41356 41504 41469 41550
rect 41515 41504 41627 41550
rect 41673 41504 41785 41550
rect 41831 41504 41943 41550
rect 41989 41504 42101 41550
rect 42147 41504 42259 41550
rect 42305 41504 42418 41550
rect 42464 41504 42576 41550
rect 42622 41504 42734 41550
rect 42780 41504 42892 41550
rect 42938 41504 43739 41550
rect 43785 41504 43790 41550
rect 40485 41501 43790 41504
rect 43842 41550 44001 41553
rect 43842 41504 43906 41550
rect 43952 41504 44001 41550
rect 43842 41501 44001 41504
rect 44053 41550 44213 41553
rect 44265 41550 44424 41553
rect 44053 41504 44071 41550
rect 44117 41504 44213 41550
rect 44282 41504 44424 41550
rect 44053 41501 44213 41504
rect 44265 41501 44424 41504
rect 44476 41501 44514 41553
rect 39492 41490 44514 41501
rect 39492 41467 42986 41490
rect 43704 41467 44514 41490
rect 39492 41015 39608 41467
rect 40215 41460 40523 41467
rect 40788 41453 42986 41467
rect 43753 41460 44514 41467
rect 44796 41587 45346 41594
rect 45584 41587 48546 41668
rect 54085 41674 54540 41751
rect 54085 41628 54223 41674
rect 54269 41634 54540 41674
rect 54269 41628 54440 41634
rect 54085 41594 54440 41628
rect 48800 41587 49982 41594
rect 50308 41587 50859 41594
rect 44796 41553 49982 41587
rect 44796 41550 44834 41553
rect 44886 41550 45045 41553
rect 45097 41550 45256 41553
rect 45308 41550 48838 41553
rect 44796 41504 44812 41550
rect 44886 41504 44925 41550
rect 44971 41504 45038 41550
rect 45097 41504 45151 41550
rect 45197 41504 45256 41550
rect 45310 41504 45619 41550
rect 45665 41504 45777 41550
rect 45823 41504 45935 41550
rect 45981 41504 46093 41550
rect 46139 41504 46251 41550
rect 46297 41504 46409 41550
rect 46455 41504 46568 41550
rect 46614 41504 46726 41550
rect 46772 41504 46884 41550
rect 46930 41504 47042 41550
rect 47088 41504 47200 41550
rect 47246 41504 47358 41550
rect 47404 41504 47516 41550
rect 47562 41504 47675 41550
rect 47721 41504 47833 41550
rect 47879 41504 47991 41550
rect 48037 41504 48149 41550
rect 48195 41504 48307 41550
rect 48353 41504 48465 41550
rect 48511 41504 48838 41550
rect 44796 41501 44834 41504
rect 44886 41501 45045 41504
rect 45097 41501 45256 41504
rect 45308 41501 48838 41504
rect 48890 41501 49048 41553
rect 49100 41501 49259 41553
rect 49311 41501 49471 41553
rect 49523 41501 49682 41553
rect 49734 41501 49892 41553
rect 49944 41501 49982 41553
rect 44796 41467 49982 41501
rect 50307 41553 50859 41587
rect 50307 41501 50346 41553
rect 50398 41550 50557 41553
rect 50609 41550 50768 41553
rect 50820 41550 50859 41553
rect 52278 41588 54440 41594
rect 54486 41588 54540 41634
rect 55927 42287 56632 42401
rect 55927 42244 56267 42287
rect 55927 42198 55961 42244
rect 56007 42241 56267 42244
rect 56313 42241 56632 42287
rect 56007 42198 56632 42241
rect 55927 42123 56632 42198
rect 55927 42081 56267 42123
rect 55927 42035 55961 42081
rect 56007 42077 56267 42081
rect 56313 42077 56632 42123
rect 56007 42035 56632 42077
rect 55927 41960 56632 42035
rect 55927 41917 56267 41960
rect 55927 41871 55961 41917
rect 56007 41914 56267 41917
rect 56313 41914 56632 41960
rect 56007 41871 56632 41914
rect 55927 41797 56632 41871
rect 55927 41754 56267 41797
rect 55927 41708 55961 41754
rect 56007 41751 56267 41754
rect 56313 41751 56632 41797
rect 56007 41708 56632 41751
rect 55927 41634 56632 41708
rect 52278 41553 54540 41588
rect 52278 41550 52316 41553
rect 52368 41550 52527 41553
rect 52579 41550 52738 41553
rect 52790 41550 52948 41553
rect 53000 41550 53159 41553
rect 53211 41550 53371 41553
rect 53423 41550 53582 41553
rect 53634 41550 53792 41553
rect 50398 41504 50467 41550
rect 50513 41504 50557 41550
rect 50617 41504 50674 41550
rect 50720 41504 50768 41550
rect 50823 41504 50880 41550
rect 50926 41504 50983 41550
rect 51029 41504 51086 41550
rect 51132 41504 51189 41550
rect 51235 41504 51292 41550
rect 51338 41504 51395 41550
rect 51441 41504 51454 41550
rect 51789 41504 51802 41550
rect 53776 41504 53792 41550
rect 50398 41501 50557 41504
rect 50609 41501 50768 41504
rect 50820 41501 50859 41504
rect 50307 41467 50859 41501
rect 44796 41460 45346 41467
rect 43362 41409 43524 41420
rect 39737 41326 39866 41355
rect 40246 41337 40362 41374
rect 43362 41363 43373 41409
rect 43513 41363 43524 41409
rect 43362 41356 43524 41363
rect 39727 41280 39740 41326
rect 39786 41315 39862 41326
rect 39827 41280 39862 41315
rect 39908 41280 39985 41326
rect 40031 41280 40108 41326
rect 40154 41280 40167 41326
rect 40246 41291 40281 41337
rect 40327 41291 40362 41337
rect 39737 41263 39775 41280
rect 39827 41263 39866 41280
rect 39737 41236 39866 41263
rect 39737 41223 39865 41236
rect 39923 41100 40085 41140
rect 39923 41048 39994 41100
rect 40046 41048 40085 41100
rect 39008 40969 39021 41015
rect 39067 40969 39144 41015
rect 39190 40969 39267 41015
rect 39313 40969 39326 41015
rect 39492 40969 39641 41015
rect 39687 40969 39730 41015
rect 39014 40937 39323 40969
rect 39492 40937 39608 40969
rect 37853 40825 38161 40830
rect 36438 40791 36953 40825
rect 37439 40791 38161 40825
rect 38658 40805 38726 40927
rect 39923 40917 40085 41048
rect 39809 40914 40085 40917
rect 39809 40906 39994 40914
rect 39809 40860 39844 40906
rect 39890 40862 39994 40906
rect 40046 40893 40085 40914
rect 40246 40893 40362 41291
rect 40718 41315 43524 41356
rect 45584 41386 48546 41467
rect 48800 41460 49982 41467
rect 50308 41460 50859 41467
rect 52278 41501 52316 41504
rect 52368 41501 52527 41504
rect 52579 41501 52738 41504
rect 52790 41501 52948 41504
rect 53000 41501 53159 41504
rect 53211 41501 53371 41504
rect 53423 41501 53582 41504
rect 53634 41501 53792 41504
rect 53844 41501 54003 41553
rect 54055 41501 54214 41553
rect 54266 41501 54540 41553
rect 52278 41466 54540 41501
rect 52278 41460 54440 41466
rect 45584 41340 45619 41386
rect 45665 41340 45777 41386
rect 45823 41340 45935 41386
rect 45981 41340 46093 41386
rect 46139 41340 46251 41386
rect 46297 41340 46409 41386
rect 46455 41340 46568 41386
rect 46614 41340 46726 41386
rect 46772 41340 46884 41386
rect 46930 41340 47042 41386
rect 47088 41340 47200 41386
rect 47246 41340 47358 41386
rect 47404 41340 47516 41386
rect 47562 41340 47675 41386
rect 47721 41340 47833 41386
rect 47879 41340 47991 41386
rect 48037 41340 48149 41386
rect 48195 41340 48307 41386
rect 48353 41340 48465 41386
rect 48511 41340 48546 41386
rect 54085 41426 54440 41460
rect 54085 41380 54223 41426
rect 54269 41420 54440 41426
rect 54486 41420 54540 41466
rect 54758 41553 55840 41594
rect 54758 41550 54855 41553
rect 54758 41504 54793 41550
rect 54839 41504 54855 41550
rect 54758 41501 54855 41504
rect 54907 41550 55066 41553
rect 54907 41504 54956 41550
rect 55002 41504 55066 41550
rect 54907 41501 55066 41504
rect 55118 41550 55278 41553
rect 55330 41550 55489 41553
rect 55164 41504 55278 41550
rect 55330 41504 55439 41550
rect 55485 41504 55489 41550
rect 55118 41501 55278 41504
rect 55330 41501 55489 41504
rect 55541 41550 55840 41553
rect 55541 41504 55599 41550
rect 55645 41504 55760 41550
rect 55806 41504 55840 41550
rect 55541 41501 55840 41504
rect 54758 41461 55840 41501
rect 55927 41588 56267 41634
rect 56313 41588 56632 41634
rect 55927 41466 56632 41588
rect 54817 41460 55579 41461
rect 54269 41380 54540 41420
rect 40718 41263 41935 41315
rect 41987 41263 43524 41315
rect 40718 41222 43524 41263
rect 44605 41280 44812 41326
rect 44858 41280 44925 41326
rect 44971 41280 45038 41326
rect 45084 41280 45151 41326
rect 45197 41280 45264 41326
rect 45310 41280 45323 41326
rect 45584 41304 48546 41340
rect 51035 41329 51343 41370
rect 51035 41326 51073 41329
rect 51125 41326 51253 41329
rect 51305 41326 51343 41329
rect 51589 41354 51657 41365
rect 44341 41214 44509 41225
rect 44341 41168 44358 41214
rect 44498 41168 44509 41214
rect 44341 41124 44509 41168
rect 42229 41084 44509 41124
rect 42229 41032 43445 41084
rect 43497 41032 44509 41084
rect 42229 40991 44509 41032
rect 44605 40893 44721 41280
rect 48905 41254 49877 41294
rect 50454 41280 50467 41326
rect 50513 41280 50571 41326
rect 50617 41280 50674 41326
rect 50720 41280 50777 41326
rect 50823 41280 50880 41326
rect 50926 41280 50983 41326
rect 51029 41280 51073 41326
rect 51132 41280 51189 41326
rect 51235 41280 51253 41326
rect 51338 41280 51395 41326
rect 51441 41280 51454 41326
rect 48905 41239 48943 41254
rect 48995 41239 49154 41254
rect 49206 41239 49365 41254
rect 49417 41239 49576 41254
rect 49628 41239 49787 41254
rect 49839 41239 49877 41254
rect 48765 41193 48778 41239
rect 48824 41193 48881 41239
rect 48927 41202 48943 41239
rect 48927 41193 48984 41202
rect 49030 41193 49087 41239
rect 49133 41202 49154 41239
rect 49133 41193 49190 41202
rect 49236 41193 49293 41239
rect 49339 41202 49365 41239
rect 49339 41193 49396 41202
rect 49442 41193 49499 41239
rect 49545 41202 49576 41239
rect 49545 41193 49602 41202
rect 49852 41193 49877 41239
rect 51035 41277 51073 41280
rect 51125 41277 51253 41280
rect 51305 41277 51343 41280
rect 51035 41237 51343 41277
rect 48557 41147 48687 41188
rect 48905 41162 49877 41193
rect 44901 41102 45241 41131
rect 44799 41056 44812 41102
rect 44858 41056 44925 41102
rect 44971 41091 45038 41102
rect 44991 41056 45038 41091
rect 45084 41056 45151 41102
rect 45197 41091 45264 41102
rect 45203 41056 45264 41091
rect 45310 41056 45323 41102
rect 48557 41095 48596 41147
rect 48648 41095 48687 41147
rect 48557 41092 48687 41095
rect 44901 41039 44939 41056
rect 44991 41039 45151 41056
rect 45203 41039 45241 41056
rect 44901 40998 45241 41039
rect 45400 40983 48379 41016
rect 45400 40937 45464 40983
rect 45604 40975 48379 40983
rect 45604 40937 46353 40975
rect 45400 40923 46353 40937
rect 46405 40923 48379 40975
rect 40046 40878 44918 40893
rect 45400 40882 48379 40923
rect 48557 40952 48622 41092
rect 48668 40952 48687 41092
rect 50262 41102 50812 41131
rect 50262 41091 50467 41102
rect 50513 41091 50571 41102
rect 49820 41015 50160 41056
rect 48765 40969 48778 41015
rect 48824 40969 48881 41015
rect 48927 40969 48984 41015
rect 49030 40969 49087 41015
rect 49133 40969 49190 41015
rect 49236 40969 49293 41015
rect 49339 40969 49396 41015
rect 49442 40969 49499 41015
rect 49545 40969 49602 41015
rect 49852 40969 50160 41015
rect 50262 41039 50300 41091
rect 50352 41056 50467 41091
rect 50563 41056 50571 41091
rect 50617 41056 50674 41102
rect 50720 41091 50777 41102
rect 50720 41056 50722 41091
rect 50352 41039 50511 41056
rect 50563 41039 50722 41056
rect 50774 41056 50777 41091
rect 50823 41056 50880 41102
rect 50926 41056 50983 41102
rect 51029 41056 51086 41102
rect 51132 41056 51189 41102
rect 51235 41056 51292 41102
rect 51338 41056 51395 41102
rect 51441 41056 51454 41102
rect 50774 41039 50812 41056
rect 50262 40998 50812 41039
rect 48557 40929 48687 40952
rect 49820 40937 50160 40969
rect 40046 40862 44812 40878
rect 39890 40860 44812 40862
rect 39809 40857 44812 40860
rect 39809 40811 43739 40857
rect 43785 40811 43906 40857
rect 43952 40811 44071 40857
rect 44117 40811 44236 40857
rect 44282 40832 44812 40857
rect 44858 40832 44925 40878
rect 44971 40832 45038 40878
rect 45084 40832 45151 40878
rect 45197 40832 45264 40878
rect 45310 40832 45323 40878
rect 48557 40877 48596 40929
rect 48648 40877 48687 40929
rect 48557 40837 48687 40877
rect 50044 40880 50160 40937
rect 51589 40932 51600 41354
rect 51646 40932 51657 41354
rect 51797 41326 52105 41363
rect 51789 41280 51802 41326
rect 53776 41280 53789 41326
rect 54085 41303 54540 41380
rect 51797 41270 51835 41280
rect 51887 41270 52015 41280
rect 52067 41270 52105 41280
rect 51797 41230 52105 41270
rect 54085 41262 54440 41303
rect 54085 41216 54223 41262
rect 54269 41257 54440 41262
rect 54486 41257 54540 41303
rect 54269 41216 54540 41257
rect 54085 41140 54540 41216
rect 54085 41124 54440 41140
rect 53585 41102 54440 41124
rect 51789 41056 51802 41102
rect 53776 41094 54440 41102
rect 54486 41094 54540 41140
rect 53776 41056 54540 41094
rect 53585 41005 54540 41056
rect 51589 40880 51657 40932
rect 54085 40977 54540 41005
rect 54085 40931 54440 40977
rect 54486 40931 54540 40977
rect 50044 40843 51657 40880
rect 51797 40878 52105 40900
rect 44282 40811 44918 40832
rect 38658 40791 39723 40805
rect 30683 40767 30855 40773
rect 30583 40727 30855 40767
rect 30901 40727 31040 40773
rect 33484 40760 34643 40789
rect 35260 40745 35273 40791
rect 35523 40745 35543 40791
rect 35626 40745 35683 40791
rect 35729 40745 35754 40791
rect 35832 40745 35889 40791
rect 35935 40745 35965 40791
rect 36038 40745 36095 40791
rect 36141 40745 36176 40791
rect 36244 40745 36301 40791
rect 36347 40745 36360 40791
rect 36438 40745 36854 40791
rect 36900 40745 36971 40791
rect 37017 40745 37088 40791
rect 37134 40745 37206 40791
rect 37252 40745 37324 40791
rect 37370 40745 37442 40791
rect 37488 40789 37909 40791
rect 37488 40745 37891 40789
rect 37955 40745 38026 40791
rect 38072 40789 38143 40791
rect 38123 40745 38143 40789
rect 38189 40745 38261 40791
rect 38307 40745 38379 40791
rect 38425 40745 38497 40791
rect 38543 40745 38556 40791
rect 38658 40745 39021 40791
rect 39067 40745 39144 40791
rect 39190 40745 39267 40791
rect 39313 40745 39641 40791
rect 39687 40745 39730 40791
rect 39809 40773 44918 40811
rect 48905 40791 49877 40831
rect 48765 40745 48778 40791
rect 48824 40745 48881 40791
rect 48927 40745 48943 40791
rect 49030 40745 49087 40791
rect 49133 40745 49154 40791
rect 49236 40745 49293 40791
rect 49339 40745 49365 40791
rect 49442 40745 49499 40791
rect 49545 40745 49576 40791
rect 49852 40745 49877 40791
rect 50044 40797 50516 40843
rect 50562 40797 50703 40843
rect 50749 40797 50890 40843
rect 50936 40797 51076 40843
rect 51122 40797 51263 40843
rect 51309 40797 51657 40843
rect 51789 40832 51802 40878
rect 53776 40832 53789 40878
rect 50044 40787 51657 40797
rect 50481 40760 51657 40787
rect 51797 40807 51835 40832
rect 51887 40807 52015 40832
rect 52067 40807 52105 40832
rect 51797 40767 52105 40807
rect 54085 40813 54540 40931
rect 54085 40773 54440 40813
rect 30583 40694 31040 40727
rect 35294 40739 35332 40745
rect 35384 40739 35543 40745
rect 35595 40739 35754 40745
rect 35806 40739 35965 40745
rect 36017 40739 36176 40745
rect 36228 40739 36266 40745
rect 34870 40694 35025 40701
rect 35294 40699 36266 40739
rect 36438 40705 36953 40745
rect 37439 40737 37891 40745
rect 37943 40737 38071 40745
rect 38123 40737 38161 40745
rect 37439 40705 38161 40737
rect 37853 40697 38161 40705
rect 27744 40601 27790 40653
rect 27842 40601 27846 40653
rect 28492 40601 28634 40653
rect 28686 40650 28845 40653
rect 28686 40604 28810 40650
rect 28686 40601 28845 40604
rect 28897 40601 29056 40653
rect 29108 40601 29196 40653
rect 27744 38853 27846 40601
rect 28492 40487 29196 40601
rect 29283 40653 30365 40694
rect 29283 40650 29582 40653
rect 29283 40604 29317 40650
rect 29363 40604 29478 40650
rect 29524 40604 29582 40650
rect 29283 40601 29582 40604
rect 29634 40650 29793 40653
rect 29845 40650 30005 40653
rect 29634 40604 29638 40650
rect 29684 40604 29793 40650
rect 29845 40604 29959 40650
rect 29634 40601 29793 40604
rect 29845 40601 30005 40604
rect 30057 40650 30216 40653
rect 30057 40604 30121 40650
rect 30167 40604 30216 40650
rect 30057 40601 30216 40604
rect 30268 40650 30365 40653
rect 30268 40604 30284 40650
rect 30330 40604 30365 40650
rect 30268 40601 30365 40604
rect 29283 40561 30365 40601
rect 30583 40653 32842 40694
rect 30583 40650 30854 40653
rect 30583 40604 30637 40650
rect 30683 40604 30854 40650
rect 30583 40601 30854 40604
rect 30906 40601 31065 40653
rect 31117 40601 31276 40653
rect 31328 40601 31486 40653
rect 31538 40601 31697 40653
rect 31749 40601 31909 40653
rect 31961 40601 32120 40653
rect 32172 40601 32330 40653
rect 32382 40601 32541 40653
rect 32593 40601 32752 40653
rect 32804 40601 32842 40653
rect 29544 40560 30306 40561
rect 30583 40560 32842 40601
rect 34717 40653 35025 40694
rect 38658 40685 39723 40745
rect 48905 40739 48943 40745
rect 48995 40739 49154 40745
rect 49206 40739 49365 40745
rect 49417 40739 49576 40745
rect 49628 40739 49787 40745
rect 49839 40739 49877 40745
rect 48905 40699 49877 40739
rect 54085 40727 54223 40773
rect 54269 40767 54440 40773
rect 54486 40767 54540 40813
rect 54269 40727 54540 40767
rect 50099 40694 50255 40701
rect 54085 40694 54540 40727
rect 55927 41420 56267 41466
rect 56313 41420 56632 41466
rect 55927 41344 56632 41420
rect 55927 41298 55961 41344
rect 56007 41303 56632 41344
rect 56007 41298 56267 41303
rect 55927 41257 56267 41298
rect 56313 41257 56632 41303
rect 55927 41181 56632 41257
rect 55927 41135 55961 41181
rect 56007 41140 56632 41181
rect 56007 41135 56267 41140
rect 55927 41094 56267 41135
rect 56313 41094 56632 41140
rect 55927 41017 56632 41094
rect 55927 40971 55961 41017
rect 56007 40977 56632 41017
rect 56007 40971 56267 40977
rect 55927 40931 56267 40971
rect 56313 40931 56632 40977
rect 55927 40854 56632 40931
rect 55927 40808 55961 40854
rect 56007 40813 56632 40854
rect 56007 40808 56267 40813
rect 55927 40767 56267 40808
rect 56313 40767 56632 40813
rect 34717 40601 34755 40653
rect 34807 40650 34935 40653
rect 34807 40604 34916 40650
rect 34807 40601 34935 40604
rect 34987 40601 35025 40653
rect 34717 40560 35025 40601
rect 50099 40653 50408 40694
rect 50099 40601 50138 40653
rect 50190 40650 50318 40653
rect 50206 40604 50318 40650
rect 50190 40601 50318 40604
rect 50370 40601 50408 40653
rect 28492 40441 28810 40487
rect 28856 40444 29196 40487
rect 28856 40441 29116 40444
rect 28492 40398 29116 40441
rect 29162 40398 29196 40444
rect 28492 40323 29196 40398
rect 28492 40277 28810 40323
rect 28856 40281 29196 40323
rect 28856 40277 29116 40281
rect 28492 40235 29116 40277
rect 29162 40235 29196 40281
rect 28492 40160 29196 40235
rect 28492 40114 28810 40160
rect 28856 40117 29196 40160
rect 28856 40114 29116 40117
rect 28492 40071 29116 40114
rect 29162 40071 29196 40117
rect 28492 39997 29196 40071
rect 28492 39951 28810 39997
rect 28856 39954 29196 39997
rect 28856 39951 29116 39954
rect 28492 39908 29116 39951
rect 29162 39908 29196 39954
rect 28492 39834 29196 39908
rect 28492 39788 28810 39834
rect 28856 39788 29196 39834
rect 30583 40527 31040 40560
rect 34870 40553 35025 40560
rect 30583 40487 30855 40527
rect 30583 40441 30637 40487
rect 30683 40481 30855 40487
rect 30901 40481 31040 40527
rect 35294 40515 36266 40555
rect 37853 40549 38161 40557
rect 35294 40509 35332 40515
rect 35384 40509 35543 40515
rect 35595 40509 35754 40515
rect 35806 40509 35965 40515
rect 36017 40509 36176 40515
rect 36228 40509 36266 40515
rect 36438 40509 36953 40549
rect 37439 40517 38161 40549
rect 37439 40509 37891 40517
rect 37943 40509 38071 40517
rect 38123 40509 38161 40517
rect 38658 40509 39723 40569
rect 50099 40560 50408 40601
rect 52278 40653 54540 40694
rect 52278 40601 52316 40653
rect 52368 40601 52527 40653
rect 52579 40601 52738 40653
rect 52790 40601 52948 40653
rect 53000 40601 53159 40653
rect 53211 40601 53371 40653
rect 53423 40601 53582 40653
rect 53634 40601 53792 40653
rect 53844 40601 54003 40653
rect 54055 40601 54214 40653
rect 54266 40650 54540 40653
rect 54266 40604 54440 40650
rect 54486 40604 54540 40650
rect 54266 40601 54540 40604
rect 52278 40560 54540 40601
rect 54758 40653 55840 40694
rect 54758 40650 54855 40653
rect 54758 40604 54793 40650
rect 54839 40604 54855 40650
rect 54758 40601 54855 40604
rect 54907 40650 55066 40653
rect 54907 40604 54956 40650
rect 55002 40604 55066 40650
rect 54907 40601 55066 40604
rect 55118 40650 55278 40653
rect 55330 40650 55489 40653
rect 55164 40604 55278 40650
rect 55330 40604 55439 40650
rect 55485 40604 55489 40650
rect 55118 40601 55278 40604
rect 55330 40601 55489 40604
rect 55541 40650 55840 40653
rect 55541 40604 55599 40650
rect 55645 40604 55760 40650
rect 55806 40604 55840 40650
rect 55541 40601 55840 40604
rect 54758 40561 55840 40601
rect 55927 40653 56632 40767
rect 57278 40653 57380 42401
rect 55927 40601 56015 40653
rect 56067 40601 56226 40653
rect 56278 40650 56437 40653
rect 56313 40604 56437 40650
rect 56278 40601 56437 40604
rect 56489 40601 56632 40653
rect 57278 40601 57281 40653
rect 57333 40601 57380 40653
rect 54817 40560 55579 40561
rect 48905 40515 49877 40555
rect 50099 40553 50255 40560
rect 48905 40509 48943 40515
rect 48995 40509 49154 40515
rect 49206 40509 49365 40515
rect 49417 40509 49576 40515
rect 49628 40509 49787 40515
rect 49839 40509 49877 40515
rect 30683 40441 31040 40481
rect 33484 40465 34643 40494
rect 30583 40364 31040 40441
rect 33019 40425 33327 40465
rect 33019 40422 33057 40425
rect 33109 40422 33237 40425
rect 33289 40422 33327 40425
rect 33484 40457 35082 40465
rect 35260 40463 35273 40509
rect 35523 40463 35543 40509
rect 35626 40463 35683 40509
rect 35729 40463 35754 40509
rect 35832 40463 35889 40509
rect 35935 40463 35965 40509
rect 36038 40463 36095 40509
rect 36141 40463 36176 40509
rect 36244 40463 36301 40509
rect 36347 40463 36360 40509
rect 36438 40463 36854 40509
rect 36900 40463 36971 40509
rect 37017 40463 37088 40509
rect 37134 40463 37206 40509
rect 37252 40463 37324 40509
rect 37370 40463 37442 40509
rect 37488 40465 37891 40509
rect 37488 40463 37909 40465
rect 37955 40463 38026 40509
rect 38123 40465 38143 40509
rect 38072 40463 38143 40465
rect 38189 40463 38261 40509
rect 38307 40463 38379 40509
rect 38425 40463 38497 40509
rect 38543 40463 38556 40509
rect 38658 40463 39021 40509
rect 39067 40463 39144 40509
rect 39190 40463 39267 40509
rect 39313 40463 39641 40509
rect 39687 40463 39730 40509
rect 31336 40376 31349 40422
rect 33323 40376 33336 40422
rect 33484 40411 33816 40457
rect 33862 40411 34002 40457
rect 34048 40411 34189 40457
rect 34235 40411 34376 40457
rect 34422 40411 34562 40457
rect 34608 40411 35082 40457
rect 35294 40423 36266 40463
rect 36438 40429 36953 40463
rect 37439 40429 38161 40463
rect 30583 40323 30855 40364
rect 30583 40277 30637 40323
rect 30683 40318 30855 40323
rect 30901 40318 31040 40364
rect 33019 40373 33057 40376
rect 33109 40373 33237 40376
rect 33289 40373 33327 40376
rect 33019 40332 33327 40373
rect 33484 40374 35082 40411
rect 30683 40277 31040 40318
rect 30583 40249 31040 40277
rect 33484 40292 33552 40374
rect 30583 40201 31493 40249
rect 30583 40160 30855 40201
rect 30583 40114 30637 40160
rect 30683 40155 30855 40160
rect 30901 40198 31493 40201
rect 30901 40155 31349 40198
rect 30683 40152 31349 40155
rect 33323 40152 33336 40198
rect 30683 40130 31493 40152
rect 30683 40114 31040 40130
rect 30583 40038 31040 40114
rect 30583 39997 30855 40038
rect 30583 39951 30637 39997
rect 30683 39992 30855 39997
rect 30901 39992 31040 40038
rect 30683 39951 31040 39992
rect 33019 39977 33327 40017
rect 33019 39974 33057 39977
rect 33109 39974 33237 39977
rect 33289 39974 33327 39977
rect 30583 39874 31040 39951
rect 31336 39928 31349 39974
rect 33323 39928 33336 39974
rect 33019 39925 33057 39928
rect 33109 39925 33237 39928
rect 33289 39925 33327 39928
rect 33019 39884 33327 39925
rect 30583 39834 30855 39874
rect 28492 39666 29196 39788
rect 28492 39620 28810 39666
rect 28856 39620 29196 39666
rect 29283 39753 30365 39794
rect 29283 39750 29582 39753
rect 29283 39704 29317 39750
rect 29363 39704 29478 39750
rect 29524 39704 29582 39750
rect 29283 39701 29582 39704
rect 29634 39750 29793 39753
rect 29845 39750 30005 39753
rect 29634 39704 29638 39750
rect 29684 39704 29793 39750
rect 29845 39704 29959 39750
rect 29634 39701 29793 39704
rect 29845 39701 30005 39704
rect 30057 39750 30216 39753
rect 30057 39704 30121 39750
rect 30167 39704 30216 39750
rect 30057 39701 30216 39704
rect 30268 39750 30365 39753
rect 30268 39704 30284 39750
rect 30330 39704 30365 39750
rect 30268 39701 30365 39704
rect 29283 39661 30365 39701
rect 30583 39788 30637 39834
rect 30683 39828 30855 39834
rect 30901 39828 31040 39874
rect 33484 39870 33495 40292
rect 33541 39870 33552 40292
rect 34964 40317 35082 40374
rect 36438 40329 36554 40429
rect 37853 40424 38161 40429
rect 38658 40449 39723 40463
rect 34964 40285 36360 40317
rect 34228 40215 34718 40256
rect 34228 40198 34267 40215
rect 34319 40198 34447 40215
rect 34499 40198 34627 40215
rect 33671 40152 33684 40198
rect 33730 40152 33787 40198
rect 33833 40152 33890 40198
rect 33936 40152 33993 40198
rect 34039 40152 34096 40198
rect 34142 40152 34199 40198
rect 34245 40163 34267 40198
rect 34245 40152 34302 40163
rect 34348 40152 34405 40198
rect 34499 40163 34508 40198
rect 34451 40152 34508 40163
rect 34554 40152 34612 40198
rect 34679 40163 34718 40215
rect 34964 40239 35273 40285
rect 35523 40239 35580 40285
rect 35626 40239 35683 40285
rect 35729 40239 35786 40285
rect 35832 40239 35889 40285
rect 35935 40239 35992 40285
rect 36038 40239 36095 40285
rect 36141 40239 36198 40285
rect 36244 40239 36301 40285
rect 36347 40239 36360 40285
rect 34964 40195 36360 40239
rect 34658 40152 34718 40163
rect 34228 40123 34718 40152
rect 36438 40189 36475 40329
rect 36521 40189 36554 40329
rect 35294 40061 36266 40095
rect 36438 40086 36554 40189
rect 36640 40329 36773 40349
rect 36640 40290 36697 40329
rect 36640 40238 36678 40290
rect 36640 40189 36697 40238
rect 36743 40189 36773 40329
rect 38658 40327 38726 40449
rect 39809 40443 44918 40481
rect 48765 40463 48778 40509
rect 48824 40463 48881 40509
rect 48927 40463 48943 40509
rect 49030 40463 49087 40509
rect 49133 40463 49154 40509
rect 49236 40463 49293 40509
rect 49339 40463 49365 40509
rect 49442 40463 49499 40509
rect 49545 40463 49576 40509
rect 49852 40463 49877 40509
rect 54085 40527 54540 40560
rect 50481 40467 51657 40494
rect 39809 40397 43739 40443
rect 43785 40397 43906 40443
rect 43952 40397 44071 40443
rect 44117 40397 44236 40443
rect 44282 40422 44918 40443
rect 48905 40423 49877 40463
rect 50044 40457 51657 40467
rect 44282 40397 44812 40422
rect 39809 40394 44812 40397
rect 39809 40348 39844 40394
rect 39890 40392 44812 40394
rect 39890 40348 39994 40392
rect 39809 40340 39994 40348
rect 40046 40376 44812 40392
rect 44858 40376 44925 40422
rect 44971 40376 45038 40422
rect 45084 40376 45151 40422
rect 45197 40376 45264 40422
rect 45310 40376 45323 40422
rect 48557 40377 48687 40417
rect 40046 40361 44918 40376
rect 40046 40340 40085 40361
rect 39809 40337 40085 40340
rect 36924 40317 37685 40324
rect 36923 40285 37931 40317
rect 36841 40239 36854 40285
rect 36900 40283 36971 40285
rect 36900 40239 36961 40283
rect 37017 40239 37088 40285
rect 37134 40283 37206 40285
rect 37134 40239 37172 40283
rect 37252 40239 37324 40285
rect 37370 40283 37442 40285
rect 37370 40239 37384 40283
rect 36923 40231 36961 40239
rect 37013 40231 37172 40239
rect 37224 40231 37384 40239
rect 37436 40239 37442 40283
rect 37488 40283 37909 40285
rect 37488 40239 37595 40283
rect 37436 40231 37595 40239
rect 37647 40239 37909 40283
rect 37955 40239 38026 40285
rect 38072 40239 38143 40285
rect 38189 40239 38261 40285
rect 38307 40239 38379 40285
rect 38425 40239 38497 40285
rect 38543 40239 38556 40285
rect 37647 40231 37931 40239
rect 36923 40198 37931 40231
rect 36923 40197 37685 40198
rect 36924 40191 37685 40197
rect 36640 40166 36773 40189
rect 38658 40187 38669 40327
rect 38715 40187 38726 40327
rect 39014 40285 39323 40317
rect 39492 40285 39608 40317
rect 39008 40239 39021 40285
rect 39067 40239 39144 40285
rect 39190 40239 39267 40285
rect 39313 40239 39326 40285
rect 39492 40239 39641 40285
rect 39687 40239 39730 40285
rect 38658 40176 38726 40187
rect 36438 40061 36953 40086
rect 37439 40083 37931 40086
rect 37439 40061 38161 40083
rect 35260 40015 35273 40061
rect 35523 40055 35580 40061
rect 35523 40015 35543 40055
rect 35626 40015 35683 40061
rect 35729 40055 35786 40061
rect 35729 40015 35754 40055
rect 35832 40015 35889 40061
rect 35935 40055 35992 40061
rect 35935 40015 35965 40055
rect 36038 40015 36095 40061
rect 36141 40055 36198 40061
rect 36141 40015 36176 40055
rect 36244 40015 36301 40061
rect 36347 40015 36360 40061
rect 36438 40015 36854 40061
rect 36900 40015 36971 40061
rect 37017 40015 37088 40061
rect 37134 40015 37206 40061
rect 37252 40015 37324 40061
rect 37370 40015 37442 40061
rect 37488 40043 37909 40061
rect 37488 40015 37891 40043
rect 37955 40015 38026 40061
rect 38072 40043 38143 40061
rect 38123 40015 38143 40043
rect 38189 40015 38261 40061
rect 38307 40015 38379 40061
rect 38425 40015 38497 40061
rect 38543 40015 38556 40061
rect 33781 39974 34089 40009
rect 35294 40003 35332 40015
rect 35384 40003 35543 40015
rect 35595 40003 35754 40015
rect 35806 40003 35965 40015
rect 36017 40003 36176 40015
rect 36228 40003 36266 40015
rect 33671 39928 33684 39974
rect 33730 39928 33787 39974
rect 33833 39969 33890 39974
rect 33871 39928 33890 39969
rect 33936 39928 33993 39974
rect 34039 39969 34096 39974
rect 34051 39928 34096 39969
rect 34142 39928 34199 39974
rect 34245 39928 34302 39974
rect 34348 39928 34405 39974
rect 34451 39928 34508 39974
rect 34554 39928 34612 39974
rect 34658 39928 34671 39974
rect 35294 39963 36266 40003
rect 36438 39966 36953 40015
rect 37439 39991 37891 40015
rect 37943 39991 38071 40015
rect 38123 39991 38161 40015
rect 37439 39966 38161 39991
rect 37853 39950 38161 39966
rect 33781 39917 33819 39928
rect 33871 39917 33999 39928
rect 34051 39917 34089 39928
rect 33781 39876 34089 39917
rect 33484 39859 33552 39870
rect 30683 39794 31040 39828
rect 30683 39788 32842 39794
rect 30583 39753 32842 39788
rect 34247 39787 35008 39794
rect 30583 39701 30854 39753
rect 30906 39701 31065 39753
rect 31117 39701 31276 39753
rect 31328 39750 31486 39753
rect 31538 39750 31697 39753
rect 31749 39750 31909 39753
rect 31961 39750 32120 39753
rect 32172 39750 32330 39753
rect 32382 39750 32541 39753
rect 32593 39750 32752 39753
rect 32804 39750 32842 39753
rect 34246 39753 35008 39787
rect 34246 39750 34284 39753
rect 34336 39750 34495 39753
rect 34547 39750 34707 39753
rect 31328 39704 31349 39750
rect 33323 39704 33336 39750
rect 33671 39704 33684 39750
rect 33730 39704 33787 39750
rect 33833 39704 33890 39750
rect 33936 39704 33993 39750
rect 34039 39704 34096 39750
rect 34142 39704 34199 39750
rect 34245 39704 34284 39750
rect 34348 39704 34405 39750
rect 34451 39704 34495 39750
rect 34554 39704 34612 39750
rect 34658 39704 34707 39750
rect 31328 39701 31486 39704
rect 31538 39701 31697 39704
rect 31749 39701 31909 39704
rect 31961 39701 32120 39704
rect 32172 39701 32330 39704
rect 32382 39701 32541 39704
rect 32593 39701 32752 39704
rect 32804 39701 32842 39704
rect 30583 39666 32842 39701
rect 34246 39701 34284 39704
rect 34336 39701 34495 39704
rect 34547 39701 34707 39704
rect 34759 39701 34918 39753
rect 34970 39701 35008 39753
rect 34246 39667 35008 39701
rect 29544 39660 30306 39661
rect 28492 39544 29196 39620
rect 28492 39503 29116 39544
rect 28492 39457 28810 39503
rect 28856 39498 29116 39503
rect 29162 39498 29196 39544
rect 28856 39457 29196 39498
rect 28492 39381 29196 39457
rect 28492 39340 29116 39381
rect 28492 39294 28810 39340
rect 28856 39335 29116 39340
rect 29162 39335 29196 39381
rect 28856 39294 29196 39335
rect 28492 39217 29196 39294
rect 28492 39177 29116 39217
rect 28492 39131 28810 39177
rect 28856 39171 29116 39177
rect 29162 39171 29196 39217
rect 28856 39131 29196 39171
rect 28492 39054 29196 39131
rect 28492 39013 29116 39054
rect 28492 38967 28810 39013
rect 28856 39008 29116 39013
rect 29162 39008 29196 39054
rect 28856 38967 29196 39008
rect 28492 38853 29196 38967
rect 30583 39620 30637 39666
rect 30683 39660 32842 39666
rect 34247 39660 35008 39667
rect 35182 39787 36364 39794
rect 35182 39753 36958 39787
rect 35182 39701 35220 39753
rect 35272 39701 35430 39753
rect 35482 39701 35641 39753
rect 35693 39701 35853 39753
rect 35905 39701 36064 39753
rect 36116 39701 36274 39753
rect 36326 39750 36958 39753
rect 36326 39704 36489 39750
rect 36723 39704 36958 39750
rect 36326 39701 36958 39704
rect 35182 39667 36958 39701
rect 37946 39753 38842 39794
rect 37946 39750 38330 39753
rect 38382 39750 38541 39753
rect 37946 39704 37957 39750
rect 38473 39704 38541 39750
rect 37946 39701 38330 39704
rect 38382 39701 38541 39704
rect 38593 39701 38752 39753
rect 38804 39701 38842 39753
rect 35182 39660 36364 39667
rect 37946 39660 38842 39701
rect 39014 39753 39323 40239
rect 39014 39701 39052 39753
rect 39104 39750 39232 39753
rect 39108 39704 39220 39750
rect 39104 39701 39232 39704
rect 39284 39701 39323 39753
rect 30683 39626 31040 39660
rect 30683 39620 30855 39626
rect 30583 39580 30855 39620
rect 30901 39580 31040 39626
rect 30583 39503 31040 39580
rect 33484 39584 33552 39595
rect 33019 39529 33327 39570
rect 33019 39526 33057 39529
rect 33109 39526 33237 39529
rect 33289 39526 33327 39529
rect 30583 39457 30637 39503
rect 30683 39462 31040 39503
rect 31336 39480 31349 39526
rect 33323 39480 33336 39526
rect 30683 39457 30855 39462
rect 30583 39416 30855 39457
rect 30901 39416 31040 39462
rect 33019 39477 33057 39480
rect 33109 39477 33237 39480
rect 33289 39477 33327 39480
rect 33019 39437 33327 39477
rect 30583 39340 31040 39416
rect 30583 39294 30637 39340
rect 30683 39324 31040 39340
rect 30683 39302 31493 39324
rect 30683 39299 31349 39302
rect 30683 39294 30855 39299
rect 30583 39253 30855 39294
rect 30901 39256 31349 39299
rect 33323 39256 33336 39302
rect 30901 39253 31493 39256
rect 30583 39205 31493 39253
rect 30583 39177 31040 39205
rect 30583 39131 30637 39177
rect 30683 39136 31040 39177
rect 30683 39131 30855 39136
rect 30583 39090 30855 39131
rect 30901 39090 31040 39136
rect 33484 39162 33495 39584
rect 33541 39162 33552 39584
rect 33781 39537 34089 39578
rect 33781 39526 33819 39537
rect 33871 39526 33999 39537
rect 34051 39526 34089 39537
rect 33671 39480 33684 39526
rect 33730 39480 33787 39526
rect 33871 39485 33890 39526
rect 33833 39480 33890 39485
rect 33936 39480 33993 39526
rect 34051 39485 34096 39526
rect 34039 39480 34096 39485
rect 34142 39480 34199 39526
rect 34245 39480 34302 39526
rect 34348 39480 34405 39526
rect 34451 39480 34508 39526
rect 34554 39480 34612 39526
rect 34658 39480 34671 39526
rect 33781 39445 34089 39480
rect 35294 39451 36266 39491
rect 37853 39488 38161 39504
rect 35294 39439 35332 39451
rect 35384 39439 35543 39451
rect 35595 39439 35754 39451
rect 35806 39439 35965 39451
rect 36017 39439 36176 39451
rect 36228 39439 36266 39451
rect 36438 39439 36953 39488
rect 37439 39463 38161 39488
rect 37439 39439 37891 39463
rect 37943 39439 38071 39463
rect 38123 39439 38161 39463
rect 35260 39393 35273 39439
rect 35523 39399 35543 39439
rect 35523 39393 35580 39399
rect 35626 39393 35683 39439
rect 35729 39399 35754 39439
rect 35729 39393 35786 39399
rect 35832 39393 35889 39439
rect 35935 39399 35965 39439
rect 35935 39393 35992 39399
rect 36038 39393 36095 39439
rect 36141 39399 36176 39439
rect 36141 39393 36198 39399
rect 36244 39393 36301 39439
rect 36347 39393 36360 39439
rect 36438 39393 36854 39439
rect 36900 39393 36971 39439
rect 37017 39393 37088 39439
rect 37134 39393 37206 39439
rect 37252 39393 37324 39439
rect 37370 39393 37442 39439
rect 37488 39411 37891 39439
rect 37488 39393 37909 39411
rect 37955 39393 38026 39439
rect 38123 39411 38143 39439
rect 38072 39393 38143 39411
rect 38189 39393 38261 39439
rect 38307 39393 38379 39439
rect 38425 39393 38497 39439
rect 38543 39393 38556 39439
rect 35294 39359 36266 39393
rect 36438 39368 36953 39393
rect 37439 39371 38161 39393
rect 37439 39368 37931 39371
rect 34228 39302 34718 39331
rect 33671 39256 33684 39302
rect 33730 39256 33787 39302
rect 33833 39256 33890 39302
rect 33936 39256 33993 39302
rect 34039 39256 34096 39302
rect 34142 39256 34199 39302
rect 34245 39291 34302 39302
rect 34245 39256 34267 39291
rect 34348 39256 34405 39302
rect 34451 39291 34508 39302
rect 34499 39256 34508 39291
rect 34554 39256 34612 39302
rect 34658 39291 34718 39302
rect 34228 39239 34267 39256
rect 34319 39239 34447 39256
rect 34499 39239 34627 39256
rect 34679 39239 34718 39291
rect 36438 39265 36554 39368
rect 34228 39198 34718 39239
rect 34964 39215 36360 39259
rect 30583 39013 31040 39090
rect 33019 39081 33327 39122
rect 33019 39078 33057 39081
rect 33109 39078 33237 39081
rect 33289 39078 33327 39081
rect 33484 39080 33552 39162
rect 34964 39169 35273 39215
rect 35523 39169 35580 39215
rect 35626 39169 35683 39215
rect 35729 39169 35786 39215
rect 35832 39169 35889 39215
rect 35935 39169 35992 39215
rect 36038 39169 36095 39215
rect 36141 39169 36198 39215
rect 36244 39169 36301 39215
rect 36347 39169 36360 39215
rect 34964 39137 36360 39169
rect 34964 39080 35082 39137
rect 31336 39032 31349 39078
rect 33323 39032 33336 39078
rect 33484 39043 35082 39080
rect 30583 38967 30637 39013
rect 30683 38973 31040 39013
rect 33019 39029 33057 39032
rect 33109 39029 33237 39032
rect 33289 39029 33327 39032
rect 33019 38989 33327 39029
rect 33484 38997 33816 39043
rect 33862 38997 34002 39043
rect 34048 38997 34189 39043
rect 34235 38997 34376 39043
rect 34422 38997 34562 39043
rect 34608 38997 35082 39043
rect 36438 39125 36475 39265
rect 36521 39125 36554 39265
rect 33484 38989 35082 38997
rect 35294 38991 36266 39031
rect 36438 39025 36554 39125
rect 36640 39265 36773 39288
rect 36640 39216 36697 39265
rect 36640 39164 36678 39216
rect 36640 39125 36697 39164
rect 36743 39125 36773 39265
rect 38658 39267 38726 39278
rect 36924 39257 37685 39263
rect 36923 39256 37685 39257
rect 36923 39223 37931 39256
rect 36923 39215 36961 39223
rect 37013 39215 37172 39223
rect 37224 39215 37384 39223
rect 36841 39169 36854 39215
rect 36900 39171 36961 39215
rect 36900 39169 36971 39171
rect 37017 39169 37088 39215
rect 37134 39171 37172 39215
rect 37134 39169 37206 39171
rect 37252 39169 37324 39215
rect 37370 39171 37384 39215
rect 37436 39215 37595 39223
rect 37436 39171 37442 39215
rect 37370 39169 37442 39171
rect 37488 39171 37595 39215
rect 37647 39215 37931 39223
rect 37647 39171 37909 39215
rect 37488 39169 37909 39171
rect 37955 39169 38026 39215
rect 38072 39169 38143 39215
rect 38189 39169 38261 39215
rect 38307 39169 38379 39215
rect 38425 39169 38497 39215
rect 38543 39169 38556 39215
rect 36923 39137 37931 39169
rect 36924 39130 37685 39137
rect 36640 39105 36773 39125
rect 38658 39127 38669 39267
rect 38715 39127 38726 39267
rect 39014 39215 39323 39701
rect 39492 39787 39608 40239
rect 39923 40206 40085 40337
rect 39923 40154 39994 40206
rect 40046 40154 40085 40206
rect 39923 40114 40085 40154
rect 39737 40018 39865 40031
rect 39737 39991 39866 40018
rect 39737 39974 39775 39991
rect 39827 39974 39866 39991
rect 39727 39928 39740 39974
rect 39827 39939 39862 39974
rect 39786 39928 39862 39939
rect 39908 39928 39985 39974
rect 40031 39928 40108 39974
rect 40154 39928 40167 39974
rect 40246 39963 40362 40361
rect 42229 40222 44509 40263
rect 42229 40170 43445 40222
rect 43497 40170 44509 40222
rect 42229 40130 44509 40170
rect 44341 40086 44509 40130
rect 44341 40040 44358 40086
rect 44498 40040 44509 40086
rect 39737 39899 39866 39928
rect 40246 39917 40281 39963
rect 40327 39917 40362 39963
rect 40246 39880 40362 39917
rect 40718 39991 43524 40032
rect 44341 40029 44509 40040
rect 40718 39939 41935 39991
rect 41987 39939 43524 39991
rect 40718 39898 43524 39939
rect 44605 39974 44721 40361
rect 45400 40331 48379 40372
rect 45400 40317 46731 40331
rect 45400 40271 45464 40317
rect 45604 40279 46731 40317
rect 46783 40279 48379 40331
rect 45604 40271 48379 40279
rect 44901 40215 45241 40256
rect 45400 40238 48379 40271
rect 48557 40325 48596 40377
rect 48648 40325 48687 40377
rect 48557 40302 48687 40325
rect 50044 40411 50516 40457
rect 50562 40411 50703 40457
rect 50749 40411 50890 40457
rect 50936 40411 51076 40457
rect 51122 40411 51263 40457
rect 51309 40411 51657 40457
rect 51797 40447 52105 40487
rect 51797 40422 51835 40447
rect 51887 40422 52015 40447
rect 52067 40422 52105 40447
rect 54085 40481 54223 40527
rect 54269 40487 54540 40527
rect 54269 40481 54440 40487
rect 54085 40441 54440 40481
rect 54486 40441 54540 40487
rect 50044 40374 51657 40411
rect 51789 40376 51802 40422
rect 53776 40376 53789 40422
rect 50044 40317 50160 40374
rect 44901 40198 44939 40215
rect 44991 40198 45151 40215
rect 45203 40198 45241 40215
rect 44799 40152 44812 40198
rect 44858 40152 44925 40198
rect 44991 40163 45038 40198
rect 44971 40152 45038 40163
rect 45084 40152 45151 40198
rect 45203 40163 45264 40198
rect 45197 40152 45264 40163
rect 45310 40152 45323 40198
rect 48557 40162 48622 40302
rect 48668 40162 48687 40302
rect 49820 40285 50160 40317
rect 48765 40239 48778 40285
rect 48824 40239 48881 40285
rect 48927 40239 48984 40285
rect 49030 40239 49087 40285
rect 49133 40239 49190 40285
rect 49236 40239 49293 40285
rect 49339 40239 49396 40285
rect 49442 40239 49499 40285
rect 49545 40239 49602 40285
rect 49852 40239 50160 40285
rect 51589 40322 51657 40374
rect 51797 40354 52105 40376
rect 49820 40198 50160 40239
rect 50262 40215 50812 40256
rect 48557 40159 48687 40162
rect 44901 40123 45241 40152
rect 48557 40107 48596 40159
rect 48648 40107 48687 40159
rect 50262 40163 50300 40215
rect 50352 40198 50511 40215
rect 50563 40198 50722 40215
rect 50352 40163 50467 40198
rect 50563 40163 50571 40198
rect 50262 40152 50467 40163
rect 50513 40152 50571 40163
rect 50617 40152 50674 40198
rect 50720 40163 50722 40198
rect 50774 40198 50812 40215
rect 50774 40163 50777 40198
rect 50720 40152 50777 40163
rect 50823 40152 50880 40198
rect 50926 40152 50983 40198
rect 51029 40152 51086 40198
rect 51132 40152 51189 40198
rect 51235 40152 51292 40198
rect 51338 40152 51395 40198
rect 51441 40152 51454 40198
rect 50262 40123 50812 40152
rect 48557 40066 48687 40107
rect 48905 40061 49877 40092
rect 48765 40015 48778 40061
rect 48824 40015 48881 40061
rect 48927 40052 48984 40061
rect 48927 40015 48943 40052
rect 49030 40015 49087 40061
rect 49133 40052 49190 40061
rect 49133 40015 49154 40052
rect 49236 40015 49293 40061
rect 49339 40052 49396 40061
rect 49339 40015 49365 40052
rect 49442 40015 49499 40061
rect 49545 40052 49602 40061
rect 49545 40015 49576 40052
rect 49852 40015 49877 40061
rect 48905 40000 48943 40015
rect 48995 40000 49154 40015
rect 49206 40000 49365 40015
rect 49417 40000 49576 40015
rect 49628 40000 49787 40015
rect 49839 40000 49877 40015
rect 44605 39928 44812 39974
rect 44858 39928 44925 39974
rect 44971 39928 45038 39974
rect 45084 39928 45151 39974
rect 45197 39928 45264 39974
rect 45310 39928 45323 39974
rect 48905 39960 49877 40000
rect 51035 39977 51343 40017
rect 51035 39974 51073 39977
rect 51125 39974 51253 39977
rect 51305 39974 51343 39977
rect 43362 39891 43524 39898
rect 43362 39845 43373 39891
rect 43513 39845 43524 39891
rect 43362 39834 43524 39845
rect 45584 39914 48546 39950
rect 50454 39928 50467 39974
rect 50513 39928 50571 39974
rect 50617 39928 50674 39974
rect 50720 39928 50777 39974
rect 50823 39928 50880 39974
rect 50926 39928 50983 39974
rect 51029 39928 51073 39974
rect 51132 39928 51189 39974
rect 51235 39928 51253 39974
rect 51338 39928 51395 39974
rect 51441 39928 51454 39974
rect 45584 39868 45619 39914
rect 45665 39868 45777 39914
rect 45823 39868 45935 39914
rect 45981 39868 46093 39914
rect 46139 39868 46251 39914
rect 46297 39868 46409 39914
rect 46455 39868 46568 39914
rect 46614 39868 46726 39914
rect 46772 39868 46884 39914
rect 46930 39868 47042 39914
rect 47088 39868 47200 39914
rect 47246 39868 47358 39914
rect 47404 39868 47516 39914
rect 47562 39868 47675 39914
rect 47721 39868 47833 39914
rect 47879 39868 47991 39914
rect 48037 39868 48149 39914
rect 48195 39868 48307 39914
rect 48353 39868 48465 39914
rect 48511 39868 48546 39914
rect 51035 39925 51073 39928
rect 51125 39925 51253 39928
rect 51305 39925 51343 39928
rect 51035 39884 51343 39925
rect 51589 39900 51600 40322
rect 51646 39900 51657 40322
rect 54085 40323 54540 40441
rect 54085 40277 54440 40323
rect 54486 40277 54540 40323
rect 54085 40249 54540 40277
rect 53585 40198 54540 40249
rect 51789 40152 51802 40198
rect 53776 40160 54540 40198
rect 53776 40152 54440 40160
rect 53585 40130 54440 40152
rect 54085 40114 54440 40130
rect 54486 40114 54540 40160
rect 54085 40038 54540 40114
rect 51797 39984 52105 40024
rect 51797 39974 51835 39984
rect 51887 39974 52015 39984
rect 52067 39974 52105 39984
rect 54085 39992 54223 40038
rect 54269 39997 54540 40038
rect 54269 39992 54440 39997
rect 51789 39928 51802 39974
rect 53776 39928 53789 39974
rect 54085 39951 54440 39992
rect 54486 39951 54540 39997
rect 51589 39889 51657 39900
rect 51797 39891 52105 39928
rect 40215 39787 40523 39794
rect 40788 39787 42986 39801
rect 43753 39787 44514 39794
rect 39492 39764 42986 39787
rect 43704 39764 44514 39787
rect 39492 39753 44514 39764
rect 39492 39750 40253 39753
rect 39492 39704 39740 39750
rect 39786 39704 39862 39750
rect 39908 39704 39985 39750
rect 40031 39704 40108 39750
rect 40154 39704 40253 39750
rect 39492 39701 40253 39704
rect 40305 39701 40433 39753
rect 40485 39750 43790 39753
rect 40485 39704 40836 39750
rect 40882 39704 40994 39750
rect 41040 39704 41152 39750
rect 41198 39704 41310 39750
rect 41356 39704 41469 39750
rect 41515 39704 41627 39750
rect 41673 39704 41785 39750
rect 41831 39704 41943 39750
rect 41989 39704 42101 39750
rect 42147 39704 42259 39750
rect 42305 39704 42418 39750
rect 42464 39704 42576 39750
rect 42622 39704 42734 39750
rect 42780 39704 42892 39750
rect 42938 39704 43739 39750
rect 43785 39704 43790 39750
rect 40485 39701 43790 39704
rect 43842 39750 44001 39753
rect 43842 39704 43906 39750
rect 43952 39704 44001 39750
rect 43842 39701 44001 39704
rect 44053 39750 44213 39753
rect 44265 39750 44424 39753
rect 44053 39704 44071 39750
rect 44117 39704 44213 39750
rect 44282 39704 44424 39750
rect 44053 39701 44213 39704
rect 44265 39701 44424 39704
rect 44476 39701 44514 39753
rect 39492 39690 44514 39701
rect 39492 39667 42986 39690
rect 43704 39667 44514 39690
rect 39492 39215 39608 39667
rect 40215 39660 40523 39667
rect 40788 39653 42986 39667
rect 43753 39660 44514 39667
rect 44796 39787 45346 39794
rect 45584 39787 48546 39868
rect 54085 39874 54540 39951
rect 54085 39828 54223 39874
rect 54269 39834 54540 39874
rect 54269 39828 54440 39834
rect 54085 39794 54440 39828
rect 48800 39787 49982 39794
rect 50308 39787 50859 39794
rect 44796 39753 49982 39787
rect 44796 39750 44834 39753
rect 44886 39750 45045 39753
rect 45097 39750 45256 39753
rect 45308 39750 48838 39753
rect 44796 39704 44812 39750
rect 44886 39704 44925 39750
rect 44971 39704 45038 39750
rect 45097 39704 45151 39750
rect 45197 39704 45256 39750
rect 45310 39704 45619 39750
rect 45665 39704 45777 39750
rect 45823 39704 45935 39750
rect 45981 39704 46093 39750
rect 46139 39704 46251 39750
rect 46297 39704 46409 39750
rect 46455 39704 46568 39750
rect 46614 39704 46726 39750
rect 46772 39704 46884 39750
rect 46930 39704 47042 39750
rect 47088 39704 47200 39750
rect 47246 39704 47358 39750
rect 47404 39704 47516 39750
rect 47562 39704 47675 39750
rect 47721 39704 47833 39750
rect 47879 39704 47991 39750
rect 48037 39704 48149 39750
rect 48195 39704 48307 39750
rect 48353 39704 48465 39750
rect 48511 39704 48838 39750
rect 44796 39701 44834 39704
rect 44886 39701 45045 39704
rect 45097 39701 45256 39704
rect 45308 39701 48838 39704
rect 48890 39701 49048 39753
rect 49100 39701 49259 39753
rect 49311 39701 49471 39753
rect 49523 39701 49682 39753
rect 49734 39701 49892 39753
rect 49944 39701 49982 39753
rect 44796 39667 49982 39701
rect 50307 39753 50859 39787
rect 50307 39701 50346 39753
rect 50398 39750 50557 39753
rect 50609 39750 50768 39753
rect 50820 39750 50859 39753
rect 52278 39788 54440 39794
rect 54486 39788 54540 39834
rect 55927 40487 56632 40601
rect 55927 40444 56267 40487
rect 55927 40398 55961 40444
rect 56007 40441 56267 40444
rect 56313 40441 56632 40487
rect 56007 40398 56632 40441
rect 55927 40323 56632 40398
rect 55927 40281 56267 40323
rect 55927 40235 55961 40281
rect 56007 40277 56267 40281
rect 56313 40277 56632 40323
rect 56007 40235 56632 40277
rect 55927 40160 56632 40235
rect 55927 40117 56267 40160
rect 55927 40071 55961 40117
rect 56007 40114 56267 40117
rect 56313 40114 56632 40160
rect 56007 40071 56632 40114
rect 55927 39997 56632 40071
rect 55927 39954 56267 39997
rect 55927 39908 55961 39954
rect 56007 39951 56267 39954
rect 56313 39951 56632 39997
rect 56007 39908 56632 39951
rect 55927 39834 56632 39908
rect 52278 39753 54540 39788
rect 52278 39750 52316 39753
rect 52368 39750 52527 39753
rect 52579 39750 52738 39753
rect 52790 39750 52948 39753
rect 53000 39750 53159 39753
rect 53211 39750 53371 39753
rect 53423 39750 53582 39753
rect 53634 39750 53792 39753
rect 50398 39704 50467 39750
rect 50513 39704 50557 39750
rect 50617 39704 50674 39750
rect 50720 39704 50768 39750
rect 50823 39704 50880 39750
rect 50926 39704 50983 39750
rect 51029 39704 51086 39750
rect 51132 39704 51189 39750
rect 51235 39704 51292 39750
rect 51338 39704 51395 39750
rect 51441 39704 51454 39750
rect 51789 39704 51802 39750
rect 53776 39704 53792 39750
rect 50398 39701 50557 39704
rect 50609 39701 50768 39704
rect 50820 39701 50859 39704
rect 50307 39667 50859 39701
rect 44796 39660 45346 39667
rect 43362 39609 43524 39620
rect 39737 39526 39866 39555
rect 40246 39537 40362 39574
rect 43362 39563 43373 39609
rect 43513 39563 43524 39609
rect 43362 39556 43524 39563
rect 39727 39480 39740 39526
rect 39786 39515 39862 39526
rect 39827 39480 39862 39515
rect 39908 39480 39985 39526
rect 40031 39480 40108 39526
rect 40154 39480 40167 39526
rect 40246 39491 40281 39537
rect 40327 39491 40362 39537
rect 39737 39463 39775 39480
rect 39827 39463 39866 39480
rect 39737 39436 39866 39463
rect 39737 39423 39865 39436
rect 39923 39300 40085 39340
rect 39923 39248 39994 39300
rect 40046 39248 40085 39300
rect 39008 39169 39021 39215
rect 39067 39169 39144 39215
rect 39190 39169 39267 39215
rect 39313 39169 39326 39215
rect 39492 39169 39641 39215
rect 39687 39169 39730 39215
rect 39014 39137 39323 39169
rect 39492 39137 39608 39169
rect 37853 39025 38161 39030
rect 36438 38991 36953 39025
rect 37439 38991 38161 39025
rect 38658 39005 38726 39127
rect 39923 39117 40085 39248
rect 39809 39114 40085 39117
rect 39809 39106 39994 39114
rect 39809 39060 39844 39106
rect 39890 39062 39994 39106
rect 40046 39093 40085 39114
rect 40246 39093 40362 39491
rect 40718 39515 43524 39556
rect 45584 39586 48546 39667
rect 48800 39660 49982 39667
rect 50308 39660 50859 39667
rect 52278 39701 52316 39704
rect 52368 39701 52527 39704
rect 52579 39701 52738 39704
rect 52790 39701 52948 39704
rect 53000 39701 53159 39704
rect 53211 39701 53371 39704
rect 53423 39701 53582 39704
rect 53634 39701 53792 39704
rect 53844 39701 54003 39753
rect 54055 39701 54214 39753
rect 54266 39701 54540 39753
rect 52278 39666 54540 39701
rect 52278 39660 54440 39666
rect 45584 39540 45619 39586
rect 45665 39540 45777 39586
rect 45823 39540 45935 39586
rect 45981 39540 46093 39586
rect 46139 39540 46251 39586
rect 46297 39540 46409 39586
rect 46455 39540 46568 39586
rect 46614 39540 46726 39586
rect 46772 39540 46884 39586
rect 46930 39540 47042 39586
rect 47088 39540 47200 39586
rect 47246 39540 47358 39586
rect 47404 39540 47516 39586
rect 47562 39540 47675 39586
rect 47721 39540 47833 39586
rect 47879 39540 47991 39586
rect 48037 39540 48149 39586
rect 48195 39540 48307 39586
rect 48353 39540 48465 39586
rect 48511 39540 48546 39586
rect 54085 39626 54440 39660
rect 54085 39580 54223 39626
rect 54269 39620 54440 39626
rect 54486 39620 54540 39666
rect 54758 39753 55840 39794
rect 54758 39750 54855 39753
rect 54758 39704 54793 39750
rect 54839 39704 54855 39750
rect 54758 39701 54855 39704
rect 54907 39750 55066 39753
rect 54907 39704 54956 39750
rect 55002 39704 55066 39750
rect 54907 39701 55066 39704
rect 55118 39750 55278 39753
rect 55330 39750 55489 39753
rect 55164 39704 55278 39750
rect 55330 39704 55439 39750
rect 55485 39704 55489 39750
rect 55118 39701 55278 39704
rect 55330 39701 55489 39704
rect 55541 39750 55840 39753
rect 55541 39704 55599 39750
rect 55645 39704 55760 39750
rect 55806 39704 55840 39750
rect 55541 39701 55840 39704
rect 54758 39661 55840 39701
rect 55927 39788 56267 39834
rect 56313 39788 56632 39834
rect 55927 39666 56632 39788
rect 54817 39660 55579 39661
rect 54269 39580 54540 39620
rect 40718 39463 41935 39515
rect 41987 39463 43524 39515
rect 40718 39422 43524 39463
rect 44605 39480 44812 39526
rect 44858 39480 44925 39526
rect 44971 39480 45038 39526
rect 45084 39480 45151 39526
rect 45197 39480 45264 39526
rect 45310 39480 45323 39526
rect 45584 39504 48546 39540
rect 51035 39529 51343 39570
rect 51035 39526 51073 39529
rect 51125 39526 51253 39529
rect 51305 39526 51343 39529
rect 51589 39554 51657 39565
rect 44341 39414 44509 39425
rect 44341 39368 44358 39414
rect 44498 39368 44509 39414
rect 44341 39324 44509 39368
rect 42229 39284 44509 39324
rect 42229 39232 43445 39284
rect 43497 39232 44509 39284
rect 42229 39191 44509 39232
rect 44605 39093 44721 39480
rect 48905 39454 49877 39494
rect 50454 39480 50467 39526
rect 50513 39480 50571 39526
rect 50617 39480 50674 39526
rect 50720 39480 50777 39526
rect 50823 39480 50880 39526
rect 50926 39480 50983 39526
rect 51029 39480 51073 39526
rect 51132 39480 51189 39526
rect 51235 39480 51253 39526
rect 51338 39480 51395 39526
rect 51441 39480 51454 39526
rect 48905 39439 48943 39454
rect 48995 39439 49154 39454
rect 49206 39439 49365 39454
rect 49417 39439 49576 39454
rect 49628 39439 49787 39454
rect 49839 39439 49877 39454
rect 48765 39393 48778 39439
rect 48824 39393 48881 39439
rect 48927 39402 48943 39439
rect 48927 39393 48984 39402
rect 49030 39393 49087 39439
rect 49133 39402 49154 39439
rect 49133 39393 49190 39402
rect 49236 39393 49293 39439
rect 49339 39402 49365 39439
rect 49339 39393 49396 39402
rect 49442 39393 49499 39439
rect 49545 39402 49576 39439
rect 49545 39393 49602 39402
rect 49852 39393 49877 39439
rect 51035 39477 51073 39480
rect 51125 39477 51253 39480
rect 51305 39477 51343 39480
rect 51035 39437 51343 39477
rect 48557 39347 48687 39388
rect 48905 39362 49877 39393
rect 44901 39302 45241 39331
rect 44799 39256 44812 39302
rect 44858 39256 44925 39302
rect 44971 39291 45038 39302
rect 44991 39256 45038 39291
rect 45084 39256 45151 39302
rect 45197 39291 45264 39302
rect 45203 39256 45264 39291
rect 45310 39256 45323 39302
rect 48557 39295 48596 39347
rect 48648 39295 48687 39347
rect 48557 39292 48687 39295
rect 44901 39239 44939 39256
rect 44991 39239 45151 39256
rect 45203 39239 45241 39256
rect 44901 39198 45241 39239
rect 45400 39183 48379 39216
rect 45400 39137 45464 39183
rect 45604 39175 48379 39183
rect 45604 39137 47108 39175
rect 45400 39123 47108 39137
rect 47160 39123 48379 39175
rect 40046 39078 44918 39093
rect 45400 39082 48379 39123
rect 48557 39152 48622 39292
rect 48668 39152 48687 39292
rect 50262 39302 50812 39331
rect 50262 39291 50467 39302
rect 50513 39291 50571 39302
rect 49820 39215 50160 39256
rect 48765 39169 48778 39215
rect 48824 39169 48881 39215
rect 48927 39169 48984 39215
rect 49030 39169 49087 39215
rect 49133 39169 49190 39215
rect 49236 39169 49293 39215
rect 49339 39169 49396 39215
rect 49442 39169 49499 39215
rect 49545 39169 49602 39215
rect 49852 39169 50160 39215
rect 50262 39239 50300 39291
rect 50352 39256 50467 39291
rect 50563 39256 50571 39291
rect 50617 39256 50674 39302
rect 50720 39291 50777 39302
rect 50720 39256 50722 39291
rect 50352 39239 50511 39256
rect 50563 39239 50722 39256
rect 50774 39256 50777 39291
rect 50823 39256 50880 39302
rect 50926 39256 50983 39302
rect 51029 39256 51086 39302
rect 51132 39256 51189 39302
rect 51235 39256 51292 39302
rect 51338 39256 51395 39302
rect 51441 39256 51454 39302
rect 50774 39239 50812 39256
rect 50262 39198 50812 39239
rect 48557 39129 48687 39152
rect 49820 39137 50160 39169
rect 40046 39062 44812 39078
rect 39890 39060 44812 39062
rect 39809 39057 44812 39060
rect 39809 39011 43739 39057
rect 43785 39011 43906 39057
rect 43952 39011 44071 39057
rect 44117 39011 44236 39057
rect 44282 39032 44812 39057
rect 44858 39032 44925 39078
rect 44971 39032 45038 39078
rect 45084 39032 45151 39078
rect 45197 39032 45264 39078
rect 45310 39032 45323 39078
rect 48557 39077 48596 39129
rect 48648 39077 48687 39129
rect 48557 39037 48687 39077
rect 50044 39080 50160 39137
rect 51589 39132 51600 39554
rect 51646 39132 51657 39554
rect 51797 39526 52105 39563
rect 51789 39480 51802 39526
rect 53776 39480 53789 39526
rect 54085 39503 54540 39580
rect 51797 39470 51835 39480
rect 51887 39470 52015 39480
rect 52067 39470 52105 39480
rect 51797 39430 52105 39470
rect 54085 39462 54440 39503
rect 54085 39416 54223 39462
rect 54269 39457 54440 39462
rect 54486 39457 54540 39503
rect 54269 39416 54540 39457
rect 54085 39340 54540 39416
rect 54085 39324 54440 39340
rect 53585 39302 54440 39324
rect 51789 39256 51802 39302
rect 53776 39294 54440 39302
rect 54486 39294 54540 39340
rect 53776 39256 54540 39294
rect 53585 39205 54540 39256
rect 51589 39080 51657 39132
rect 54085 39177 54540 39205
rect 54085 39131 54440 39177
rect 54486 39131 54540 39177
rect 50044 39043 51657 39080
rect 51797 39078 52105 39100
rect 44282 39011 44918 39032
rect 38658 38991 39723 39005
rect 30683 38967 30855 38973
rect 30583 38927 30855 38967
rect 30901 38927 31040 38973
rect 33484 38960 34643 38989
rect 35260 38945 35273 38991
rect 35523 38945 35543 38991
rect 35626 38945 35683 38991
rect 35729 38945 35754 38991
rect 35832 38945 35889 38991
rect 35935 38945 35965 38991
rect 36038 38945 36095 38991
rect 36141 38945 36176 38991
rect 36244 38945 36301 38991
rect 36347 38945 36360 38991
rect 36438 38945 36854 38991
rect 36900 38945 36971 38991
rect 37017 38945 37088 38991
rect 37134 38945 37206 38991
rect 37252 38945 37324 38991
rect 37370 38945 37442 38991
rect 37488 38989 37909 38991
rect 37488 38945 37891 38989
rect 37955 38945 38026 38991
rect 38072 38989 38143 38991
rect 38123 38945 38143 38989
rect 38189 38945 38261 38991
rect 38307 38945 38379 38991
rect 38425 38945 38497 38991
rect 38543 38945 38556 38991
rect 38658 38945 39021 38991
rect 39067 38945 39144 38991
rect 39190 38945 39267 38991
rect 39313 38945 39641 38991
rect 39687 38945 39730 38991
rect 39809 38973 44918 39011
rect 48905 38991 49877 39031
rect 48765 38945 48778 38991
rect 48824 38945 48881 38991
rect 48927 38945 48943 38991
rect 49030 38945 49087 38991
rect 49133 38945 49154 38991
rect 49236 38945 49293 38991
rect 49339 38945 49365 38991
rect 49442 38945 49499 38991
rect 49545 38945 49576 38991
rect 49852 38945 49877 38991
rect 50044 38997 50516 39043
rect 50562 38997 50703 39043
rect 50749 38997 50890 39043
rect 50936 38997 51076 39043
rect 51122 38997 51263 39043
rect 51309 38997 51657 39043
rect 51789 39032 51802 39078
rect 53776 39032 53789 39078
rect 50044 38987 51657 38997
rect 50481 38960 51657 38987
rect 51797 39007 51835 39032
rect 51887 39007 52015 39032
rect 52067 39007 52105 39032
rect 51797 38967 52105 39007
rect 54085 39013 54540 39131
rect 54085 38973 54440 39013
rect 30583 38894 31040 38927
rect 35294 38939 35332 38945
rect 35384 38939 35543 38945
rect 35595 38939 35754 38945
rect 35806 38939 35965 38945
rect 36017 38939 36176 38945
rect 36228 38939 36266 38945
rect 34870 38894 35025 38901
rect 35294 38899 36266 38939
rect 36438 38905 36953 38945
rect 37439 38937 37891 38945
rect 37943 38937 38071 38945
rect 38123 38937 38161 38945
rect 37439 38905 38161 38937
rect 37853 38897 38161 38905
rect 27744 38801 27790 38853
rect 27842 38801 27846 38853
rect 28492 38801 28634 38853
rect 28686 38850 28845 38853
rect 28686 38804 28810 38850
rect 28686 38801 28845 38804
rect 28897 38801 29056 38853
rect 29108 38801 29196 38853
rect 27744 37053 27846 38801
rect 28492 38687 29196 38801
rect 29283 38853 30365 38894
rect 29283 38850 29582 38853
rect 29283 38804 29317 38850
rect 29363 38804 29478 38850
rect 29524 38804 29582 38850
rect 29283 38801 29582 38804
rect 29634 38850 29793 38853
rect 29845 38850 30005 38853
rect 29634 38804 29638 38850
rect 29684 38804 29793 38850
rect 29845 38804 29959 38850
rect 29634 38801 29793 38804
rect 29845 38801 30005 38804
rect 30057 38850 30216 38853
rect 30057 38804 30121 38850
rect 30167 38804 30216 38850
rect 30057 38801 30216 38804
rect 30268 38850 30365 38853
rect 30268 38804 30284 38850
rect 30330 38804 30365 38850
rect 30268 38801 30365 38804
rect 29283 38761 30365 38801
rect 30583 38853 32842 38894
rect 30583 38850 30854 38853
rect 30583 38804 30637 38850
rect 30683 38804 30854 38850
rect 30583 38801 30854 38804
rect 30906 38801 31065 38853
rect 31117 38801 31276 38853
rect 31328 38801 31486 38853
rect 31538 38801 31697 38853
rect 31749 38801 31909 38853
rect 31961 38801 32120 38853
rect 32172 38801 32330 38853
rect 32382 38801 32541 38853
rect 32593 38801 32752 38853
rect 32804 38801 32842 38853
rect 29544 38760 30306 38761
rect 30583 38760 32842 38801
rect 34717 38853 35025 38894
rect 38658 38885 39723 38945
rect 48905 38939 48943 38945
rect 48995 38939 49154 38945
rect 49206 38939 49365 38945
rect 49417 38939 49576 38945
rect 49628 38939 49787 38945
rect 49839 38939 49877 38945
rect 48905 38899 49877 38939
rect 54085 38927 54223 38973
rect 54269 38967 54440 38973
rect 54486 38967 54540 39013
rect 54269 38927 54540 38967
rect 50099 38894 50255 38901
rect 54085 38894 54540 38927
rect 55927 39620 56267 39666
rect 56313 39620 56632 39666
rect 55927 39544 56632 39620
rect 55927 39498 55961 39544
rect 56007 39503 56632 39544
rect 56007 39498 56267 39503
rect 55927 39457 56267 39498
rect 56313 39457 56632 39503
rect 55927 39381 56632 39457
rect 55927 39335 55961 39381
rect 56007 39340 56632 39381
rect 56007 39335 56267 39340
rect 55927 39294 56267 39335
rect 56313 39294 56632 39340
rect 55927 39217 56632 39294
rect 55927 39171 55961 39217
rect 56007 39177 56632 39217
rect 56007 39171 56267 39177
rect 55927 39131 56267 39171
rect 56313 39131 56632 39177
rect 55927 39054 56632 39131
rect 55927 39008 55961 39054
rect 56007 39013 56632 39054
rect 56007 39008 56267 39013
rect 55927 38967 56267 39008
rect 56313 38967 56632 39013
rect 34717 38801 34755 38853
rect 34807 38850 34935 38853
rect 34807 38804 34916 38850
rect 34807 38801 34935 38804
rect 34987 38801 35025 38853
rect 34717 38760 35025 38801
rect 50099 38853 50408 38894
rect 50099 38801 50138 38853
rect 50190 38850 50318 38853
rect 50206 38804 50318 38850
rect 50190 38801 50318 38804
rect 50370 38801 50408 38853
rect 28492 38641 28810 38687
rect 28856 38644 29196 38687
rect 28856 38641 29116 38644
rect 28492 38598 29116 38641
rect 29162 38598 29196 38644
rect 28492 38523 29196 38598
rect 28492 38477 28810 38523
rect 28856 38481 29196 38523
rect 28856 38477 29116 38481
rect 28492 38435 29116 38477
rect 29162 38435 29196 38481
rect 28492 38360 29196 38435
rect 28492 38314 28810 38360
rect 28856 38317 29196 38360
rect 28856 38314 29116 38317
rect 28492 38271 29116 38314
rect 29162 38271 29196 38317
rect 28492 38197 29196 38271
rect 28492 38151 28810 38197
rect 28856 38154 29196 38197
rect 28856 38151 29116 38154
rect 28492 38108 29116 38151
rect 29162 38108 29196 38154
rect 28492 38034 29196 38108
rect 28492 37988 28810 38034
rect 28856 37988 29196 38034
rect 30583 38727 31040 38760
rect 34870 38753 35025 38760
rect 30583 38687 30855 38727
rect 30583 38641 30637 38687
rect 30683 38681 30855 38687
rect 30901 38681 31040 38727
rect 35294 38715 36266 38755
rect 37853 38749 38161 38757
rect 35294 38709 35332 38715
rect 35384 38709 35543 38715
rect 35595 38709 35754 38715
rect 35806 38709 35965 38715
rect 36017 38709 36176 38715
rect 36228 38709 36266 38715
rect 36438 38709 36953 38749
rect 37439 38717 38161 38749
rect 37439 38709 37891 38717
rect 37943 38709 38071 38717
rect 38123 38709 38161 38717
rect 38658 38709 39723 38769
rect 50099 38760 50408 38801
rect 52278 38853 54540 38894
rect 52278 38801 52316 38853
rect 52368 38801 52527 38853
rect 52579 38801 52738 38853
rect 52790 38801 52948 38853
rect 53000 38801 53159 38853
rect 53211 38801 53371 38853
rect 53423 38801 53582 38853
rect 53634 38801 53792 38853
rect 53844 38801 54003 38853
rect 54055 38801 54214 38853
rect 54266 38850 54540 38853
rect 54266 38804 54440 38850
rect 54486 38804 54540 38850
rect 54266 38801 54540 38804
rect 52278 38760 54540 38801
rect 54758 38853 55840 38894
rect 54758 38850 54855 38853
rect 54758 38804 54793 38850
rect 54839 38804 54855 38850
rect 54758 38801 54855 38804
rect 54907 38850 55066 38853
rect 54907 38804 54956 38850
rect 55002 38804 55066 38850
rect 54907 38801 55066 38804
rect 55118 38850 55278 38853
rect 55330 38850 55489 38853
rect 55164 38804 55278 38850
rect 55330 38804 55439 38850
rect 55485 38804 55489 38850
rect 55118 38801 55278 38804
rect 55330 38801 55489 38804
rect 55541 38850 55840 38853
rect 55541 38804 55599 38850
rect 55645 38804 55760 38850
rect 55806 38804 55840 38850
rect 55541 38801 55840 38804
rect 54758 38761 55840 38801
rect 55927 38853 56632 38967
rect 57278 38853 57380 40601
rect 55927 38801 56015 38853
rect 56067 38801 56226 38853
rect 56278 38850 56437 38853
rect 56313 38804 56437 38850
rect 56278 38801 56437 38804
rect 56489 38801 56632 38853
rect 57278 38801 57281 38853
rect 57333 38801 57380 38853
rect 54817 38760 55579 38761
rect 48905 38715 49877 38755
rect 50099 38753 50255 38760
rect 48905 38709 48943 38715
rect 48995 38709 49154 38715
rect 49206 38709 49365 38715
rect 49417 38709 49576 38715
rect 49628 38709 49787 38715
rect 49839 38709 49877 38715
rect 30683 38641 31040 38681
rect 33484 38665 34643 38694
rect 30583 38564 31040 38641
rect 33019 38625 33327 38665
rect 33019 38622 33057 38625
rect 33109 38622 33237 38625
rect 33289 38622 33327 38625
rect 33484 38657 35082 38665
rect 35260 38663 35273 38709
rect 35523 38663 35543 38709
rect 35626 38663 35683 38709
rect 35729 38663 35754 38709
rect 35832 38663 35889 38709
rect 35935 38663 35965 38709
rect 36038 38663 36095 38709
rect 36141 38663 36176 38709
rect 36244 38663 36301 38709
rect 36347 38663 36360 38709
rect 36438 38663 36854 38709
rect 36900 38663 36971 38709
rect 37017 38663 37088 38709
rect 37134 38663 37206 38709
rect 37252 38663 37324 38709
rect 37370 38663 37442 38709
rect 37488 38665 37891 38709
rect 37488 38663 37909 38665
rect 37955 38663 38026 38709
rect 38123 38665 38143 38709
rect 38072 38663 38143 38665
rect 38189 38663 38261 38709
rect 38307 38663 38379 38709
rect 38425 38663 38497 38709
rect 38543 38663 38556 38709
rect 38658 38663 39021 38709
rect 39067 38663 39144 38709
rect 39190 38663 39267 38709
rect 39313 38663 39641 38709
rect 39687 38663 39730 38709
rect 31336 38576 31349 38622
rect 33323 38576 33336 38622
rect 33484 38611 33816 38657
rect 33862 38611 34002 38657
rect 34048 38611 34189 38657
rect 34235 38611 34376 38657
rect 34422 38611 34562 38657
rect 34608 38611 35082 38657
rect 35294 38623 36266 38663
rect 36438 38629 36953 38663
rect 37439 38629 38161 38663
rect 30583 38523 30855 38564
rect 30583 38477 30637 38523
rect 30683 38518 30855 38523
rect 30901 38518 31040 38564
rect 33019 38573 33057 38576
rect 33109 38573 33237 38576
rect 33289 38573 33327 38576
rect 33019 38532 33327 38573
rect 33484 38574 35082 38611
rect 30683 38477 31040 38518
rect 30583 38449 31040 38477
rect 33484 38492 33552 38574
rect 30583 38401 31493 38449
rect 30583 38360 30855 38401
rect 30583 38314 30637 38360
rect 30683 38355 30855 38360
rect 30901 38398 31493 38401
rect 30901 38355 31349 38398
rect 30683 38352 31349 38355
rect 33323 38352 33336 38398
rect 30683 38330 31493 38352
rect 30683 38314 31040 38330
rect 30583 38238 31040 38314
rect 30583 38197 30855 38238
rect 30583 38151 30637 38197
rect 30683 38192 30855 38197
rect 30901 38192 31040 38238
rect 30683 38151 31040 38192
rect 33019 38177 33327 38217
rect 33019 38174 33057 38177
rect 33109 38174 33237 38177
rect 33289 38174 33327 38177
rect 30583 38074 31040 38151
rect 31336 38128 31349 38174
rect 33323 38128 33336 38174
rect 33019 38125 33057 38128
rect 33109 38125 33237 38128
rect 33289 38125 33327 38128
rect 33019 38084 33327 38125
rect 30583 38034 30855 38074
rect 28492 37866 29196 37988
rect 28492 37820 28810 37866
rect 28856 37820 29196 37866
rect 29283 37953 30365 37994
rect 29283 37950 29582 37953
rect 29283 37904 29317 37950
rect 29363 37904 29478 37950
rect 29524 37904 29582 37950
rect 29283 37901 29582 37904
rect 29634 37950 29793 37953
rect 29845 37950 30005 37953
rect 29634 37904 29638 37950
rect 29684 37904 29793 37950
rect 29845 37904 29959 37950
rect 29634 37901 29793 37904
rect 29845 37901 30005 37904
rect 30057 37950 30216 37953
rect 30057 37904 30121 37950
rect 30167 37904 30216 37950
rect 30057 37901 30216 37904
rect 30268 37950 30365 37953
rect 30268 37904 30284 37950
rect 30330 37904 30365 37950
rect 30268 37901 30365 37904
rect 29283 37861 30365 37901
rect 30583 37988 30637 38034
rect 30683 38028 30855 38034
rect 30901 38028 31040 38074
rect 33484 38070 33495 38492
rect 33541 38070 33552 38492
rect 34964 38517 35082 38574
rect 36438 38529 36554 38629
rect 37853 38624 38161 38629
rect 38658 38649 39723 38663
rect 34964 38485 36360 38517
rect 34228 38415 34718 38456
rect 34228 38398 34267 38415
rect 34319 38398 34447 38415
rect 34499 38398 34627 38415
rect 33671 38352 33684 38398
rect 33730 38352 33787 38398
rect 33833 38352 33890 38398
rect 33936 38352 33993 38398
rect 34039 38352 34096 38398
rect 34142 38352 34199 38398
rect 34245 38363 34267 38398
rect 34245 38352 34302 38363
rect 34348 38352 34405 38398
rect 34499 38363 34508 38398
rect 34451 38352 34508 38363
rect 34554 38352 34612 38398
rect 34679 38363 34718 38415
rect 34964 38439 35273 38485
rect 35523 38439 35580 38485
rect 35626 38439 35683 38485
rect 35729 38439 35786 38485
rect 35832 38439 35889 38485
rect 35935 38439 35992 38485
rect 36038 38439 36095 38485
rect 36141 38439 36198 38485
rect 36244 38439 36301 38485
rect 36347 38439 36360 38485
rect 34964 38395 36360 38439
rect 34658 38352 34718 38363
rect 34228 38323 34718 38352
rect 36438 38389 36475 38529
rect 36521 38389 36554 38529
rect 35294 38261 36266 38295
rect 36438 38286 36554 38389
rect 36640 38529 36773 38549
rect 36640 38490 36697 38529
rect 36640 38438 36678 38490
rect 36640 38389 36697 38438
rect 36743 38389 36773 38529
rect 38658 38527 38726 38649
rect 39809 38643 44918 38681
rect 48765 38663 48778 38709
rect 48824 38663 48881 38709
rect 48927 38663 48943 38709
rect 49030 38663 49087 38709
rect 49133 38663 49154 38709
rect 49236 38663 49293 38709
rect 49339 38663 49365 38709
rect 49442 38663 49499 38709
rect 49545 38663 49576 38709
rect 49852 38663 49877 38709
rect 54085 38727 54540 38760
rect 50481 38667 51657 38694
rect 39809 38597 43739 38643
rect 43785 38597 43906 38643
rect 43952 38597 44071 38643
rect 44117 38597 44236 38643
rect 44282 38622 44918 38643
rect 48905 38623 49877 38663
rect 50044 38657 51657 38667
rect 44282 38597 44812 38622
rect 39809 38594 44812 38597
rect 39809 38548 39844 38594
rect 39890 38592 44812 38594
rect 39890 38548 39994 38592
rect 39809 38540 39994 38548
rect 40046 38576 44812 38592
rect 44858 38576 44925 38622
rect 44971 38576 45038 38622
rect 45084 38576 45151 38622
rect 45197 38576 45264 38622
rect 45310 38576 45323 38622
rect 48557 38577 48687 38617
rect 40046 38561 44918 38576
rect 40046 38540 40085 38561
rect 39809 38537 40085 38540
rect 36924 38517 37685 38524
rect 36923 38485 37931 38517
rect 36841 38439 36854 38485
rect 36900 38483 36971 38485
rect 36900 38439 36961 38483
rect 37017 38439 37088 38485
rect 37134 38483 37206 38485
rect 37134 38439 37172 38483
rect 37252 38439 37324 38485
rect 37370 38483 37442 38485
rect 37370 38439 37384 38483
rect 36923 38431 36961 38439
rect 37013 38431 37172 38439
rect 37224 38431 37384 38439
rect 37436 38439 37442 38483
rect 37488 38483 37909 38485
rect 37488 38439 37595 38483
rect 37436 38431 37595 38439
rect 37647 38439 37909 38483
rect 37955 38439 38026 38485
rect 38072 38439 38143 38485
rect 38189 38439 38261 38485
rect 38307 38439 38379 38485
rect 38425 38439 38497 38485
rect 38543 38439 38556 38485
rect 37647 38431 37931 38439
rect 36923 38398 37931 38431
rect 36923 38397 37685 38398
rect 36924 38391 37685 38397
rect 36640 38366 36773 38389
rect 38658 38387 38669 38527
rect 38715 38387 38726 38527
rect 39014 38485 39323 38517
rect 39492 38485 39608 38517
rect 39008 38439 39021 38485
rect 39067 38439 39144 38485
rect 39190 38439 39267 38485
rect 39313 38439 39326 38485
rect 39492 38439 39641 38485
rect 39687 38439 39730 38485
rect 38658 38376 38726 38387
rect 36438 38261 36953 38286
rect 37439 38283 37931 38286
rect 37439 38261 38161 38283
rect 35260 38215 35273 38261
rect 35523 38255 35580 38261
rect 35523 38215 35543 38255
rect 35626 38215 35683 38261
rect 35729 38255 35786 38261
rect 35729 38215 35754 38255
rect 35832 38215 35889 38261
rect 35935 38255 35992 38261
rect 35935 38215 35965 38255
rect 36038 38215 36095 38261
rect 36141 38255 36198 38261
rect 36141 38215 36176 38255
rect 36244 38215 36301 38261
rect 36347 38215 36360 38261
rect 36438 38215 36854 38261
rect 36900 38215 36971 38261
rect 37017 38215 37088 38261
rect 37134 38215 37206 38261
rect 37252 38215 37324 38261
rect 37370 38215 37442 38261
rect 37488 38243 37909 38261
rect 37488 38215 37891 38243
rect 37955 38215 38026 38261
rect 38072 38243 38143 38261
rect 38123 38215 38143 38243
rect 38189 38215 38261 38261
rect 38307 38215 38379 38261
rect 38425 38215 38497 38261
rect 38543 38215 38556 38261
rect 33781 38174 34089 38209
rect 35294 38203 35332 38215
rect 35384 38203 35543 38215
rect 35595 38203 35754 38215
rect 35806 38203 35965 38215
rect 36017 38203 36176 38215
rect 36228 38203 36266 38215
rect 33671 38128 33684 38174
rect 33730 38128 33787 38174
rect 33833 38169 33890 38174
rect 33871 38128 33890 38169
rect 33936 38128 33993 38174
rect 34039 38169 34096 38174
rect 34051 38128 34096 38169
rect 34142 38128 34199 38174
rect 34245 38128 34302 38174
rect 34348 38128 34405 38174
rect 34451 38128 34508 38174
rect 34554 38128 34612 38174
rect 34658 38128 34671 38174
rect 35294 38163 36266 38203
rect 36438 38166 36953 38215
rect 37439 38191 37891 38215
rect 37943 38191 38071 38215
rect 38123 38191 38161 38215
rect 37439 38166 38161 38191
rect 37853 38150 38161 38166
rect 33781 38117 33819 38128
rect 33871 38117 33999 38128
rect 34051 38117 34089 38128
rect 33781 38076 34089 38117
rect 33484 38059 33552 38070
rect 30683 37994 31040 38028
rect 30683 37988 32842 37994
rect 30583 37953 32842 37988
rect 34247 37987 35008 37994
rect 30583 37901 30854 37953
rect 30906 37901 31065 37953
rect 31117 37901 31276 37953
rect 31328 37950 31486 37953
rect 31538 37950 31697 37953
rect 31749 37950 31909 37953
rect 31961 37950 32120 37953
rect 32172 37950 32330 37953
rect 32382 37950 32541 37953
rect 32593 37950 32752 37953
rect 32804 37950 32842 37953
rect 34246 37953 35008 37987
rect 34246 37950 34284 37953
rect 34336 37950 34495 37953
rect 34547 37950 34707 37953
rect 31328 37904 31349 37950
rect 33323 37904 33336 37950
rect 33671 37904 33684 37950
rect 33730 37904 33787 37950
rect 33833 37904 33890 37950
rect 33936 37904 33993 37950
rect 34039 37904 34096 37950
rect 34142 37904 34199 37950
rect 34245 37904 34284 37950
rect 34348 37904 34405 37950
rect 34451 37904 34495 37950
rect 34554 37904 34612 37950
rect 34658 37904 34707 37950
rect 31328 37901 31486 37904
rect 31538 37901 31697 37904
rect 31749 37901 31909 37904
rect 31961 37901 32120 37904
rect 32172 37901 32330 37904
rect 32382 37901 32541 37904
rect 32593 37901 32752 37904
rect 32804 37901 32842 37904
rect 30583 37866 32842 37901
rect 34246 37901 34284 37904
rect 34336 37901 34495 37904
rect 34547 37901 34707 37904
rect 34759 37901 34918 37953
rect 34970 37901 35008 37953
rect 34246 37867 35008 37901
rect 29544 37860 30306 37861
rect 28492 37744 29196 37820
rect 28492 37703 29116 37744
rect 28492 37657 28810 37703
rect 28856 37698 29116 37703
rect 29162 37698 29196 37744
rect 28856 37657 29196 37698
rect 28492 37581 29196 37657
rect 28492 37540 29116 37581
rect 28492 37494 28810 37540
rect 28856 37535 29116 37540
rect 29162 37535 29196 37581
rect 28856 37494 29196 37535
rect 28492 37417 29196 37494
rect 28492 37377 29116 37417
rect 28492 37331 28810 37377
rect 28856 37371 29116 37377
rect 29162 37371 29196 37417
rect 28856 37331 29196 37371
rect 28492 37254 29196 37331
rect 28492 37213 29116 37254
rect 28492 37167 28810 37213
rect 28856 37208 29116 37213
rect 29162 37208 29196 37254
rect 28856 37167 29196 37208
rect 28492 37053 29196 37167
rect 30583 37820 30637 37866
rect 30683 37860 32842 37866
rect 34247 37860 35008 37867
rect 35182 37987 36364 37994
rect 35182 37953 36958 37987
rect 35182 37901 35220 37953
rect 35272 37901 35430 37953
rect 35482 37901 35641 37953
rect 35693 37901 35853 37953
rect 35905 37901 36064 37953
rect 36116 37901 36274 37953
rect 36326 37950 36958 37953
rect 36326 37904 36489 37950
rect 36723 37904 36958 37950
rect 36326 37901 36958 37904
rect 35182 37867 36958 37901
rect 37946 37953 38842 37994
rect 37946 37950 38330 37953
rect 38382 37950 38541 37953
rect 37946 37904 37957 37950
rect 38473 37904 38541 37950
rect 37946 37901 38330 37904
rect 38382 37901 38541 37904
rect 38593 37901 38752 37953
rect 38804 37901 38842 37953
rect 35182 37860 36364 37867
rect 37946 37860 38842 37901
rect 39014 37953 39323 38439
rect 39014 37901 39052 37953
rect 39104 37950 39232 37953
rect 39108 37904 39220 37950
rect 39104 37901 39232 37904
rect 39284 37901 39323 37953
rect 30683 37826 31040 37860
rect 30683 37820 30855 37826
rect 30583 37780 30855 37820
rect 30901 37780 31040 37826
rect 30583 37703 31040 37780
rect 33484 37784 33552 37795
rect 33019 37729 33327 37770
rect 33019 37726 33057 37729
rect 33109 37726 33237 37729
rect 33289 37726 33327 37729
rect 30583 37657 30637 37703
rect 30683 37662 31040 37703
rect 31336 37680 31349 37726
rect 33323 37680 33336 37726
rect 30683 37657 30855 37662
rect 30583 37616 30855 37657
rect 30901 37616 31040 37662
rect 33019 37677 33057 37680
rect 33109 37677 33237 37680
rect 33289 37677 33327 37680
rect 33019 37637 33327 37677
rect 30583 37540 31040 37616
rect 30583 37494 30637 37540
rect 30683 37524 31040 37540
rect 30683 37502 31493 37524
rect 30683 37499 31349 37502
rect 30683 37494 30855 37499
rect 30583 37453 30855 37494
rect 30901 37456 31349 37499
rect 33323 37456 33336 37502
rect 30901 37453 31493 37456
rect 30583 37405 31493 37453
rect 30583 37377 31040 37405
rect 30583 37331 30637 37377
rect 30683 37336 31040 37377
rect 30683 37331 30855 37336
rect 30583 37290 30855 37331
rect 30901 37290 31040 37336
rect 33484 37362 33495 37784
rect 33541 37362 33552 37784
rect 33781 37737 34089 37778
rect 33781 37726 33819 37737
rect 33871 37726 33999 37737
rect 34051 37726 34089 37737
rect 33671 37680 33684 37726
rect 33730 37680 33787 37726
rect 33871 37685 33890 37726
rect 33833 37680 33890 37685
rect 33936 37680 33993 37726
rect 34051 37685 34096 37726
rect 34039 37680 34096 37685
rect 34142 37680 34199 37726
rect 34245 37680 34302 37726
rect 34348 37680 34405 37726
rect 34451 37680 34508 37726
rect 34554 37680 34612 37726
rect 34658 37680 34671 37726
rect 33781 37645 34089 37680
rect 35294 37651 36266 37691
rect 37853 37688 38161 37704
rect 35294 37639 35332 37651
rect 35384 37639 35543 37651
rect 35595 37639 35754 37651
rect 35806 37639 35965 37651
rect 36017 37639 36176 37651
rect 36228 37639 36266 37651
rect 36438 37639 36953 37688
rect 37439 37663 38161 37688
rect 37439 37639 37891 37663
rect 37943 37639 38071 37663
rect 38123 37639 38161 37663
rect 35260 37593 35273 37639
rect 35523 37599 35543 37639
rect 35523 37593 35580 37599
rect 35626 37593 35683 37639
rect 35729 37599 35754 37639
rect 35729 37593 35786 37599
rect 35832 37593 35889 37639
rect 35935 37599 35965 37639
rect 35935 37593 35992 37599
rect 36038 37593 36095 37639
rect 36141 37599 36176 37639
rect 36141 37593 36198 37599
rect 36244 37593 36301 37639
rect 36347 37593 36360 37639
rect 36438 37593 36854 37639
rect 36900 37593 36971 37639
rect 37017 37593 37088 37639
rect 37134 37593 37206 37639
rect 37252 37593 37324 37639
rect 37370 37593 37442 37639
rect 37488 37611 37891 37639
rect 37488 37593 37909 37611
rect 37955 37593 38026 37639
rect 38123 37611 38143 37639
rect 38072 37593 38143 37611
rect 38189 37593 38261 37639
rect 38307 37593 38379 37639
rect 38425 37593 38497 37639
rect 38543 37593 38556 37639
rect 35294 37559 36266 37593
rect 36438 37568 36953 37593
rect 37439 37571 38161 37593
rect 37439 37568 37931 37571
rect 34228 37502 34718 37531
rect 33671 37456 33684 37502
rect 33730 37456 33787 37502
rect 33833 37456 33890 37502
rect 33936 37456 33993 37502
rect 34039 37456 34096 37502
rect 34142 37456 34199 37502
rect 34245 37491 34302 37502
rect 34245 37456 34267 37491
rect 34348 37456 34405 37502
rect 34451 37491 34508 37502
rect 34499 37456 34508 37491
rect 34554 37456 34612 37502
rect 34658 37491 34718 37502
rect 34228 37439 34267 37456
rect 34319 37439 34447 37456
rect 34499 37439 34627 37456
rect 34679 37439 34718 37491
rect 36438 37465 36554 37568
rect 34228 37398 34718 37439
rect 34964 37415 36360 37459
rect 30583 37213 31040 37290
rect 33019 37281 33327 37322
rect 33019 37278 33057 37281
rect 33109 37278 33237 37281
rect 33289 37278 33327 37281
rect 33484 37280 33552 37362
rect 34964 37369 35273 37415
rect 35523 37369 35580 37415
rect 35626 37369 35683 37415
rect 35729 37369 35786 37415
rect 35832 37369 35889 37415
rect 35935 37369 35992 37415
rect 36038 37369 36095 37415
rect 36141 37369 36198 37415
rect 36244 37369 36301 37415
rect 36347 37369 36360 37415
rect 34964 37337 36360 37369
rect 34964 37280 35082 37337
rect 31336 37232 31349 37278
rect 33323 37232 33336 37278
rect 33484 37243 35082 37280
rect 30583 37167 30637 37213
rect 30683 37173 31040 37213
rect 33019 37229 33057 37232
rect 33109 37229 33237 37232
rect 33289 37229 33327 37232
rect 33019 37189 33327 37229
rect 33484 37197 33816 37243
rect 33862 37197 34002 37243
rect 34048 37197 34189 37243
rect 34235 37197 34376 37243
rect 34422 37197 34562 37243
rect 34608 37197 35082 37243
rect 36438 37325 36475 37465
rect 36521 37325 36554 37465
rect 33484 37189 35082 37197
rect 35294 37191 36266 37231
rect 36438 37225 36554 37325
rect 36640 37465 36773 37488
rect 36640 37416 36697 37465
rect 36640 37364 36678 37416
rect 36640 37325 36697 37364
rect 36743 37325 36773 37465
rect 38658 37467 38726 37478
rect 36924 37457 37685 37463
rect 36923 37456 37685 37457
rect 36923 37423 37931 37456
rect 36923 37415 36961 37423
rect 37013 37415 37172 37423
rect 37224 37415 37384 37423
rect 36841 37369 36854 37415
rect 36900 37371 36961 37415
rect 36900 37369 36971 37371
rect 37017 37369 37088 37415
rect 37134 37371 37172 37415
rect 37134 37369 37206 37371
rect 37252 37369 37324 37415
rect 37370 37371 37384 37415
rect 37436 37415 37595 37423
rect 37436 37371 37442 37415
rect 37370 37369 37442 37371
rect 37488 37371 37595 37415
rect 37647 37415 37931 37423
rect 37647 37371 37909 37415
rect 37488 37369 37909 37371
rect 37955 37369 38026 37415
rect 38072 37369 38143 37415
rect 38189 37369 38261 37415
rect 38307 37369 38379 37415
rect 38425 37369 38497 37415
rect 38543 37369 38556 37415
rect 36923 37337 37931 37369
rect 36924 37330 37685 37337
rect 36640 37305 36773 37325
rect 38658 37327 38669 37467
rect 38715 37327 38726 37467
rect 39014 37415 39323 37901
rect 39492 37987 39608 38439
rect 39923 38406 40085 38537
rect 39923 38354 39994 38406
rect 40046 38354 40085 38406
rect 39923 38314 40085 38354
rect 39737 38218 39865 38231
rect 39737 38191 39866 38218
rect 39737 38174 39775 38191
rect 39827 38174 39866 38191
rect 39727 38128 39740 38174
rect 39827 38139 39862 38174
rect 39786 38128 39862 38139
rect 39908 38128 39985 38174
rect 40031 38128 40108 38174
rect 40154 38128 40167 38174
rect 40246 38163 40362 38561
rect 42229 38422 44509 38463
rect 42229 38370 43445 38422
rect 43497 38370 44509 38422
rect 42229 38330 44509 38370
rect 44341 38286 44509 38330
rect 44341 38240 44358 38286
rect 44498 38240 44509 38286
rect 39737 38099 39866 38128
rect 40246 38117 40281 38163
rect 40327 38117 40362 38163
rect 40246 38080 40362 38117
rect 40718 38191 43524 38232
rect 44341 38229 44509 38240
rect 40718 38139 41935 38191
rect 41987 38139 43524 38191
rect 40718 38098 43524 38139
rect 44605 38174 44721 38561
rect 45400 38531 48379 38572
rect 45400 38517 47486 38531
rect 45400 38471 45464 38517
rect 45604 38479 47486 38517
rect 47538 38479 48379 38531
rect 45604 38471 48379 38479
rect 44901 38415 45241 38456
rect 45400 38438 48379 38471
rect 48557 38525 48596 38577
rect 48648 38525 48687 38577
rect 48557 38502 48687 38525
rect 50044 38611 50516 38657
rect 50562 38611 50703 38657
rect 50749 38611 50890 38657
rect 50936 38611 51076 38657
rect 51122 38611 51263 38657
rect 51309 38611 51657 38657
rect 51797 38647 52105 38687
rect 51797 38622 51835 38647
rect 51887 38622 52015 38647
rect 52067 38622 52105 38647
rect 54085 38681 54223 38727
rect 54269 38687 54540 38727
rect 54269 38681 54440 38687
rect 54085 38641 54440 38681
rect 54486 38641 54540 38687
rect 50044 38574 51657 38611
rect 51789 38576 51802 38622
rect 53776 38576 53789 38622
rect 50044 38517 50160 38574
rect 44901 38398 44939 38415
rect 44991 38398 45151 38415
rect 45203 38398 45241 38415
rect 44799 38352 44812 38398
rect 44858 38352 44925 38398
rect 44991 38363 45038 38398
rect 44971 38352 45038 38363
rect 45084 38352 45151 38398
rect 45203 38363 45264 38398
rect 45197 38352 45264 38363
rect 45310 38352 45323 38398
rect 48557 38362 48622 38502
rect 48668 38362 48687 38502
rect 49820 38485 50160 38517
rect 48765 38439 48778 38485
rect 48824 38439 48881 38485
rect 48927 38439 48984 38485
rect 49030 38439 49087 38485
rect 49133 38439 49190 38485
rect 49236 38439 49293 38485
rect 49339 38439 49396 38485
rect 49442 38439 49499 38485
rect 49545 38439 49602 38485
rect 49852 38439 50160 38485
rect 51589 38522 51657 38574
rect 51797 38554 52105 38576
rect 49820 38398 50160 38439
rect 50262 38415 50812 38456
rect 48557 38359 48687 38362
rect 44901 38323 45241 38352
rect 48557 38307 48596 38359
rect 48648 38307 48687 38359
rect 50262 38363 50300 38415
rect 50352 38398 50511 38415
rect 50563 38398 50722 38415
rect 50352 38363 50467 38398
rect 50563 38363 50571 38398
rect 50262 38352 50467 38363
rect 50513 38352 50571 38363
rect 50617 38352 50674 38398
rect 50720 38363 50722 38398
rect 50774 38398 50812 38415
rect 50774 38363 50777 38398
rect 50720 38352 50777 38363
rect 50823 38352 50880 38398
rect 50926 38352 50983 38398
rect 51029 38352 51086 38398
rect 51132 38352 51189 38398
rect 51235 38352 51292 38398
rect 51338 38352 51395 38398
rect 51441 38352 51454 38398
rect 50262 38323 50812 38352
rect 48557 38266 48687 38307
rect 48905 38261 49877 38292
rect 48765 38215 48778 38261
rect 48824 38215 48881 38261
rect 48927 38252 48984 38261
rect 48927 38215 48943 38252
rect 49030 38215 49087 38261
rect 49133 38252 49190 38261
rect 49133 38215 49154 38252
rect 49236 38215 49293 38261
rect 49339 38252 49396 38261
rect 49339 38215 49365 38252
rect 49442 38215 49499 38261
rect 49545 38252 49602 38261
rect 49545 38215 49576 38252
rect 49852 38215 49877 38261
rect 48905 38200 48943 38215
rect 48995 38200 49154 38215
rect 49206 38200 49365 38215
rect 49417 38200 49576 38215
rect 49628 38200 49787 38215
rect 49839 38200 49877 38215
rect 44605 38128 44812 38174
rect 44858 38128 44925 38174
rect 44971 38128 45038 38174
rect 45084 38128 45151 38174
rect 45197 38128 45264 38174
rect 45310 38128 45323 38174
rect 48905 38160 49877 38200
rect 51035 38177 51343 38217
rect 51035 38174 51073 38177
rect 51125 38174 51253 38177
rect 51305 38174 51343 38177
rect 43362 38091 43524 38098
rect 43362 38045 43373 38091
rect 43513 38045 43524 38091
rect 43362 38034 43524 38045
rect 45584 38114 48546 38150
rect 50454 38128 50467 38174
rect 50513 38128 50571 38174
rect 50617 38128 50674 38174
rect 50720 38128 50777 38174
rect 50823 38128 50880 38174
rect 50926 38128 50983 38174
rect 51029 38128 51073 38174
rect 51132 38128 51189 38174
rect 51235 38128 51253 38174
rect 51338 38128 51395 38174
rect 51441 38128 51454 38174
rect 45584 38068 45619 38114
rect 45665 38068 45777 38114
rect 45823 38068 45935 38114
rect 45981 38068 46093 38114
rect 46139 38068 46251 38114
rect 46297 38068 46409 38114
rect 46455 38068 46568 38114
rect 46614 38068 46726 38114
rect 46772 38068 46884 38114
rect 46930 38068 47042 38114
rect 47088 38068 47200 38114
rect 47246 38068 47358 38114
rect 47404 38068 47516 38114
rect 47562 38068 47675 38114
rect 47721 38068 47833 38114
rect 47879 38068 47991 38114
rect 48037 38068 48149 38114
rect 48195 38068 48307 38114
rect 48353 38068 48465 38114
rect 48511 38068 48546 38114
rect 51035 38125 51073 38128
rect 51125 38125 51253 38128
rect 51305 38125 51343 38128
rect 51035 38084 51343 38125
rect 51589 38100 51600 38522
rect 51646 38100 51657 38522
rect 54085 38523 54540 38641
rect 54085 38477 54440 38523
rect 54486 38477 54540 38523
rect 54085 38449 54540 38477
rect 53585 38398 54540 38449
rect 51789 38352 51802 38398
rect 53776 38360 54540 38398
rect 53776 38352 54440 38360
rect 53585 38330 54440 38352
rect 54085 38314 54440 38330
rect 54486 38314 54540 38360
rect 54085 38238 54540 38314
rect 51797 38184 52105 38224
rect 51797 38174 51835 38184
rect 51887 38174 52015 38184
rect 52067 38174 52105 38184
rect 54085 38192 54223 38238
rect 54269 38197 54540 38238
rect 54269 38192 54440 38197
rect 51789 38128 51802 38174
rect 53776 38128 53789 38174
rect 54085 38151 54440 38192
rect 54486 38151 54540 38197
rect 51589 38089 51657 38100
rect 51797 38091 52105 38128
rect 40215 37987 40523 37994
rect 40788 37987 42986 38001
rect 43753 37987 44514 37994
rect 39492 37964 42986 37987
rect 43704 37964 44514 37987
rect 39492 37953 44514 37964
rect 39492 37950 40253 37953
rect 39492 37904 39740 37950
rect 39786 37904 39862 37950
rect 39908 37904 39985 37950
rect 40031 37904 40108 37950
rect 40154 37904 40253 37950
rect 39492 37901 40253 37904
rect 40305 37901 40433 37953
rect 40485 37950 43790 37953
rect 40485 37904 40836 37950
rect 40882 37904 40994 37950
rect 41040 37904 41152 37950
rect 41198 37904 41310 37950
rect 41356 37904 41469 37950
rect 41515 37904 41627 37950
rect 41673 37904 41785 37950
rect 41831 37904 41943 37950
rect 41989 37904 42101 37950
rect 42147 37904 42259 37950
rect 42305 37904 42418 37950
rect 42464 37904 42576 37950
rect 42622 37904 42734 37950
rect 42780 37904 42892 37950
rect 42938 37904 43739 37950
rect 43785 37904 43790 37950
rect 40485 37901 43790 37904
rect 43842 37950 44001 37953
rect 43842 37904 43906 37950
rect 43952 37904 44001 37950
rect 43842 37901 44001 37904
rect 44053 37950 44213 37953
rect 44265 37950 44424 37953
rect 44053 37904 44071 37950
rect 44117 37904 44213 37950
rect 44282 37904 44424 37950
rect 44053 37901 44213 37904
rect 44265 37901 44424 37904
rect 44476 37901 44514 37953
rect 39492 37890 44514 37901
rect 39492 37867 42986 37890
rect 43704 37867 44514 37890
rect 39492 37415 39608 37867
rect 40215 37860 40523 37867
rect 40788 37853 42986 37867
rect 43753 37860 44514 37867
rect 44796 37987 45346 37994
rect 45584 37987 48546 38068
rect 54085 38074 54540 38151
rect 54085 38028 54223 38074
rect 54269 38034 54540 38074
rect 54269 38028 54440 38034
rect 54085 37994 54440 38028
rect 48800 37987 49982 37994
rect 50308 37987 50859 37994
rect 44796 37953 49982 37987
rect 44796 37950 44834 37953
rect 44886 37950 45045 37953
rect 45097 37950 45256 37953
rect 45308 37950 48838 37953
rect 44796 37904 44812 37950
rect 44886 37904 44925 37950
rect 44971 37904 45038 37950
rect 45097 37904 45151 37950
rect 45197 37904 45256 37950
rect 45310 37904 45619 37950
rect 45665 37904 45777 37950
rect 45823 37904 45935 37950
rect 45981 37904 46093 37950
rect 46139 37904 46251 37950
rect 46297 37904 46409 37950
rect 46455 37904 46568 37950
rect 46614 37904 46726 37950
rect 46772 37904 46884 37950
rect 46930 37904 47042 37950
rect 47088 37904 47200 37950
rect 47246 37904 47358 37950
rect 47404 37904 47516 37950
rect 47562 37904 47675 37950
rect 47721 37904 47833 37950
rect 47879 37904 47991 37950
rect 48037 37904 48149 37950
rect 48195 37904 48307 37950
rect 48353 37904 48465 37950
rect 48511 37904 48838 37950
rect 44796 37901 44834 37904
rect 44886 37901 45045 37904
rect 45097 37901 45256 37904
rect 45308 37901 48838 37904
rect 48890 37901 49048 37953
rect 49100 37901 49259 37953
rect 49311 37901 49471 37953
rect 49523 37901 49682 37953
rect 49734 37901 49892 37953
rect 49944 37901 49982 37953
rect 44796 37867 49982 37901
rect 50307 37953 50859 37987
rect 50307 37901 50346 37953
rect 50398 37950 50557 37953
rect 50609 37950 50768 37953
rect 50820 37950 50859 37953
rect 52278 37988 54440 37994
rect 54486 37988 54540 38034
rect 55927 38687 56632 38801
rect 55927 38644 56267 38687
rect 55927 38598 55961 38644
rect 56007 38641 56267 38644
rect 56313 38641 56632 38687
rect 56007 38598 56632 38641
rect 55927 38523 56632 38598
rect 55927 38481 56267 38523
rect 55927 38435 55961 38481
rect 56007 38477 56267 38481
rect 56313 38477 56632 38523
rect 56007 38435 56632 38477
rect 55927 38360 56632 38435
rect 55927 38317 56267 38360
rect 55927 38271 55961 38317
rect 56007 38314 56267 38317
rect 56313 38314 56632 38360
rect 56007 38271 56632 38314
rect 55927 38197 56632 38271
rect 55927 38154 56267 38197
rect 55927 38108 55961 38154
rect 56007 38151 56267 38154
rect 56313 38151 56632 38197
rect 56007 38108 56632 38151
rect 55927 38034 56632 38108
rect 52278 37953 54540 37988
rect 52278 37950 52316 37953
rect 52368 37950 52527 37953
rect 52579 37950 52738 37953
rect 52790 37950 52948 37953
rect 53000 37950 53159 37953
rect 53211 37950 53371 37953
rect 53423 37950 53582 37953
rect 53634 37950 53792 37953
rect 50398 37904 50467 37950
rect 50513 37904 50557 37950
rect 50617 37904 50674 37950
rect 50720 37904 50768 37950
rect 50823 37904 50880 37950
rect 50926 37904 50983 37950
rect 51029 37904 51086 37950
rect 51132 37904 51189 37950
rect 51235 37904 51292 37950
rect 51338 37904 51395 37950
rect 51441 37904 51454 37950
rect 51789 37904 51802 37950
rect 53776 37904 53792 37950
rect 50398 37901 50557 37904
rect 50609 37901 50768 37904
rect 50820 37901 50859 37904
rect 50307 37867 50859 37901
rect 44796 37860 45346 37867
rect 43362 37809 43524 37820
rect 39737 37726 39866 37755
rect 40246 37737 40362 37774
rect 43362 37763 43373 37809
rect 43513 37763 43524 37809
rect 43362 37756 43524 37763
rect 39727 37680 39740 37726
rect 39786 37715 39862 37726
rect 39827 37680 39862 37715
rect 39908 37680 39985 37726
rect 40031 37680 40108 37726
rect 40154 37680 40167 37726
rect 40246 37691 40281 37737
rect 40327 37691 40362 37737
rect 39737 37663 39775 37680
rect 39827 37663 39866 37680
rect 39737 37636 39866 37663
rect 39737 37623 39865 37636
rect 39923 37500 40085 37540
rect 39923 37448 39994 37500
rect 40046 37448 40085 37500
rect 39008 37369 39021 37415
rect 39067 37369 39144 37415
rect 39190 37369 39267 37415
rect 39313 37369 39326 37415
rect 39492 37369 39641 37415
rect 39687 37369 39730 37415
rect 39014 37337 39323 37369
rect 39492 37337 39608 37369
rect 37853 37225 38161 37230
rect 36438 37191 36953 37225
rect 37439 37191 38161 37225
rect 38658 37205 38726 37327
rect 39923 37317 40085 37448
rect 39809 37314 40085 37317
rect 39809 37306 39994 37314
rect 39809 37260 39844 37306
rect 39890 37262 39994 37306
rect 40046 37293 40085 37314
rect 40246 37293 40362 37691
rect 40718 37715 43524 37756
rect 45584 37786 48546 37867
rect 48800 37860 49982 37867
rect 50308 37860 50859 37867
rect 52278 37901 52316 37904
rect 52368 37901 52527 37904
rect 52579 37901 52738 37904
rect 52790 37901 52948 37904
rect 53000 37901 53159 37904
rect 53211 37901 53371 37904
rect 53423 37901 53582 37904
rect 53634 37901 53792 37904
rect 53844 37901 54003 37953
rect 54055 37901 54214 37953
rect 54266 37901 54540 37953
rect 52278 37866 54540 37901
rect 52278 37860 54440 37866
rect 45584 37740 45619 37786
rect 45665 37740 45777 37786
rect 45823 37740 45935 37786
rect 45981 37740 46093 37786
rect 46139 37740 46251 37786
rect 46297 37740 46409 37786
rect 46455 37740 46568 37786
rect 46614 37740 46726 37786
rect 46772 37740 46884 37786
rect 46930 37740 47042 37786
rect 47088 37740 47200 37786
rect 47246 37740 47358 37786
rect 47404 37740 47516 37786
rect 47562 37740 47675 37786
rect 47721 37740 47833 37786
rect 47879 37740 47991 37786
rect 48037 37740 48149 37786
rect 48195 37740 48307 37786
rect 48353 37740 48465 37786
rect 48511 37740 48546 37786
rect 54085 37826 54440 37860
rect 54085 37780 54223 37826
rect 54269 37820 54440 37826
rect 54486 37820 54540 37866
rect 54758 37953 55840 37994
rect 54758 37950 54855 37953
rect 54758 37904 54793 37950
rect 54839 37904 54855 37950
rect 54758 37901 54855 37904
rect 54907 37950 55066 37953
rect 54907 37904 54956 37950
rect 55002 37904 55066 37950
rect 54907 37901 55066 37904
rect 55118 37950 55278 37953
rect 55330 37950 55489 37953
rect 55164 37904 55278 37950
rect 55330 37904 55439 37950
rect 55485 37904 55489 37950
rect 55118 37901 55278 37904
rect 55330 37901 55489 37904
rect 55541 37950 55840 37953
rect 55541 37904 55599 37950
rect 55645 37904 55760 37950
rect 55806 37904 55840 37950
rect 55541 37901 55840 37904
rect 54758 37861 55840 37901
rect 55927 37988 56267 38034
rect 56313 37988 56632 38034
rect 55927 37866 56632 37988
rect 54817 37860 55579 37861
rect 54269 37780 54540 37820
rect 40718 37663 41935 37715
rect 41987 37663 43524 37715
rect 40718 37622 43524 37663
rect 44605 37680 44812 37726
rect 44858 37680 44925 37726
rect 44971 37680 45038 37726
rect 45084 37680 45151 37726
rect 45197 37680 45264 37726
rect 45310 37680 45323 37726
rect 45584 37704 48546 37740
rect 51035 37729 51343 37770
rect 51035 37726 51073 37729
rect 51125 37726 51253 37729
rect 51305 37726 51343 37729
rect 51589 37754 51657 37765
rect 44341 37614 44509 37625
rect 44341 37568 44358 37614
rect 44498 37568 44509 37614
rect 44341 37524 44509 37568
rect 42229 37484 44509 37524
rect 42229 37432 43445 37484
rect 43497 37432 44509 37484
rect 42229 37391 44509 37432
rect 44605 37293 44721 37680
rect 48905 37654 49877 37694
rect 50454 37680 50467 37726
rect 50513 37680 50571 37726
rect 50617 37680 50674 37726
rect 50720 37680 50777 37726
rect 50823 37680 50880 37726
rect 50926 37680 50983 37726
rect 51029 37680 51073 37726
rect 51132 37680 51189 37726
rect 51235 37680 51253 37726
rect 51338 37680 51395 37726
rect 51441 37680 51454 37726
rect 48905 37639 48943 37654
rect 48995 37639 49154 37654
rect 49206 37639 49365 37654
rect 49417 37639 49576 37654
rect 49628 37639 49787 37654
rect 49839 37639 49877 37654
rect 48765 37593 48778 37639
rect 48824 37593 48881 37639
rect 48927 37602 48943 37639
rect 48927 37593 48984 37602
rect 49030 37593 49087 37639
rect 49133 37602 49154 37639
rect 49133 37593 49190 37602
rect 49236 37593 49293 37639
rect 49339 37602 49365 37639
rect 49339 37593 49396 37602
rect 49442 37593 49499 37639
rect 49545 37602 49576 37639
rect 49545 37593 49602 37602
rect 49852 37593 49877 37639
rect 51035 37677 51073 37680
rect 51125 37677 51253 37680
rect 51305 37677 51343 37680
rect 51035 37637 51343 37677
rect 48557 37547 48687 37588
rect 48905 37562 49877 37593
rect 44901 37502 45241 37531
rect 44799 37456 44812 37502
rect 44858 37456 44925 37502
rect 44971 37491 45038 37502
rect 44991 37456 45038 37491
rect 45084 37456 45151 37502
rect 45197 37491 45264 37502
rect 45203 37456 45264 37491
rect 45310 37456 45323 37502
rect 48557 37495 48596 37547
rect 48648 37495 48687 37547
rect 48557 37492 48687 37495
rect 44901 37439 44939 37456
rect 44991 37439 45151 37456
rect 45203 37439 45241 37456
rect 44901 37398 45241 37439
rect 45400 37383 48379 37416
rect 45400 37337 45464 37383
rect 45604 37375 48379 37383
rect 45604 37337 47864 37375
rect 45400 37323 47864 37337
rect 47916 37323 48379 37375
rect 40046 37278 44918 37293
rect 45400 37282 48379 37323
rect 48557 37352 48622 37492
rect 48668 37352 48687 37492
rect 50262 37502 50812 37531
rect 50262 37491 50467 37502
rect 50513 37491 50571 37502
rect 49820 37415 50160 37456
rect 48765 37369 48778 37415
rect 48824 37369 48881 37415
rect 48927 37369 48984 37415
rect 49030 37369 49087 37415
rect 49133 37369 49190 37415
rect 49236 37369 49293 37415
rect 49339 37369 49396 37415
rect 49442 37369 49499 37415
rect 49545 37369 49602 37415
rect 49852 37369 50160 37415
rect 50262 37439 50300 37491
rect 50352 37456 50467 37491
rect 50563 37456 50571 37491
rect 50617 37456 50674 37502
rect 50720 37491 50777 37502
rect 50720 37456 50722 37491
rect 50352 37439 50511 37456
rect 50563 37439 50722 37456
rect 50774 37456 50777 37491
rect 50823 37456 50880 37502
rect 50926 37456 50983 37502
rect 51029 37456 51086 37502
rect 51132 37456 51189 37502
rect 51235 37456 51292 37502
rect 51338 37456 51395 37502
rect 51441 37456 51454 37502
rect 50774 37439 50812 37456
rect 50262 37398 50812 37439
rect 48557 37329 48687 37352
rect 49820 37337 50160 37369
rect 40046 37262 44812 37278
rect 39890 37260 44812 37262
rect 39809 37257 44812 37260
rect 39809 37211 43739 37257
rect 43785 37211 43906 37257
rect 43952 37211 44071 37257
rect 44117 37211 44236 37257
rect 44282 37232 44812 37257
rect 44858 37232 44925 37278
rect 44971 37232 45038 37278
rect 45084 37232 45151 37278
rect 45197 37232 45264 37278
rect 45310 37232 45323 37278
rect 48557 37277 48596 37329
rect 48648 37277 48687 37329
rect 48557 37237 48687 37277
rect 50044 37280 50160 37337
rect 51589 37332 51600 37754
rect 51646 37332 51657 37754
rect 51797 37726 52105 37763
rect 51789 37680 51802 37726
rect 53776 37680 53789 37726
rect 54085 37703 54540 37780
rect 51797 37670 51835 37680
rect 51887 37670 52015 37680
rect 52067 37670 52105 37680
rect 51797 37630 52105 37670
rect 54085 37662 54440 37703
rect 54085 37616 54223 37662
rect 54269 37657 54440 37662
rect 54486 37657 54540 37703
rect 54269 37616 54540 37657
rect 54085 37540 54540 37616
rect 54085 37524 54440 37540
rect 53585 37502 54440 37524
rect 51789 37456 51802 37502
rect 53776 37494 54440 37502
rect 54486 37494 54540 37540
rect 53776 37456 54540 37494
rect 53585 37405 54540 37456
rect 51589 37280 51657 37332
rect 54085 37377 54540 37405
rect 54085 37331 54440 37377
rect 54486 37331 54540 37377
rect 50044 37243 51657 37280
rect 51797 37278 52105 37300
rect 44282 37211 44918 37232
rect 38658 37191 39723 37205
rect 30683 37167 30855 37173
rect 30583 37127 30855 37167
rect 30901 37127 31040 37173
rect 33484 37160 34643 37189
rect 35260 37145 35273 37191
rect 35523 37145 35543 37191
rect 35626 37145 35683 37191
rect 35729 37145 35754 37191
rect 35832 37145 35889 37191
rect 35935 37145 35965 37191
rect 36038 37145 36095 37191
rect 36141 37145 36176 37191
rect 36244 37145 36301 37191
rect 36347 37145 36360 37191
rect 36438 37145 36854 37191
rect 36900 37145 36971 37191
rect 37017 37145 37088 37191
rect 37134 37145 37206 37191
rect 37252 37145 37324 37191
rect 37370 37145 37442 37191
rect 37488 37189 37909 37191
rect 37488 37145 37891 37189
rect 37955 37145 38026 37191
rect 38072 37189 38143 37191
rect 38123 37145 38143 37189
rect 38189 37145 38261 37191
rect 38307 37145 38379 37191
rect 38425 37145 38497 37191
rect 38543 37145 38556 37191
rect 38658 37145 39021 37191
rect 39067 37145 39144 37191
rect 39190 37145 39267 37191
rect 39313 37145 39641 37191
rect 39687 37145 39730 37191
rect 39809 37173 44918 37211
rect 48905 37191 49877 37231
rect 48765 37145 48778 37191
rect 48824 37145 48881 37191
rect 48927 37145 48943 37191
rect 49030 37145 49087 37191
rect 49133 37145 49154 37191
rect 49236 37145 49293 37191
rect 49339 37145 49365 37191
rect 49442 37145 49499 37191
rect 49545 37145 49576 37191
rect 49852 37145 49877 37191
rect 50044 37197 50516 37243
rect 50562 37197 50703 37243
rect 50749 37197 50890 37243
rect 50936 37197 51076 37243
rect 51122 37197 51263 37243
rect 51309 37197 51657 37243
rect 51789 37232 51802 37278
rect 53776 37232 53789 37278
rect 50044 37187 51657 37197
rect 50481 37160 51657 37187
rect 51797 37207 51835 37232
rect 51887 37207 52015 37232
rect 52067 37207 52105 37232
rect 51797 37167 52105 37207
rect 54085 37213 54540 37331
rect 54085 37173 54440 37213
rect 30583 37094 31040 37127
rect 35294 37139 35332 37145
rect 35384 37139 35543 37145
rect 35595 37139 35754 37145
rect 35806 37139 35965 37145
rect 36017 37139 36176 37145
rect 36228 37139 36266 37145
rect 34870 37094 35025 37101
rect 35294 37099 36266 37139
rect 36438 37105 36953 37145
rect 37439 37137 37891 37145
rect 37943 37137 38071 37145
rect 38123 37137 38161 37145
rect 37439 37105 38161 37137
rect 37853 37097 38161 37105
rect 27744 37001 27790 37053
rect 27842 37001 27846 37053
rect 28492 37001 28634 37053
rect 28686 37050 28845 37053
rect 28686 37004 28810 37050
rect 28686 37001 28845 37004
rect 28897 37001 29056 37053
rect 29108 37001 29196 37053
rect 27744 35996 27846 37001
rect 28492 36887 29196 37001
rect 29283 37053 30365 37094
rect 29283 37050 29582 37053
rect 29283 37004 29317 37050
rect 29363 37004 29478 37050
rect 29524 37004 29582 37050
rect 29283 37001 29582 37004
rect 29634 37050 29793 37053
rect 29845 37050 30005 37053
rect 29634 37004 29638 37050
rect 29684 37004 29793 37050
rect 29845 37004 29959 37050
rect 29634 37001 29793 37004
rect 29845 37001 30005 37004
rect 30057 37050 30216 37053
rect 30057 37004 30121 37050
rect 30167 37004 30216 37050
rect 30057 37001 30216 37004
rect 30268 37050 30365 37053
rect 30268 37004 30284 37050
rect 30330 37004 30365 37050
rect 30268 37001 30365 37004
rect 29283 36961 30365 37001
rect 30583 37053 32842 37094
rect 30583 37050 30854 37053
rect 30583 37004 30637 37050
rect 30683 37004 30854 37050
rect 30583 37001 30854 37004
rect 30906 37001 31065 37053
rect 31117 37001 31276 37053
rect 31328 37001 31486 37053
rect 31538 37001 31697 37053
rect 31749 37001 31909 37053
rect 31961 37001 32120 37053
rect 32172 37001 32330 37053
rect 32382 37001 32541 37053
rect 32593 37001 32752 37053
rect 32804 37001 32842 37053
rect 29544 36960 30306 36961
rect 30583 36960 32842 37001
rect 34717 37053 35025 37094
rect 38658 37085 39723 37145
rect 48905 37139 48943 37145
rect 48995 37139 49154 37145
rect 49206 37139 49365 37145
rect 49417 37139 49576 37145
rect 49628 37139 49787 37145
rect 49839 37139 49877 37145
rect 48905 37099 49877 37139
rect 54085 37127 54223 37173
rect 54269 37167 54440 37173
rect 54486 37167 54540 37213
rect 54269 37127 54540 37167
rect 50099 37094 50255 37101
rect 54085 37094 54540 37127
rect 55927 37820 56267 37866
rect 56313 37820 56632 37866
rect 55927 37744 56632 37820
rect 55927 37698 55961 37744
rect 56007 37703 56632 37744
rect 56007 37698 56267 37703
rect 55927 37657 56267 37698
rect 56313 37657 56632 37703
rect 55927 37581 56632 37657
rect 55927 37535 55961 37581
rect 56007 37540 56632 37581
rect 56007 37535 56267 37540
rect 55927 37494 56267 37535
rect 56313 37494 56632 37540
rect 55927 37417 56632 37494
rect 55927 37371 55961 37417
rect 56007 37377 56632 37417
rect 56007 37371 56267 37377
rect 55927 37331 56267 37371
rect 56313 37331 56632 37377
rect 55927 37254 56632 37331
rect 55927 37208 55961 37254
rect 56007 37213 56632 37254
rect 56007 37208 56267 37213
rect 55927 37167 56267 37208
rect 56313 37167 56632 37213
rect 34717 37001 34755 37053
rect 34807 37050 34935 37053
rect 34807 37004 34916 37050
rect 34807 37001 34935 37004
rect 34987 37001 35025 37053
rect 34717 36960 35025 37001
rect 50099 37053 50408 37094
rect 50099 37001 50138 37053
rect 50190 37050 50318 37053
rect 50206 37004 50318 37050
rect 50190 37001 50318 37004
rect 50370 37001 50408 37053
rect 28492 36841 28810 36887
rect 28856 36844 29196 36887
rect 28856 36841 29116 36844
rect 28492 36798 29116 36841
rect 29162 36798 29196 36844
rect 28492 36723 29196 36798
rect 28492 36677 28810 36723
rect 28856 36681 29196 36723
rect 28856 36677 29116 36681
rect 28492 36635 29116 36677
rect 29162 36635 29196 36681
rect 28492 36560 29196 36635
rect 28492 36514 28810 36560
rect 28856 36517 29196 36560
rect 28856 36514 29116 36517
rect 28492 36471 29116 36514
rect 29162 36471 29196 36517
rect 28492 36397 29196 36471
rect 28492 36351 28810 36397
rect 28856 36354 29196 36397
rect 28856 36351 29116 36354
rect 28492 36308 29116 36351
rect 29162 36308 29196 36354
rect 28492 36234 29196 36308
rect 28492 36188 28810 36234
rect 28856 36188 29196 36234
rect 30583 36927 31040 36960
rect 34870 36953 35025 36960
rect 30583 36887 30855 36927
rect 30583 36841 30637 36887
rect 30683 36881 30855 36887
rect 30901 36881 31040 36927
rect 35294 36915 36266 36955
rect 37853 36949 38161 36957
rect 35294 36909 35332 36915
rect 35384 36909 35543 36915
rect 35595 36909 35754 36915
rect 35806 36909 35965 36915
rect 36017 36909 36176 36915
rect 36228 36909 36266 36915
rect 36438 36909 36953 36949
rect 37439 36917 38161 36949
rect 37439 36909 37891 36917
rect 37943 36909 38071 36917
rect 38123 36909 38161 36917
rect 38658 36909 39723 36969
rect 50099 36960 50408 37001
rect 52278 37053 54540 37094
rect 52278 37001 52316 37053
rect 52368 37001 52527 37053
rect 52579 37001 52738 37053
rect 52790 37001 52948 37053
rect 53000 37001 53159 37053
rect 53211 37001 53371 37053
rect 53423 37001 53582 37053
rect 53634 37001 53792 37053
rect 53844 37001 54003 37053
rect 54055 37001 54214 37053
rect 54266 37050 54540 37053
rect 54266 37004 54440 37050
rect 54486 37004 54540 37050
rect 54266 37001 54540 37004
rect 52278 36960 54540 37001
rect 54758 37053 55840 37094
rect 54758 37050 54855 37053
rect 54758 37004 54793 37050
rect 54839 37004 54855 37050
rect 54758 37001 54855 37004
rect 54907 37050 55066 37053
rect 54907 37004 54956 37050
rect 55002 37004 55066 37050
rect 54907 37001 55066 37004
rect 55118 37050 55278 37053
rect 55330 37050 55489 37053
rect 55164 37004 55278 37050
rect 55330 37004 55439 37050
rect 55485 37004 55489 37050
rect 55118 37001 55278 37004
rect 55330 37001 55489 37004
rect 55541 37050 55840 37053
rect 55541 37004 55599 37050
rect 55645 37004 55760 37050
rect 55806 37004 55840 37050
rect 55541 37001 55840 37004
rect 54758 36961 55840 37001
rect 55927 37053 56632 37167
rect 57278 37053 57380 38801
rect 55927 37001 56015 37053
rect 56067 37001 56226 37053
rect 56278 37050 56437 37053
rect 56313 37004 56437 37050
rect 56278 37001 56437 37004
rect 56489 37001 56632 37053
rect 57278 37001 57281 37053
rect 57333 37001 57380 37053
rect 54817 36960 55579 36961
rect 48905 36915 49877 36955
rect 50099 36953 50255 36960
rect 48905 36909 48943 36915
rect 48995 36909 49154 36915
rect 49206 36909 49365 36915
rect 49417 36909 49576 36915
rect 49628 36909 49787 36915
rect 49839 36909 49877 36915
rect 30683 36841 31040 36881
rect 33484 36865 34643 36894
rect 30583 36764 31040 36841
rect 33019 36825 33327 36865
rect 33019 36822 33057 36825
rect 33109 36822 33237 36825
rect 33289 36822 33327 36825
rect 33484 36857 35082 36865
rect 35260 36863 35273 36909
rect 35523 36863 35543 36909
rect 35626 36863 35683 36909
rect 35729 36863 35754 36909
rect 35832 36863 35889 36909
rect 35935 36863 35965 36909
rect 36038 36863 36095 36909
rect 36141 36863 36176 36909
rect 36244 36863 36301 36909
rect 36347 36863 36360 36909
rect 36438 36863 36854 36909
rect 36900 36863 36971 36909
rect 37017 36863 37088 36909
rect 37134 36863 37206 36909
rect 37252 36863 37324 36909
rect 37370 36863 37442 36909
rect 37488 36865 37891 36909
rect 37488 36863 37909 36865
rect 37955 36863 38026 36909
rect 38123 36865 38143 36909
rect 38072 36863 38143 36865
rect 38189 36863 38261 36909
rect 38307 36863 38379 36909
rect 38425 36863 38497 36909
rect 38543 36863 38556 36909
rect 38658 36863 39021 36909
rect 39067 36863 39144 36909
rect 39190 36863 39267 36909
rect 39313 36863 39641 36909
rect 39687 36863 39730 36909
rect 31336 36776 31349 36822
rect 33323 36776 33336 36822
rect 33484 36811 33816 36857
rect 33862 36811 34002 36857
rect 34048 36811 34189 36857
rect 34235 36811 34376 36857
rect 34422 36811 34562 36857
rect 34608 36811 35082 36857
rect 35294 36823 36266 36863
rect 36438 36829 36953 36863
rect 37439 36829 38161 36863
rect 30583 36723 30855 36764
rect 30583 36677 30637 36723
rect 30683 36718 30855 36723
rect 30901 36718 31040 36764
rect 33019 36773 33057 36776
rect 33109 36773 33237 36776
rect 33289 36773 33327 36776
rect 33019 36732 33327 36773
rect 33484 36774 35082 36811
rect 30683 36677 31040 36718
rect 30583 36649 31040 36677
rect 33484 36692 33552 36774
rect 30583 36601 31493 36649
rect 30583 36560 30855 36601
rect 30583 36514 30637 36560
rect 30683 36555 30855 36560
rect 30901 36598 31493 36601
rect 30901 36555 31349 36598
rect 30683 36552 31349 36555
rect 33323 36552 33336 36598
rect 30683 36530 31493 36552
rect 30683 36514 31040 36530
rect 30583 36438 31040 36514
rect 30583 36397 30855 36438
rect 30583 36351 30637 36397
rect 30683 36392 30855 36397
rect 30901 36392 31040 36438
rect 30683 36351 31040 36392
rect 33019 36377 33327 36417
rect 33019 36374 33057 36377
rect 33109 36374 33237 36377
rect 33289 36374 33327 36377
rect 30583 36274 31040 36351
rect 31336 36328 31349 36374
rect 33323 36328 33336 36374
rect 33019 36325 33057 36328
rect 33109 36325 33237 36328
rect 33289 36325 33327 36328
rect 33019 36284 33327 36325
rect 30583 36234 30855 36274
rect 28492 36027 29196 36188
rect 29283 36153 30365 36194
rect 29283 36150 29582 36153
rect 29283 36104 29317 36150
rect 29363 36104 29478 36150
rect 29524 36104 29582 36150
rect 29283 36101 29582 36104
rect 29634 36150 29793 36153
rect 29845 36150 30005 36153
rect 29634 36104 29638 36150
rect 29684 36104 29793 36150
rect 29845 36104 29959 36150
rect 29634 36101 29793 36104
rect 29845 36101 30005 36104
rect 30057 36150 30216 36153
rect 30057 36104 30121 36150
rect 30167 36104 30216 36150
rect 30057 36101 30216 36104
rect 30268 36150 30365 36153
rect 30268 36104 30284 36150
rect 30330 36104 30365 36150
rect 30268 36101 30365 36104
rect 29283 36061 30365 36101
rect 30583 36188 30637 36234
rect 30683 36228 30855 36234
rect 30901 36228 31040 36274
rect 33484 36270 33495 36692
rect 33541 36270 33552 36692
rect 34964 36717 35082 36774
rect 36438 36729 36554 36829
rect 37853 36824 38161 36829
rect 38658 36849 39723 36863
rect 34964 36685 36360 36717
rect 34228 36615 34718 36656
rect 34228 36598 34267 36615
rect 34319 36598 34447 36615
rect 34499 36598 34627 36615
rect 33671 36552 33684 36598
rect 33730 36552 33787 36598
rect 33833 36552 33890 36598
rect 33936 36552 33993 36598
rect 34039 36552 34096 36598
rect 34142 36552 34199 36598
rect 34245 36563 34267 36598
rect 34245 36552 34302 36563
rect 34348 36552 34405 36598
rect 34499 36563 34508 36598
rect 34451 36552 34508 36563
rect 34554 36552 34612 36598
rect 34679 36563 34718 36615
rect 34964 36639 35273 36685
rect 35523 36639 35580 36685
rect 35626 36639 35683 36685
rect 35729 36639 35786 36685
rect 35832 36639 35889 36685
rect 35935 36639 35992 36685
rect 36038 36639 36095 36685
rect 36141 36639 36198 36685
rect 36244 36639 36301 36685
rect 36347 36639 36360 36685
rect 34964 36595 36360 36639
rect 34658 36552 34718 36563
rect 34228 36523 34718 36552
rect 36438 36589 36475 36729
rect 36521 36589 36554 36729
rect 35294 36461 36266 36495
rect 36438 36486 36554 36589
rect 36640 36729 36773 36749
rect 36640 36690 36697 36729
rect 36640 36638 36678 36690
rect 36640 36589 36697 36638
rect 36743 36589 36773 36729
rect 38658 36727 38726 36849
rect 39809 36843 44918 36881
rect 48765 36863 48778 36909
rect 48824 36863 48881 36909
rect 48927 36863 48943 36909
rect 49030 36863 49087 36909
rect 49133 36863 49154 36909
rect 49236 36863 49293 36909
rect 49339 36863 49365 36909
rect 49442 36863 49499 36909
rect 49545 36863 49576 36909
rect 49852 36863 49877 36909
rect 54085 36927 54540 36960
rect 50481 36867 51657 36894
rect 39809 36797 43739 36843
rect 43785 36797 43906 36843
rect 43952 36797 44071 36843
rect 44117 36797 44236 36843
rect 44282 36822 44918 36843
rect 48905 36823 49877 36863
rect 50044 36857 51657 36867
rect 44282 36797 44812 36822
rect 39809 36794 44812 36797
rect 39809 36748 39844 36794
rect 39890 36792 44812 36794
rect 39890 36748 39994 36792
rect 39809 36740 39994 36748
rect 40046 36776 44812 36792
rect 44858 36776 44925 36822
rect 44971 36776 45038 36822
rect 45084 36776 45151 36822
rect 45197 36776 45264 36822
rect 45310 36776 45323 36822
rect 48557 36777 48687 36817
rect 40046 36761 44918 36776
rect 40046 36740 40085 36761
rect 39809 36737 40085 36740
rect 36924 36717 37685 36724
rect 36923 36685 37931 36717
rect 36841 36639 36854 36685
rect 36900 36683 36971 36685
rect 36900 36639 36961 36683
rect 37017 36639 37088 36685
rect 37134 36683 37206 36685
rect 37134 36639 37172 36683
rect 37252 36639 37324 36685
rect 37370 36683 37442 36685
rect 37370 36639 37384 36683
rect 36923 36631 36961 36639
rect 37013 36631 37172 36639
rect 37224 36631 37384 36639
rect 37436 36639 37442 36683
rect 37488 36683 37909 36685
rect 37488 36639 37595 36683
rect 37436 36631 37595 36639
rect 37647 36639 37909 36683
rect 37955 36639 38026 36685
rect 38072 36639 38143 36685
rect 38189 36639 38261 36685
rect 38307 36639 38379 36685
rect 38425 36639 38497 36685
rect 38543 36639 38556 36685
rect 37647 36631 37931 36639
rect 36923 36598 37931 36631
rect 36923 36597 37685 36598
rect 36924 36591 37685 36597
rect 36640 36566 36773 36589
rect 38658 36587 38669 36727
rect 38715 36587 38726 36727
rect 39014 36685 39323 36717
rect 39492 36685 39608 36717
rect 39008 36639 39021 36685
rect 39067 36639 39144 36685
rect 39190 36639 39267 36685
rect 39313 36639 39326 36685
rect 39492 36639 39641 36685
rect 39687 36639 39730 36685
rect 38658 36576 38726 36587
rect 36438 36461 36953 36486
rect 37439 36483 37931 36486
rect 37439 36461 38161 36483
rect 35260 36415 35273 36461
rect 35523 36455 35580 36461
rect 35523 36415 35543 36455
rect 35626 36415 35683 36461
rect 35729 36455 35786 36461
rect 35729 36415 35754 36455
rect 35832 36415 35889 36461
rect 35935 36455 35992 36461
rect 35935 36415 35965 36455
rect 36038 36415 36095 36461
rect 36141 36455 36198 36461
rect 36141 36415 36176 36455
rect 36244 36415 36301 36461
rect 36347 36415 36360 36461
rect 36438 36415 36854 36461
rect 36900 36415 36971 36461
rect 37017 36415 37088 36461
rect 37134 36415 37206 36461
rect 37252 36415 37324 36461
rect 37370 36415 37442 36461
rect 37488 36443 37909 36461
rect 37488 36415 37891 36443
rect 37955 36415 38026 36461
rect 38072 36443 38143 36461
rect 38123 36415 38143 36443
rect 38189 36415 38261 36461
rect 38307 36415 38379 36461
rect 38425 36415 38497 36461
rect 38543 36415 38556 36461
rect 33781 36374 34089 36409
rect 35294 36403 35332 36415
rect 35384 36403 35543 36415
rect 35595 36403 35754 36415
rect 35806 36403 35965 36415
rect 36017 36403 36176 36415
rect 36228 36403 36266 36415
rect 33671 36328 33684 36374
rect 33730 36328 33787 36374
rect 33833 36369 33890 36374
rect 33871 36328 33890 36369
rect 33936 36328 33993 36374
rect 34039 36369 34096 36374
rect 34051 36328 34096 36369
rect 34142 36328 34199 36374
rect 34245 36328 34302 36374
rect 34348 36328 34405 36374
rect 34451 36328 34508 36374
rect 34554 36328 34612 36374
rect 34658 36328 34671 36374
rect 35294 36363 36266 36403
rect 36438 36366 36953 36415
rect 37439 36391 37891 36415
rect 37943 36391 38071 36415
rect 38123 36391 38161 36415
rect 37439 36366 38161 36391
rect 37853 36350 38161 36366
rect 33781 36317 33819 36328
rect 33871 36317 33999 36328
rect 34051 36317 34089 36328
rect 33781 36276 34089 36317
rect 33484 36259 33552 36270
rect 30683 36194 31040 36228
rect 30683 36188 32842 36194
rect 30583 36153 32842 36188
rect 34247 36187 35008 36194
rect 30583 36101 30854 36153
rect 30906 36101 31065 36153
rect 31117 36101 31276 36153
rect 31328 36150 31486 36153
rect 31538 36150 31697 36153
rect 31749 36150 31909 36153
rect 31961 36150 32120 36153
rect 32172 36150 32330 36153
rect 32382 36150 32541 36153
rect 32593 36150 32752 36153
rect 32804 36150 32842 36153
rect 34246 36153 35008 36187
rect 34246 36150 34284 36153
rect 34336 36150 34495 36153
rect 34547 36150 34707 36153
rect 31328 36104 31349 36150
rect 33323 36104 33336 36150
rect 33671 36104 33684 36150
rect 33730 36104 33787 36150
rect 33833 36104 33890 36150
rect 33936 36104 33993 36150
rect 34039 36104 34096 36150
rect 34142 36104 34199 36150
rect 34245 36104 34284 36150
rect 34348 36104 34405 36150
rect 34451 36104 34495 36150
rect 34554 36104 34612 36150
rect 34658 36104 34707 36150
rect 31328 36101 31486 36104
rect 31538 36101 31697 36104
rect 31749 36101 31909 36104
rect 31961 36101 32120 36104
rect 32172 36101 32330 36104
rect 32382 36101 32541 36104
rect 32593 36101 32752 36104
rect 32804 36101 32842 36104
rect 30583 36061 32842 36101
rect 34246 36101 34284 36104
rect 34336 36101 34495 36104
rect 34547 36101 34707 36104
rect 34759 36101 34918 36153
rect 34970 36101 35008 36153
rect 34246 36067 35008 36101
rect 34247 36061 35008 36067
rect 35182 36187 36364 36194
rect 35182 36153 36958 36187
rect 35182 36101 35220 36153
rect 35272 36101 35430 36153
rect 35482 36101 35641 36153
rect 35693 36101 35853 36153
rect 35905 36101 36064 36153
rect 36116 36101 36274 36153
rect 36326 36150 36958 36153
rect 36326 36104 36489 36150
rect 36723 36104 36958 36150
rect 36326 36101 36958 36104
rect 35182 36067 36958 36101
rect 37946 36153 38842 36194
rect 37946 36150 38330 36153
rect 38382 36150 38541 36153
rect 37946 36104 37957 36150
rect 38473 36104 38541 36150
rect 37946 36101 38330 36104
rect 38382 36101 38541 36104
rect 38593 36101 38752 36153
rect 38804 36101 38842 36153
rect 29544 36060 30306 36061
rect 30748 36060 32842 36061
rect 35182 36060 36364 36067
rect 37946 36061 38842 36101
rect 39014 36153 39323 36639
rect 39014 36101 39052 36153
rect 39104 36150 39232 36153
rect 39108 36104 39220 36150
rect 39104 36101 39232 36104
rect 39284 36101 39323 36153
rect 39014 36067 39323 36101
rect 39492 36187 39608 36639
rect 39923 36606 40085 36737
rect 39923 36554 39994 36606
rect 40046 36554 40085 36606
rect 39923 36514 40085 36554
rect 39737 36418 39865 36431
rect 39737 36391 39866 36418
rect 39737 36374 39775 36391
rect 39827 36374 39866 36391
rect 39727 36328 39740 36374
rect 39827 36339 39862 36374
rect 39786 36328 39862 36339
rect 39908 36328 39985 36374
rect 40031 36328 40108 36374
rect 40154 36328 40167 36374
rect 40246 36363 40362 36761
rect 42229 36622 44509 36663
rect 42229 36570 43445 36622
rect 43497 36570 44509 36622
rect 42229 36530 44509 36570
rect 44341 36486 44509 36530
rect 44341 36440 44358 36486
rect 44498 36440 44509 36486
rect 39737 36299 39866 36328
rect 40246 36317 40281 36363
rect 40327 36317 40362 36363
rect 40246 36280 40362 36317
rect 40718 36391 43524 36432
rect 44341 36429 44509 36440
rect 40718 36339 41935 36391
rect 41987 36339 43524 36391
rect 40718 36298 43524 36339
rect 44605 36374 44721 36761
rect 45400 36731 48379 36772
rect 45400 36717 48241 36731
rect 45400 36671 45464 36717
rect 45604 36679 48241 36717
rect 48293 36679 48379 36731
rect 45604 36671 48379 36679
rect 44901 36615 45241 36656
rect 45400 36638 48379 36671
rect 48557 36725 48596 36777
rect 48648 36725 48687 36777
rect 48557 36702 48687 36725
rect 50044 36811 50516 36857
rect 50562 36811 50703 36857
rect 50749 36811 50890 36857
rect 50936 36811 51076 36857
rect 51122 36811 51263 36857
rect 51309 36811 51657 36857
rect 51797 36847 52105 36887
rect 51797 36822 51835 36847
rect 51887 36822 52015 36847
rect 52067 36822 52105 36847
rect 54085 36881 54223 36927
rect 54269 36887 54540 36927
rect 54269 36881 54440 36887
rect 54085 36841 54440 36881
rect 54486 36841 54540 36887
rect 50044 36774 51657 36811
rect 51789 36776 51802 36822
rect 53776 36776 53789 36822
rect 50044 36717 50160 36774
rect 44901 36598 44939 36615
rect 44991 36598 45151 36615
rect 45203 36598 45241 36615
rect 44799 36552 44812 36598
rect 44858 36552 44925 36598
rect 44991 36563 45038 36598
rect 44971 36552 45038 36563
rect 45084 36552 45151 36598
rect 45203 36563 45264 36598
rect 45197 36552 45264 36563
rect 45310 36552 45323 36598
rect 48557 36562 48622 36702
rect 48668 36562 48687 36702
rect 49820 36685 50160 36717
rect 48765 36639 48778 36685
rect 48824 36639 48881 36685
rect 48927 36639 48984 36685
rect 49030 36639 49087 36685
rect 49133 36639 49190 36685
rect 49236 36639 49293 36685
rect 49339 36639 49396 36685
rect 49442 36639 49499 36685
rect 49545 36639 49602 36685
rect 49852 36639 50160 36685
rect 51589 36722 51657 36774
rect 51797 36754 52105 36776
rect 49820 36598 50160 36639
rect 50262 36615 50812 36656
rect 48557 36559 48687 36562
rect 44901 36523 45241 36552
rect 48557 36507 48596 36559
rect 48648 36507 48687 36559
rect 50262 36563 50300 36615
rect 50352 36598 50511 36615
rect 50563 36598 50722 36615
rect 50352 36563 50467 36598
rect 50563 36563 50571 36598
rect 50262 36552 50467 36563
rect 50513 36552 50571 36563
rect 50617 36552 50674 36598
rect 50720 36563 50722 36598
rect 50774 36598 50812 36615
rect 50774 36563 50777 36598
rect 50720 36552 50777 36563
rect 50823 36552 50880 36598
rect 50926 36552 50983 36598
rect 51029 36552 51086 36598
rect 51132 36552 51189 36598
rect 51235 36552 51292 36598
rect 51338 36552 51395 36598
rect 51441 36552 51454 36598
rect 50262 36523 50812 36552
rect 48557 36466 48687 36507
rect 48905 36461 49877 36492
rect 48765 36415 48778 36461
rect 48824 36415 48881 36461
rect 48927 36452 48984 36461
rect 48927 36415 48943 36452
rect 49030 36415 49087 36461
rect 49133 36452 49190 36461
rect 49133 36415 49154 36452
rect 49236 36415 49293 36461
rect 49339 36452 49396 36461
rect 49339 36415 49365 36452
rect 49442 36415 49499 36461
rect 49545 36452 49602 36461
rect 49545 36415 49576 36452
rect 49852 36415 49877 36461
rect 48905 36400 48943 36415
rect 48995 36400 49154 36415
rect 49206 36400 49365 36415
rect 49417 36400 49576 36415
rect 49628 36400 49787 36415
rect 49839 36400 49877 36415
rect 44605 36328 44812 36374
rect 44858 36328 44925 36374
rect 44971 36328 45038 36374
rect 45084 36328 45151 36374
rect 45197 36328 45264 36374
rect 45310 36328 45323 36374
rect 48905 36360 49877 36400
rect 51035 36377 51343 36417
rect 51035 36374 51073 36377
rect 51125 36374 51253 36377
rect 51305 36374 51343 36377
rect 43362 36291 43524 36298
rect 43362 36245 43373 36291
rect 43513 36245 43524 36291
rect 43362 36234 43524 36245
rect 45584 36314 48546 36350
rect 50454 36328 50467 36374
rect 50513 36328 50571 36374
rect 50617 36328 50674 36374
rect 50720 36328 50777 36374
rect 50823 36328 50880 36374
rect 50926 36328 50983 36374
rect 51029 36328 51073 36374
rect 51132 36328 51189 36374
rect 51235 36328 51253 36374
rect 51338 36328 51395 36374
rect 51441 36328 51454 36374
rect 45584 36268 45619 36314
rect 45665 36268 45777 36314
rect 45823 36268 45935 36314
rect 45981 36268 46093 36314
rect 46139 36268 46251 36314
rect 46297 36268 46409 36314
rect 46455 36268 46568 36314
rect 46614 36268 46726 36314
rect 46772 36268 46884 36314
rect 46930 36268 47042 36314
rect 47088 36268 47200 36314
rect 47246 36268 47358 36314
rect 47404 36268 47516 36314
rect 47562 36268 47675 36314
rect 47721 36268 47833 36314
rect 47879 36268 47991 36314
rect 48037 36268 48149 36314
rect 48195 36268 48307 36314
rect 48353 36268 48465 36314
rect 48511 36268 48546 36314
rect 51035 36325 51073 36328
rect 51125 36325 51253 36328
rect 51305 36325 51343 36328
rect 51035 36284 51343 36325
rect 51589 36300 51600 36722
rect 51646 36300 51657 36722
rect 54085 36723 54540 36841
rect 54085 36677 54440 36723
rect 54486 36677 54540 36723
rect 54085 36649 54540 36677
rect 53585 36598 54540 36649
rect 51789 36552 51802 36598
rect 53776 36560 54540 36598
rect 53776 36552 54440 36560
rect 53585 36530 54440 36552
rect 54085 36514 54440 36530
rect 54486 36514 54540 36560
rect 54085 36438 54540 36514
rect 51797 36384 52105 36424
rect 51797 36374 51835 36384
rect 51887 36374 52015 36384
rect 52067 36374 52105 36384
rect 54085 36392 54223 36438
rect 54269 36397 54540 36438
rect 54269 36392 54440 36397
rect 51789 36328 51802 36374
rect 53776 36328 53789 36374
rect 54085 36351 54440 36392
rect 54486 36351 54540 36397
rect 51589 36289 51657 36300
rect 51797 36291 52105 36328
rect 40215 36187 40523 36193
rect 40788 36187 42986 36201
rect 43753 36187 44514 36194
rect 39492 36164 42986 36187
rect 43704 36164 44514 36187
rect 39492 36153 44514 36164
rect 39492 36150 40253 36153
rect 39492 36104 39740 36150
rect 39786 36104 39862 36150
rect 39908 36104 39985 36150
rect 40031 36104 40108 36150
rect 40154 36104 40253 36150
rect 39492 36101 40253 36104
rect 40305 36101 40433 36153
rect 40485 36150 43790 36153
rect 40485 36104 40836 36150
rect 40882 36104 40994 36150
rect 41040 36104 41152 36150
rect 41198 36104 41310 36150
rect 41356 36104 41469 36150
rect 41515 36104 41627 36150
rect 41673 36104 41785 36150
rect 41831 36104 41943 36150
rect 41989 36104 42101 36150
rect 42147 36104 42259 36150
rect 42305 36104 42418 36150
rect 42464 36104 42576 36150
rect 42622 36104 42734 36150
rect 42780 36104 42892 36150
rect 42938 36104 43739 36150
rect 43785 36104 43790 36150
rect 40485 36101 43790 36104
rect 43842 36150 44001 36153
rect 43842 36104 43906 36150
rect 43952 36104 44001 36150
rect 43842 36101 44001 36104
rect 44053 36150 44213 36153
rect 44265 36150 44424 36153
rect 44053 36104 44071 36150
rect 44117 36104 44213 36150
rect 44282 36104 44424 36150
rect 44053 36101 44213 36104
rect 44265 36101 44424 36104
rect 44476 36101 44514 36153
rect 39492 36090 44514 36101
rect 39492 36067 42986 36090
rect 43704 36067 44514 36090
rect 37946 36060 38324 36061
rect 39014 36060 39322 36067
rect 40215 36060 40523 36067
rect 40788 36053 42986 36067
rect 43753 36061 44514 36067
rect 44796 36187 45346 36194
rect 45584 36187 48546 36268
rect 54085 36274 54540 36351
rect 54085 36228 54223 36274
rect 54269 36234 54540 36274
rect 54269 36228 54440 36234
rect 54085 36194 54440 36228
rect 48800 36187 49982 36194
rect 50308 36187 50859 36194
rect 44796 36153 49982 36187
rect 44796 36150 44834 36153
rect 44886 36150 45045 36153
rect 45097 36150 45256 36153
rect 45308 36150 48838 36153
rect 44796 36104 44812 36150
rect 44886 36104 44925 36150
rect 44971 36104 45038 36150
rect 45097 36104 45151 36150
rect 45197 36104 45256 36150
rect 45310 36104 45619 36150
rect 45665 36104 45777 36150
rect 45823 36104 45935 36150
rect 45981 36104 46093 36150
rect 46139 36104 46251 36150
rect 46297 36104 46409 36150
rect 46455 36104 46568 36150
rect 46614 36104 46726 36150
rect 46772 36104 46884 36150
rect 46930 36104 47042 36150
rect 47088 36104 47200 36150
rect 47246 36104 47358 36150
rect 47404 36104 47516 36150
rect 47562 36104 47675 36150
rect 47721 36104 47833 36150
rect 47879 36104 47991 36150
rect 48037 36104 48149 36150
rect 48195 36104 48307 36150
rect 48353 36104 48465 36150
rect 48511 36104 48838 36150
rect 44796 36101 44834 36104
rect 44886 36101 45045 36104
rect 45097 36101 45256 36104
rect 45308 36101 48838 36104
rect 48890 36101 49048 36153
rect 49100 36101 49259 36153
rect 49311 36101 49471 36153
rect 49523 36101 49682 36153
rect 49734 36101 49892 36153
rect 49944 36101 49982 36153
rect 44796 36067 49982 36101
rect 50307 36153 50859 36187
rect 50307 36101 50346 36153
rect 50398 36150 50557 36153
rect 50609 36150 50768 36153
rect 50820 36150 50859 36153
rect 52278 36188 54440 36194
rect 54486 36188 54540 36234
rect 55927 36887 56632 37001
rect 55927 36844 56267 36887
rect 55927 36798 55961 36844
rect 56007 36841 56267 36844
rect 56313 36841 56632 36887
rect 56007 36798 56632 36841
rect 55927 36723 56632 36798
rect 55927 36681 56267 36723
rect 55927 36635 55961 36681
rect 56007 36677 56267 36681
rect 56313 36677 56632 36723
rect 56007 36635 56632 36677
rect 55927 36560 56632 36635
rect 55927 36517 56267 36560
rect 55927 36471 55961 36517
rect 56007 36514 56267 36517
rect 56313 36514 56632 36560
rect 56007 36471 56632 36514
rect 55927 36397 56632 36471
rect 55927 36354 56267 36397
rect 55927 36308 55961 36354
rect 56007 36351 56267 36354
rect 56313 36351 56632 36397
rect 56007 36308 56632 36351
rect 55927 36234 56632 36308
rect 52278 36153 54540 36188
rect 52278 36150 52316 36153
rect 52368 36150 52527 36153
rect 52579 36150 52738 36153
rect 52790 36150 52948 36153
rect 53000 36150 53159 36153
rect 53211 36150 53371 36153
rect 53423 36150 53582 36153
rect 53634 36150 53792 36153
rect 50398 36104 50467 36150
rect 50513 36104 50557 36150
rect 50617 36104 50674 36150
rect 50720 36104 50768 36150
rect 50823 36104 50880 36150
rect 50926 36104 50983 36150
rect 51029 36104 51086 36150
rect 51132 36104 51189 36150
rect 51235 36104 51292 36150
rect 51338 36104 51395 36150
rect 51441 36104 51454 36150
rect 51789 36104 51802 36150
rect 53776 36104 53792 36150
rect 50398 36101 50557 36104
rect 50609 36101 50768 36104
rect 50820 36101 50859 36104
rect 50307 36067 50859 36101
rect 44796 36061 45346 36067
rect 48800 36060 49982 36067
rect 50308 36060 50859 36067
rect 52278 36101 52316 36104
rect 52368 36101 52527 36104
rect 52579 36101 52738 36104
rect 52790 36101 52948 36104
rect 53000 36101 53159 36104
rect 53211 36101 53371 36104
rect 53423 36101 53582 36104
rect 53634 36101 53792 36104
rect 53844 36101 54003 36153
rect 54055 36101 54214 36153
rect 54266 36101 54540 36153
rect 52278 36061 54540 36101
rect 54758 36153 55840 36194
rect 54758 36150 54855 36153
rect 54758 36104 54793 36150
rect 54839 36104 54855 36150
rect 54758 36101 54855 36104
rect 54907 36150 55066 36153
rect 54907 36104 54956 36150
rect 55002 36104 55066 36150
rect 54907 36101 55066 36104
rect 55118 36150 55278 36153
rect 55330 36150 55489 36153
rect 55164 36104 55278 36150
rect 55330 36104 55439 36150
rect 55485 36104 55489 36150
rect 55118 36101 55278 36104
rect 55330 36101 55489 36104
rect 55541 36150 55840 36153
rect 55541 36104 55599 36150
rect 55645 36104 55760 36150
rect 55806 36104 55840 36150
rect 55541 36101 55840 36104
rect 54758 36061 55840 36101
rect 55927 36188 56267 36234
rect 56313 36188 56632 36234
rect 52278 36060 54377 36061
rect 54817 36060 55579 36061
rect 55927 36027 56632 36188
rect 28492 35996 28891 36027
rect 27744 35985 28891 35996
rect 56621 35996 56632 36027
rect 57278 35996 57380 37001
rect 27744 34938 27828 35985
rect 56621 35977 57380 35996
rect 27387 34909 27449 34938
rect 24369 34886 27449 34909
rect 27749 34886 27828 34938
rect 24369 34848 27498 34886
rect 24369 34796 25400 34848
rect 25452 34796 25524 34848
rect 25576 34796 25648 34848
rect 25700 34796 25772 34848
rect 25824 34796 25896 34848
rect 25948 34814 27498 34848
rect 27744 34814 27828 34886
rect 25948 34796 27449 34814
rect 24369 34762 27449 34796
rect 27749 34762 27828 34814
rect 24369 34739 27498 34762
rect 25388 34724 25960 34739
rect 25388 34672 25400 34724
rect 25452 34672 25524 34724
rect 25576 34672 25648 34724
rect 25700 34672 25772 34724
rect 25824 34672 25896 34724
rect 25948 34672 25960 34724
rect 25388 34660 25960 34672
rect 27387 34690 27498 34739
rect 27744 34690 27828 34762
rect 27387 34638 27449 34690
rect 27749 34638 27828 34690
rect 27387 34566 27498 34638
rect 27744 34613 27828 34638
rect 57295 34613 57380 35977
rect 27744 34602 57380 34613
rect 27744 34566 27846 34602
rect 27387 34514 27449 34566
rect 27749 34514 27846 34566
rect 26772 33432 27214 33519
rect 26772 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27214 33432
rect 26772 33215 27214 33380
rect 26772 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27214 33215
rect 26772 32997 27214 33163
rect 26772 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27214 32997
rect 26772 32779 27214 32945
rect 26772 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27214 32779
rect 26772 32562 27214 32727
rect 26772 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27214 32562
rect 26772 32344 27214 32510
rect 26772 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27214 32344
rect 26772 32127 27214 32292
rect 26772 32075 26861 32127
rect 26913 32075 27073 32127
rect 27125 32075 27214 32127
rect 26772 31909 27214 32075
rect 26772 31857 26861 31909
rect 26913 31857 27073 31909
rect 27125 31857 27214 31909
rect 26772 31691 27214 31857
rect 26772 31639 26861 31691
rect 26913 31639 27073 31691
rect 27125 31639 27214 31691
rect 26772 31474 27214 31639
rect 26772 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27214 31474
rect 26772 31256 27214 31422
rect 26772 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27214 31256
rect 26772 31038 27214 31204
rect 26772 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27214 31038
rect 26772 30821 27214 30986
rect 26772 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27214 30821
rect 26772 30603 27214 30769
rect 26772 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27214 30603
rect 26772 30386 27214 30551
rect 26772 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27214 30386
rect 26772 30168 27214 30334
rect 26772 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27214 30168
rect 26772 29950 27214 30116
rect 26772 29898 26861 29950
rect 26913 29898 27073 29950
rect 27125 29898 27214 29950
rect 26772 29733 27214 29898
rect 26772 29681 26861 29733
rect 26913 29681 27073 29733
rect 27125 29681 27214 29733
rect 26772 29515 27214 29681
rect 26772 29463 26861 29515
rect 26913 29463 27073 29515
rect 27125 29463 27214 29515
rect 26772 29297 27214 29463
rect 26772 29245 26861 29297
rect 26913 29245 27073 29297
rect 27125 29245 27214 29297
rect 26772 29080 27214 29245
rect 26772 29028 26861 29080
rect 26913 29028 27073 29080
rect 27125 29028 27214 29080
rect 26772 28862 27214 29028
rect 26772 28810 26861 28862
rect 26913 28810 27073 28862
rect 27125 28810 27214 28862
rect 26772 28644 27214 28810
rect 26772 28592 26861 28644
rect 26913 28592 27073 28644
rect 27125 28592 27214 28644
rect 26772 28427 27214 28592
rect 26772 28375 26861 28427
rect 26913 28375 27073 28427
rect 27125 28375 27214 28427
rect 26772 28209 27214 28375
rect 26772 28157 26861 28209
rect 26913 28157 27073 28209
rect 27125 28157 27214 28209
rect 26772 27992 27214 28157
rect 26772 27940 26861 27992
rect 26913 27940 27073 27992
rect 27125 27940 27214 27992
rect 26772 27774 27214 27940
rect 26772 27722 26861 27774
rect 26913 27722 27073 27774
rect 27125 27722 27214 27774
rect 26772 27556 27214 27722
rect 26772 27504 26861 27556
rect 26913 27504 27073 27556
rect 27125 27504 27214 27556
rect 26772 27339 27214 27504
rect 26772 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27214 27339
rect 26772 27121 27214 27287
rect 26772 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27214 27121
rect 26772 26903 27214 27069
rect 26772 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27214 26903
rect 26772 26686 27214 26851
rect 26772 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27214 26686
rect 26772 26468 27214 26634
rect 26772 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27214 26468
rect 26772 26250 27214 26416
rect 26772 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27214 26250
rect 26772 26033 27214 26198
rect 26772 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27214 26033
rect 26772 25815 27214 25981
rect 26772 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27214 25815
rect 26772 25598 27214 25763
rect 26772 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27214 25598
rect 26772 25380 27214 25546
rect 26772 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27214 25380
rect 26772 25162 27214 25328
rect 26772 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27214 25162
rect 26772 24945 27214 25110
rect 26772 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27214 24945
rect 26772 24727 27214 24893
rect 26772 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27214 24727
rect 26772 24509 27214 24675
rect 26772 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27214 24509
rect 26772 24292 27214 24457
rect 26772 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27214 24292
rect 26772 24074 27214 24240
rect 26772 24022 26861 24074
rect 26913 24022 27073 24074
rect 27125 24022 27214 24074
rect 26772 23857 27214 24022
rect 26772 23805 26861 23857
rect 26913 23805 27073 23857
rect 27125 23805 27214 23857
rect 26772 23639 27214 23805
rect 26772 23587 26861 23639
rect 26913 23587 27073 23639
rect 27125 23587 27214 23639
rect 26772 23421 27214 23587
rect 26772 23369 26861 23421
rect 26913 23369 27073 23421
rect 27125 23369 27214 23421
rect 26772 23204 27214 23369
rect 26772 23152 26861 23204
rect 26913 23152 27073 23204
rect 27125 23152 27214 23204
rect 26772 22986 27214 23152
rect 26772 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27214 22986
rect 26772 22768 27214 22934
rect 26772 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27214 22768
rect 26772 22551 27214 22716
rect 26772 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27214 22551
rect 26772 22333 27214 22499
rect 26772 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27214 22333
rect 26772 22115 27214 22281
rect 26772 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27214 22115
rect 26772 21898 27214 22063
rect 26772 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27214 21898
rect 26772 21680 27214 21846
rect 26772 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27214 21680
rect 26772 21463 27214 21628
rect 26772 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27214 21463
rect 26772 21245 27214 21411
rect 26772 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27214 21245
rect 26772 21027 27214 21193
rect 26772 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27214 21027
rect 26772 20810 27214 20975
rect 26772 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27214 20810
rect 26772 20592 27214 20758
rect 26772 20540 26861 20592
rect 26913 20540 27073 20592
rect 27125 20540 27214 20592
rect 26772 20374 27214 20540
rect 26772 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27214 20374
rect 26772 20157 27214 20322
rect 26772 20105 26861 20157
rect 26913 20105 27073 20157
rect 27125 20105 27214 20157
rect 26772 19939 27214 20105
rect 26772 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27214 19939
rect 26772 19722 27214 19887
rect 26772 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27214 19722
rect 26772 19504 27214 19670
rect 26772 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27214 19504
rect 26772 19286 27214 19452
rect 26772 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27214 19286
rect 26772 19068 27214 19234
rect 26772 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27214 19068
rect 26772 18851 27214 19016
rect 26772 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27214 18851
rect 26772 18633 27214 18799
rect 26772 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27214 18633
rect 26772 18416 27214 18581
rect 26772 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27214 18416
rect 26772 18198 27214 18364
rect 26772 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27214 18198
rect 26772 17980 27214 18146
rect 26772 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27214 17980
rect 26772 17763 27214 17928
rect 26772 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27214 17763
rect 26772 17545 27214 17711
rect 26772 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27214 17545
rect 26772 17327 27214 17493
rect 26772 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27214 17327
rect 26772 17110 27214 17275
rect 26772 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27214 17110
rect 26772 16892 27214 17058
rect 26772 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27214 16892
rect 26772 16675 27214 16840
rect 26772 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27214 16675
rect 26772 16457 27214 16623
rect 26772 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27214 16457
rect 26772 16239 27214 16405
rect 26772 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27214 16239
rect 26772 16022 27214 16187
rect 26772 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27214 16022
rect 26772 15804 27214 15970
rect 26772 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27214 15804
rect 26772 15586 27214 15752
rect 26772 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27214 15586
rect 26772 15369 27214 15534
rect 26772 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27214 15369
rect 26772 15151 27214 15317
rect 26772 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27214 15151
rect 26772 14933 27214 15099
rect 26772 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27214 14933
rect 26772 14716 27214 14881
rect 26772 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27214 14716
rect 26772 14498 27214 14664
rect 26772 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27214 14498
rect 26772 14281 27214 14446
rect 26772 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27214 14281
rect 26772 14063 27214 14229
rect 26772 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27214 14063
rect 26772 13845 27214 14011
rect 26772 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27214 13845
rect 26772 13628 27214 13793
rect 26772 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27214 13628
rect 26772 13410 27214 13576
rect 26772 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27214 13410
rect 26772 13192 27214 13358
rect 26772 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27214 13192
rect 26772 12975 27214 13140
rect 26772 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27214 12975
rect 26772 12757 27214 12923
rect 26772 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27214 12757
rect 26772 12540 27214 12705
rect 26772 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27214 12540
rect 26772 12322 27214 12488
rect 26772 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27214 12322
rect 26772 12104 27214 12270
rect 26772 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27214 12104
rect 26772 11887 27214 12052
rect 26772 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27214 11887
rect 26772 11669 27214 11835
rect 26772 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27214 11669
rect 26772 11451 27214 11617
rect 26772 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27214 11451
rect 26772 11234 27214 11399
rect 26772 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27214 11234
rect 26772 11016 27214 11182
rect 26772 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27214 11016
rect 26772 10798 27214 10964
rect 26772 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27214 10798
rect 26772 10581 27214 10746
rect 26772 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27214 10581
rect 26772 10363 27214 10529
rect 26772 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27214 10363
rect 26772 10146 27214 10311
rect 26772 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27214 10146
rect 26772 9928 27214 10094
rect 26772 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27214 9928
rect 26772 9710 27214 9876
rect 26772 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27214 9710
rect 26772 9493 27214 9658
rect 26772 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27214 9493
rect 26772 9275 27214 9441
rect 26772 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27214 9275
rect 26772 9057 27214 9223
rect 26772 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27214 9057
rect 26772 8840 27214 9005
rect 26772 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27214 8840
rect 26772 8622 27214 8788
rect 26772 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27214 8622
rect 26772 8404 27214 8570
rect 26772 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27214 8404
rect 26772 8187 27214 8352
rect 26772 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27214 8187
rect 26772 7969 27214 8135
rect 26772 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27214 7969
rect 26772 7752 27214 7917
rect 26772 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27214 7752
rect 26772 7534 27214 7700
rect 26772 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27214 7534
rect 26772 7316 27214 7482
rect 26772 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27214 7316
rect 26772 7099 27214 7264
rect 26772 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27214 7099
rect 26772 6881 27214 7047
rect 26772 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27214 6881
rect 26772 6663 27214 6829
rect 26772 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27214 6663
rect 26772 6446 27214 6611
rect 26772 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27214 6446
rect 26772 6228 27214 6394
rect 26772 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27214 6228
rect 26772 6011 27214 6176
rect 26772 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27214 6011
rect 26772 5793 27214 5959
rect 26772 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27214 5793
rect 26772 5575 27214 5741
rect 26772 5523 26861 5575
rect 26913 5523 27073 5575
rect 27125 5523 27214 5575
rect 26772 5358 27214 5523
rect 26772 5306 26861 5358
rect 26913 5306 27073 5358
rect 27125 5306 27214 5358
rect 26772 4587 27214 5306
rect 26772 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27214 4587
rect 26772 4370 27214 4535
rect 26772 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27214 4370
rect 26772 4152 27214 4318
rect 26772 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27214 4152
rect 26772 3934 27214 4100
rect 26772 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27214 3934
rect 26772 3717 27214 3882
rect 26772 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27214 3717
rect 26772 1777 27214 3665
rect 27387 33432 27498 34514
rect 27744 34256 27846 34514
rect 57292 34256 57380 34602
rect 27744 34245 57380 34256
rect 27387 33380 27476 33432
rect 27387 33215 27498 33380
rect 27387 33163 27476 33215
rect 27387 32997 27498 33163
rect 27387 32945 27476 32997
rect 27387 32779 27498 32945
rect 27387 32727 27476 32779
rect 27387 32562 27498 32727
rect 27387 32510 27476 32562
rect 27387 32344 27498 32510
rect 27387 32292 27476 32344
rect 27387 32127 27498 32292
rect 27387 32075 27476 32127
rect 27387 31909 27498 32075
rect 27387 31857 27476 31909
rect 27387 31691 27498 31857
rect 27387 31639 27476 31691
rect 27387 31474 27498 31639
rect 27387 31422 27476 31474
rect 27387 31256 27498 31422
rect 27387 31204 27476 31256
rect 27387 31038 27498 31204
rect 27387 30986 27476 31038
rect 27387 30821 27498 30986
rect 27387 30769 27476 30821
rect 27387 30603 27498 30769
rect 27387 30551 27476 30603
rect 27387 30386 27498 30551
rect 27387 30334 27476 30386
rect 27387 30168 27498 30334
rect 27387 30116 27476 30168
rect 27387 29950 27498 30116
rect 27387 29898 27476 29950
rect 27387 29733 27498 29898
rect 27387 29681 27476 29733
rect 27387 29515 27498 29681
rect 27387 29463 27476 29515
rect 27387 29297 27498 29463
rect 27387 29245 27476 29297
rect 27387 29080 27498 29245
rect 27387 29028 27476 29080
rect 27387 28862 27498 29028
rect 27387 28810 27476 28862
rect 27387 28644 27498 28810
rect 27387 28592 27476 28644
rect 27387 28427 27498 28592
rect 27387 28375 27476 28427
rect 27387 28209 27498 28375
rect 27387 28157 27476 28209
rect 27387 27992 27498 28157
rect 27387 27940 27476 27992
rect 27387 27774 27498 27940
rect 27387 27722 27476 27774
rect 27387 27556 27498 27722
rect 27387 27504 27476 27556
rect 27387 27339 27498 27504
rect 27387 27287 27476 27339
rect 27387 27121 27498 27287
rect 27387 27069 27476 27121
rect 27387 26903 27498 27069
rect 27387 26851 27476 26903
rect 27387 26686 27498 26851
rect 27387 26634 27476 26686
rect 27387 26468 27498 26634
rect 27387 26416 27476 26468
rect 27387 26250 27498 26416
rect 27387 26198 27476 26250
rect 27387 26033 27498 26198
rect 27387 25981 27476 26033
rect 27387 25815 27498 25981
rect 27387 25763 27476 25815
rect 27387 25598 27498 25763
rect 27387 25546 27476 25598
rect 27387 25380 27498 25546
rect 27387 25328 27476 25380
rect 27387 25162 27498 25328
rect 27387 25110 27476 25162
rect 27387 24945 27498 25110
rect 27387 24893 27476 24945
rect 27387 24727 27498 24893
rect 27387 24675 27476 24727
rect 27387 24509 27498 24675
rect 27387 24457 27476 24509
rect 27387 24292 27498 24457
rect 27387 24240 27476 24292
rect 27387 24074 27498 24240
rect 27387 24022 27476 24074
rect 27387 23857 27498 24022
rect 27387 23805 27476 23857
rect 27387 23639 27498 23805
rect 27387 23587 27476 23639
rect 27387 23421 27498 23587
rect 27387 23369 27476 23421
rect 27387 23204 27498 23369
rect 27387 23152 27476 23204
rect 27387 22986 27498 23152
rect 27387 22934 27476 22986
rect 27387 22768 27498 22934
rect 27387 22716 27476 22768
rect 27387 22551 27498 22716
rect 27387 22499 27476 22551
rect 27387 22333 27498 22499
rect 27387 22281 27476 22333
rect 27387 22115 27498 22281
rect 27387 22063 27476 22115
rect 27387 21898 27498 22063
rect 27387 21846 27476 21898
rect 27387 21680 27498 21846
rect 27387 21628 27476 21680
rect 27387 21463 27498 21628
rect 27387 21411 27476 21463
rect 27387 21245 27498 21411
rect 27387 21193 27476 21245
rect 27387 21027 27498 21193
rect 27387 20975 27476 21027
rect 27387 20810 27498 20975
rect 27387 20758 27476 20810
rect 27387 20592 27498 20758
rect 27387 20540 27476 20592
rect 27387 20374 27498 20540
rect 27387 20322 27476 20374
rect 27387 20157 27498 20322
rect 27387 20105 27476 20157
rect 27387 19939 27498 20105
rect 27387 19887 27476 19939
rect 27387 19722 27498 19887
rect 27387 19670 27476 19722
rect 27387 19504 27498 19670
rect 27387 19452 27476 19504
rect 27387 19286 27498 19452
rect 27387 19234 27476 19286
rect 27387 19068 27498 19234
rect 27387 19016 27476 19068
rect 27387 18851 27498 19016
rect 27387 18799 27476 18851
rect 27387 18633 27498 18799
rect 27387 18581 27476 18633
rect 27387 18416 27498 18581
rect 27387 18364 27476 18416
rect 27387 18198 27498 18364
rect 27387 18146 27476 18198
rect 27387 17980 27498 18146
rect 27387 17928 27476 17980
rect 27387 17763 27498 17928
rect 27387 17711 27476 17763
rect 27387 17545 27498 17711
rect 27387 17493 27476 17545
rect 27387 17327 27498 17493
rect 27387 17275 27476 17327
rect 27387 17110 27498 17275
rect 27387 17058 27476 17110
rect 27387 16892 27498 17058
rect 27387 16840 27476 16892
rect 27387 16675 27498 16840
rect 27387 16623 27476 16675
rect 27387 16457 27498 16623
rect 27387 16405 27476 16457
rect 27387 16239 27498 16405
rect 27387 16187 27476 16239
rect 27387 16022 27498 16187
rect 27387 15970 27476 16022
rect 27387 15804 27498 15970
rect 27387 15752 27476 15804
rect 27387 15586 27498 15752
rect 27387 15534 27476 15586
rect 27387 15369 27498 15534
rect 27387 15317 27476 15369
rect 27387 15151 27498 15317
rect 27387 15099 27476 15151
rect 27387 14933 27498 15099
rect 27387 14881 27476 14933
rect 27387 14716 27498 14881
rect 27387 14664 27476 14716
rect 27387 14498 27498 14664
rect 27387 14446 27476 14498
rect 27387 14281 27498 14446
rect 27387 14229 27476 14281
rect 27387 14063 27498 14229
rect 27387 14011 27476 14063
rect 27387 13845 27498 14011
rect 27387 13793 27476 13845
rect 27387 13628 27498 13793
rect 27387 13576 27476 13628
rect 27387 13410 27498 13576
rect 27387 13358 27476 13410
rect 27387 13192 27498 13358
rect 27387 13140 27476 13192
rect 27387 12975 27498 13140
rect 27387 12923 27476 12975
rect 27387 12757 27498 12923
rect 27387 12705 27476 12757
rect 27387 12540 27498 12705
rect 27387 12488 27476 12540
rect 27387 12322 27498 12488
rect 27387 12270 27476 12322
rect 27387 12104 27498 12270
rect 27387 12052 27476 12104
rect 27387 11887 27498 12052
rect 27387 11835 27476 11887
rect 27387 11669 27498 11835
rect 27387 11617 27476 11669
rect 27387 11451 27498 11617
rect 27387 11399 27476 11451
rect 27387 11234 27498 11399
rect 27387 11182 27476 11234
rect 27387 11016 27498 11182
rect 27387 10964 27476 11016
rect 27387 10798 27498 10964
rect 27387 10746 27476 10798
rect 27387 10581 27498 10746
rect 27387 10529 27476 10581
rect 27387 10363 27498 10529
rect 27387 10311 27476 10363
rect 27387 10146 27498 10311
rect 27387 10094 27476 10146
rect 27387 9928 27498 10094
rect 27387 9876 27476 9928
rect 27387 9710 27498 9876
rect 27387 9658 27476 9710
rect 27387 9493 27498 9658
rect 27387 9441 27476 9493
rect 27387 9275 27498 9441
rect 27387 9223 27476 9275
rect 27387 9057 27498 9223
rect 27387 9005 27476 9057
rect 27387 8840 27498 9005
rect 27387 8788 27476 8840
rect 27387 8622 27498 8788
rect 27387 8570 27476 8622
rect 27387 8404 27498 8570
rect 27387 8352 27476 8404
rect 27387 8187 27498 8352
rect 27387 8135 27476 8187
rect 27387 7969 27498 8135
rect 27387 7917 27476 7969
rect 27387 7752 27498 7917
rect 27387 7700 27476 7752
rect 27387 7534 27498 7700
rect 27387 7482 27476 7534
rect 27387 7316 27498 7482
rect 27387 7264 27476 7316
rect 27387 7099 27498 7264
rect 27387 7047 27476 7099
rect 27387 6881 27498 7047
rect 27387 6829 27476 6881
rect 27387 6663 27498 6829
rect 27387 6611 27476 6663
rect 27387 6446 27498 6611
rect 27387 6394 27476 6446
rect 27387 6228 27498 6394
rect 27387 6176 27476 6228
rect 27387 6011 27498 6176
rect 27387 5959 27476 6011
rect 27387 5793 27498 5959
rect 27387 5741 27476 5793
rect 27387 5575 27498 5741
rect 27387 5523 27476 5575
rect 27387 5358 27498 5523
rect 27387 5306 27476 5358
rect 27387 4587 27498 5306
rect 27387 4535 27476 4587
rect 27387 4370 27498 4535
rect 27387 4318 27476 4370
rect 27387 4152 27498 4318
rect 27387 4100 27476 4152
rect 27387 3934 27498 4100
rect 27387 3882 27476 3934
rect 27387 3717 27498 3882
rect 27387 3665 27476 3717
rect 2562 1689 2742 1701
rect 2562 1637 2574 1689
rect 2730 1637 2742 1689
rect 2562 1625 2742 1637
rect 12627 1689 12807 1701
rect 12627 1637 12639 1689
rect 12795 1637 12807 1689
rect 12627 1625 12807 1637
rect 13077 1689 13257 1701
rect 13077 1637 13089 1689
rect 13245 1637 13257 1689
rect 13077 1625 13257 1637
rect 23427 1689 23607 1701
rect 23427 1637 23439 1689
rect 23595 1637 23607 1689
rect 23427 1625 23607 1637
rect 27387 1282 27498 3665
rect 717 1117 27498 1282
rect 27744 1925 27828 34245
rect 49896 6349 50076 6361
rect 49896 6347 49908 6349
rect 49728 6301 49908 6347
rect 49896 6297 49908 6301
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 51642 5199 51822 5211
rect 51642 5196 51654 5199
rect 49963 5150 51654 5196
rect 51642 5147 51654 5150
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 50834 3890 56586 3901
rect 28628 3869 40180 3880
rect 28628 3823 28639 3869
rect 28685 3823 28755 3869
rect 28801 3823 28871 3869
rect 28917 3823 28987 3869
rect 29033 3823 29103 3869
rect 29149 3823 29219 3869
rect 29265 3823 29335 3869
rect 29381 3823 29451 3869
rect 29497 3823 29567 3869
rect 29613 3823 29683 3869
rect 29729 3823 29799 3869
rect 29845 3823 29915 3869
rect 29961 3823 30031 3869
rect 30077 3823 30147 3869
rect 30193 3823 30263 3869
rect 30309 3823 30379 3869
rect 30425 3823 30495 3869
rect 30541 3823 30611 3869
rect 30657 3823 30727 3869
rect 30773 3823 30843 3869
rect 30889 3823 30959 3869
rect 31005 3823 31075 3869
rect 31121 3823 31191 3869
rect 31237 3823 31307 3869
rect 31353 3823 31423 3869
rect 31469 3823 31539 3869
rect 31585 3823 31655 3869
rect 31701 3823 31771 3869
rect 31817 3823 31887 3869
rect 31933 3823 32003 3869
rect 32049 3823 32119 3869
rect 32165 3823 32235 3869
rect 32281 3823 32351 3869
rect 32397 3823 32467 3869
rect 32513 3823 32583 3869
rect 32629 3823 32699 3869
rect 32745 3823 32815 3869
rect 32861 3823 32931 3869
rect 32977 3823 33047 3869
rect 33093 3823 33163 3869
rect 33209 3823 33279 3869
rect 33325 3823 33395 3869
rect 33441 3823 33511 3869
rect 33557 3823 33627 3869
rect 33673 3823 33743 3869
rect 33789 3823 33859 3869
rect 33905 3823 33975 3869
rect 34021 3823 34091 3869
rect 34137 3823 34207 3869
rect 34253 3823 34323 3869
rect 34369 3823 34439 3869
rect 34485 3823 34555 3869
rect 34601 3823 34671 3869
rect 34717 3823 34787 3869
rect 34833 3823 34903 3869
rect 34949 3823 35019 3869
rect 35065 3823 35135 3869
rect 35181 3823 35251 3869
rect 35297 3823 35367 3869
rect 35413 3823 35483 3869
rect 35529 3823 35599 3869
rect 35645 3823 35715 3869
rect 35761 3823 35831 3869
rect 35877 3823 35947 3869
rect 35993 3823 36063 3869
rect 36109 3823 36179 3869
rect 36225 3823 36295 3869
rect 36341 3823 36411 3869
rect 36457 3823 36527 3869
rect 36573 3823 36643 3869
rect 36689 3823 36759 3869
rect 36805 3823 36875 3869
rect 36921 3823 36991 3869
rect 37037 3823 37107 3869
rect 37153 3823 37223 3869
rect 37269 3823 37339 3869
rect 37385 3823 37455 3869
rect 37501 3823 37571 3869
rect 37617 3823 37687 3869
rect 37733 3823 37803 3869
rect 37849 3823 37919 3869
rect 37965 3823 38035 3869
rect 38081 3823 38151 3869
rect 38197 3823 38267 3869
rect 38313 3823 38383 3869
rect 38429 3823 38499 3869
rect 38545 3823 38615 3869
rect 38661 3823 38731 3869
rect 38777 3823 38847 3869
rect 38893 3823 38963 3869
rect 39009 3823 39079 3869
rect 39125 3823 39195 3869
rect 39241 3823 39311 3869
rect 39357 3823 39427 3869
rect 39473 3823 39543 3869
rect 39589 3823 39659 3869
rect 39705 3823 39775 3869
rect 39821 3823 39891 3869
rect 39937 3823 40007 3869
rect 40053 3823 40123 3869
rect 40169 3823 40180 3869
rect 28628 3753 40180 3823
rect 28628 3707 28639 3753
rect 28685 3707 28755 3753
rect 28801 3707 28871 3753
rect 28917 3707 28987 3753
rect 29033 3707 29103 3753
rect 29149 3707 29219 3753
rect 29265 3707 29335 3753
rect 29381 3707 29451 3753
rect 29497 3707 29567 3753
rect 29613 3707 29683 3753
rect 29729 3707 29799 3753
rect 29845 3707 29915 3753
rect 29961 3707 30031 3753
rect 30077 3707 30147 3753
rect 30193 3707 30263 3753
rect 30309 3707 30379 3753
rect 30425 3707 30495 3753
rect 30541 3707 30611 3753
rect 30657 3707 30727 3753
rect 30773 3707 30843 3753
rect 30889 3707 30959 3753
rect 31005 3707 31075 3753
rect 31121 3707 31191 3753
rect 31237 3707 31307 3753
rect 31353 3707 31423 3753
rect 31469 3707 31539 3753
rect 31585 3707 31655 3753
rect 31701 3707 31771 3753
rect 31817 3707 31887 3753
rect 31933 3707 32003 3753
rect 32049 3707 32119 3753
rect 32165 3707 32235 3753
rect 32281 3707 32351 3753
rect 32397 3707 32467 3753
rect 32513 3707 32583 3753
rect 32629 3707 32699 3753
rect 32745 3707 32815 3753
rect 32861 3707 32931 3753
rect 32977 3707 33047 3753
rect 33093 3707 33163 3753
rect 33209 3707 33279 3753
rect 33325 3707 33395 3753
rect 33441 3707 33511 3753
rect 33557 3707 33627 3753
rect 33673 3707 33743 3753
rect 33789 3707 33859 3753
rect 33905 3707 33975 3753
rect 34021 3707 34091 3753
rect 34137 3707 34207 3753
rect 34253 3707 34323 3753
rect 34369 3707 34439 3753
rect 34485 3707 34555 3753
rect 34601 3707 34671 3753
rect 34717 3707 34787 3753
rect 34833 3707 34903 3753
rect 34949 3707 35019 3753
rect 35065 3707 35135 3753
rect 35181 3707 35251 3753
rect 35297 3707 35367 3753
rect 35413 3707 35483 3753
rect 35529 3707 35599 3753
rect 35645 3707 35715 3753
rect 35761 3707 35831 3753
rect 35877 3707 35947 3753
rect 35993 3707 36063 3753
rect 36109 3707 36179 3753
rect 36225 3707 36295 3753
rect 36341 3707 36411 3753
rect 36457 3707 36527 3753
rect 36573 3707 36643 3753
rect 36689 3707 36759 3753
rect 36805 3707 36875 3753
rect 36921 3707 36991 3753
rect 37037 3707 37107 3753
rect 37153 3707 37223 3753
rect 37269 3707 37339 3753
rect 37385 3707 37455 3753
rect 37501 3707 37571 3753
rect 37617 3707 37687 3753
rect 37733 3707 37803 3753
rect 37849 3707 37919 3753
rect 37965 3707 38035 3753
rect 38081 3707 38151 3753
rect 38197 3707 38267 3753
rect 38313 3707 38383 3753
rect 38429 3707 38499 3753
rect 38545 3707 38615 3753
rect 38661 3707 38731 3753
rect 38777 3707 38847 3753
rect 38893 3707 38963 3753
rect 39009 3707 39079 3753
rect 39125 3707 39195 3753
rect 39241 3707 39311 3753
rect 39357 3707 39427 3753
rect 39473 3707 39543 3753
rect 39589 3707 39659 3753
rect 39705 3707 39775 3753
rect 39821 3707 39891 3753
rect 39937 3707 40007 3753
rect 40053 3707 40123 3753
rect 40169 3707 40180 3753
rect 28628 3637 40180 3707
rect 28628 3591 28639 3637
rect 28685 3591 28755 3637
rect 28801 3591 28871 3637
rect 28917 3591 28987 3637
rect 29033 3591 29103 3637
rect 29149 3591 29219 3637
rect 29265 3591 29335 3637
rect 29381 3591 29451 3637
rect 29497 3591 29567 3637
rect 29613 3591 29683 3637
rect 29729 3591 29799 3637
rect 29845 3591 29915 3637
rect 29961 3591 30031 3637
rect 30077 3591 30147 3637
rect 30193 3591 30263 3637
rect 30309 3591 30379 3637
rect 30425 3591 30495 3637
rect 30541 3591 30611 3637
rect 30657 3591 30727 3637
rect 30773 3591 30843 3637
rect 30889 3591 30959 3637
rect 31005 3591 31075 3637
rect 31121 3591 31191 3637
rect 31237 3591 31307 3637
rect 31353 3591 31423 3637
rect 31469 3591 31539 3637
rect 31585 3591 31655 3637
rect 31701 3591 31771 3637
rect 31817 3591 31887 3637
rect 31933 3591 32003 3637
rect 32049 3591 32119 3637
rect 32165 3591 32235 3637
rect 32281 3591 32351 3637
rect 32397 3591 32467 3637
rect 32513 3591 32583 3637
rect 32629 3591 32699 3637
rect 32745 3591 32815 3637
rect 32861 3591 32931 3637
rect 32977 3591 33047 3637
rect 33093 3591 33163 3637
rect 33209 3591 33279 3637
rect 33325 3591 33395 3637
rect 33441 3591 33511 3637
rect 33557 3591 33627 3637
rect 33673 3591 33743 3637
rect 33789 3591 33859 3637
rect 33905 3591 33975 3637
rect 34021 3591 34091 3637
rect 34137 3591 34207 3637
rect 34253 3591 34323 3637
rect 34369 3591 34439 3637
rect 34485 3591 34555 3637
rect 34601 3591 34671 3637
rect 34717 3591 34787 3637
rect 34833 3591 34903 3637
rect 34949 3591 35019 3637
rect 35065 3591 35135 3637
rect 35181 3591 35251 3637
rect 35297 3591 35367 3637
rect 35413 3591 35483 3637
rect 35529 3591 35599 3637
rect 35645 3591 35715 3637
rect 35761 3591 35831 3637
rect 35877 3591 35947 3637
rect 35993 3591 36063 3637
rect 36109 3591 36179 3637
rect 36225 3591 36295 3637
rect 36341 3591 36411 3637
rect 36457 3591 36527 3637
rect 36573 3591 36643 3637
rect 36689 3591 36759 3637
rect 36805 3591 36875 3637
rect 36921 3591 36991 3637
rect 37037 3591 37107 3637
rect 37153 3591 37223 3637
rect 37269 3591 37339 3637
rect 37385 3591 37455 3637
rect 37501 3591 37571 3637
rect 37617 3591 37687 3637
rect 37733 3591 37803 3637
rect 37849 3591 37919 3637
rect 37965 3591 38035 3637
rect 38081 3591 38151 3637
rect 38197 3591 38267 3637
rect 38313 3591 38383 3637
rect 38429 3591 38499 3637
rect 38545 3591 38615 3637
rect 38661 3591 38731 3637
rect 38777 3591 38847 3637
rect 38893 3591 38963 3637
rect 39009 3591 39079 3637
rect 39125 3591 39195 3637
rect 39241 3591 39311 3637
rect 39357 3591 39427 3637
rect 39473 3591 39543 3637
rect 39589 3591 39659 3637
rect 39705 3591 39775 3637
rect 39821 3591 39891 3637
rect 39937 3591 40007 3637
rect 40053 3591 40123 3637
rect 40169 3591 40180 3637
rect 28628 3521 40180 3591
rect 28628 3475 28639 3521
rect 28685 3475 28755 3521
rect 28801 3475 28871 3521
rect 28917 3475 28987 3521
rect 29033 3475 29103 3521
rect 29149 3475 29219 3521
rect 29265 3475 29335 3521
rect 29381 3475 29451 3521
rect 29497 3475 29567 3521
rect 29613 3475 29683 3521
rect 29729 3475 29799 3521
rect 29845 3475 29915 3521
rect 29961 3475 30031 3521
rect 30077 3475 30147 3521
rect 30193 3475 30263 3521
rect 30309 3475 30379 3521
rect 30425 3475 30495 3521
rect 30541 3475 30611 3521
rect 30657 3475 30727 3521
rect 30773 3475 30843 3521
rect 30889 3475 30959 3521
rect 31005 3475 31075 3521
rect 31121 3475 31191 3521
rect 31237 3475 31307 3521
rect 31353 3475 31423 3521
rect 31469 3475 31539 3521
rect 31585 3475 31655 3521
rect 31701 3475 31771 3521
rect 31817 3475 31887 3521
rect 31933 3475 32003 3521
rect 32049 3475 32119 3521
rect 32165 3475 32235 3521
rect 32281 3475 32351 3521
rect 32397 3475 32467 3521
rect 32513 3475 32583 3521
rect 32629 3475 32699 3521
rect 32745 3475 32815 3521
rect 32861 3475 32931 3521
rect 32977 3475 33047 3521
rect 33093 3475 33163 3521
rect 33209 3475 33279 3521
rect 33325 3475 33395 3521
rect 33441 3475 33511 3521
rect 33557 3475 33627 3521
rect 33673 3475 33743 3521
rect 33789 3475 33859 3521
rect 33905 3475 33975 3521
rect 34021 3475 34091 3521
rect 34137 3475 34207 3521
rect 34253 3475 34323 3521
rect 34369 3475 34439 3521
rect 34485 3475 34555 3521
rect 34601 3475 34671 3521
rect 34717 3475 34787 3521
rect 34833 3475 34903 3521
rect 34949 3475 35019 3521
rect 35065 3475 35135 3521
rect 35181 3475 35251 3521
rect 35297 3475 35367 3521
rect 35413 3475 35483 3521
rect 35529 3475 35599 3521
rect 35645 3475 35715 3521
rect 35761 3475 35831 3521
rect 35877 3475 35947 3521
rect 35993 3475 36063 3521
rect 36109 3475 36179 3521
rect 36225 3475 36295 3521
rect 36341 3475 36411 3521
rect 36457 3475 36527 3521
rect 36573 3475 36643 3521
rect 36689 3475 36759 3521
rect 36805 3475 36875 3521
rect 36921 3475 36991 3521
rect 37037 3475 37107 3521
rect 37153 3475 37223 3521
rect 37269 3475 37339 3521
rect 37385 3475 37455 3521
rect 37501 3475 37571 3521
rect 37617 3475 37687 3521
rect 37733 3475 37803 3521
rect 37849 3475 37919 3521
rect 37965 3475 38035 3521
rect 38081 3475 38151 3521
rect 38197 3475 38267 3521
rect 38313 3475 38383 3521
rect 38429 3475 38499 3521
rect 38545 3475 38615 3521
rect 38661 3475 38731 3521
rect 38777 3475 38847 3521
rect 38893 3475 38963 3521
rect 39009 3475 39079 3521
rect 39125 3475 39195 3521
rect 39241 3475 39311 3521
rect 39357 3475 39427 3521
rect 39473 3475 39543 3521
rect 39589 3475 39659 3521
rect 39705 3475 39775 3521
rect 39821 3475 39891 3521
rect 39937 3475 40007 3521
rect 40053 3475 40123 3521
rect 40169 3475 40180 3521
rect 28628 3405 40180 3475
rect 28628 3359 28639 3405
rect 28685 3359 28755 3405
rect 28801 3359 28871 3405
rect 28917 3359 28987 3405
rect 29033 3359 29103 3405
rect 29149 3359 29219 3405
rect 29265 3359 29335 3405
rect 29381 3359 29451 3405
rect 29497 3359 29567 3405
rect 29613 3359 29683 3405
rect 29729 3359 29799 3405
rect 29845 3359 29915 3405
rect 29961 3359 30031 3405
rect 30077 3359 30147 3405
rect 30193 3359 30263 3405
rect 30309 3359 30379 3405
rect 30425 3359 30495 3405
rect 30541 3359 30611 3405
rect 30657 3359 30727 3405
rect 30773 3359 30843 3405
rect 30889 3359 30959 3405
rect 31005 3359 31075 3405
rect 31121 3359 31191 3405
rect 31237 3359 31307 3405
rect 31353 3359 31423 3405
rect 31469 3359 31539 3405
rect 31585 3359 31655 3405
rect 31701 3359 31771 3405
rect 31817 3359 31887 3405
rect 31933 3359 32003 3405
rect 32049 3359 32119 3405
rect 32165 3359 32235 3405
rect 32281 3359 32351 3405
rect 32397 3359 32467 3405
rect 32513 3359 32583 3405
rect 32629 3359 32699 3405
rect 32745 3359 32815 3405
rect 32861 3359 32931 3405
rect 32977 3359 33047 3405
rect 33093 3359 33163 3405
rect 33209 3359 33279 3405
rect 33325 3359 33395 3405
rect 33441 3359 33511 3405
rect 33557 3359 33627 3405
rect 33673 3359 33743 3405
rect 33789 3359 33859 3405
rect 33905 3359 33975 3405
rect 34021 3359 34091 3405
rect 34137 3359 34207 3405
rect 34253 3359 34323 3405
rect 34369 3359 34439 3405
rect 34485 3359 34555 3405
rect 34601 3359 34671 3405
rect 34717 3359 34787 3405
rect 34833 3359 34903 3405
rect 34949 3359 35019 3405
rect 35065 3359 35135 3405
rect 35181 3359 35251 3405
rect 35297 3359 35367 3405
rect 35413 3359 35483 3405
rect 35529 3359 35599 3405
rect 35645 3359 35715 3405
rect 35761 3359 35831 3405
rect 35877 3359 35947 3405
rect 35993 3359 36063 3405
rect 36109 3359 36179 3405
rect 36225 3359 36295 3405
rect 36341 3359 36411 3405
rect 36457 3359 36527 3405
rect 36573 3359 36643 3405
rect 36689 3359 36759 3405
rect 36805 3359 36875 3405
rect 36921 3359 36991 3405
rect 37037 3359 37107 3405
rect 37153 3359 37223 3405
rect 37269 3359 37339 3405
rect 37385 3359 37455 3405
rect 37501 3359 37571 3405
rect 37617 3359 37687 3405
rect 37733 3359 37803 3405
rect 37849 3359 37919 3405
rect 37965 3359 38035 3405
rect 38081 3359 38151 3405
rect 38197 3359 38267 3405
rect 38313 3359 38383 3405
rect 38429 3359 38499 3405
rect 38545 3359 38615 3405
rect 38661 3359 38731 3405
rect 38777 3359 38847 3405
rect 38893 3359 38963 3405
rect 39009 3359 39079 3405
rect 39125 3359 39195 3405
rect 39241 3359 39311 3405
rect 39357 3359 39427 3405
rect 39473 3359 39543 3405
rect 39589 3359 39659 3405
rect 39705 3359 39775 3405
rect 39821 3359 39891 3405
rect 39937 3359 40007 3405
rect 40053 3359 40123 3405
rect 40169 3359 40180 3405
rect 28628 3289 40180 3359
rect 50834 3844 50845 3890
rect 50891 3844 50961 3890
rect 51007 3844 51077 3890
rect 51123 3844 51193 3890
rect 51239 3844 51309 3890
rect 51355 3844 51425 3890
rect 51471 3844 51541 3890
rect 51587 3844 51657 3890
rect 51703 3844 51773 3890
rect 51819 3844 51889 3890
rect 51935 3844 52005 3890
rect 52051 3844 52121 3890
rect 52167 3844 52237 3890
rect 52283 3844 52353 3890
rect 52399 3844 52469 3890
rect 52515 3844 52585 3890
rect 52631 3844 52701 3890
rect 52747 3844 52817 3890
rect 52863 3844 52933 3890
rect 52979 3844 53049 3890
rect 53095 3844 53165 3890
rect 53211 3844 53281 3890
rect 53327 3844 53397 3890
rect 53443 3844 53513 3890
rect 53559 3844 53629 3890
rect 53675 3844 53745 3890
rect 53791 3844 53861 3890
rect 53907 3844 53977 3890
rect 54023 3844 54093 3890
rect 54139 3844 54209 3890
rect 54255 3844 54325 3890
rect 54371 3844 54441 3890
rect 54487 3844 54557 3890
rect 54603 3844 54673 3890
rect 54719 3844 54789 3890
rect 54835 3844 54905 3890
rect 54951 3844 55021 3890
rect 55067 3844 55137 3890
rect 55183 3844 55253 3890
rect 55299 3844 55369 3890
rect 55415 3844 55485 3890
rect 55531 3844 55601 3890
rect 55647 3844 55717 3890
rect 55763 3844 55833 3890
rect 55879 3844 55949 3890
rect 55995 3844 56065 3890
rect 56111 3844 56181 3890
rect 56227 3844 56297 3890
rect 56343 3844 56413 3890
rect 56459 3844 56529 3890
rect 56575 3844 56586 3890
rect 50834 3774 56586 3844
rect 50834 3728 50845 3774
rect 50891 3728 50961 3774
rect 51007 3728 51077 3774
rect 51123 3728 51193 3774
rect 51239 3728 51309 3774
rect 51355 3728 51425 3774
rect 51471 3728 51541 3774
rect 51587 3728 51657 3774
rect 51703 3728 51773 3774
rect 51819 3728 51889 3774
rect 51935 3728 52005 3774
rect 52051 3728 52121 3774
rect 52167 3728 52237 3774
rect 52283 3728 52353 3774
rect 52399 3728 52469 3774
rect 52515 3728 52585 3774
rect 52631 3728 52701 3774
rect 52747 3728 52817 3774
rect 52863 3728 52933 3774
rect 52979 3728 53049 3774
rect 53095 3728 53165 3774
rect 53211 3728 53281 3774
rect 53327 3728 53397 3774
rect 53443 3728 53513 3774
rect 53559 3728 53629 3774
rect 53675 3728 53745 3774
rect 53791 3728 53861 3774
rect 53907 3728 53977 3774
rect 54023 3728 54093 3774
rect 54139 3728 54209 3774
rect 54255 3728 54325 3774
rect 54371 3728 54441 3774
rect 54487 3728 54557 3774
rect 54603 3728 54673 3774
rect 54719 3728 54789 3774
rect 54835 3728 54905 3774
rect 54951 3728 55021 3774
rect 55067 3728 55137 3774
rect 55183 3728 55253 3774
rect 55299 3728 55369 3774
rect 55415 3728 55485 3774
rect 55531 3728 55601 3774
rect 55647 3728 55717 3774
rect 55763 3728 55833 3774
rect 55879 3728 55949 3774
rect 55995 3728 56065 3774
rect 56111 3728 56181 3774
rect 56227 3728 56297 3774
rect 56343 3728 56413 3774
rect 56459 3728 56529 3774
rect 56575 3728 56586 3774
rect 50834 3658 56586 3728
rect 50834 3612 50845 3658
rect 50891 3612 50961 3658
rect 51007 3612 51077 3658
rect 51123 3612 51193 3658
rect 51239 3612 51309 3658
rect 51355 3612 51425 3658
rect 51471 3612 51541 3658
rect 51587 3612 51657 3658
rect 51703 3612 51773 3658
rect 51819 3612 51889 3658
rect 51935 3612 52005 3658
rect 52051 3612 52121 3658
rect 52167 3612 52237 3658
rect 52283 3612 52353 3658
rect 52399 3612 52469 3658
rect 52515 3612 52585 3658
rect 52631 3612 52701 3658
rect 52747 3612 52817 3658
rect 52863 3612 52933 3658
rect 52979 3612 53049 3658
rect 53095 3612 53165 3658
rect 53211 3612 53281 3658
rect 53327 3612 53397 3658
rect 53443 3612 53513 3658
rect 53559 3612 53629 3658
rect 53675 3612 53745 3658
rect 53791 3612 53861 3658
rect 53907 3612 53977 3658
rect 54023 3612 54093 3658
rect 54139 3612 54209 3658
rect 54255 3612 54325 3658
rect 54371 3612 54441 3658
rect 54487 3612 54557 3658
rect 54603 3612 54673 3658
rect 54719 3612 54789 3658
rect 54835 3612 54905 3658
rect 54951 3612 55021 3658
rect 55067 3612 55137 3658
rect 55183 3612 55253 3658
rect 55299 3612 55369 3658
rect 55415 3612 55485 3658
rect 55531 3612 55601 3658
rect 55647 3612 55717 3658
rect 55763 3612 55833 3658
rect 55879 3612 55949 3658
rect 55995 3612 56065 3658
rect 56111 3612 56181 3658
rect 56227 3612 56297 3658
rect 56343 3612 56413 3658
rect 56459 3612 56529 3658
rect 56575 3612 56586 3658
rect 50834 3542 56586 3612
rect 50834 3496 50845 3542
rect 50891 3496 50961 3542
rect 51007 3496 51077 3542
rect 51123 3496 51193 3542
rect 51239 3496 51309 3542
rect 51355 3496 51425 3542
rect 51471 3496 51541 3542
rect 51587 3496 51657 3542
rect 51703 3496 51773 3542
rect 51819 3496 51889 3542
rect 51935 3496 52005 3542
rect 52051 3496 52121 3542
rect 52167 3496 52237 3542
rect 52283 3496 52353 3542
rect 52399 3496 52469 3542
rect 52515 3496 52585 3542
rect 52631 3496 52701 3542
rect 52747 3496 52817 3542
rect 52863 3496 52933 3542
rect 52979 3496 53049 3542
rect 53095 3496 53165 3542
rect 53211 3496 53281 3542
rect 53327 3496 53397 3542
rect 53443 3496 53513 3542
rect 53559 3496 53629 3542
rect 53675 3496 53745 3542
rect 53791 3496 53861 3542
rect 53907 3496 53977 3542
rect 54023 3496 54093 3542
rect 54139 3496 54209 3542
rect 54255 3496 54325 3542
rect 54371 3496 54441 3542
rect 54487 3496 54557 3542
rect 54603 3496 54673 3542
rect 54719 3496 54789 3542
rect 54835 3496 54905 3542
rect 54951 3496 55021 3542
rect 55067 3496 55137 3542
rect 55183 3496 55253 3542
rect 55299 3496 55369 3542
rect 55415 3496 55485 3542
rect 55531 3496 55601 3542
rect 55647 3496 55717 3542
rect 55763 3496 55833 3542
rect 55879 3496 55949 3542
rect 55995 3496 56065 3542
rect 56111 3496 56181 3542
rect 56227 3496 56297 3542
rect 56343 3496 56413 3542
rect 56459 3496 56529 3542
rect 56575 3496 56586 3542
rect 50834 3426 56586 3496
rect 50834 3380 50845 3426
rect 50891 3380 50961 3426
rect 51007 3380 51077 3426
rect 51123 3380 51193 3426
rect 51239 3380 51309 3426
rect 51355 3380 51425 3426
rect 51471 3380 51541 3426
rect 51587 3380 51657 3426
rect 51703 3380 51773 3426
rect 51819 3380 51889 3426
rect 51935 3380 52005 3426
rect 52051 3380 52121 3426
rect 52167 3380 52237 3426
rect 52283 3380 52353 3426
rect 52399 3380 52469 3426
rect 52515 3380 52585 3426
rect 52631 3380 52701 3426
rect 52747 3380 52817 3426
rect 52863 3380 52933 3426
rect 52979 3380 53049 3426
rect 53095 3380 53165 3426
rect 53211 3380 53281 3426
rect 53327 3380 53397 3426
rect 53443 3380 53513 3426
rect 53559 3380 53629 3426
rect 53675 3380 53745 3426
rect 53791 3380 53861 3426
rect 53907 3380 53977 3426
rect 54023 3380 54093 3426
rect 54139 3380 54209 3426
rect 54255 3380 54325 3426
rect 54371 3380 54441 3426
rect 54487 3380 54557 3426
rect 54603 3380 54673 3426
rect 54719 3380 54789 3426
rect 54835 3380 54905 3426
rect 54951 3380 55021 3426
rect 55067 3380 55137 3426
rect 55183 3380 55253 3426
rect 55299 3380 55369 3426
rect 55415 3380 55485 3426
rect 55531 3380 55601 3426
rect 55647 3380 55717 3426
rect 55763 3380 55833 3426
rect 55879 3380 55949 3426
rect 55995 3380 56065 3426
rect 56111 3380 56181 3426
rect 56227 3380 56297 3426
rect 56343 3380 56413 3426
rect 56459 3380 56529 3426
rect 56575 3380 56586 3426
rect 50834 3310 56586 3380
rect 28628 3243 28639 3289
rect 28685 3243 28755 3289
rect 28801 3243 28871 3289
rect 28917 3243 28987 3289
rect 29033 3243 29103 3289
rect 29149 3243 29219 3289
rect 29265 3243 29335 3289
rect 29381 3243 29451 3289
rect 29497 3243 29567 3289
rect 29613 3243 29683 3289
rect 29729 3243 29799 3289
rect 29845 3243 29915 3289
rect 29961 3243 30031 3289
rect 30077 3243 30147 3289
rect 30193 3243 30263 3289
rect 30309 3243 30379 3289
rect 30425 3243 30495 3289
rect 30541 3243 30611 3289
rect 30657 3243 30727 3289
rect 30773 3243 30843 3289
rect 30889 3243 30959 3289
rect 31005 3243 31075 3289
rect 31121 3243 31191 3289
rect 31237 3243 31307 3289
rect 31353 3243 31423 3289
rect 31469 3243 31539 3289
rect 31585 3243 31655 3289
rect 31701 3243 31771 3289
rect 31817 3243 31887 3289
rect 31933 3243 32003 3289
rect 32049 3243 32119 3289
rect 32165 3243 32235 3289
rect 32281 3243 32351 3289
rect 32397 3243 32467 3289
rect 32513 3243 32583 3289
rect 32629 3243 32699 3289
rect 32745 3243 32815 3289
rect 32861 3243 32931 3289
rect 32977 3243 33047 3289
rect 33093 3243 33163 3289
rect 33209 3243 33279 3289
rect 33325 3243 33395 3289
rect 33441 3243 33511 3289
rect 33557 3243 33627 3289
rect 33673 3243 33743 3289
rect 33789 3243 33859 3289
rect 33905 3243 33975 3289
rect 34021 3243 34091 3289
rect 34137 3243 34207 3289
rect 34253 3243 34323 3289
rect 34369 3243 34439 3289
rect 34485 3243 34555 3289
rect 34601 3243 34671 3289
rect 34717 3243 34787 3289
rect 34833 3243 34903 3289
rect 34949 3243 35019 3289
rect 35065 3243 35135 3289
rect 35181 3243 35251 3289
rect 35297 3243 35367 3289
rect 35413 3243 35483 3289
rect 35529 3243 35599 3289
rect 35645 3243 35715 3289
rect 35761 3243 35831 3289
rect 35877 3243 35947 3289
rect 35993 3243 36063 3289
rect 36109 3243 36179 3289
rect 36225 3243 36295 3289
rect 36341 3243 36411 3289
rect 36457 3243 36527 3289
rect 36573 3243 36643 3289
rect 36689 3243 36759 3289
rect 36805 3243 36875 3289
rect 36921 3243 36991 3289
rect 37037 3243 37107 3289
rect 37153 3243 37223 3289
rect 37269 3243 37339 3289
rect 37385 3243 37455 3289
rect 37501 3243 37571 3289
rect 37617 3243 37687 3289
rect 37733 3243 37803 3289
rect 37849 3243 37919 3289
rect 37965 3243 38035 3289
rect 38081 3243 38151 3289
rect 38197 3243 38267 3289
rect 38313 3243 38383 3289
rect 38429 3243 38499 3289
rect 38545 3243 38615 3289
rect 38661 3243 38731 3289
rect 38777 3243 38847 3289
rect 38893 3243 38963 3289
rect 39009 3243 39079 3289
rect 39125 3243 39195 3289
rect 39241 3243 39311 3289
rect 39357 3243 39427 3289
rect 39473 3243 39543 3289
rect 39589 3243 39659 3289
rect 39705 3243 39775 3289
rect 39821 3243 39891 3289
rect 39937 3243 40007 3289
rect 40053 3243 40123 3289
rect 40169 3243 40180 3289
rect 28628 3173 40180 3243
rect 40611 3282 40791 3294
rect 40611 3230 40623 3282
rect 40779 3230 40791 3282
rect 40611 3218 40791 3230
rect 50834 3264 50845 3310
rect 50891 3264 50961 3310
rect 51007 3264 51077 3310
rect 51123 3264 51193 3310
rect 51239 3264 51309 3310
rect 51355 3264 51425 3310
rect 51471 3264 51541 3310
rect 51587 3264 51657 3310
rect 51703 3264 51773 3310
rect 51819 3264 51889 3310
rect 51935 3264 52005 3310
rect 52051 3264 52121 3310
rect 52167 3264 52237 3310
rect 52283 3264 52353 3310
rect 52399 3264 52469 3310
rect 52515 3264 52585 3310
rect 52631 3264 52701 3310
rect 52747 3264 52817 3310
rect 52863 3264 52933 3310
rect 52979 3264 53049 3310
rect 53095 3264 53165 3310
rect 53211 3264 53281 3310
rect 53327 3264 53397 3310
rect 53443 3264 53513 3310
rect 53559 3264 53629 3310
rect 53675 3264 53745 3310
rect 53791 3264 53861 3310
rect 53907 3264 53977 3310
rect 54023 3264 54093 3310
rect 54139 3264 54209 3310
rect 54255 3264 54325 3310
rect 54371 3264 54441 3310
rect 54487 3264 54557 3310
rect 54603 3264 54673 3310
rect 54719 3264 54789 3310
rect 54835 3264 54905 3310
rect 54951 3264 55021 3310
rect 55067 3264 55137 3310
rect 55183 3264 55253 3310
rect 55299 3264 55369 3310
rect 55415 3264 55485 3310
rect 55531 3264 55601 3310
rect 55647 3264 55717 3310
rect 55763 3264 55833 3310
rect 55879 3264 55949 3310
rect 55995 3264 56065 3310
rect 56111 3264 56181 3310
rect 56227 3264 56297 3310
rect 56343 3264 56413 3310
rect 56459 3264 56529 3310
rect 56575 3264 56586 3310
rect 28628 3127 28639 3173
rect 28685 3127 28755 3173
rect 28801 3127 28871 3173
rect 28917 3127 28987 3173
rect 29033 3127 29103 3173
rect 29149 3127 29219 3173
rect 29265 3127 29335 3173
rect 29381 3127 29451 3173
rect 29497 3127 29567 3173
rect 29613 3127 29683 3173
rect 29729 3127 29799 3173
rect 29845 3127 29915 3173
rect 29961 3127 30031 3173
rect 30077 3127 30147 3173
rect 30193 3127 30263 3173
rect 30309 3127 30379 3173
rect 30425 3127 30495 3173
rect 30541 3127 30611 3173
rect 30657 3127 30727 3173
rect 30773 3127 30843 3173
rect 30889 3127 30959 3173
rect 31005 3127 31075 3173
rect 31121 3127 31191 3173
rect 31237 3127 31307 3173
rect 31353 3127 31423 3173
rect 31469 3127 31539 3173
rect 31585 3127 31655 3173
rect 31701 3127 31771 3173
rect 31817 3127 31887 3173
rect 31933 3127 32003 3173
rect 32049 3127 32119 3173
rect 32165 3127 32235 3173
rect 32281 3127 32351 3173
rect 32397 3127 32467 3173
rect 32513 3127 32583 3173
rect 32629 3127 32699 3173
rect 32745 3127 32815 3173
rect 32861 3127 32931 3173
rect 32977 3127 33047 3173
rect 33093 3127 33163 3173
rect 33209 3127 33279 3173
rect 33325 3127 33395 3173
rect 33441 3127 33511 3173
rect 33557 3127 33627 3173
rect 33673 3127 33743 3173
rect 33789 3127 33859 3173
rect 33905 3127 33975 3173
rect 34021 3127 34091 3173
rect 34137 3127 34207 3173
rect 34253 3127 34323 3173
rect 34369 3127 34439 3173
rect 34485 3127 34555 3173
rect 34601 3127 34671 3173
rect 34717 3127 34787 3173
rect 34833 3127 34903 3173
rect 34949 3127 35019 3173
rect 35065 3127 35135 3173
rect 35181 3127 35251 3173
rect 35297 3127 35367 3173
rect 35413 3127 35483 3173
rect 35529 3127 35599 3173
rect 35645 3127 35715 3173
rect 35761 3127 35831 3173
rect 35877 3127 35947 3173
rect 35993 3127 36063 3173
rect 36109 3127 36179 3173
rect 36225 3127 36295 3173
rect 36341 3127 36411 3173
rect 36457 3127 36527 3173
rect 36573 3127 36643 3173
rect 36689 3127 36759 3173
rect 36805 3127 36875 3173
rect 36921 3127 36991 3173
rect 37037 3127 37107 3173
rect 37153 3127 37223 3173
rect 37269 3127 37339 3173
rect 37385 3127 37455 3173
rect 37501 3127 37571 3173
rect 37617 3127 37687 3173
rect 37733 3127 37803 3173
rect 37849 3127 37919 3173
rect 37965 3127 38035 3173
rect 38081 3127 38151 3173
rect 38197 3127 38267 3173
rect 38313 3127 38383 3173
rect 38429 3127 38499 3173
rect 38545 3127 38615 3173
rect 38661 3127 38731 3173
rect 38777 3127 38847 3173
rect 38893 3127 38963 3173
rect 39009 3127 39079 3173
rect 39125 3127 39195 3173
rect 39241 3127 39311 3173
rect 39357 3127 39427 3173
rect 39473 3127 39543 3173
rect 39589 3127 39659 3173
rect 39705 3127 39775 3173
rect 39821 3127 39891 3173
rect 39937 3127 40007 3173
rect 40053 3127 40123 3173
rect 40169 3127 40180 3173
rect 28628 3057 40180 3127
rect 28628 3011 28639 3057
rect 28685 3011 28755 3057
rect 28801 3011 28871 3057
rect 28917 3011 28987 3057
rect 29033 3011 29103 3057
rect 29149 3011 29219 3057
rect 29265 3011 29335 3057
rect 29381 3011 29451 3057
rect 29497 3011 29567 3057
rect 29613 3011 29683 3057
rect 29729 3011 29799 3057
rect 29845 3011 29915 3057
rect 29961 3011 30031 3057
rect 30077 3011 30147 3057
rect 30193 3011 30263 3057
rect 30309 3011 30379 3057
rect 30425 3011 30495 3057
rect 30541 3011 30611 3057
rect 30657 3011 30727 3057
rect 30773 3011 30843 3057
rect 30889 3011 30959 3057
rect 31005 3011 31075 3057
rect 31121 3011 31191 3057
rect 31237 3011 31307 3057
rect 31353 3011 31423 3057
rect 31469 3011 31539 3057
rect 31585 3011 31655 3057
rect 31701 3011 31771 3057
rect 31817 3011 31887 3057
rect 31933 3011 32003 3057
rect 32049 3011 32119 3057
rect 32165 3011 32235 3057
rect 32281 3011 32351 3057
rect 32397 3011 32467 3057
rect 32513 3011 32583 3057
rect 32629 3011 32699 3057
rect 32745 3011 32815 3057
rect 32861 3011 32931 3057
rect 32977 3011 33047 3057
rect 33093 3011 33163 3057
rect 33209 3011 33279 3057
rect 33325 3011 33395 3057
rect 33441 3011 33511 3057
rect 33557 3011 33627 3057
rect 33673 3011 33743 3057
rect 33789 3011 33859 3057
rect 33905 3011 33975 3057
rect 34021 3011 34091 3057
rect 34137 3011 34207 3057
rect 34253 3011 34323 3057
rect 34369 3011 34439 3057
rect 34485 3011 34555 3057
rect 34601 3011 34671 3057
rect 34717 3011 34787 3057
rect 34833 3011 34903 3057
rect 34949 3011 35019 3057
rect 35065 3011 35135 3057
rect 35181 3011 35251 3057
rect 35297 3011 35367 3057
rect 35413 3011 35483 3057
rect 35529 3011 35599 3057
rect 35645 3011 35715 3057
rect 35761 3011 35831 3057
rect 35877 3011 35947 3057
rect 35993 3011 36063 3057
rect 36109 3011 36179 3057
rect 36225 3011 36295 3057
rect 36341 3011 36411 3057
rect 36457 3011 36527 3057
rect 36573 3011 36643 3057
rect 36689 3011 36759 3057
rect 36805 3011 36875 3057
rect 36921 3011 36991 3057
rect 37037 3011 37107 3057
rect 37153 3011 37223 3057
rect 37269 3011 37339 3057
rect 37385 3011 37455 3057
rect 37501 3011 37571 3057
rect 37617 3011 37687 3057
rect 37733 3011 37803 3057
rect 37849 3011 37919 3057
rect 37965 3011 38035 3057
rect 38081 3011 38151 3057
rect 38197 3011 38267 3057
rect 38313 3011 38383 3057
rect 38429 3011 38499 3057
rect 38545 3011 38615 3057
rect 38661 3011 38731 3057
rect 38777 3011 38847 3057
rect 38893 3011 38963 3057
rect 39009 3011 39079 3057
rect 39125 3011 39195 3057
rect 39241 3011 39311 3057
rect 39357 3011 39427 3057
rect 39473 3011 39543 3057
rect 39589 3011 39659 3057
rect 39705 3011 39775 3057
rect 39821 3011 39891 3057
rect 39937 3011 40007 3057
rect 40053 3011 40123 3057
rect 40169 3011 40180 3057
rect 28628 2941 40180 3011
rect 28628 2895 28639 2941
rect 28685 2895 28755 2941
rect 28801 2895 28871 2941
rect 28917 2895 28987 2941
rect 29033 2895 29103 2941
rect 29149 2895 29219 2941
rect 29265 2895 29335 2941
rect 29381 2895 29451 2941
rect 29497 2895 29567 2941
rect 29613 2895 29683 2941
rect 29729 2895 29799 2941
rect 29845 2895 29915 2941
rect 29961 2895 30031 2941
rect 30077 2895 30147 2941
rect 30193 2895 30263 2941
rect 30309 2895 30379 2941
rect 30425 2895 30495 2941
rect 30541 2895 30611 2941
rect 30657 2895 30727 2941
rect 30773 2895 30843 2941
rect 30889 2895 30959 2941
rect 31005 2895 31075 2941
rect 31121 2895 31191 2941
rect 31237 2895 31307 2941
rect 31353 2895 31423 2941
rect 31469 2895 31539 2941
rect 31585 2895 31655 2941
rect 31701 2895 31771 2941
rect 31817 2895 31887 2941
rect 31933 2895 32003 2941
rect 32049 2895 32119 2941
rect 32165 2895 32235 2941
rect 32281 2895 32351 2941
rect 32397 2895 32467 2941
rect 32513 2895 32583 2941
rect 32629 2895 32699 2941
rect 32745 2895 32815 2941
rect 32861 2895 32931 2941
rect 32977 2895 33047 2941
rect 33093 2895 33163 2941
rect 33209 2895 33279 2941
rect 33325 2895 33395 2941
rect 33441 2895 33511 2941
rect 33557 2895 33627 2941
rect 33673 2895 33743 2941
rect 33789 2895 33859 2941
rect 33905 2895 33975 2941
rect 34021 2895 34091 2941
rect 34137 2895 34207 2941
rect 34253 2895 34323 2941
rect 34369 2895 34439 2941
rect 34485 2895 34555 2941
rect 34601 2895 34671 2941
rect 34717 2895 34787 2941
rect 34833 2895 34903 2941
rect 34949 2895 35019 2941
rect 35065 2895 35135 2941
rect 35181 2895 35251 2941
rect 35297 2895 35367 2941
rect 35413 2895 35483 2941
rect 35529 2895 35599 2941
rect 35645 2895 35715 2941
rect 35761 2895 35831 2941
rect 35877 2895 35947 2941
rect 35993 2895 36063 2941
rect 36109 2895 36179 2941
rect 36225 2895 36295 2941
rect 36341 2895 36411 2941
rect 36457 2895 36527 2941
rect 36573 2895 36643 2941
rect 36689 2895 36759 2941
rect 36805 2895 36875 2941
rect 36921 2895 36991 2941
rect 37037 2895 37107 2941
rect 37153 2895 37223 2941
rect 37269 2895 37339 2941
rect 37385 2895 37455 2941
rect 37501 2895 37571 2941
rect 37617 2895 37687 2941
rect 37733 2895 37803 2941
rect 37849 2895 37919 2941
rect 37965 2895 38035 2941
rect 38081 2895 38151 2941
rect 38197 2895 38267 2941
rect 38313 2895 38383 2941
rect 38429 2895 38499 2941
rect 38545 2895 38615 2941
rect 38661 2895 38731 2941
rect 38777 2895 38847 2941
rect 38893 2895 38963 2941
rect 39009 2895 39079 2941
rect 39125 2895 39195 2941
rect 39241 2895 39311 2941
rect 39357 2895 39427 2941
rect 39473 2895 39543 2941
rect 39589 2895 39659 2941
rect 39705 2895 39775 2941
rect 39821 2895 39891 2941
rect 39937 2895 40007 2941
rect 40053 2895 40123 2941
rect 40169 2895 40180 2941
rect 28628 2825 40180 2895
rect 28628 2779 28639 2825
rect 28685 2779 28755 2825
rect 28801 2779 28871 2825
rect 28917 2779 28987 2825
rect 29033 2779 29103 2825
rect 29149 2779 29219 2825
rect 29265 2779 29335 2825
rect 29381 2779 29451 2825
rect 29497 2779 29567 2825
rect 29613 2779 29683 2825
rect 29729 2779 29799 2825
rect 29845 2779 29915 2825
rect 29961 2779 30031 2825
rect 30077 2779 30147 2825
rect 30193 2779 30263 2825
rect 30309 2779 30379 2825
rect 30425 2779 30495 2825
rect 30541 2779 30611 2825
rect 30657 2779 30727 2825
rect 30773 2779 30843 2825
rect 30889 2779 30959 2825
rect 31005 2779 31075 2825
rect 31121 2779 31191 2825
rect 31237 2779 31307 2825
rect 31353 2779 31423 2825
rect 31469 2779 31539 2825
rect 31585 2779 31655 2825
rect 31701 2779 31771 2825
rect 31817 2779 31887 2825
rect 31933 2779 32003 2825
rect 32049 2779 32119 2825
rect 32165 2779 32235 2825
rect 32281 2779 32351 2825
rect 32397 2779 32467 2825
rect 32513 2779 32583 2825
rect 32629 2779 32699 2825
rect 32745 2779 32815 2825
rect 32861 2779 32931 2825
rect 32977 2779 33047 2825
rect 33093 2779 33163 2825
rect 33209 2779 33279 2825
rect 33325 2779 33395 2825
rect 33441 2779 33511 2825
rect 33557 2779 33627 2825
rect 33673 2779 33743 2825
rect 33789 2779 33859 2825
rect 33905 2779 33975 2825
rect 34021 2779 34091 2825
rect 34137 2779 34207 2825
rect 34253 2779 34323 2825
rect 34369 2779 34439 2825
rect 34485 2779 34555 2825
rect 34601 2779 34671 2825
rect 34717 2779 34787 2825
rect 34833 2779 34903 2825
rect 34949 2779 35019 2825
rect 35065 2779 35135 2825
rect 35181 2779 35251 2825
rect 35297 2779 35367 2825
rect 35413 2779 35483 2825
rect 35529 2779 35599 2825
rect 35645 2779 35715 2825
rect 35761 2779 35831 2825
rect 35877 2779 35947 2825
rect 35993 2779 36063 2825
rect 36109 2779 36179 2825
rect 36225 2779 36295 2825
rect 36341 2779 36411 2825
rect 36457 2779 36527 2825
rect 36573 2779 36643 2825
rect 36689 2779 36759 2825
rect 36805 2779 36875 2825
rect 36921 2779 36991 2825
rect 37037 2779 37107 2825
rect 37153 2779 37223 2825
rect 37269 2779 37339 2825
rect 37385 2779 37455 2825
rect 37501 2779 37571 2825
rect 37617 2779 37687 2825
rect 37733 2779 37803 2825
rect 37849 2779 37919 2825
rect 37965 2779 38035 2825
rect 38081 2779 38151 2825
rect 38197 2779 38267 2825
rect 38313 2779 38383 2825
rect 38429 2779 38499 2825
rect 38545 2779 38615 2825
rect 38661 2779 38731 2825
rect 38777 2779 38847 2825
rect 38893 2779 38963 2825
rect 39009 2779 39079 2825
rect 39125 2779 39195 2825
rect 39241 2779 39311 2825
rect 39357 2779 39427 2825
rect 39473 2779 39543 2825
rect 39589 2779 39659 2825
rect 39705 2779 39775 2825
rect 39821 2779 39891 2825
rect 39937 2779 40007 2825
rect 40053 2779 40123 2825
rect 40169 2779 40180 2825
rect 28628 2709 40180 2779
rect 28628 2663 28639 2709
rect 28685 2663 28755 2709
rect 28801 2663 28871 2709
rect 28917 2663 28987 2709
rect 29033 2663 29103 2709
rect 29149 2663 29219 2709
rect 29265 2663 29335 2709
rect 29381 2663 29451 2709
rect 29497 2663 29567 2709
rect 29613 2663 29683 2709
rect 29729 2663 29799 2709
rect 29845 2663 29915 2709
rect 29961 2663 30031 2709
rect 30077 2663 30147 2709
rect 30193 2663 30263 2709
rect 30309 2663 30379 2709
rect 30425 2663 30495 2709
rect 30541 2663 30611 2709
rect 30657 2663 30727 2709
rect 30773 2663 30843 2709
rect 30889 2663 30959 2709
rect 31005 2663 31075 2709
rect 31121 2663 31191 2709
rect 31237 2663 31307 2709
rect 31353 2663 31423 2709
rect 31469 2663 31539 2709
rect 31585 2663 31655 2709
rect 31701 2663 31771 2709
rect 31817 2663 31887 2709
rect 31933 2663 32003 2709
rect 32049 2663 32119 2709
rect 32165 2663 32235 2709
rect 32281 2663 32351 2709
rect 32397 2663 32467 2709
rect 32513 2663 32583 2709
rect 32629 2663 32699 2709
rect 32745 2663 32815 2709
rect 32861 2663 32931 2709
rect 32977 2663 33047 2709
rect 33093 2663 33163 2709
rect 33209 2663 33279 2709
rect 33325 2663 33395 2709
rect 33441 2663 33511 2709
rect 33557 2663 33627 2709
rect 33673 2663 33743 2709
rect 33789 2663 33859 2709
rect 33905 2663 33975 2709
rect 34021 2663 34091 2709
rect 34137 2663 34207 2709
rect 34253 2663 34323 2709
rect 34369 2663 34439 2709
rect 34485 2663 34555 2709
rect 34601 2663 34671 2709
rect 34717 2663 34787 2709
rect 34833 2663 34903 2709
rect 34949 2663 35019 2709
rect 35065 2663 35135 2709
rect 35181 2663 35251 2709
rect 35297 2663 35367 2709
rect 35413 2663 35483 2709
rect 35529 2663 35599 2709
rect 35645 2663 35715 2709
rect 35761 2663 35831 2709
rect 35877 2663 35947 2709
rect 35993 2663 36063 2709
rect 36109 2663 36179 2709
rect 36225 2663 36295 2709
rect 36341 2663 36411 2709
rect 36457 2663 36527 2709
rect 36573 2663 36643 2709
rect 36689 2663 36759 2709
rect 36805 2663 36875 2709
rect 36921 2663 36991 2709
rect 37037 2663 37107 2709
rect 37153 2663 37223 2709
rect 37269 2663 37339 2709
rect 37385 2663 37455 2709
rect 37501 2663 37571 2709
rect 37617 2663 37687 2709
rect 37733 2663 37803 2709
rect 37849 2663 37919 2709
rect 37965 2663 38035 2709
rect 38081 2663 38151 2709
rect 38197 2663 38267 2709
rect 38313 2663 38383 2709
rect 38429 2663 38499 2709
rect 38545 2663 38615 2709
rect 38661 2663 38731 2709
rect 38777 2663 38847 2709
rect 38893 2663 38963 2709
rect 39009 2663 39079 2709
rect 39125 2663 39195 2709
rect 39241 2663 39311 2709
rect 39357 2663 39427 2709
rect 39473 2663 39543 2709
rect 39589 2663 39659 2709
rect 39705 2663 39775 2709
rect 39821 2663 39891 2709
rect 39937 2663 40007 2709
rect 40053 2663 40123 2709
rect 40169 2663 40180 2709
rect 28628 2593 40180 2663
rect 28628 2547 28639 2593
rect 28685 2547 28755 2593
rect 28801 2547 28871 2593
rect 28917 2547 28987 2593
rect 29033 2547 29103 2593
rect 29149 2547 29219 2593
rect 29265 2547 29335 2593
rect 29381 2547 29451 2593
rect 29497 2547 29567 2593
rect 29613 2547 29683 2593
rect 29729 2547 29799 2593
rect 29845 2547 29915 2593
rect 29961 2547 30031 2593
rect 30077 2547 30147 2593
rect 30193 2547 30263 2593
rect 30309 2547 30379 2593
rect 30425 2547 30495 2593
rect 30541 2547 30611 2593
rect 30657 2547 30727 2593
rect 30773 2547 30843 2593
rect 30889 2547 30959 2593
rect 31005 2547 31075 2593
rect 31121 2547 31191 2593
rect 31237 2547 31307 2593
rect 31353 2547 31423 2593
rect 31469 2547 31539 2593
rect 31585 2547 31655 2593
rect 31701 2547 31771 2593
rect 31817 2547 31887 2593
rect 31933 2547 32003 2593
rect 32049 2547 32119 2593
rect 32165 2547 32235 2593
rect 32281 2547 32351 2593
rect 32397 2547 32467 2593
rect 32513 2547 32583 2593
rect 32629 2547 32699 2593
rect 32745 2547 32815 2593
rect 32861 2547 32931 2593
rect 32977 2547 33047 2593
rect 33093 2547 33163 2593
rect 33209 2547 33279 2593
rect 33325 2547 33395 2593
rect 33441 2547 33511 2593
rect 33557 2547 33627 2593
rect 33673 2547 33743 2593
rect 33789 2547 33859 2593
rect 33905 2547 33975 2593
rect 34021 2547 34091 2593
rect 34137 2547 34207 2593
rect 34253 2547 34323 2593
rect 34369 2547 34439 2593
rect 34485 2547 34555 2593
rect 34601 2547 34671 2593
rect 34717 2547 34787 2593
rect 34833 2547 34903 2593
rect 34949 2547 35019 2593
rect 35065 2547 35135 2593
rect 35181 2547 35251 2593
rect 35297 2547 35367 2593
rect 35413 2547 35483 2593
rect 35529 2547 35599 2593
rect 35645 2547 35715 2593
rect 35761 2547 35831 2593
rect 35877 2547 35947 2593
rect 35993 2547 36063 2593
rect 36109 2547 36179 2593
rect 36225 2547 36295 2593
rect 36341 2547 36411 2593
rect 36457 2547 36527 2593
rect 36573 2547 36643 2593
rect 36689 2547 36759 2593
rect 36805 2547 36875 2593
rect 36921 2547 36991 2593
rect 37037 2547 37107 2593
rect 37153 2547 37223 2593
rect 37269 2547 37339 2593
rect 37385 2547 37455 2593
rect 37501 2547 37571 2593
rect 37617 2547 37687 2593
rect 37733 2547 37803 2593
rect 37849 2547 37919 2593
rect 37965 2547 38035 2593
rect 38081 2547 38151 2593
rect 38197 2547 38267 2593
rect 38313 2547 38383 2593
rect 38429 2547 38499 2593
rect 38545 2547 38615 2593
rect 38661 2547 38731 2593
rect 38777 2547 38847 2593
rect 38893 2547 38963 2593
rect 39009 2547 39079 2593
rect 39125 2547 39195 2593
rect 39241 2547 39311 2593
rect 39357 2547 39427 2593
rect 39473 2547 39543 2593
rect 39589 2547 39659 2593
rect 39705 2547 39775 2593
rect 39821 2547 39891 2593
rect 39937 2547 40007 2593
rect 40053 2547 40123 2593
rect 40169 2547 40180 2593
rect 28628 2477 40180 2547
rect 28628 2431 28639 2477
rect 28685 2431 28755 2477
rect 28801 2431 28871 2477
rect 28917 2431 28987 2477
rect 29033 2431 29103 2477
rect 29149 2431 29219 2477
rect 29265 2431 29335 2477
rect 29381 2431 29451 2477
rect 29497 2431 29567 2477
rect 29613 2431 29683 2477
rect 29729 2431 29799 2477
rect 29845 2431 29915 2477
rect 29961 2431 30031 2477
rect 30077 2431 30147 2477
rect 30193 2431 30263 2477
rect 30309 2431 30379 2477
rect 30425 2431 30495 2477
rect 30541 2431 30611 2477
rect 30657 2431 30727 2477
rect 30773 2431 30843 2477
rect 30889 2431 30959 2477
rect 31005 2431 31075 2477
rect 31121 2431 31191 2477
rect 31237 2431 31307 2477
rect 31353 2431 31423 2477
rect 31469 2431 31539 2477
rect 31585 2431 31655 2477
rect 31701 2431 31771 2477
rect 31817 2431 31887 2477
rect 31933 2431 32003 2477
rect 32049 2431 32119 2477
rect 32165 2431 32235 2477
rect 32281 2431 32351 2477
rect 32397 2431 32467 2477
rect 32513 2431 32583 2477
rect 32629 2431 32699 2477
rect 32745 2431 32815 2477
rect 32861 2431 32931 2477
rect 32977 2431 33047 2477
rect 33093 2431 33163 2477
rect 33209 2431 33279 2477
rect 33325 2431 33395 2477
rect 33441 2431 33511 2477
rect 33557 2431 33627 2477
rect 33673 2431 33743 2477
rect 33789 2431 33859 2477
rect 33905 2431 33975 2477
rect 34021 2431 34091 2477
rect 34137 2431 34207 2477
rect 34253 2431 34323 2477
rect 34369 2431 34439 2477
rect 34485 2431 34555 2477
rect 34601 2431 34671 2477
rect 34717 2431 34787 2477
rect 34833 2431 34903 2477
rect 34949 2431 35019 2477
rect 35065 2431 35135 2477
rect 35181 2431 35251 2477
rect 35297 2431 35367 2477
rect 35413 2431 35483 2477
rect 35529 2431 35599 2477
rect 35645 2431 35715 2477
rect 35761 2431 35831 2477
rect 35877 2431 35947 2477
rect 35993 2431 36063 2477
rect 36109 2431 36179 2477
rect 36225 2431 36295 2477
rect 36341 2431 36411 2477
rect 36457 2431 36527 2477
rect 36573 2431 36643 2477
rect 36689 2431 36759 2477
rect 36805 2431 36875 2477
rect 36921 2431 36991 2477
rect 37037 2431 37107 2477
rect 37153 2431 37223 2477
rect 37269 2431 37339 2477
rect 37385 2431 37455 2477
rect 37501 2431 37571 2477
rect 37617 2431 37687 2477
rect 37733 2431 37803 2477
rect 37849 2431 37919 2477
rect 37965 2431 38035 2477
rect 38081 2431 38151 2477
rect 38197 2431 38267 2477
rect 38313 2431 38383 2477
rect 38429 2431 38499 2477
rect 38545 2431 38615 2477
rect 38661 2431 38731 2477
rect 38777 2431 38847 2477
rect 38893 2431 38963 2477
rect 39009 2431 39079 2477
rect 39125 2431 39195 2477
rect 39241 2431 39311 2477
rect 39357 2431 39427 2477
rect 39473 2431 39543 2477
rect 39589 2431 39659 2477
rect 39705 2431 39775 2477
rect 39821 2431 39891 2477
rect 39937 2431 40007 2477
rect 40053 2431 40123 2477
rect 40169 2431 40180 2477
rect 28628 2361 40180 2431
rect 28628 2315 28639 2361
rect 28685 2315 28755 2361
rect 28801 2315 28871 2361
rect 28917 2315 28987 2361
rect 29033 2315 29103 2361
rect 29149 2315 29219 2361
rect 29265 2315 29335 2361
rect 29381 2315 29451 2361
rect 29497 2315 29567 2361
rect 29613 2315 29683 2361
rect 29729 2315 29799 2361
rect 29845 2315 29915 2361
rect 29961 2315 30031 2361
rect 30077 2315 30147 2361
rect 30193 2315 30263 2361
rect 30309 2315 30379 2361
rect 30425 2315 30495 2361
rect 30541 2315 30611 2361
rect 30657 2315 30727 2361
rect 30773 2315 30843 2361
rect 30889 2315 30959 2361
rect 31005 2315 31075 2361
rect 31121 2315 31191 2361
rect 31237 2315 31307 2361
rect 31353 2315 31423 2361
rect 31469 2315 31539 2361
rect 31585 2315 31655 2361
rect 31701 2315 31771 2361
rect 31817 2315 31887 2361
rect 31933 2315 32003 2361
rect 32049 2315 32119 2361
rect 32165 2315 32235 2361
rect 32281 2315 32351 2361
rect 32397 2315 32467 2361
rect 32513 2315 32583 2361
rect 32629 2315 32699 2361
rect 32745 2315 32815 2361
rect 32861 2315 32931 2361
rect 32977 2315 33047 2361
rect 33093 2315 33163 2361
rect 33209 2315 33279 2361
rect 33325 2315 33395 2361
rect 33441 2315 33511 2361
rect 33557 2315 33627 2361
rect 33673 2315 33743 2361
rect 33789 2315 33859 2361
rect 33905 2315 33975 2361
rect 34021 2315 34091 2361
rect 34137 2315 34207 2361
rect 34253 2315 34323 2361
rect 34369 2315 34439 2361
rect 34485 2315 34555 2361
rect 34601 2315 34671 2361
rect 34717 2315 34787 2361
rect 34833 2315 34903 2361
rect 34949 2315 35019 2361
rect 35065 2315 35135 2361
rect 35181 2315 35251 2361
rect 35297 2315 35367 2361
rect 35413 2315 35483 2361
rect 35529 2315 35599 2361
rect 35645 2315 35715 2361
rect 35761 2315 35831 2361
rect 35877 2315 35947 2361
rect 35993 2315 36063 2361
rect 36109 2315 36179 2361
rect 36225 2315 36295 2361
rect 36341 2315 36411 2361
rect 36457 2315 36527 2361
rect 36573 2315 36643 2361
rect 36689 2315 36759 2361
rect 36805 2315 36875 2361
rect 36921 2315 36991 2361
rect 37037 2315 37107 2361
rect 37153 2315 37223 2361
rect 37269 2315 37339 2361
rect 37385 2315 37455 2361
rect 37501 2315 37571 2361
rect 37617 2315 37687 2361
rect 37733 2315 37803 2361
rect 37849 2315 37919 2361
rect 37965 2315 38035 2361
rect 38081 2315 38151 2361
rect 38197 2315 38267 2361
rect 38313 2315 38383 2361
rect 38429 2315 38499 2361
rect 38545 2315 38615 2361
rect 38661 2315 38731 2361
rect 38777 2315 38847 2361
rect 38893 2315 38963 2361
rect 39009 2315 39079 2361
rect 39125 2315 39195 2361
rect 39241 2315 39311 2361
rect 39357 2315 39427 2361
rect 39473 2315 39543 2361
rect 39589 2315 39659 2361
rect 39705 2315 39775 2361
rect 39821 2315 39891 2361
rect 39937 2315 40007 2361
rect 40053 2315 40123 2361
rect 40169 2315 40180 2361
rect 28628 2245 40180 2315
rect 28628 2199 28639 2245
rect 28685 2199 28755 2245
rect 28801 2199 28871 2245
rect 28917 2199 28987 2245
rect 29033 2199 29103 2245
rect 29149 2199 29219 2245
rect 29265 2199 29335 2245
rect 29381 2199 29451 2245
rect 29497 2199 29567 2245
rect 29613 2199 29683 2245
rect 29729 2199 29799 2245
rect 29845 2199 29915 2245
rect 29961 2199 30031 2245
rect 30077 2199 30147 2245
rect 30193 2199 30263 2245
rect 30309 2199 30379 2245
rect 30425 2199 30495 2245
rect 30541 2199 30611 2245
rect 30657 2199 30727 2245
rect 30773 2199 30843 2245
rect 30889 2199 30959 2245
rect 31005 2199 31075 2245
rect 31121 2199 31191 2245
rect 31237 2199 31307 2245
rect 31353 2199 31423 2245
rect 31469 2199 31539 2245
rect 31585 2199 31655 2245
rect 31701 2199 31771 2245
rect 31817 2199 31887 2245
rect 31933 2199 32003 2245
rect 32049 2199 32119 2245
rect 32165 2199 32235 2245
rect 32281 2199 32351 2245
rect 32397 2199 32467 2245
rect 32513 2199 32583 2245
rect 32629 2199 32699 2245
rect 32745 2199 32815 2245
rect 32861 2199 32931 2245
rect 32977 2199 33047 2245
rect 33093 2199 33163 2245
rect 33209 2199 33279 2245
rect 33325 2199 33395 2245
rect 33441 2199 33511 2245
rect 33557 2199 33627 2245
rect 33673 2199 33743 2245
rect 33789 2199 33859 2245
rect 33905 2199 33975 2245
rect 34021 2199 34091 2245
rect 34137 2199 34207 2245
rect 34253 2199 34323 2245
rect 34369 2199 34439 2245
rect 34485 2199 34555 2245
rect 34601 2199 34671 2245
rect 34717 2199 34787 2245
rect 34833 2199 34903 2245
rect 34949 2199 35019 2245
rect 35065 2199 35135 2245
rect 35181 2199 35251 2245
rect 35297 2199 35367 2245
rect 35413 2199 35483 2245
rect 35529 2199 35599 2245
rect 35645 2199 35715 2245
rect 35761 2199 35831 2245
rect 35877 2199 35947 2245
rect 35993 2199 36063 2245
rect 36109 2199 36179 2245
rect 36225 2199 36295 2245
rect 36341 2199 36411 2245
rect 36457 2199 36527 2245
rect 36573 2199 36643 2245
rect 36689 2199 36759 2245
rect 36805 2199 36875 2245
rect 36921 2199 36991 2245
rect 37037 2199 37107 2245
rect 37153 2199 37223 2245
rect 37269 2199 37339 2245
rect 37385 2199 37455 2245
rect 37501 2199 37571 2245
rect 37617 2199 37687 2245
rect 37733 2199 37803 2245
rect 37849 2199 37919 2245
rect 37965 2199 38035 2245
rect 38081 2199 38151 2245
rect 38197 2199 38267 2245
rect 38313 2199 38383 2245
rect 38429 2199 38499 2245
rect 38545 2199 38615 2245
rect 38661 2199 38731 2245
rect 38777 2199 38847 2245
rect 38893 2199 38963 2245
rect 39009 2199 39079 2245
rect 39125 2199 39195 2245
rect 39241 2199 39311 2245
rect 39357 2199 39427 2245
rect 39473 2199 39543 2245
rect 39589 2199 39659 2245
rect 39705 2199 39775 2245
rect 39821 2199 39891 2245
rect 39937 2199 40007 2245
rect 40053 2199 40123 2245
rect 40169 2199 40180 2245
rect 28628 2129 40180 2199
rect 28628 2083 28639 2129
rect 28685 2083 28755 2129
rect 28801 2083 28871 2129
rect 28917 2083 28987 2129
rect 29033 2083 29103 2129
rect 29149 2083 29219 2129
rect 29265 2083 29335 2129
rect 29381 2083 29451 2129
rect 29497 2083 29567 2129
rect 29613 2083 29683 2129
rect 29729 2083 29799 2129
rect 29845 2083 29915 2129
rect 29961 2083 30031 2129
rect 30077 2083 30147 2129
rect 30193 2083 30263 2129
rect 30309 2083 30379 2129
rect 30425 2083 30495 2129
rect 30541 2083 30611 2129
rect 30657 2083 30727 2129
rect 30773 2083 30843 2129
rect 30889 2083 30959 2129
rect 31005 2083 31075 2129
rect 31121 2083 31191 2129
rect 31237 2083 31307 2129
rect 31353 2083 31423 2129
rect 31469 2083 31539 2129
rect 31585 2083 31655 2129
rect 31701 2083 31771 2129
rect 31817 2083 31887 2129
rect 31933 2083 32003 2129
rect 32049 2083 32119 2129
rect 32165 2083 32235 2129
rect 32281 2083 32351 2129
rect 32397 2083 32467 2129
rect 32513 2083 32583 2129
rect 32629 2083 32699 2129
rect 32745 2083 32815 2129
rect 32861 2083 32931 2129
rect 32977 2083 33047 2129
rect 33093 2083 33163 2129
rect 33209 2083 33279 2129
rect 33325 2083 33395 2129
rect 33441 2083 33511 2129
rect 33557 2083 33627 2129
rect 33673 2083 33743 2129
rect 33789 2083 33859 2129
rect 33905 2083 33975 2129
rect 34021 2083 34091 2129
rect 34137 2083 34207 2129
rect 34253 2083 34323 2129
rect 34369 2083 34439 2129
rect 34485 2083 34555 2129
rect 34601 2083 34671 2129
rect 34717 2083 34787 2129
rect 34833 2083 34903 2129
rect 34949 2083 35019 2129
rect 35065 2083 35135 2129
rect 35181 2083 35251 2129
rect 35297 2083 35367 2129
rect 35413 2083 35483 2129
rect 35529 2083 35599 2129
rect 35645 2083 35715 2129
rect 35761 2083 35831 2129
rect 35877 2083 35947 2129
rect 35993 2083 36063 2129
rect 36109 2083 36179 2129
rect 36225 2083 36295 2129
rect 36341 2083 36411 2129
rect 36457 2083 36527 2129
rect 36573 2083 36643 2129
rect 36689 2083 36759 2129
rect 36805 2083 36875 2129
rect 36921 2083 36991 2129
rect 37037 2083 37107 2129
rect 37153 2083 37223 2129
rect 37269 2083 37339 2129
rect 37385 2083 37455 2129
rect 37501 2083 37571 2129
rect 37617 2083 37687 2129
rect 37733 2083 37803 2129
rect 37849 2083 37919 2129
rect 37965 2083 38035 2129
rect 38081 2083 38151 2129
rect 38197 2083 38267 2129
rect 38313 2083 38383 2129
rect 38429 2083 38499 2129
rect 38545 2083 38615 2129
rect 38661 2083 38731 2129
rect 38777 2083 38847 2129
rect 38893 2083 38963 2129
rect 39009 2083 39079 2129
rect 39125 2083 39195 2129
rect 39241 2083 39311 2129
rect 39357 2083 39427 2129
rect 39473 2083 39543 2129
rect 39589 2083 39659 2129
rect 39705 2083 39775 2129
rect 39821 2083 39891 2129
rect 39937 2083 40007 2129
rect 40053 2083 40123 2129
rect 40169 2083 40180 2129
rect 28628 2013 40180 2083
rect 28628 1967 28639 2013
rect 28685 1967 28755 2013
rect 28801 1967 28871 2013
rect 28917 1967 28987 2013
rect 29033 1967 29103 2013
rect 29149 1967 29219 2013
rect 29265 1967 29335 2013
rect 29381 1967 29451 2013
rect 29497 1967 29567 2013
rect 29613 1967 29683 2013
rect 29729 1967 29799 2013
rect 29845 1967 29915 2013
rect 29961 1967 30031 2013
rect 30077 1967 30147 2013
rect 30193 1967 30263 2013
rect 30309 1967 30379 2013
rect 30425 1967 30495 2013
rect 30541 1967 30611 2013
rect 30657 1967 30727 2013
rect 30773 1967 30843 2013
rect 30889 1967 30959 2013
rect 31005 1967 31075 2013
rect 31121 1967 31191 2013
rect 31237 1967 31307 2013
rect 31353 1967 31423 2013
rect 31469 1967 31539 2013
rect 31585 1967 31655 2013
rect 31701 1967 31771 2013
rect 31817 1967 31887 2013
rect 31933 1967 32003 2013
rect 32049 1967 32119 2013
rect 32165 1967 32235 2013
rect 32281 1967 32351 2013
rect 32397 1967 32467 2013
rect 32513 1967 32583 2013
rect 32629 1967 32699 2013
rect 32745 1967 32815 2013
rect 32861 1967 32931 2013
rect 32977 1967 33047 2013
rect 33093 1967 33163 2013
rect 33209 1967 33279 2013
rect 33325 1967 33395 2013
rect 33441 1967 33511 2013
rect 33557 1967 33627 2013
rect 33673 1967 33743 2013
rect 33789 1967 33859 2013
rect 33905 1967 33975 2013
rect 34021 1967 34091 2013
rect 34137 1967 34207 2013
rect 34253 1967 34323 2013
rect 34369 1967 34439 2013
rect 34485 1967 34555 2013
rect 34601 1967 34671 2013
rect 34717 1967 34787 2013
rect 34833 1967 34903 2013
rect 34949 1967 35019 2013
rect 35065 1967 35135 2013
rect 35181 1967 35251 2013
rect 35297 1967 35367 2013
rect 35413 1967 35483 2013
rect 35529 1967 35599 2013
rect 35645 1967 35715 2013
rect 35761 1967 35831 2013
rect 35877 1967 35947 2013
rect 35993 1967 36063 2013
rect 36109 1967 36179 2013
rect 36225 1967 36295 2013
rect 36341 1967 36411 2013
rect 36457 1967 36527 2013
rect 36573 1967 36643 2013
rect 36689 1967 36759 2013
rect 36805 1967 36875 2013
rect 36921 1967 36991 2013
rect 37037 1967 37107 2013
rect 37153 1967 37223 2013
rect 37269 1967 37339 2013
rect 37385 1967 37455 2013
rect 37501 1967 37571 2013
rect 37617 1967 37687 2013
rect 37733 1967 37803 2013
rect 37849 1967 37919 2013
rect 37965 1967 38035 2013
rect 38081 1967 38151 2013
rect 38197 1967 38267 2013
rect 38313 1967 38383 2013
rect 38429 1967 38499 2013
rect 38545 1967 38615 2013
rect 38661 1967 38731 2013
rect 38777 1967 38847 2013
rect 38893 1967 38963 2013
rect 39009 1967 39079 2013
rect 39125 1967 39195 2013
rect 39241 1967 39311 2013
rect 39357 1967 39427 2013
rect 39473 1967 39543 2013
rect 39589 1967 39659 2013
rect 39705 1967 39775 2013
rect 39821 1967 39891 2013
rect 39937 1967 40007 2013
rect 40053 1967 40123 2013
rect 40169 1967 40180 2013
rect 28628 1925 40180 1967
rect 50834 3194 56586 3264
rect 50834 3148 50845 3194
rect 50891 3148 50961 3194
rect 51007 3148 51077 3194
rect 51123 3148 51193 3194
rect 51239 3148 51309 3194
rect 51355 3148 51425 3194
rect 51471 3148 51541 3194
rect 51587 3148 51657 3194
rect 51703 3148 51773 3194
rect 51819 3148 51889 3194
rect 51935 3148 52005 3194
rect 52051 3148 52121 3194
rect 52167 3148 52237 3194
rect 52283 3148 52353 3194
rect 52399 3148 52469 3194
rect 52515 3148 52585 3194
rect 52631 3148 52701 3194
rect 52747 3148 52817 3194
rect 52863 3148 52933 3194
rect 52979 3148 53049 3194
rect 53095 3148 53165 3194
rect 53211 3148 53281 3194
rect 53327 3148 53397 3194
rect 53443 3148 53513 3194
rect 53559 3148 53629 3194
rect 53675 3148 53745 3194
rect 53791 3148 53861 3194
rect 53907 3148 53977 3194
rect 54023 3148 54093 3194
rect 54139 3148 54209 3194
rect 54255 3148 54325 3194
rect 54371 3148 54441 3194
rect 54487 3148 54557 3194
rect 54603 3148 54673 3194
rect 54719 3148 54789 3194
rect 54835 3148 54905 3194
rect 54951 3148 55021 3194
rect 55067 3148 55137 3194
rect 55183 3148 55253 3194
rect 55299 3148 55369 3194
rect 55415 3148 55485 3194
rect 55531 3148 55601 3194
rect 55647 3148 55717 3194
rect 55763 3148 55833 3194
rect 55879 3148 55949 3194
rect 55995 3148 56065 3194
rect 56111 3148 56181 3194
rect 56227 3148 56297 3194
rect 56343 3148 56413 3194
rect 56459 3148 56529 3194
rect 56575 3148 56586 3194
rect 50834 3078 56586 3148
rect 50834 3032 50845 3078
rect 50891 3032 50961 3078
rect 51007 3032 51077 3078
rect 51123 3032 51193 3078
rect 51239 3032 51309 3078
rect 51355 3032 51425 3078
rect 51471 3032 51541 3078
rect 51587 3032 51657 3078
rect 51703 3032 51773 3078
rect 51819 3032 51889 3078
rect 51935 3032 52005 3078
rect 52051 3032 52121 3078
rect 52167 3032 52237 3078
rect 52283 3032 52353 3078
rect 52399 3032 52469 3078
rect 52515 3032 52585 3078
rect 52631 3032 52701 3078
rect 52747 3032 52817 3078
rect 52863 3032 52933 3078
rect 52979 3032 53049 3078
rect 53095 3032 53165 3078
rect 53211 3032 53281 3078
rect 53327 3032 53397 3078
rect 53443 3032 53513 3078
rect 53559 3032 53629 3078
rect 53675 3032 53745 3078
rect 53791 3032 53861 3078
rect 53907 3032 53977 3078
rect 54023 3032 54093 3078
rect 54139 3032 54209 3078
rect 54255 3032 54325 3078
rect 54371 3032 54441 3078
rect 54487 3032 54557 3078
rect 54603 3032 54673 3078
rect 54719 3032 54789 3078
rect 54835 3032 54905 3078
rect 54951 3032 55021 3078
rect 55067 3032 55137 3078
rect 55183 3032 55253 3078
rect 55299 3032 55369 3078
rect 55415 3032 55485 3078
rect 55531 3032 55601 3078
rect 55647 3032 55717 3078
rect 55763 3032 55833 3078
rect 55879 3032 55949 3078
rect 55995 3032 56065 3078
rect 56111 3032 56181 3078
rect 56227 3032 56297 3078
rect 56343 3032 56413 3078
rect 56459 3032 56529 3078
rect 56575 3032 56586 3078
rect 50834 2962 56586 3032
rect 50834 2916 50845 2962
rect 50891 2916 50961 2962
rect 51007 2916 51077 2962
rect 51123 2916 51193 2962
rect 51239 2916 51309 2962
rect 51355 2916 51425 2962
rect 51471 2916 51541 2962
rect 51587 2916 51657 2962
rect 51703 2916 51773 2962
rect 51819 2916 51889 2962
rect 51935 2916 52005 2962
rect 52051 2916 52121 2962
rect 52167 2916 52237 2962
rect 52283 2916 52353 2962
rect 52399 2916 52469 2962
rect 52515 2916 52585 2962
rect 52631 2916 52701 2962
rect 52747 2916 52817 2962
rect 52863 2916 52933 2962
rect 52979 2916 53049 2962
rect 53095 2916 53165 2962
rect 53211 2916 53281 2962
rect 53327 2916 53397 2962
rect 53443 2916 53513 2962
rect 53559 2916 53629 2962
rect 53675 2916 53745 2962
rect 53791 2916 53861 2962
rect 53907 2916 53977 2962
rect 54023 2916 54093 2962
rect 54139 2916 54209 2962
rect 54255 2916 54325 2962
rect 54371 2916 54441 2962
rect 54487 2916 54557 2962
rect 54603 2916 54673 2962
rect 54719 2916 54789 2962
rect 54835 2916 54905 2962
rect 54951 2916 55021 2962
rect 55067 2916 55137 2962
rect 55183 2916 55253 2962
rect 55299 2916 55369 2962
rect 55415 2916 55485 2962
rect 55531 2916 55601 2962
rect 55647 2916 55717 2962
rect 55763 2916 55833 2962
rect 55879 2916 55949 2962
rect 55995 2916 56065 2962
rect 56111 2916 56181 2962
rect 56227 2916 56297 2962
rect 56343 2916 56413 2962
rect 56459 2916 56529 2962
rect 56575 2916 56586 2962
rect 50834 2846 56586 2916
rect 50834 2800 50845 2846
rect 50891 2800 50961 2846
rect 51007 2800 51077 2846
rect 51123 2800 51193 2846
rect 51239 2800 51309 2846
rect 51355 2800 51425 2846
rect 51471 2800 51541 2846
rect 51587 2800 51657 2846
rect 51703 2800 51773 2846
rect 51819 2800 51889 2846
rect 51935 2800 52005 2846
rect 52051 2800 52121 2846
rect 52167 2800 52237 2846
rect 52283 2800 52353 2846
rect 52399 2800 52469 2846
rect 52515 2800 52585 2846
rect 52631 2800 52701 2846
rect 52747 2800 52817 2846
rect 52863 2800 52933 2846
rect 52979 2800 53049 2846
rect 53095 2800 53165 2846
rect 53211 2800 53281 2846
rect 53327 2800 53397 2846
rect 53443 2800 53513 2846
rect 53559 2800 53629 2846
rect 53675 2800 53745 2846
rect 53791 2800 53861 2846
rect 53907 2800 53977 2846
rect 54023 2800 54093 2846
rect 54139 2800 54209 2846
rect 54255 2800 54325 2846
rect 54371 2800 54441 2846
rect 54487 2800 54557 2846
rect 54603 2800 54673 2846
rect 54719 2800 54789 2846
rect 54835 2800 54905 2846
rect 54951 2800 55021 2846
rect 55067 2800 55137 2846
rect 55183 2800 55253 2846
rect 55299 2800 55369 2846
rect 55415 2800 55485 2846
rect 55531 2800 55601 2846
rect 55647 2800 55717 2846
rect 55763 2800 55833 2846
rect 55879 2800 55949 2846
rect 55995 2800 56065 2846
rect 56111 2800 56181 2846
rect 56227 2800 56297 2846
rect 56343 2800 56413 2846
rect 56459 2800 56529 2846
rect 56575 2800 56586 2846
rect 50834 2730 56586 2800
rect 50834 2684 50845 2730
rect 50891 2684 50961 2730
rect 51007 2684 51077 2730
rect 51123 2684 51193 2730
rect 51239 2684 51309 2730
rect 51355 2684 51425 2730
rect 51471 2684 51541 2730
rect 51587 2684 51657 2730
rect 51703 2684 51773 2730
rect 51819 2684 51889 2730
rect 51935 2684 52005 2730
rect 52051 2684 52121 2730
rect 52167 2684 52237 2730
rect 52283 2684 52353 2730
rect 52399 2684 52469 2730
rect 52515 2684 52585 2730
rect 52631 2684 52701 2730
rect 52747 2684 52817 2730
rect 52863 2684 52933 2730
rect 52979 2684 53049 2730
rect 53095 2684 53165 2730
rect 53211 2684 53281 2730
rect 53327 2684 53397 2730
rect 53443 2684 53513 2730
rect 53559 2684 53629 2730
rect 53675 2684 53745 2730
rect 53791 2684 53861 2730
rect 53907 2684 53977 2730
rect 54023 2684 54093 2730
rect 54139 2684 54209 2730
rect 54255 2684 54325 2730
rect 54371 2684 54441 2730
rect 54487 2684 54557 2730
rect 54603 2684 54673 2730
rect 54719 2684 54789 2730
rect 54835 2684 54905 2730
rect 54951 2684 55021 2730
rect 55067 2684 55137 2730
rect 55183 2684 55253 2730
rect 55299 2684 55369 2730
rect 55415 2684 55485 2730
rect 55531 2684 55601 2730
rect 55647 2684 55717 2730
rect 55763 2684 55833 2730
rect 55879 2684 55949 2730
rect 55995 2684 56065 2730
rect 56111 2684 56181 2730
rect 56227 2684 56297 2730
rect 56343 2684 56413 2730
rect 56459 2684 56529 2730
rect 56575 2684 56586 2730
rect 50834 2614 56586 2684
rect 50834 2568 50845 2614
rect 50891 2568 50961 2614
rect 51007 2568 51077 2614
rect 51123 2568 51193 2614
rect 51239 2568 51309 2614
rect 51355 2568 51425 2614
rect 51471 2568 51541 2614
rect 51587 2568 51657 2614
rect 51703 2568 51773 2614
rect 51819 2568 51889 2614
rect 51935 2568 52005 2614
rect 52051 2568 52121 2614
rect 52167 2568 52237 2614
rect 52283 2568 52353 2614
rect 52399 2568 52469 2614
rect 52515 2568 52585 2614
rect 52631 2568 52701 2614
rect 52747 2568 52817 2614
rect 52863 2568 52933 2614
rect 52979 2568 53049 2614
rect 53095 2568 53165 2614
rect 53211 2568 53281 2614
rect 53327 2568 53397 2614
rect 53443 2568 53513 2614
rect 53559 2568 53629 2614
rect 53675 2568 53745 2614
rect 53791 2568 53861 2614
rect 53907 2568 53977 2614
rect 54023 2568 54093 2614
rect 54139 2568 54209 2614
rect 54255 2568 54325 2614
rect 54371 2568 54441 2614
rect 54487 2568 54557 2614
rect 54603 2568 54673 2614
rect 54719 2568 54789 2614
rect 54835 2568 54905 2614
rect 54951 2568 55021 2614
rect 55067 2568 55137 2614
rect 55183 2568 55253 2614
rect 55299 2568 55369 2614
rect 55415 2568 55485 2614
rect 55531 2568 55601 2614
rect 55647 2568 55717 2614
rect 55763 2568 55833 2614
rect 55879 2568 55949 2614
rect 55995 2568 56065 2614
rect 56111 2568 56181 2614
rect 56227 2568 56297 2614
rect 56343 2568 56413 2614
rect 56459 2568 56529 2614
rect 56575 2568 56586 2614
rect 50834 2498 56586 2568
rect 50834 2452 50845 2498
rect 50891 2452 50961 2498
rect 51007 2452 51077 2498
rect 51123 2452 51193 2498
rect 51239 2452 51309 2498
rect 51355 2452 51425 2498
rect 51471 2452 51541 2498
rect 51587 2452 51657 2498
rect 51703 2452 51773 2498
rect 51819 2452 51889 2498
rect 51935 2452 52005 2498
rect 52051 2452 52121 2498
rect 52167 2452 52237 2498
rect 52283 2452 52353 2498
rect 52399 2452 52469 2498
rect 52515 2452 52585 2498
rect 52631 2452 52701 2498
rect 52747 2452 52817 2498
rect 52863 2452 52933 2498
rect 52979 2452 53049 2498
rect 53095 2452 53165 2498
rect 53211 2452 53281 2498
rect 53327 2452 53397 2498
rect 53443 2452 53513 2498
rect 53559 2452 53629 2498
rect 53675 2452 53745 2498
rect 53791 2452 53861 2498
rect 53907 2452 53977 2498
rect 54023 2452 54093 2498
rect 54139 2452 54209 2498
rect 54255 2452 54325 2498
rect 54371 2452 54441 2498
rect 54487 2452 54557 2498
rect 54603 2452 54673 2498
rect 54719 2452 54789 2498
rect 54835 2452 54905 2498
rect 54951 2452 55021 2498
rect 55067 2452 55137 2498
rect 55183 2452 55253 2498
rect 55299 2452 55369 2498
rect 55415 2452 55485 2498
rect 55531 2452 55601 2498
rect 55647 2452 55717 2498
rect 55763 2452 55833 2498
rect 55879 2452 55949 2498
rect 55995 2452 56065 2498
rect 56111 2452 56181 2498
rect 56227 2452 56297 2498
rect 56343 2452 56413 2498
rect 56459 2452 56529 2498
rect 56575 2452 56586 2498
rect 50834 2382 56586 2452
rect 50834 2336 50845 2382
rect 50891 2336 50961 2382
rect 51007 2336 51077 2382
rect 51123 2336 51193 2382
rect 51239 2336 51309 2382
rect 51355 2336 51425 2382
rect 51471 2336 51541 2382
rect 51587 2336 51657 2382
rect 51703 2336 51773 2382
rect 51819 2336 51889 2382
rect 51935 2336 52005 2382
rect 52051 2336 52121 2382
rect 52167 2336 52237 2382
rect 52283 2336 52353 2382
rect 52399 2336 52469 2382
rect 52515 2336 52585 2382
rect 52631 2336 52701 2382
rect 52747 2336 52817 2382
rect 52863 2336 52933 2382
rect 52979 2336 53049 2382
rect 53095 2336 53165 2382
rect 53211 2336 53281 2382
rect 53327 2336 53397 2382
rect 53443 2336 53513 2382
rect 53559 2336 53629 2382
rect 53675 2336 53745 2382
rect 53791 2336 53861 2382
rect 53907 2336 53977 2382
rect 54023 2336 54093 2382
rect 54139 2336 54209 2382
rect 54255 2336 54325 2382
rect 54371 2336 54441 2382
rect 54487 2336 54557 2382
rect 54603 2336 54673 2382
rect 54719 2336 54789 2382
rect 54835 2336 54905 2382
rect 54951 2336 55021 2382
rect 55067 2336 55137 2382
rect 55183 2336 55253 2382
rect 55299 2336 55369 2382
rect 55415 2336 55485 2382
rect 55531 2336 55601 2382
rect 55647 2336 55717 2382
rect 55763 2336 55833 2382
rect 55879 2336 55949 2382
rect 55995 2336 56065 2382
rect 56111 2336 56181 2382
rect 56227 2336 56297 2382
rect 56343 2336 56413 2382
rect 56459 2336 56529 2382
rect 56575 2336 56586 2382
rect 50834 2266 56586 2336
rect 50834 2220 50845 2266
rect 50891 2220 50961 2266
rect 51007 2220 51077 2266
rect 51123 2220 51193 2266
rect 51239 2220 51309 2266
rect 51355 2220 51425 2266
rect 51471 2220 51541 2266
rect 51587 2220 51657 2266
rect 51703 2220 51773 2266
rect 51819 2220 51889 2266
rect 51935 2220 52005 2266
rect 52051 2220 52121 2266
rect 52167 2220 52237 2266
rect 52283 2220 52353 2266
rect 52399 2220 52469 2266
rect 52515 2220 52585 2266
rect 52631 2220 52701 2266
rect 52747 2220 52817 2266
rect 52863 2220 52933 2266
rect 52979 2220 53049 2266
rect 53095 2220 53165 2266
rect 53211 2220 53281 2266
rect 53327 2220 53397 2266
rect 53443 2220 53513 2266
rect 53559 2220 53629 2266
rect 53675 2220 53745 2266
rect 53791 2220 53861 2266
rect 53907 2220 53977 2266
rect 54023 2220 54093 2266
rect 54139 2220 54209 2266
rect 54255 2220 54325 2266
rect 54371 2220 54441 2266
rect 54487 2220 54557 2266
rect 54603 2220 54673 2266
rect 54719 2220 54789 2266
rect 54835 2220 54905 2266
rect 54951 2220 55021 2266
rect 55067 2220 55137 2266
rect 55183 2220 55253 2266
rect 55299 2220 55369 2266
rect 55415 2220 55485 2266
rect 55531 2220 55601 2266
rect 55647 2220 55717 2266
rect 55763 2220 55833 2266
rect 55879 2220 55949 2266
rect 55995 2220 56065 2266
rect 56111 2220 56181 2266
rect 56227 2220 56297 2266
rect 56343 2220 56413 2266
rect 56459 2220 56529 2266
rect 56575 2220 56586 2266
rect 50834 2150 56586 2220
rect 50834 2104 50845 2150
rect 50891 2104 50961 2150
rect 51007 2104 51077 2150
rect 51123 2104 51193 2150
rect 51239 2104 51309 2150
rect 51355 2104 51425 2150
rect 51471 2104 51541 2150
rect 51587 2104 51657 2150
rect 51703 2104 51773 2150
rect 51819 2104 51889 2150
rect 51935 2104 52005 2150
rect 52051 2104 52121 2150
rect 52167 2104 52237 2150
rect 52283 2104 52353 2150
rect 52399 2104 52469 2150
rect 52515 2104 52585 2150
rect 52631 2104 52701 2150
rect 52747 2104 52817 2150
rect 52863 2104 52933 2150
rect 52979 2104 53049 2150
rect 53095 2104 53165 2150
rect 53211 2104 53281 2150
rect 53327 2104 53397 2150
rect 53443 2104 53513 2150
rect 53559 2104 53629 2150
rect 53675 2104 53745 2150
rect 53791 2104 53861 2150
rect 53907 2104 53977 2150
rect 54023 2104 54093 2150
rect 54139 2104 54209 2150
rect 54255 2104 54325 2150
rect 54371 2104 54441 2150
rect 54487 2104 54557 2150
rect 54603 2104 54673 2150
rect 54719 2104 54789 2150
rect 54835 2104 54905 2150
rect 54951 2104 55021 2150
rect 55067 2104 55137 2150
rect 55183 2104 55253 2150
rect 55299 2104 55369 2150
rect 55415 2104 55485 2150
rect 55531 2104 55601 2150
rect 55647 2104 55717 2150
rect 55763 2104 55833 2150
rect 55879 2104 55949 2150
rect 55995 2104 56065 2150
rect 56111 2104 56181 2150
rect 56227 2104 56297 2150
rect 56343 2104 56413 2150
rect 56459 2104 56529 2150
rect 56575 2104 56586 2150
rect 50834 2034 56586 2104
rect 50834 1988 50845 2034
rect 50891 1988 50961 2034
rect 51007 1988 51077 2034
rect 51123 1988 51193 2034
rect 51239 1988 51309 2034
rect 51355 1988 51425 2034
rect 51471 1988 51541 2034
rect 51587 1988 51657 2034
rect 51703 1988 51773 2034
rect 51819 1988 51889 2034
rect 51935 1988 52005 2034
rect 52051 1988 52121 2034
rect 52167 1988 52237 2034
rect 52283 1988 52353 2034
rect 52399 1988 52469 2034
rect 52515 1988 52585 2034
rect 52631 1988 52701 2034
rect 52747 1988 52817 2034
rect 52863 1988 52933 2034
rect 52979 1988 53049 2034
rect 53095 1988 53165 2034
rect 53211 1988 53281 2034
rect 53327 1988 53397 2034
rect 53443 1988 53513 2034
rect 53559 1988 53629 2034
rect 53675 1988 53745 2034
rect 53791 1988 53861 2034
rect 53907 1988 53977 2034
rect 54023 1988 54093 2034
rect 54139 1988 54209 2034
rect 54255 1988 54325 2034
rect 54371 1988 54441 2034
rect 54487 1988 54557 2034
rect 54603 1988 54673 2034
rect 54719 1988 54789 2034
rect 54835 1988 54905 2034
rect 54951 1988 55021 2034
rect 55067 1988 55137 2034
rect 55183 1988 55253 2034
rect 55299 1988 55369 2034
rect 55415 1988 55485 2034
rect 55531 1988 55601 2034
rect 55647 1988 55717 2034
rect 55763 1988 55833 2034
rect 55879 1988 55949 2034
rect 55995 1988 56065 2034
rect 56111 1988 56181 2034
rect 56227 1988 56297 2034
rect 56343 1988 56413 2034
rect 56459 1988 56529 2034
rect 56575 1988 56586 2034
rect 50834 1925 56586 1988
rect 57295 1925 57380 34245
rect 57626 45294 85733 45463
rect 57626 4587 57737 45294
rect 58790 44338 59517 45294
rect 58790 44286 58814 44338
rect 58866 44286 58938 44338
rect 58990 44286 59062 44338
rect 59114 44286 59186 44338
rect 59238 44286 59310 44338
rect 59362 44286 59434 44338
rect 59486 44286 59517 44338
rect 58790 44214 59517 44286
rect 58790 44162 58814 44214
rect 58866 44162 58938 44214
rect 58990 44162 59062 44214
rect 59114 44162 59186 44214
rect 59238 44162 59310 44214
rect 59362 44162 59434 44214
rect 59486 44162 59517 44214
rect 58790 44076 59517 44162
rect 84435 40526 84966 40726
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 84369 35126 85151 35326
rect 57909 33432 58351 33519
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33215 58351 33380
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 32997 58351 33163
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32779 58351 32945
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32562 58351 32727
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32344 58351 32510
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32075 57998 32127
rect 58050 32075 58210 32127
rect 58262 32075 58351 32127
rect 57909 31909 58351 32075
rect 83398 32048 83834 32122
rect 57909 31857 57998 31909
rect 58050 31857 58210 31909
rect 58262 31857 58351 31909
rect 57909 31691 58351 31857
rect 57909 31639 57998 31691
rect 58050 31639 58210 31691
rect 58262 31639 58351 31691
rect 57909 31474 58351 31639
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29950 58351 30116
rect 57909 29898 57998 29950
rect 58050 29898 58210 29950
rect 58262 29898 58351 29950
rect 57909 29733 58351 29898
rect 57909 29681 57998 29733
rect 58050 29681 58210 29733
rect 58262 29681 58351 29733
rect 57909 29515 58351 29681
rect 57909 29463 57998 29515
rect 58050 29463 58210 29515
rect 58262 29463 58351 29515
rect 57909 29297 58351 29463
rect 57909 29245 57998 29297
rect 58050 29245 58210 29297
rect 58262 29245 58351 29297
rect 57909 29080 58351 29245
rect 57909 29028 57998 29080
rect 58050 29028 58210 29080
rect 58262 29028 58351 29080
rect 57909 28862 58351 29028
rect 57909 28810 57998 28862
rect 58050 28810 58210 28862
rect 58262 28810 58351 28862
rect 57909 28644 58351 28810
rect 57909 28592 57998 28644
rect 58050 28592 58210 28644
rect 58262 28592 58351 28644
rect 57909 28427 58351 28592
rect 57909 28375 57998 28427
rect 58050 28375 58210 28427
rect 58262 28375 58351 28427
rect 57909 28209 58351 28375
rect 57909 28157 57998 28209
rect 58050 28157 58210 28209
rect 58262 28157 58351 28209
rect 57909 27992 58351 28157
rect 57909 27940 57998 27992
rect 58050 27940 58210 27992
rect 58262 27940 58351 27992
rect 57909 27774 58351 27940
rect 57909 27722 57998 27774
rect 58050 27722 58210 27774
rect 58262 27722 58351 27774
rect 57909 27556 58351 27722
rect 57909 27504 57998 27556
rect 58050 27504 58210 27556
rect 58262 27504 58351 27556
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24074 58351 24240
rect 57909 24022 57998 24074
rect 58050 24022 58210 24074
rect 58262 24022 58351 24074
rect 57909 23857 58351 24022
rect 57909 23805 57998 23857
rect 58050 23805 58210 23857
rect 58262 23805 58351 23857
rect 57909 23639 58351 23805
rect 57909 23587 57998 23639
rect 58050 23587 58210 23639
rect 58262 23587 58351 23639
rect 57909 23421 58351 23587
rect 57909 23369 57998 23421
rect 58050 23369 58210 23421
rect 58262 23369 58351 23421
rect 57909 23204 58351 23369
rect 57909 23152 57998 23204
rect 58050 23152 58210 23204
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20540 58210 20592
rect 58262 20540 58351 20592
rect 57909 20374 58351 20540
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20157 58351 20322
rect 57909 20105 57998 20157
rect 58050 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 19939 58351 20105
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13628 58351 13793
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13410 58351 13576
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13192 58351 13358
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 12975 58351 13140
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12757 58351 12923
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12540 58351 12705
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12322 58351 12488
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12104 58351 12270
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 11887 58351 12052
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11669 58351 11835
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9275 58351 9441
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9057 58351 9223
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8840 58351 9005
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8622 58351 8788
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8404 58351 8570
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8187 58351 8352
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5523 57998 5575
rect 58050 5523 58210 5575
rect 58262 5523 58351 5575
rect 57909 5358 58351 5523
rect 57909 5306 57998 5358
rect 58050 5306 58210 5358
rect 58262 5306 58351 5358
rect 57909 5220 58351 5306
rect 57647 4535 57737 4587
rect 57626 4370 57737 4535
rect 57647 4318 57737 4370
rect 57626 4152 57737 4318
rect 57647 4100 57737 4152
rect 57626 3934 57737 4100
rect 57647 3882 57737 3934
rect 57626 3717 57737 3882
rect 57647 3665 57737 3717
rect 27744 1918 57380 1925
rect 27744 1897 50845 1918
rect 27744 1851 28639 1897
rect 28685 1851 28755 1897
rect 28801 1851 28871 1897
rect 28917 1851 28987 1897
rect 29033 1851 29103 1897
rect 29149 1851 29219 1897
rect 29265 1851 29335 1897
rect 29381 1851 29451 1897
rect 29497 1851 29567 1897
rect 29613 1851 29683 1897
rect 29729 1851 29799 1897
rect 29845 1851 29915 1897
rect 29961 1851 30031 1897
rect 30077 1851 30147 1897
rect 30193 1851 30263 1897
rect 30309 1851 30379 1897
rect 30425 1851 30495 1897
rect 30541 1851 30611 1897
rect 30657 1851 30727 1897
rect 30773 1851 30843 1897
rect 30889 1851 30959 1897
rect 31005 1851 31075 1897
rect 31121 1851 31191 1897
rect 31237 1851 31307 1897
rect 31353 1851 31423 1897
rect 31469 1851 31539 1897
rect 31585 1851 31655 1897
rect 31701 1851 31771 1897
rect 31817 1851 31887 1897
rect 31933 1851 32003 1897
rect 32049 1851 32119 1897
rect 32165 1851 32235 1897
rect 32281 1851 32351 1897
rect 32397 1851 32467 1897
rect 32513 1851 32583 1897
rect 32629 1851 32699 1897
rect 32745 1851 32815 1897
rect 32861 1851 32931 1897
rect 32977 1851 33047 1897
rect 33093 1851 33163 1897
rect 33209 1851 33279 1897
rect 33325 1851 33395 1897
rect 33441 1851 33511 1897
rect 33557 1851 33627 1897
rect 33673 1851 33743 1897
rect 33789 1851 33859 1897
rect 33905 1851 33975 1897
rect 34021 1851 34091 1897
rect 34137 1851 34207 1897
rect 34253 1851 34323 1897
rect 34369 1851 34439 1897
rect 34485 1851 34555 1897
rect 34601 1851 34671 1897
rect 34717 1851 34787 1897
rect 34833 1851 34903 1897
rect 34949 1851 35019 1897
rect 35065 1851 35135 1897
rect 35181 1851 35251 1897
rect 35297 1851 35367 1897
rect 35413 1851 35483 1897
rect 35529 1851 35599 1897
rect 35645 1851 35715 1897
rect 35761 1851 35831 1897
rect 35877 1851 35947 1897
rect 35993 1851 36063 1897
rect 36109 1851 36179 1897
rect 36225 1851 36295 1897
rect 36341 1851 36411 1897
rect 36457 1851 36527 1897
rect 36573 1851 36643 1897
rect 36689 1851 36759 1897
rect 36805 1851 36875 1897
rect 36921 1851 36991 1897
rect 37037 1851 37107 1897
rect 37153 1851 37223 1897
rect 37269 1851 37339 1897
rect 37385 1851 37455 1897
rect 37501 1851 37571 1897
rect 37617 1851 37687 1897
rect 37733 1851 37803 1897
rect 37849 1851 37919 1897
rect 37965 1851 38035 1897
rect 38081 1851 38151 1897
rect 38197 1851 38267 1897
rect 38313 1851 38383 1897
rect 38429 1851 38499 1897
rect 38545 1851 38615 1897
rect 38661 1851 38731 1897
rect 38777 1851 38847 1897
rect 38893 1851 38963 1897
rect 39009 1851 39079 1897
rect 39125 1851 39195 1897
rect 39241 1851 39311 1897
rect 39357 1851 39427 1897
rect 39473 1851 39543 1897
rect 39589 1851 39659 1897
rect 39705 1851 39775 1897
rect 39821 1851 39891 1897
rect 39937 1851 40007 1897
rect 40053 1851 40123 1897
rect 40169 1872 50845 1897
rect 50891 1872 50961 1918
rect 51007 1872 51077 1918
rect 51123 1872 51193 1918
rect 51239 1872 51309 1918
rect 51355 1872 51425 1918
rect 51471 1872 51541 1918
rect 51587 1872 51657 1918
rect 51703 1872 51773 1918
rect 51819 1872 51889 1918
rect 51935 1872 52005 1918
rect 52051 1872 52121 1918
rect 52167 1872 52237 1918
rect 52283 1872 52353 1918
rect 52399 1872 52469 1918
rect 52515 1872 52585 1918
rect 52631 1872 52701 1918
rect 52747 1872 52817 1918
rect 52863 1872 52933 1918
rect 52979 1872 53049 1918
rect 53095 1872 53165 1918
rect 53211 1872 53281 1918
rect 53327 1872 53397 1918
rect 53443 1872 53513 1918
rect 53559 1872 53629 1918
rect 53675 1872 53745 1918
rect 53791 1872 53861 1918
rect 53907 1872 53977 1918
rect 54023 1872 54093 1918
rect 54139 1872 54209 1918
rect 54255 1872 54325 1918
rect 54371 1872 54441 1918
rect 54487 1872 54557 1918
rect 54603 1872 54673 1918
rect 54719 1872 54789 1918
rect 54835 1872 54905 1918
rect 54951 1872 55021 1918
rect 55067 1872 55137 1918
rect 55183 1872 55253 1918
rect 55299 1872 55369 1918
rect 55415 1872 55485 1918
rect 55531 1872 55601 1918
rect 55647 1872 55717 1918
rect 55763 1872 55833 1918
rect 55879 1872 55949 1918
rect 55995 1872 56065 1918
rect 56111 1872 56181 1918
rect 56227 1872 56297 1918
rect 56343 1872 56413 1918
rect 56459 1872 56529 1918
rect 56575 1872 57380 1918
rect 40169 1851 57380 1872
rect 27744 1802 57380 1851
rect 27744 1781 50845 1802
rect 27744 1735 28639 1781
rect 28685 1735 28755 1781
rect 28801 1735 28871 1781
rect 28917 1735 28987 1781
rect 29033 1735 29103 1781
rect 29149 1735 29219 1781
rect 29265 1735 29335 1781
rect 29381 1735 29451 1781
rect 29497 1735 29567 1781
rect 29613 1735 29683 1781
rect 29729 1735 29799 1781
rect 29845 1735 29915 1781
rect 29961 1735 30031 1781
rect 30077 1735 30147 1781
rect 30193 1735 30263 1781
rect 30309 1735 30379 1781
rect 30425 1735 30495 1781
rect 30541 1735 30611 1781
rect 30657 1735 30727 1781
rect 30773 1735 30843 1781
rect 30889 1735 30959 1781
rect 31005 1735 31075 1781
rect 31121 1735 31191 1781
rect 31237 1735 31307 1781
rect 31353 1735 31423 1781
rect 31469 1735 31539 1781
rect 31585 1735 31655 1781
rect 31701 1735 31771 1781
rect 31817 1735 31887 1781
rect 31933 1735 32003 1781
rect 32049 1735 32119 1781
rect 32165 1735 32235 1781
rect 32281 1735 32351 1781
rect 32397 1735 32467 1781
rect 32513 1735 32583 1781
rect 32629 1735 32699 1781
rect 32745 1735 32815 1781
rect 32861 1735 32931 1781
rect 32977 1735 33047 1781
rect 33093 1735 33163 1781
rect 33209 1735 33279 1781
rect 33325 1735 33395 1781
rect 33441 1735 33511 1781
rect 33557 1735 33627 1781
rect 33673 1735 33743 1781
rect 33789 1735 33859 1781
rect 33905 1735 33975 1781
rect 34021 1735 34091 1781
rect 34137 1735 34207 1781
rect 34253 1735 34323 1781
rect 34369 1735 34439 1781
rect 34485 1735 34555 1781
rect 34601 1735 34671 1781
rect 34717 1735 34787 1781
rect 34833 1735 34903 1781
rect 34949 1735 35019 1781
rect 35065 1735 35135 1781
rect 35181 1735 35251 1781
rect 35297 1735 35367 1781
rect 35413 1735 35483 1781
rect 35529 1735 35599 1781
rect 35645 1735 35715 1781
rect 35761 1735 35831 1781
rect 35877 1735 35947 1781
rect 35993 1735 36063 1781
rect 36109 1735 36179 1781
rect 36225 1735 36295 1781
rect 36341 1735 36411 1781
rect 36457 1735 36527 1781
rect 36573 1735 36643 1781
rect 36689 1735 36759 1781
rect 36805 1735 36875 1781
rect 36921 1735 36991 1781
rect 37037 1735 37107 1781
rect 37153 1735 37223 1781
rect 37269 1735 37339 1781
rect 37385 1735 37455 1781
rect 37501 1735 37571 1781
rect 37617 1735 37687 1781
rect 37733 1735 37803 1781
rect 37849 1735 37919 1781
rect 37965 1735 38035 1781
rect 38081 1735 38151 1781
rect 38197 1735 38267 1781
rect 38313 1735 38383 1781
rect 38429 1735 38499 1781
rect 38545 1735 38615 1781
rect 38661 1735 38731 1781
rect 38777 1735 38847 1781
rect 38893 1735 38963 1781
rect 39009 1735 39079 1781
rect 39125 1735 39195 1781
rect 39241 1735 39311 1781
rect 39357 1735 39427 1781
rect 39473 1735 39543 1781
rect 39589 1735 39659 1781
rect 39705 1735 39775 1781
rect 39821 1735 39891 1781
rect 39937 1735 40007 1781
rect 40053 1735 40123 1781
rect 40169 1756 50845 1781
rect 50891 1756 50961 1802
rect 51007 1756 51077 1802
rect 51123 1756 51193 1802
rect 51239 1756 51309 1802
rect 51355 1756 51425 1802
rect 51471 1756 51541 1802
rect 51587 1756 51657 1802
rect 51703 1756 51773 1802
rect 51819 1756 51889 1802
rect 51935 1756 52005 1802
rect 52051 1756 52121 1802
rect 52167 1756 52237 1802
rect 52283 1756 52353 1802
rect 52399 1756 52469 1802
rect 52515 1756 52585 1802
rect 52631 1756 52701 1802
rect 52747 1756 52817 1802
rect 52863 1756 52933 1802
rect 52979 1756 53049 1802
rect 53095 1756 53165 1802
rect 53211 1756 53281 1802
rect 53327 1756 53397 1802
rect 53443 1756 53513 1802
rect 53559 1756 53629 1802
rect 53675 1756 53745 1802
rect 53791 1756 53861 1802
rect 53907 1756 53977 1802
rect 54023 1756 54093 1802
rect 54139 1756 54209 1802
rect 54255 1756 54325 1802
rect 54371 1756 54441 1802
rect 54487 1756 54557 1802
rect 54603 1756 54673 1802
rect 54719 1756 54789 1802
rect 54835 1756 54905 1802
rect 54951 1756 55021 1802
rect 55067 1756 55137 1802
rect 55183 1756 55253 1802
rect 55299 1756 55369 1802
rect 55415 1756 55485 1802
rect 55531 1756 55601 1802
rect 55647 1756 55717 1802
rect 55763 1756 55833 1802
rect 55879 1756 55949 1802
rect 55995 1756 56065 1802
rect 56111 1756 56181 1802
rect 56227 1756 56297 1802
rect 56343 1756 56413 1802
rect 56459 1756 56529 1802
rect 56575 1756 57380 1802
rect 40169 1735 57380 1756
rect 27744 1686 57380 1735
rect 27744 1665 50845 1686
rect 27744 1619 28639 1665
rect 28685 1619 28755 1665
rect 28801 1619 28871 1665
rect 28917 1619 28987 1665
rect 29033 1619 29103 1665
rect 29149 1619 29219 1665
rect 29265 1619 29335 1665
rect 29381 1619 29451 1665
rect 29497 1619 29567 1665
rect 29613 1619 29683 1665
rect 29729 1619 29799 1665
rect 29845 1619 29915 1665
rect 29961 1619 30031 1665
rect 30077 1619 30147 1665
rect 30193 1619 30263 1665
rect 30309 1619 30379 1665
rect 30425 1619 30495 1665
rect 30541 1619 30611 1665
rect 30657 1619 30727 1665
rect 30773 1619 30843 1665
rect 30889 1619 30959 1665
rect 31005 1619 31075 1665
rect 31121 1619 31191 1665
rect 31237 1619 31307 1665
rect 31353 1619 31423 1665
rect 31469 1619 31539 1665
rect 31585 1619 31655 1665
rect 31701 1619 31771 1665
rect 31817 1619 31887 1665
rect 31933 1619 32003 1665
rect 32049 1619 32119 1665
rect 32165 1619 32235 1665
rect 32281 1619 32351 1665
rect 32397 1619 32467 1665
rect 32513 1619 32583 1665
rect 32629 1619 32699 1665
rect 32745 1619 32815 1665
rect 32861 1619 32931 1665
rect 32977 1619 33047 1665
rect 33093 1619 33163 1665
rect 33209 1619 33279 1665
rect 33325 1619 33395 1665
rect 33441 1619 33511 1665
rect 33557 1619 33627 1665
rect 33673 1619 33743 1665
rect 33789 1619 33859 1665
rect 33905 1619 33975 1665
rect 34021 1619 34091 1665
rect 34137 1619 34207 1665
rect 34253 1619 34323 1665
rect 34369 1619 34439 1665
rect 34485 1619 34555 1665
rect 34601 1619 34671 1665
rect 34717 1619 34787 1665
rect 34833 1619 34903 1665
rect 34949 1619 35019 1665
rect 35065 1619 35135 1665
rect 35181 1619 35251 1665
rect 35297 1619 35367 1665
rect 35413 1619 35483 1665
rect 35529 1619 35599 1665
rect 35645 1619 35715 1665
rect 35761 1619 35831 1665
rect 35877 1619 35947 1665
rect 35993 1619 36063 1665
rect 36109 1619 36179 1665
rect 36225 1619 36295 1665
rect 36341 1619 36411 1665
rect 36457 1619 36527 1665
rect 36573 1619 36643 1665
rect 36689 1619 36759 1665
rect 36805 1619 36875 1665
rect 36921 1619 36991 1665
rect 37037 1619 37107 1665
rect 37153 1619 37223 1665
rect 37269 1619 37339 1665
rect 37385 1619 37455 1665
rect 37501 1619 37571 1665
rect 37617 1619 37687 1665
rect 37733 1619 37803 1665
rect 37849 1619 37919 1665
rect 37965 1619 38035 1665
rect 38081 1619 38151 1665
rect 38197 1619 38267 1665
rect 38313 1619 38383 1665
rect 38429 1619 38499 1665
rect 38545 1619 38615 1665
rect 38661 1619 38731 1665
rect 38777 1619 38847 1665
rect 38893 1619 38963 1665
rect 39009 1619 39079 1665
rect 39125 1619 39195 1665
rect 39241 1619 39311 1665
rect 39357 1619 39427 1665
rect 39473 1619 39543 1665
rect 39589 1619 39659 1665
rect 39705 1619 39775 1665
rect 39821 1619 39891 1665
rect 39937 1619 40007 1665
rect 40053 1619 40123 1665
rect 40169 1640 50845 1665
rect 50891 1640 50961 1686
rect 51007 1640 51077 1686
rect 51123 1640 51193 1686
rect 51239 1640 51309 1686
rect 51355 1640 51425 1686
rect 51471 1640 51541 1686
rect 51587 1640 51657 1686
rect 51703 1640 51773 1686
rect 51819 1640 51889 1686
rect 51935 1640 52005 1686
rect 52051 1640 52121 1686
rect 52167 1640 52237 1686
rect 52283 1640 52353 1686
rect 52399 1640 52469 1686
rect 52515 1640 52585 1686
rect 52631 1640 52701 1686
rect 52747 1640 52817 1686
rect 52863 1640 52933 1686
rect 52979 1640 53049 1686
rect 53095 1640 53165 1686
rect 53211 1640 53281 1686
rect 53327 1640 53397 1686
rect 53443 1640 53513 1686
rect 53559 1640 53629 1686
rect 53675 1640 53745 1686
rect 53791 1640 53861 1686
rect 53907 1640 53977 1686
rect 54023 1640 54093 1686
rect 54139 1640 54209 1686
rect 54255 1640 54325 1686
rect 54371 1640 54441 1686
rect 54487 1640 54557 1686
rect 54603 1640 54673 1686
rect 54719 1640 54789 1686
rect 54835 1640 54905 1686
rect 54951 1640 55021 1686
rect 55067 1640 55137 1686
rect 55183 1640 55253 1686
rect 55299 1640 55369 1686
rect 55415 1640 55485 1686
rect 55531 1640 55601 1686
rect 55647 1640 55717 1686
rect 55763 1640 55833 1686
rect 55879 1640 55949 1686
rect 55995 1640 56065 1686
rect 56111 1640 56181 1686
rect 56227 1640 56297 1686
rect 56343 1640 56413 1686
rect 56459 1640 56529 1686
rect 56575 1640 57380 1686
rect 40169 1619 57380 1640
rect 27744 1570 57380 1619
rect 27744 1549 50845 1570
rect 27744 1503 28639 1549
rect 28685 1503 28755 1549
rect 28801 1503 28871 1549
rect 28917 1503 28987 1549
rect 29033 1503 29103 1549
rect 29149 1503 29219 1549
rect 29265 1503 29335 1549
rect 29381 1503 29451 1549
rect 29497 1503 29567 1549
rect 29613 1503 29683 1549
rect 29729 1503 29799 1549
rect 29845 1503 29915 1549
rect 29961 1503 30031 1549
rect 30077 1503 30147 1549
rect 30193 1503 30263 1549
rect 30309 1503 30379 1549
rect 30425 1503 30495 1549
rect 30541 1503 30611 1549
rect 30657 1503 30727 1549
rect 30773 1503 30843 1549
rect 30889 1503 30959 1549
rect 31005 1503 31075 1549
rect 31121 1503 31191 1549
rect 31237 1503 31307 1549
rect 31353 1503 31423 1549
rect 31469 1503 31539 1549
rect 31585 1503 31655 1549
rect 31701 1503 31771 1549
rect 31817 1503 31887 1549
rect 31933 1503 32003 1549
rect 32049 1503 32119 1549
rect 32165 1503 32235 1549
rect 32281 1503 32351 1549
rect 32397 1503 32467 1549
rect 32513 1503 32583 1549
rect 32629 1503 32699 1549
rect 32745 1503 32815 1549
rect 32861 1503 32931 1549
rect 32977 1503 33047 1549
rect 33093 1503 33163 1549
rect 33209 1503 33279 1549
rect 33325 1503 33395 1549
rect 33441 1503 33511 1549
rect 33557 1503 33627 1549
rect 33673 1503 33743 1549
rect 33789 1503 33859 1549
rect 33905 1503 33975 1549
rect 34021 1503 34091 1549
rect 34137 1503 34207 1549
rect 34253 1503 34323 1549
rect 34369 1503 34439 1549
rect 34485 1503 34555 1549
rect 34601 1503 34671 1549
rect 34717 1503 34787 1549
rect 34833 1503 34903 1549
rect 34949 1503 35019 1549
rect 35065 1503 35135 1549
rect 35181 1503 35251 1549
rect 35297 1503 35367 1549
rect 35413 1503 35483 1549
rect 35529 1503 35599 1549
rect 35645 1503 35715 1549
rect 35761 1503 35831 1549
rect 35877 1503 35947 1549
rect 35993 1503 36063 1549
rect 36109 1503 36179 1549
rect 36225 1503 36295 1549
rect 36341 1503 36411 1549
rect 36457 1503 36527 1549
rect 36573 1503 36643 1549
rect 36689 1503 36759 1549
rect 36805 1503 36875 1549
rect 36921 1503 36991 1549
rect 37037 1503 37107 1549
rect 37153 1503 37223 1549
rect 37269 1503 37339 1549
rect 37385 1503 37455 1549
rect 37501 1503 37571 1549
rect 37617 1503 37687 1549
rect 37733 1503 37803 1549
rect 37849 1503 37919 1549
rect 37965 1503 38035 1549
rect 38081 1503 38151 1549
rect 38197 1503 38267 1549
rect 38313 1503 38383 1549
rect 38429 1503 38499 1549
rect 38545 1503 38615 1549
rect 38661 1503 38731 1549
rect 38777 1503 38847 1549
rect 38893 1503 38963 1549
rect 39009 1503 39079 1549
rect 39125 1503 39195 1549
rect 39241 1503 39311 1549
rect 39357 1503 39427 1549
rect 39473 1503 39543 1549
rect 39589 1503 39659 1549
rect 39705 1503 39775 1549
rect 39821 1503 39891 1549
rect 39937 1503 40007 1549
rect 40053 1503 40123 1549
rect 40169 1524 50845 1549
rect 50891 1524 50961 1570
rect 51007 1524 51077 1570
rect 51123 1524 51193 1570
rect 51239 1524 51309 1570
rect 51355 1524 51425 1570
rect 51471 1524 51541 1570
rect 51587 1524 51657 1570
rect 51703 1524 51773 1570
rect 51819 1524 51889 1570
rect 51935 1524 52005 1570
rect 52051 1524 52121 1570
rect 52167 1524 52237 1570
rect 52283 1524 52353 1570
rect 52399 1524 52469 1570
rect 52515 1524 52585 1570
rect 52631 1524 52701 1570
rect 52747 1524 52817 1570
rect 52863 1524 52933 1570
rect 52979 1524 53049 1570
rect 53095 1524 53165 1570
rect 53211 1524 53281 1570
rect 53327 1524 53397 1570
rect 53443 1524 53513 1570
rect 53559 1524 53629 1570
rect 53675 1524 53745 1570
rect 53791 1524 53861 1570
rect 53907 1524 53977 1570
rect 54023 1524 54093 1570
rect 54139 1524 54209 1570
rect 54255 1524 54325 1570
rect 54371 1524 54441 1570
rect 54487 1524 54557 1570
rect 54603 1524 54673 1570
rect 54719 1524 54789 1570
rect 54835 1524 54905 1570
rect 54951 1524 55021 1570
rect 55067 1524 55137 1570
rect 55183 1524 55253 1570
rect 55299 1524 55369 1570
rect 55415 1524 55485 1570
rect 55531 1524 55601 1570
rect 55647 1524 55717 1570
rect 55763 1524 55833 1570
rect 55879 1524 55949 1570
rect 55995 1524 56065 1570
rect 56111 1524 56181 1570
rect 56227 1524 56297 1570
rect 56343 1524 56413 1570
rect 56459 1524 56529 1570
rect 56575 1524 57380 1570
rect 40169 1503 57380 1524
rect 27744 1454 57380 1503
rect 27744 1433 50845 1454
rect 27744 1387 28639 1433
rect 28685 1387 28755 1433
rect 28801 1387 28871 1433
rect 28917 1387 28987 1433
rect 29033 1387 29103 1433
rect 29149 1387 29219 1433
rect 29265 1387 29335 1433
rect 29381 1387 29451 1433
rect 29497 1387 29567 1433
rect 29613 1387 29683 1433
rect 29729 1387 29799 1433
rect 29845 1387 29915 1433
rect 29961 1387 30031 1433
rect 30077 1387 30147 1433
rect 30193 1387 30263 1433
rect 30309 1387 30379 1433
rect 30425 1387 30495 1433
rect 30541 1387 30611 1433
rect 30657 1387 30727 1433
rect 30773 1387 30843 1433
rect 30889 1387 30959 1433
rect 31005 1387 31075 1433
rect 31121 1387 31191 1433
rect 31237 1387 31307 1433
rect 31353 1387 31423 1433
rect 31469 1387 31539 1433
rect 31585 1387 31655 1433
rect 31701 1387 31771 1433
rect 31817 1387 31887 1433
rect 31933 1387 32003 1433
rect 32049 1387 32119 1433
rect 32165 1387 32235 1433
rect 32281 1387 32351 1433
rect 32397 1387 32467 1433
rect 32513 1387 32583 1433
rect 32629 1387 32699 1433
rect 32745 1387 32815 1433
rect 32861 1387 32931 1433
rect 32977 1387 33047 1433
rect 33093 1387 33163 1433
rect 33209 1387 33279 1433
rect 33325 1387 33395 1433
rect 33441 1387 33511 1433
rect 33557 1387 33627 1433
rect 33673 1387 33743 1433
rect 33789 1387 33859 1433
rect 33905 1387 33975 1433
rect 34021 1387 34091 1433
rect 34137 1387 34207 1433
rect 34253 1387 34323 1433
rect 34369 1387 34439 1433
rect 34485 1387 34555 1433
rect 34601 1387 34671 1433
rect 34717 1387 34787 1433
rect 34833 1387 34903 1433
rect 34949 1387 35019 1433
rect 35065 1387 35135 1433
rect 35181 1387 35251 1433
rect 35297 1387 35367 1433
rect 35413 1387 35483 1433
rect 35529 1387 35599 1433
rect 35645 1387 35715 1433
rect 35761 1387 35831 1433
rect 35877 1387 35947 1433
rect 35993 1387 36063 1433
rect 36109 1387 36179 1433
rect 36225 1387 36295 1433
rect 36341 1387 36411 1433
rect 36457 1387 36527 1433
rect 36573 1387 36643 1433
rect 36689 1387 36759 1433
rect 36805 1387 36875 1433
rect 36921 1387 36991 1433
rect 37037 1387 37107 1433
rect 37153 1387 37223 1433
rect 37269 1387 37339 1433
rect 37385 1387 37455 1433
rect 37501 1387 37571 1433
rect 37617 1387 37687 1433
rect 37733 1387 37803 1433
rect 37849 1387 37919 1433
rect 37965 1387 38035 1433
rect 38081 1387 38151 1433
rect 38197 1387 38267 1433
rect 38313 1387 38383 1433
rect 38429 1387 38499 1433
rect 38545 1387 38615 1433
rect 38661 1387 38731 1433
rect 38777 1387 38847 1433
rect 38893 1387 38963 1433
rect 39009 1387 39079 1433
rect 39125 1387 39195 1433
rect 39241 1387 39311 1433
rect 39357 1387 39427 1433
rect 39473 1387 39543 1433
rect 39589 1387 39659 1433
rect 39705 1387 39775 1433
rect 39821 1387 39891 1433
rect 39937 1387 40007 1433
rect 40053 1387 40123 1433
rect 40169 1408 50845 1433
rect 50891 1408 50961 1454
rect 51007 1408 51077 1454
rect 51123 1408 51193 1454
rect 51239 1408 51309 1454
rect 51355 1408 51425 1454
rect 51471 1408 51541 1454
rect 51587 1408 51657 1454
rect 51703 1408 51773 1454
rect 51819 1408 51889 1454
rect 51935 1408 52005 1454
rect 52051 1408 52121 1454
rect 52167 1408 52237 1454
rect 52283 1408 52353 1454
rect 52399 1408 52469 1454
rect 52515 1408 52585 1454
rect 52631 1408 52701 1454
rect 52747 1408 52817 1454
rect 52863 1408 52933 1454
rect 52979 1408 53049 1454
rect 53095 1408 53165 1454
rect 53211 1408 53281 1454
rect 53327 1408 53397 1454
rect 53443 1408 53513 1454
rect 53559 1408 53629 1454
rect 53675 1408 53745 1454
rect 53791 1408 53861 1454
rect 53907 1408 53977 1454
rect 54023 1408 54093 1454
rect 54139 1408 54209 1454
rect 54255 1408 54325 1454
rect 54371 1408 54441 1454
rect 54487 1408 54557 1454
rect 54603 1408 54673 1454
rect 54719 1408 54789 1454
rect 54835 1408 54905 1454
rect 54951 1408 55021 1454
rect 55067 1408 55137 1454
rect 55183 1408 55253 1454
rect 55299 1408 55369 1454
rect 55415 1408 55485 1454
rect 55531 1408 55601 1454
rect 55647 1408 55717 1454
rect 55763 1408 55833 1454
rect 55879 1408 55949 1454
rect 55995 1408 56065 1454
rect 56111 1408 56181 1454
rect 56227 1408 56297 1454
rect 56343 1408 56413 1454
rect 56459 1408 56529 1454
rect 56575 1408 57380 1454
rect 40169 1387 57380 1408
rect 27744 1338 57380 1387
rect 27744 1317 50845 1338
rect 27744 1271 28639 1317
rect 28685 1271 28755 1317
rect 28801 1271 28871 1317
rect 28917 1271 28987 1317
rect 29033 1271 29103 1317
rect 29149 1271 29219 1317
rect 29265 1271 29335 1317
rect 29381 1271 29451 1317
rect 29497 1271 29567 1317
rect 29613 1271 29683 1317
rect 29729 1271 29799 1317
rect 29845 1271 29915 1317
rect 29961 1271 30031 1317
rect 30077 1271 30147 1317
rect 30193 1271 30263 1317
rect 30309 1271 30379 1317
rect 30425 1271 30495 1317
rect 30541 1271 30611 1317
rect 30657 1271 30727 1317
rect 30773 1271 30843 1317
rect 30889 1271 30959 1317
rect 31005 1271 31075 1317
rect 31121 1271 31191 1317
rect 31237 1271 31307 1317
rect 31353 1271 31423 1317
rect 31469 1271 31539 1317
rect 31585 1271 31655 1317
rect 31701 1271 31771 1317
rect 31817 1271 31887 1317
rect 31933 1271 32003 1317
rect 32049 1271 32119 1317
rect 32165 1271 32235 1317
rect 32281 1271 32351 1317
rect 32397 1271 32467 1317
rect 32513 1271 32583 1317
rect 32629 1271 32699 1317
rect 32745 1271 32815 1317
rect 32861 1271 32931 1317
rect 32977 1271 33047 1317
rect 33093 1271 33163 1317
rect 33209 1271 33279 1317
rect 33325 1271 33395 1317
rect 33441 1271 33511 1317
rect 33557 1271 33627 1317
rect 33673 1271 33743 1317
rect 33789 1271 33859 1317
rect 33905 1271 33975 1317
rect 34021 1271 34091 1317
rect 34137 1271 34207 1317
rect 34253 1271 34323 1317
rect 34369 1271 34439 1317
rect 34485 1271 34555 1317
rect 34601 1271 34671 1317
rect 34717 1271 34787 1317
rect 34833 1271 34903 1317
rect 34949 1271 35019 1317
rect 35065 1271 35135 1317
rect 35181 1271 35251 1317
rect 35297 1271 35367 1317
rect 35413 1271 35483 1317
rect 35529 1271 35599 1317
rect 35645 1271 35715 1317
rect 35761 1271 35831 1317
rect 35877 1271 35947 1317
rect 35993 1271 36063 1317
rect 36109 1271 36179 1317
rect 36225 1271 36295 1317
rect 36341 1271 36411 1317
rect 36457 1271 36527 1317
rect 36573 1271 36643 1317
rect 36689 1271 36759 1317
rect 36805 1271 36875 1317
rect 36921 1271 36991 1317
rect 37037 1271 37107 1317
rect 37153 1271 37223 1317
rect 37269 1271 37339 1317
rect 37385 1271 37455 1317
rect 37501 1271 37571 1317
rect 37617 1271 37687 1317
rect 37733 1271 37803 1317
rect 37849 1271 37919 1317
rect 37965 1271 38035 1317
rect 38081 1271 38151 1317
rect 38197 1271 38267 1317
rect 38313 1271 38383 1317
rect 38429 1271 38499 1317
rect 38545 1271 38615 1317
rect 38661 1271 38731 1317
rect 38777 1271 38847 1317
rect 38893 1271 38963 1317
rect 39009 1271 39079 1317
rect 39125 1271 39195 1317
rect 39241 1271 39311 1317
rect 39357 1271 39427 1317
rect 39473 1271 39543 1317
rect 39589 1271 39659 1317
rect 39705 1271 39775 1317
rect 39821 1271 39891 1317
rect 39937 1271 40007 1317
rect 40053 1271 40123 1317
rect 40169 1292 50845 1317
rect 50891 1292 50961 1338
rect 51007 1292 51077 1338
rect 51123 1292 51193 1338
rect 51239 1292 51309 1338
rect 51355 1292 51425 1338
rect 51471 1292 51541 1338
rect 51587 1292 51657 1338
rect 51703 1292 51773 1338
rect 51819 1292 51889 1338
rect 51935 1292 52005 1338
rect 52051 1292 52121 1338
rect 52167 1292 52237 1338
rect 52283 1292 52353 1338
rect 52399 1292 52469 1338
rect 52515 1292 52585 1338
rect 52631 1292 52701 1338
rect 52747 1292 52817 1338
rect 52863 1292 52933 1338
rect 52979 1292 53049 1338
rect 53095 1292 53165 1338
rect 53211 1292 53281 1338
rect 53327 1292 53397 1338
rect 53443 1292 53513 1338
rect 53559 1292 53629 1338
rect 53675 1292 53745 1338
rect 53791 1292 53861 1338
rect 53907 1292 53977 1338
rect 54023 1292 54093 1338
rect 54139 1292 54209 1338
rect 54255 1292 54325 1338
rect 54371 1292 54441 1338
rect 54487 1292 54557 1338
rect 54603 1292 54673 1338
rect 54719 1292 54789 1338
rect 54835 1292 54905 1338
rect 54951 1292 55021 1338
rect 55067 1292 55137 1338
rect 55183 1292 55253 1338
rect 55299 1292 55369 1338
rect 55415 1292 55485 1338
rect 55531 1292 55601 1338
rect 55647 1292 55717 1338
rect 55763 1292 55833 1338
rect 55879 1292 55949 1338
rect 55995 1292 56065 1338
rect 56111 1292 56181 1338
rect 56227 1292 56297 1338
rect 56343 1292 56413 1338
rect 56459 1292 56529 1338
rect 56575 1292 57380 1338
rect 40169 1271 57380 1292
rect 27744 1222 57380 1271
rect 27744 1201 50845 1222
rect 27744 1155 28639 1201
rect 28685 1155 28755 1201
rect 28801 1155 28871 1201
rect 28917 1155 28987 1201
rect 29033 1155 29103 1201
rect 29149 1155 29219 1201
rect 29265 1155 29335 1201
rect 29381 1155 29451 1201
rect 29497 1155 29567 1201
rect 29613 1155 29683 1201
rect 29729 1155 29799 1201
rect 29845 1155 29915 1201
rect 29961 1155 30031 1201
rect 30077 1155 30147 1201
rect 30193 1155 30263 1201
rect 30309 1155 30379 1201
rect 30425 1155 30495 1201
rect 30541 1155 30611 1201
rect 30657 1155 30727 1201
rect 30773 1155 30843 1201
rect 30889 1155 30959 1201
rect 31005 1155 31075 1201
rect 31121 1155 31191 1201
rect 31237 1155 31307 1201
rect 31353 1155 31423 1201
rect 31469 1155 31539 1201
rect 31585 1155 31655 1201
rect 31701 1155 31771 1201
rect 31817 1155 31887 1201
rect 31933 1155 32003 1201
rect 32049 1155 32119 1201
rect 32165 1155 32235 1201
rect 32281 1155 32351 1201
rect 32397 1155 32467 1201
rect 32513 1155 32583 1201
rect 32629 1155 32699 1201
rect 32745 1155 32815 1201
rect 32861 1155 32931 1201
rect 32977 1155 33047 1201
rect 33093 1155 33163 1201
rect 33209 1155 33279 1201
rect 33325 1155 33395 1201
rect 33441 1155 33511 1201
rect 33557 1155 33627 1201
rect 33673 1155 33743 1201
rect 33789 1155 33859 1201
rect 33905 1155 33975 1201
rect 34021 1155 34091 1201
rect 34137 1155 34207 1201
rect 34253 1155 34323 1201
rect 34369 1155 34439 1201
rect 34485 1155 34555 1201
rect 34601 1155 34671 1201
rect 34717 1155 34787 1201
rect 34833 1155 34903 1201
rect 34949 1155 35019 1201
rect 35065 1155 35135 1201
rect 35181 1155 35251 1201
rect 35297 1155 35367 1201
rect 35413 1155 35483 1201
rect 35529 1155 35599 1201
rect 35645 1155 35715 1201
rect 35761 1155 35831 1201
rect 35877 1155 35947 1201
rect 35993 1155 36063 1201
rect 36109 1155 36179 1201
rect 36225 1155 36295 1201
rect 36341 1155 36411 1201
rect 36457 1155 36527 1201
rect 36573 1155 36643 1201
rect 36689 1155 36759 1201
rect 36805 1155 36875 1201
rect 36921 1155 36991 1201
rect 37037 1155 37107 1201
rect 37153 1155 37223 1201
rect 37269 1155 37339 1201
rect 37385 1155 37455 1201
rect 37501 1155 37571 1201
rect 37617 1155 37687 1201
rect 37733 1155 37803 1201
rect 37849 1155 37919 1201
rect 37965 1155 38035 1201
rect 38081 1155 38151 1201
rect 38197 1155 38267 1201
rect 38313 1155 38383 1201
rect 38429 1155 38499 1201
rect 38545 1155 38615 1201
rect 38661 1155 38731 1201
rect 38777 1155 38847 1201
rect 38893 1155 38963 1201
rect 39009 1155 39079 1201
rect 39125 1155 39195 1201
rect 39241 1155 39311 1201
rect 39357 1155 39427 1201
rect 39473 1155 39543 1201
rect 39589 1155 39659 1201
rect 39705 1155 39775 1201
rect 39821 1155 39891 1201
rect 39937 1155 40007 1201
rect 40053 1155 40123 1201
rect 40169 1176 50845 1201
rect 50891 1176 50961 1222
rect 51007 1176 51077 1222
rect 51123 1176 51193 1222
rect 51239 1176 51309 1222
rect 51355 1176 51425 1222
rect 51471 1176 51541 1222
rect 51587 1176 51657 1222
rect 51703 1176 51773 1222
rect 51819 1176 51889 1222
rect 51935 1176 52005 1222
rect 52051 1176 52121 1222
rect 52167 1176 52237 1222
rect 52283 1176 52353 1222
rect 52399 1176 52469 1222
rect 52515 1176 52585 1222
rect 52631 1176 52701 1222
rect 52747 1176 52817 1222
rect 52863 1176 52933 1222
rect 52979 1176 53049 1222
rect 53095 1176 53165 1222
rect 53211 1176 53281 1222
rect 53327 1176 53397 1222
rect 53443 1176 53513 1222
rect 53559 1176 53629 1222
rect 53675 1176 53745 1222
rect 53791 1176 53861 1222
rect 53907 1176 53977 1222
rect 54023 1176 54093 1222
rect 54139 1176 54209 1222
rect 54255 1176 54325 1222
rect 54371 1176 54441 1222
rect 54487 1176 54557 1222
rect 54603 1176 54673 1222
rect 54719 1176 54789 1222
rect 54835 1176 54905 1222
rect 54951 1176 55021 1222
rect 55067 1176 55137 1222
rect 55183 1176 55253 1222
rect 55299 1176 55369 1222
rect 55415 1176 55485 1222
rect 55531 1176 55601 1222
rect 55647 1176 55717 1222
rect 55763 1176 55833 1222
rect 55879 1176 55949 1222
rect 55995 1176 56065 1222
rect 56111 1176 56181 1222
rect 56227 1176 56297 1222
rect 56343 1176 56413 1222
rect 56459 1176 56529 1222
rect 56575 1176 57380 1222
rect 40169 1155 57380 1176
rect 27744 1117 57380 1155
rect 57626 1282 57737 3665
rect 57909 4587 58351 4728
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4370 58351 4535
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4152 58351 4318
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57909 1777 58351 3665
rect 62138 1689 62318 1701
rect 62138 1637 62150 1689
rect 62306 1637 62318 1689
rect 62138 1625 62318 1637
rect 72203 1689 72383 1701
rect 72203 1637 72215 1689
rect 72371 1637 72383 1689
rect 72203 1625 72383 1637
rect 72653 1689 72833 1701
rect 72653 1637 72665 1689
rect 72821 1637 72833 1689
rect 72653 1625 72833 1637
rect 82718 1689 82898 1701
rect 82718 1637 82730 1689
rect 82886 1637 82898 1689
rect 82718 1625 82898 1637
rect 85722 1282 85733 45294
rect 57626 1117 85733 1282
rect 86079 1117 86090 45563
rect 282 1023 86090 1117
rect 282 1015 48668 1023
rect 282 969 371 1015
rect 417 969 495 1015
rect 541 969 619 1015
rect 665 969 743 1015
rect 789 969 867 1015
rect 913 969 991 1015
rect 1037 969 1115 1015
rect 1161 969 1239 1015
rect 1285 969 1363 1015
rect 1409 969 1487 1015
rect 1533 969 1611 1015
rect 1657 969 1735 1015
rect 1781 969 1859 1015
rect 1905 969 1983 1015
rect 2029 969 2107 1015
rect 2153 969 2231 1015
rect 2277 969 2355 1015
rect 2401 969 2479 1015
rect 2525 969 2603 1015
rect 2649 969 2727 1015
rect 2773 969 2851 1015
rect 2897 969 2975 1015
rect 3021 969 3099 1015
rect 3145 969 3223 1015
rect 3269 969 3347 1015
rect 3393 969 3471 1015
rect 3517 969 3595 1015
rect 3641 969 3719 1015
rect 3765 969 3843 1015
rect 3889 969 3967 1015
rect 4013 969 4091 1015
rect 4137 969 4215 1015
rect 4261 969 4339 1015
rect 4385 969 4463 1015
rect 4509 969 4587 1015
rect 4633 969 4711 1015
rect 4757 969 4835 1015
rect 4881 969 4959 1015
rect 5005 969 5083 1015
rect 5129 969 5207 1015
rect 5253 969 5331 1015
rect 5377 969 5455 1015
rect 5501 969 5579 1015
rect 5625 969 5703 1015
rect 5749 969 5827 1015
rect 5873 969 5951 1015
rect 5997 969 6075 1015
rect 6121 969 6199 1015
rect 6245 969 6323 1015
rect 6369 969 6447 1015
rect 6493 969 6571 1015
rect 6617 969 6695 1015
rect 6741 969 6819 1015
rect 6865 969 6943 1015
rect 6989 969 7067 1015
rect 7113 969 7191 1015
rect 7237 969 7315 1015
rect 7361 969 7439 1015
rect 7485 969 7563 1015
rect 7609 969 7687 1015
rect 7733 969 7811 1015
rect 7857 969 7935 1015
rect 7981 969 8059 1015
rect 8105 969 8183 1015
rect 8229 969 8307 1015
rect 8353 969 8431 1015
rect 8477 969 8555 1015
rect 8601 969 8679 1015
rect 8725 969 8803 1015
rect 8849 969 8927 1015
rect 8973 969 9051 1015
rect 9097 969 9175 1015
rect 9221 969 9299 1015
rect 9345 969 9423 1015
rect 9469 969 9547 1015
rect 9593 969 9671 1015
rect 9717 969 9795 1015
rect 9841 969 9919 1015
rect 9965 969 10043 1015
rect 10089 969 10167 1015
rect 10213 969 10291 1015
rect 10337 969 10415 1015
rect 10461 969 10539 1015
rect 10585 969 10663 1015
rect 10709 969 10787 1015
rect 10833 969 10911 1015
rect 10957 969 11035 1015
rect 11081 969 11159 1015
rect 11205 969 11283 1015
rect 11329 969 11407 1015
rect 11453 969 11531 1015
rect 11577 969 11655 1015
rect 11701 969 11779 1015
rect 11825 969 11903 1015
rect 11949 969 12027 1015
rect 12073 969 12151 1015
rect 12197 969 12275 1015
rect 12321 969 12399 1015
rect 12445 969 12523 1015
rect 12569 969 12647 1015
rect 12693 969 12771 1015
rect 12817 969 12895 1015
rect 12941 969 13019 1015
rect 13065 969 13143 1015
rect 13189 969 13267 1015
rect 13313 969 13391 1015
rect 13437 969 13515 1015
rect 13561 969 13639 1015
rect 13685 969 13763 1015
rect 13809 969 13887 1015
rect 13933 969 14011 1015
rect 14057 969 14135 1015
rect 14181 969 14259 1015
rect 14305 969 14383 1015
rect 14429 969 14507 1015
rect 14553 969 14631 1015
rect 14677 969 14755 1015
rect 14801 969 14879 1015
rect 14925 969 15003 1015
rect 15049 969 15127 1015
rect 15173 969 15251 1015
rect 15297 969 15375 1015
rect 15421 969 15499 1015
rect 15545 969 15623 1015
rect 15669 969 15747 1015
rect 15793 969 15871 1015
rect 15917 969 15995 1015
rect 16041 969 16119 1015
rect 16165 969 16243 1015
rect 16289 969 16367 1015
rect 16413 969 16491 1015
rect 16537 969 16615 1015
rect 16661 969 16739 1015
rect 16785 969 16863 1015
rect 16909 969 16987 1015
rect 17033 969 17111 1015
rect 17157 969 17235 1015
rect 17281 969 17359 1015
rect 17405 969 17483 1015
rect 17529 969 17607 1015
rect 17653 969 17731 1015
rect 17777 969 17855 1015
rect 17901 969 17979 1015
rect 18025 969 18103 1015
rect 18149 969 18227 1015
rect 18273 969 18351 1015
rect 18397 969 18475 1015
rect 18521 969 18599 1015
rect 18645 969 18723 1015
rect 18769 969 18847 1015
rect 18893 969 18971 1015
rect 19017 969 19095 1015
rect 19141 969 19219 1015
rect 19265 969 19343 1015
rect 19389 969 19467 1015
rect 19513 969 19591 1015
rect 19637 969 19715 1015
rect 19761 969 19839 1015
rect 19885 969 19963 1015
rect 20009 969 20087 1015
rect 20133 969 20211 1015
rect 20257 969 20335 1015
rect 20381 969 20459 1015
rect 20505 969 20583 1015
rect 20629 969 20707 1015
rect 20753 969 20831 1015
rect 20877 969 20955 1015
rect 21001 969 21079 1015
rect 21125 969 21203 1015
rect 21249 969 21327 1015
rect 21373 969 21451 1015
rect 21497 969 21575 1015
rect 21621 969 21699 1015
rect 21745 969 21823 1015
rect 21869 969 21947 1015
rect 21993 969 22071 1015
rect 22117 969 22195 1015
rect 22241 969 22319 1015
rect 22365 969 22443 1015
rect 22489 969 22567 1015
rect 22613 969 22691 1015
rect 22737 969 22815 1015
rect 22861 969 22939 1015
rect 22985 969 23063 1015
rect 23109 969 23187 1015
rect 23233 969 23311 1015
rect 23357 969 23435 1015
rect 23481 969 23559 1015
rect 23605 969 23683 1015
rect 23729 969 23807 1015
rect 23853 969 23931 1015
rect 23977 969 24055 1015
rect 24101 969 24179 1015
rect 24225 969 24303 1015
rect 24349 969 24427 1015
rect 24473 969 24551 1015
rect 24597 969 24675 1015
rect 24721 969 24799 1015
rect 24845 969 24923 1015
rect 24969 969 25047 1015
rect 25093 969 25171 1015
rect 25217 969 25295 1015
rect 25341 969 25419 1015
rect 25465 969 25543 1015
rect 25589 969 25667 1015
rect 25713 969 25791 1015
rect 25837 969 25915 1015
rect 25961 969 26039 1015
rect 26085 969 26163 1015
rect 26209 969 26287 1015
rect 26333 969 26411 1015
rect 26457 969 26535 1015
rect 26581 969 26659 1015
rect 26705 969 26783 1015
rect 26829 969 26907 1015
rect 26953 969 27031 1015
rect 27077 969 27155 1015
rect 27201 969 27279 1015
rect 27325 969 27403 1015
rect 27449 969 27527 1015
rect 27573 969 27651 1015
rect 27697 969 27775 1015
rect 27821 969 27899 1015
rect 27945 969 28023 1015
rect 28069 969 28147 1015
rect 28193 969 28271 1015
rect 28317 969 28395 1015
rect 28441 969 28519 1015
rect 28565 969 28643 1015
rect 28689 969 28767 1015
rect 28813 969 28891 1015
rect 28937 969 29015 1015
rect 29061 969 29139 1015
rect 29185 969 29263 1015
rect 29309 969 29387 1015
rect 29433 969 29511 1015
rect 29557 969 29635 1015
rect 29681 969 29759 1015
rect 29805 969 29883 1015
rect 29929 969 30007 1015
rect 30053 969 30131 1015
rect 30177 969 30255 1015
rect 30301 969 30379 1015
rect 30425 969 30503 1015
rect 30549 969 30627 1015
rect 30673 969 30751 1015
rect 30797 969 30875 1015
rect 30921 969 30999 1015
rect 31045 969 31123 1015
rect 31169 969 31247 1015
rect 31293 969 31371 1015
rect 31417 969 31495 1015
rect 31541 969 31619 1015
rect 31665 969 31743 1015
rect 31789 969 31867 1015
rect 31913 969 31991 1015
rect 32037 969 32115 1015
rect 32161 969 32239 1015
rect 32285 969 32363 1015
rect 32409 969 32487 1015
rect 32533 969 32611 1015
rect 32657 969 32735 1015
rect 32781 969 32859 1015
rect 32905 969 32983 1015
rect 33029 969 33107 1015
rect 33153 969 33231 1015
rect 33277 969 33355 1015
rect 33401 969 33479 1015
rect 33525 969 33603 1015
rect 33649 969 33727 1015
rect 33773 969 33851 1015
rect 33897 969 33975 1015
rect 34021 969 34099 1015
rect 34145 969 34223 1015
rect 34269 969 34347 1015
rect 34393 969 34471 1015
rect 34517 969 34595 1015
rect 34641 969 34719 1015
rect 34765 969 34843 1015
rect 34889 969 34967 1015
rect 35013 969 35091 1015
rect 35137 969 35215 1015
rect 35261 969 35339 1015
rect 35385 969 35463 1015
rect 35509 969 35587 1015
rect 35633 969 35711 1015
rect 35757 969 35835 1015
rect 35881 969 35959 1015
rect 36005 969 36083 1015
rect 36129 969 36207 1015
rect 36253 969 36331 1015
rect 36377 969 36455 1015
rect 36501 969 36579 1015
rect 36625 969 36703 1015
rect 36749 969 36827 1015
rect 36873 969 36951 1015
rect 36997 969 37075 1015
rect 37121 969 37199 1015
rect 37245 969 37323 1015
rect 37369 969 37447 1015
rect 37493 969 37571 1015
rect 37617 969 37695 1015
rect 37741 969 37819 1015
rect 37865 969 37943 1015
rect 37989 969 38067 1015
rect 38113 969 38191 1015
rect 38237 969 38315 1015
rect 38361 969 38439 1015
rect 38485 969 38563 1015
rect 38609 969 38687 1015
rect 38733 969 38811 1015
rect 38857 969 38935 1015
rect 38981 969 39059 1015
rect 39105 969 39183 1015
rect 39229 969 39307 1015
rect 39353 969 39431 1015
rect 39477 969 39555 1015
rect 39601 969 39679 1015
rect 39725 969 39803 1015
rect 39849 969 39927 1015
rect 39973 969 40051 1015
rect 40097 969 40175 1015
rect 40221 969 40299 1015
rect 40345 969 40423 1015
rect 40469 969 40547 1015
rect 40593 969 40671 1015
rect 40717 969 40795 1015
rect 40841 969 40919 1015
rect 40965 969 41043 1015
rect 41089 969 41167 1015
rect 41213 969 41291 1015
rect 41337 969 41415 1015
rect 41461 969 41539 1015
rect 41585 969 41663 1015
rect 41709 969 41787 1015
rect 41833 969 41911 1015
rect 41957 969 42035 1015
rect 42081 969 42159 1015
rect 42205 969 42283 1015
rect 42329 969 42407 1015
rect 42453 969 42531 1015
rect 42577 969 42655 1015
rect 42701 969 42779 1015
rect 42825 969 42903 1015
rect 42949 969 43027 1015
rect 43073 969 43151 1015
rect 43197 969 43275 1015
rect 43321 969 43399 1015
rect 43445 969 43523 1015
rect 43569 969 43647 1015
rect 43693 969 43771 1015
rect 43817 969 43895 1015
rect 43941 969 44019 1015
rect 44065 969 44143 1015
rect 44189 969 44267 1015
rect 44313 969 44391 1015
rect 44437 969 44515 1015
rect 44561 969 44639 1015
rect 44685 969 44763 1015
rect 44809 969 44887 1015
rect 44933 969 45011 1015
rect 45057 969 45135 1015
rect 45181 969 45259 1015
rect 45305 969 45383 1015
rect 45429 969 45507 1015
rect 45553 969 45631 1015
rect 45677 969 45755 1015
rect 45801 969 45879 1015
rect 45925 969 46003 1015
rect 46049 969 46127 1015
rect 46173 969 46251 1015
rect 46297 969 46375 1015
rect 46421 969 46499 1015
rect 46545 969 46623 1015
rect 46669 969 46747 1015
rect 46793 969 46871 1015
rect 46917 969 46995 1015
rect 47041 969 47119 1015
rect 47165 969 47243 1015
rect 47289 969 47367 1015
rect 47413 969 47491 1015
rect 47537 969 47615 1015
rect 47661 969 47739 1015
rect 47785 969 47863 1015
rect 47909 969 47987 1015
rect 48033 969 48111 1015
rect 48157 969 48235 1015
rect 48281 969 48359 1015
rect 48405 969 48483 1015
rect 48529 969 48607 1015
rect 48653 971 48668 1015
rect 48720 1015 48792 1023
rect 48720 971 48731 1015
rect 48653 969 48731 971
rect 48777 971 48792 1015
rect 48844 1015 48916 1023
rect 48844 971 48855 1015
rect 48777 969 48855 971
rect 48901 971 48916 1015
rect 48968 1015 86090 1023
rect 48968 971 48979 1015
rect 48901 969 48979 971
rect 49025 969 49103 1015
rect 49149 969 49227 1015
rect 49273 969 49351 1015
rect 49397 969 49475 1015
rect 49521 969 49599 1015
rect 49645 969 49723 1015
rect 49769 969 49847 1015
rect 49893 969 49971 1015
rect 50017 969 50095 1015
rect 50141 969 50219 1015
rect 50265 969 50343 1015
rect 50389 969 50467 1015
rect 50513 969 50591 1015
rect 50637 969 50715 1015
rect 50761 969 50839 1015
rect 50885 969 50963 1015
rect 51009 969 51087 1015
rect 51133 969 51211 1015
rect 51257 969 51335 1015
rect 51381 969 51459 1015
rect 51505 969 51583 1015
rect 51629 969 51707 1015
rect 51753 969 51831 1015
rect 51877 969 51955 1015
rect 52001 969 52079 1015
rect 52125 969 52203 1015
rect 52249 969 52327 1015
rect 52373 969 52451 1015
rect 52497 969 52575 1015
rect 52621 969 52699 1015
rect 52745 969 52823 1015
rect 52869 969 52947 1015
rect 52993 969 53071 1015
rect 53117 969 53195 1015
rect 53241 969 53319 1015
rect 53365 969 53443 1015
rect 53489 969 53567 1015
rect 53613 969 53691 1015
rect 53737 969 53815 1015
rect 53861 1006 53939 1015
rect 53861 969 53907 1006
rect 53985 969 54063 1015
rect 54109 969 54187 1015
rect 54233 969 54311 1015
rect 54357 969 54435 1015
rect 54481 969 54559 1015
rect 54605 969 54683 1015
rect 54729 969 54807 1015
rect 54853 969 54931 1015
rect 54977 969 55055 1015
rect 55101 969 55179 1015
rect 55225 969 55303 1015
rect 55349 969 55427 1015
rect 55473 969 55551 1015
rect 55597 969 55675 1015
rect 55721 969 55799 1015
rect 55845 969 55923 1015
rect 55969 969 56047 1015
rect 56093 969 56171 1015
rect 56217 969 56295 1015
rect 56341 969 56419 1015
rect 56465 969 56543 1015
rect 56589 969 56667 1015
rect 56713 969 56791 1015
rect 56837 969 56915 1015
rect 56961 969 57039 1015
rect 57085 969 57163 1015
rect 57209 969 57287 1015
rect 57333 969 57411 1015
rect 57457 969 57535 1015
rect 57581 969 57659 1015
rect 57705 969 57783 1015
rect 57829 969 57907 1015
rect 57953 969 58031 1015
rect 58077 969 58155 1015
rect 58201 969 58279 1015
rect 58325 969 58403 1015
rect 58449 969 58527 1015
rect 58573 969 58651 1015
rect 58697 969 58775 1015
rect 58821 969 58899 1015
rect 58945 969 59023 1015
rect 59069 969 59147 1015
rect 59193 969 59271 1015
rect 59317 969 59395 1015
rect 59441 969 59519 1015
rect 59565 969 59643 1015
rect 59689 969 59767 1015
rect 59813 969 59891 1015
rect 59937 969 60015 1015
rect 60061 969 60139 1015
rect 60185 969 60263 1015
rect 60309 969 60387 1015
rect 60433 969 60511 1015
rect 60557 969 60635 1015
rect 60681 969 60759 1015
rect 60805 969 60883 1015
rect 60929 969 61007 1015
rect 61053 969 61131 1015
rect 61177 969 61255 1015
rect 61301 969 61379 1015
rect 61425 969 61503 1015
rect 61549 969 61627 1015
rect 61673 969 61751 1015
rect 61797 969 61875 1015
rect 61921 969 61999 1015
rect 62045 969 62123 1015
rect 62169 969 62247 1015
rect 62293 969 62371 1015
rect 62417 969 62495 1015
rect 62541 969 62619 1015
rect 62665 969 62743 1015
rect 62789 969 62867 1015
rect 62913 969 62991 1015
rect 63037 969 63115 1015
rect 63161 969 63239 1015
rect 63285 969 63363 1015
rect 63409 969 63487 1015
rect 63533 969 63611 1015
rect 63657 969 63735 1015
rect 63781 969 63859 1015
rect 63905 969 63983 1015
rect 64029 969 64107 1015
rect 64153 969 64231 1015
rect 64277 969 64355 1015
rect 64401 969 64479 1015
rect 64525 969 64603 1015
rect 64649 969 64727 1015
rect 64773 969 64851 1015
rect 64897 969 64975 1015
rect 65021 969 65099 1015
rect 65145 969 65223 1015
rect 65269 969 65347 1015
rect 65393 969 65471 1015
rect 65517 969 65595 1015
rect 65641 969 65719 1015
rect 65765 969 65843 1015
rect 65889 969 65967 1015
rect 66013 969 66091 1015
rect 66137 969 66215 1015
rect 66261 969 66339 1015
rect 66385 969 66463 1015
rect 66509 969 66587 1015
rect 66633 969 66711 1015
rect 66757 969 66835 1015
rect 66881 969 66959 1015
rect 67005 969 67083 1015
rect 67129 969 67207 1015
rect 67253 969 67331 1015
rect 67377 969 67455 1015
rect 67501 969 67579 1015
rect 67625 969 67703 1015
rect 67749 969 67827 1015
rect 67873 969 67951 1015
rect 67997 969 68075 1015
rect 68121 969 68199 1015
rect 68245 969 68323 1015
rect 68369 969 68447 1015
rect 68493 969 68571 1015
rect 68617 969 68695 1015
rect 68741 969 68819 1015
rect 68865 969 68943 1015
rect 68989 969 69067 1015
rect 69113 969 69191 1015
rect 69237 969 69315 1015
rect 69361 969 69439 1015
rect 69485 969 69563 1015
rect 69609 969 69687 1015
rect 69733 969 69811 1015
rect 69857 969 69935 1015
rect 69981 969 70059 1015
rect 70105 969 70183 1015
rect 70229 969 70307 1015
rect 70353 969 70431 1015
rect 70477 969 70555 1015
rect 70601 969 70679 1015
rect 70725 969 70803 1015
rect 70849 969 70927 1015
rect 70973 969 71051 1015
rect 71097 969 71175 1015
rect 71221 969 71299 1015
rect 71345 969 71423 1015
rect 71469 969 71547 1015
rect 71593 969 71671 1015
rect 71717 969 71795 1015
rect 71841 969 71919 1015
rect 71965 969 72043 1015
rect 72089 969 72167 1015
rect 72213 969 72291 1015
rect 72337 969 72415 1015
rect 72461 969 72539 1015
rect 72585 969 72663 1015
rect 72709 969 72787 1015
rect 72833 969 72911 1015
rect 72957 969 73035 1015
rect 73081 969 73159 1015
rect 73205 969 73283 1015
rect 73329 969 73407 1015
rect 73453 969 73531 1015
rect 73577 969 73655 1015
rect 73701 969 73779 1015
rect 73825 969 73903 1015
rect 73949 969 74027 1015
rect 74073 969 74151 1015
rect 74197 969 74275 1015
rect 74321 969 74399 1015
rect 74445 969 74523 1015
rect 74569 969 74647 1015
rect 74693 969 74771 1015
rect 74817 969 74895 1015
rect 74941 969 75019 1015
rect 75065 969 75143 1015
rect 75189 969 75267 1015
rect 75313 969 75391 1015
rect 75437 969 75515 1015
rect 75561 969 75639 1015
rect 75685 969 75763 1015
rect 75809 969 75887 1015
rect 75933 969 76011 1015
rect 76057 969 76135 1015
rect 76181 969 76259 1015
rect 76305 969 76383 1015
rect 76429 969 76507 1015
rect 76553 969 76631 1015
rect 76677 969 76755 1015
rect 76801 969 76879 1015
rect 76925 969 77003 1015
rect 77049 969 77127 1015
rect 77173 969 77251 1015
rect 77297 969 77375 1015
rect 77421 969 77499 1015
rect 77545 969 77623 1015
rect 77669 969 77747 1015
rect 77793 969 77871 1015
rect 77917 969 77995 1015
rect 78041 969 78119 1015
rect 78165 969 78243 1015
rect 78289 969 78367 1015
rect 78413 969 78491 1015
rect 78537 969 78615 1015
rect 78661 969 78739 1015
rect 78785 969 78863 1015
rect 78909 969 78987 1015
rect 79033 969 79111 1015
rect 79157 969 79235 1015
rect 79281 969 79359 1015
rect 79405 969 79483 1015
rect 79529 969 79607 1015
rect 79653 969 79731 1015
rect 79777 969 79855 1015
rect 79901 969 79979 1015
rect 80025 969 80103 1015
rect 80149 969 80227 1015
rect 80273 969 80351 1015
rect 80397 969 80475 1015
rect 80521 969 80599 1015
rect 80645 969 80723 1015
rect 80769 969 80847 1015
rect 80893 969 80971 1015
rect 81017 969 81095 1015
rect 81141 969 81219 1015
rect 81265 969 81343 1015
rect 81389 969 81467 1015
rect 81513 969 81591 1015
rect 81637 969 81715 1015
rect 81761 969 81839 1015
rect 81885 969 81963 1015
rect 82009 969 82087 1015
rect 82133 969 82211 1015
rect 82257 969 82335 1015
rect 82381 969 82459 1015
rect 82505 969 82583 1015
rect 82629 969 82707 1015
rect 82753 969 82831 1015
rect 82877 969 82955 1015
rect 83001 969 83079 1015
rect 83125 969 83203 1015
rect 83249 969 83327 1015
rect 83373 969 83451 1015
rect 83497 969 83575 1015
rect 83621 969 83699 1015
rect 83745 969 83823 1015
rect 83869 969 83947 1015
rect 83993 969 84071 1015
rect 84117 969 84195 1015
rect 84241 969 84319 1015
rect 84365 969 84443 1015
rect 84489 969 84567 1015
rect 84613 969 84691 1015
rect 84737 969 84815 1015
rect 84861 969 84939 1015
rect 84985 969 85063 1015
rect 85109 969 85187 1015
rect 85233 969 85311 1015
rect 85357 969 85435 1015
rect 85481 969 85559 1015
rect 85605 969 85683 1015
rect 85729 969 85807 1015
rect 85853 969 85931 1015
rect 85977 969 86090 1015
rect 282 914 53907 969
rect 282 891 29090 914
rect 29142 891 29787 914
rect 29839 899 53907 914
rect 29839 891 48668 899
rect 282 845 371 891
rect 417 845 495 891
rect 541 845 619 891
rect 665 845 743 891
rect 789 845 867 891
rect 913 845 991 891
rect 1037 845 1115 891
rect 1161 845 1239 891
rect 1285 845 1363 891
rect 1409 845 1487 891
rect 1533 845 1611 891
rect 1657 845 1735 891
rect 1781 845 1859 891
rect 1905 845 1983 891
rect 2029 845 2107 891
rect 2153 845 2231 891
rect 2277 845 2355 891
rect 2401 845 2479 891
rect 2525 845 2603 891
rect 2649 845 2727 891
rect 2773 845 2851 891
rect 2897 845 2975 891
rect 3021 845 3099 891
rect 3145 845 3223 891
rect 3269 845 3347 891
rect 3393 845 3471 891
rect 3517 845 3595 891
rect 3641 845 3719 891
rect 3765 845 3843 891
rect 3889 845 3967 891
rect 4013 845 4091 891
rect 4137 845 4215 891
rect 4261 845 4339 891
rect 4385 845 4463 891
rect 4509 845 4587 891
rect 4633 845 4711 891
rect 4757 845 4835 891
rect 4881 845 4959 891
rect 5005 845 5083 891
rect 5129 845 5207 891
rect 5253 845 5331 891
rect 5377 845 5455 891
rect 5501 845 5579 891
rect 5625 845 5703 891
rect 5749 845 5827 891
rect 5873 845 5951 891
rect 5997 845 6075 891
rect 6121 845 6199 891
rect 6245 845 6323 891
rect 6369 845 6447 891
rect 6493 845 6571 891
rect 6617 845 6695 891
rect 6741 845 6819 891
rect 6865 845 6943 891
rect 6989 845 7067 891
rect 7113 845 7191 891
rect 7237 845 7315 891
rect 7361 845 7439 891
rect 7485 845 7563 891
rect 7609 845 7687 891
rect 7733 845 7811 891
rect 7857 845 7935 891
rect 7981 845 8059 891
rect 8105 845 8183 891
rect 8229 845 8307 891
rect 8353 845 8431 891
rect 8477 845 8555 891
rect 8601 845 8679 891
rect 8725 845 8803 891
rect 8849 845 8927 891
rect 8973 845 9051 891
rect 9097 845 9175 891
rect 9221 845 9299 891
rect 9345 845 9423 891
rect 9469 845 9547 891
rect 9593 845 9671 891
rect 9717 845 9795 891
rect 9841 845 9919 891
rect 9965 845 10043 891
rect 10089 845 10167 891
rect 10213 845 10291 891
rect 10337 845 10415 891
rect 10461 845 10539 891
rect 10585 845 10663 891
rect 10709 845 10787 891
rect 10833 845 10911 891
rect 10957 845 11035 891
rect 11081 845 11159 891
rect 11205 845 11283 891
rect 11329 845 11407 891
rect 11453 845 11531 891
rect 11577 845 11655 891
rect 11701 845 11779 891
rect 11825 845 11903 891
rect 11949 845 12027 891
rect 12073 845 12151 891
rect 12197 845 12275 891
rect 12321 845 12399 891
rect 12445 845 12523 891
rect 12569 845 12647 891
rect 12693 845 12771 891
rect 12817 845 12895 891
rect 12941 845 13019 891
rect 13065 845 13143 891
rect 13189 845 13267 891
rect 13313 845 13391 891
rect 13437 845 13515 891
rect 13561 845 13639 891
rect 13685 845 13763 891
rect 13809 845 13887 891
rect 13933 845 14011 891
rect 14057 845 14135 891
rect 14181 845 14259 891
rect 14305 845 14383 891
rect 14429 845 14507 891
rect 14553 845 14631 891
rect 14677 845 14755 891
rect 14801 845 14879 891
rect 14925 845 15003 891
rect 15049 845 15127 891
rect 15173 845 15251 891
rect 15297 845 15375 891
rect 15421 845 15499 891
rect 15545 845 15623 891
rect 15669 845 15747 891
rect 15793 845 15871 891
rect 15917 845 15995 891
rect 16041 845 16119 891
rect 16165 845 16243 891
rect 16289 845 16367 891
rect 16413 845 16491 891
rect 16537 845 16615 891
rect 16661 845 16739 891
rect 16785 845 16863 891
rect 16909 845 16987 891
rect 17033 845 17111 891
rect 17157 845 17235 891
rect 17281 845 17359 891
rect 17405 845 17483 891
rect 17529 845 17607 891
rect 17653 845 17731 891
rect 17777 845 17855 891
rect 17901 845 17979 891
rect 18025 845 18103 891
rect 18149 845 18227 891
rect 18273 845 18351 891
rect 18397 845 18475 891
rect 18521 845 18599 891
rect 18645 845 18723 891
rect 18769 845 18847 891
rect 18893 845 18971 891
rect 19017 845 19095 891
rect 19141 845 19219 891
rect 19265 845 19343 891
rect 19389 845 19467 891
rect 19513 845 19591 891
rect 19637 845 19715 891
rect 19761 845 19839 891
rect 19885 845 19963 891
rect 20009 845 20087 891
rect 20133 845 20211 891
rect 20257 845 20335 891
rect 20381 845 20459 891
rect 20505 845 20583 891
rect 20629 845 20707 891
rect 20753 845 20831 891
rect 20877 845 20955 891
rect 21001 845 21079 891
rect 21125 845 21203 891
rect 21249 845 21327 891
rect 21373 845 21451 891
rect 21497 845 21575 891
rect 21621 845 21699 891
rect 21745 845 21823 891
rect 21869 845 21947 891
rect 21993 845 22071 891
rect 22117 845 22195 891
rect 22241 845 22319 891
rect 22365 845 22443 891
rect 22489 845 22567 891
rect 22613 845 22691 891
rect 22737 845 22815 891
rect 22861 845 22939 891
rect 22985 845 23063 891
rect 23109 845 23187 891
rect 23233 845 23311 891
rect 23357 845 23435 891
rect 23481 845 23559 891
rect 23605 845 23683 891
rect 23729 845 23807 891
rect 23853 845 23931 891
rect 23977 845 24055 891
rect 24101 845 24179 891
rect 24225 845 24303 891
rect 24349 845 24427 891
rect 24473 845 24551 891
rect 24597 845 24675 891
rect 24721 845 24799 891
rect 24845 845 24923 891
rect 24969 845 25047 891
rect 25093 845 25171 891
rect 25217 845 25295 891
rect 25341 845 25419 891
rect 25465 845 25543 891
rect 25589 845 25667 891
rect 25713 845 25791 891
rect 25837 845 25915 891
rect 25961 845 26039 891
rect 26085 845 26163 891
rect 26209 845 26287 891
rect 26333 845 26411 891
rect 26457 845 26535 891
rect 26581 845 26659 891
rect 26705 845 26783 891
rect 26829 845 26907 891
rect 26953 845 27031 891
rect 27077 845 27155 891
rect 27201 845 27279 891
rect 27325 845 27403 891
rect 27449 845 27527 891
rect 27573 845 27651 891
rect 27697 845 27775 891
rect 27821 845 27899 891
rect 27945 845 28023 891
rect 28069 845 28147 891
rect 28193 845 28271 891
rect 28317 845 28395 891
rect 28441 845 28519 891
rect 28565 845 28643 891
rect 28689 845 28767 891
rect 28813 845 28891 891
rect 28937 845 29015 891
rect 29061 845 29090 891
rect 29185 845 29263 891
rect 29309 845 29387 891
rect 29433 845 29511 891
rect 29557 845 29635 891
rect 29681 845 29759 891
rect 29839 845 29883 891
rect 29929 845 30007 891
rect 30053 845 30131 891
rect 30177 845 30255 891
rect 30301 845 30379 891
rect 30425 845 30503 891
rect 30549 845 30627 891
rect 30673 845 30751 891
rect 30797 845 30875 891
rect 30921 845 30999 891
rect 31045 845 31123 891
rect 31169 845 31247 891
rect 31293 845 31371 891
rect 31417 845 31495 891
rect 31541 845 31619 891
rect 31665 845 31743 891
rect 31789 845 31867 891
rect 31913 845 31991 891
rect 32037 845 32115 891
rect 32161 845 32239 891
rect 32285 845 32363 891
rect 32409 845 32487 891
rect 32533 845 32611 891
rect 32657 845 32735 891
rect 32781 845 32859 891
rect 32905 845 32983 891
rect 33029 845 33107 891
rect 33153 845 33231 891
rect 33277 845 33355 891
rect 33401 845 33479 891
rect 33525 845 33603 891
rect 33649 845 33727 891
rect 33773 845 33851 891
rect 33897 845 33975 891
rect 34021 845 34099 891
rect 34145 845 34223 891
rect 34269 845 34347 891
rect 34393 845 34471 891
rect 34517 845 34595 891
rect 34641 845 34719 891
rect 34765 845 34843 891
rect 34889 845 34967 891
rect 35013 845 35091 891
rect 35137 845 35215 891
rect 35261 845 35339 891
rect 35385 845 35463 891
rect 35509 845 35587 891
rect 35633 845 35711 891
rect 35757 845 35835 891
rect 35881 845 35959 891
rect 36005 845 36083 891
rect 36129 845 36207 891
rect 36253 845 36331 891
rect 36377 845 36455 891
rect 36501 845 36579 891
rect 36625 845 36703 891
rect 36749 845 36827 891
rect 36873 845 36951 891
rect 36997 845 37075 891
rect 37121 845 37199 891
rect 37245 845 37323 891
rect 37369 845 37447 891
rect 37493 845 37571 891
rect 37617 845 37695 891
rect 37741 845 37819 891
rect 37865 845 37943 891
rect 37989 845 38067 891
rect 38113 845 38191 891
rect 38237 845 38315 891
rect 38361 845 38439 891
rect 38485 845 38563 891
rect 38609 845 38687 891
rect 38733 845 38811 891
rect 38857 845 38935 891
rect 38981 845 39059 891
rect 39105 845 39183 891
rect 39229 845 39307 891
rect 39353 845 39431 891
rect 39477 845 39555 891
rect 39601 845 39679 891
rect 39725 845 39803 891
rect 39849 845 39927 891
rect 39973 845 40051 891
rect 40097 845 40175 891
rect 40221 845 40299 891
rect 40345 845 40423 891
rect 40469 845 40547 891
rect 40593 845 40671 891
rect 40717 845 40795 891
rect 40841 845 40919 891
rect 40965 845 41043 891
rect 41089 845 41167 891
rect 41213 845 41291 891
rect 41337 845 41415 891
rect 41461 845 41539 891
rect 41585 845 41663 891
rect 41709 845 41787 891
rect 41833 845 41911 891
rect 41957 845 42035 891
rect 42081 845 42159 891
rect 42205 845 42283 891
rect 42329 845 42407 891
rect 42453 845 42531 891
rect 42577 845 42655 891
rect 42701 845 42779 891
rect 42825 845 42903 891
rect 42949 845 43027 891
rect 43073 845 43151 891
rect 43197 845 43275 891
rect 43321 845 43399 891
rect 43445 845 43523 891
rect 43569 845 43647 891
rect 43693 845 43771 891
rect 43817 845 43895 891
rect 43941 845 44019 891
rect 44065 845 44143 891
rect 44189 845 44267 891
rect 44313 845 44391 891
rect 44437 845 44515 891
rect 44561 845 44639 891
rect 44685 845 44763 891
rect 44809 845 44887 891
rect 44933 845 45011 891
rect 45057 845 45135 891
rect 45181 845 45259 891
rect 45305 845 45383 891
rect 45429 845 45507 891
rect 45553 845 45631 891
rect 45677 845 45755 891
rect 45801 845 45879 891
rect 45925 845 46003 891
rect 46049 845 46127 891
rect 46173 845 46251 891
rect 46297 845 46375 891
rect 46421 845 46499 891
rect 46545 845 46623 891
rect 46669 845 46747 891
rect 46793 845 46871 891
rect 46917 845 46995 891
rect 47041 845 47119 891
rect 47165 845 47243 891
rect 47289 845 47367 891
rect 47413 845 47491 891
rect 47537 845 47615 891
rect 47661 845 47739 891
rect 47785 845 47863 891
rect 47909 845 47987 891
rect 48033 845 48111 891
rect 48157 845 48235 891
rect 48281 845 48359 891
rect 48405 845 48483 891
rect 48529 845 48607 891
rect 48653 847 48668 891
rect 48720 891 48792 899
rect 48720 847 48731 891
rect 48653 845 48731 847
rect 48777 847 48792 891
rect 48844 891 48916 899
rect 48844 847 48855 891
rect 48777 845 48855 847
rect 48901 847 48916 891
rect 48968 891 53907 899
rect 53959 891 86090 969
rect 48968 847 48979 891
rect 48901 845 48979 847
rect 49025 845 49103 891
rect 49149 845 49227 891
rect 49273 845 49351 891
rect 49397 845 49475 891
rect 49521 845 49599 891
rect 49645 845 49723 891
rect 49769 845 49847 891
rect 49893 845 49971 891
rect 50017 845 50095 891
rect 50141 845 50219 891
rect 50265 845 50343 891
rect 50389 845 50467 891
rect 50513 845 50591 891
rect 50637 845 50715 891
rect 50761 845 50839 891
rect 50885 845 50963 891
rect 51009 845 51087 891
rect 51133 845 51211 891
rect 51257 845 51335 891
rect 51381 845 51459 891
rect 51505 845 51583 891
rect 51629 845 51707 891
rect 51753 845 51831 891
rect 51877 845 51955 891
rect 52001 845 52079 891
rect 52125 845 52203 891
rect 52249 845 52327 891
rect 52373 845 52451 891
rect 52497 845 52575 891
rect 52621 845 52699 891
rect 52745 845 52823 891
rect 52869 845 52947 891
rect 52993 845 53071 891
rect 53117 845 53195 891
rect 53241 845 53319 891
rect 53365 845 53443 891
rect 53489 845 53567 891
rect 53613 845 53691 891
rect 53737 845 53815 891
rect 53861 845 53907 891
rect 53985 845 54063 891
rect 54109 845 54187 891
rect 54233 845 54311 891
rect 54357 845 54435 891
rect 54481 845 54559 891
rect 54605 845 54683 891
rect 54729 845 54807 891
rect 54853 845 54931 891
rect 54977 845 55055 891
rect 55101 845 55179 891
rect 55225 845 55303 891
rect 55349 845 55427 891
rect 55473 845 55551 891
rect 55597 845 55675 891
rect 55721 845 55799 891
rect 55845 845 55923 891
rect 55969 845 56047 891
rect 56093 845 56171 891
rect 56217 845 56295 891
rect 56341 845 56419 891
rect 56465 845 56543 891
rect 56589 845 56667 891
rect 56713 845 56791 891
rect 56837 845 56915 891
rect 56961 845 57039 891
rect 57085 845 57163 891
rect 57209 845 57287 891
rect 57333 845 57411 891
rect 57457 845 57535 891
rect 57581 845 57659 891
rect 57705 845 57783 891
rect 57829 845 57907 891
rect 57953 845 58031 891
rect 58077 845 58155 891
rect 58201 845 58279 891
rect 58325 845 58403 891
rect 58449 845 58527 891
rect 58573 845 58651 891
rect 58697 845 58775 891
rect 58821 845 58899 891
rect 58945 845 59023 891
rect 59069 845 59147 891
rect 59193 845 59271 891
rect 59317 845 59395 891
rect 59441 845 59519 891
rect 59565 845 59643 891
rect 59689 845 59767 891
rect 59813 845 59891 891
rect 59937 845 60015 891
rect 60061 845 60139 891
rect 60185 845 60263 891
rect 60309 845 60387 891
rect 60433 845 60511 891
rect 60557 845 60635 891
rect 60681 845 60759 891
rect 60805 845 60883 891
rect 60929 845 61007 891
rect 61053 845 61131 891
rect 61177 845 61255 891
rect 61301 845 61379 891
rect 61425 845 61503 891
rect 61549 845 61627 891
rect 61673 845 61751 891
rect 61797 845 61875 891
rect 61921 845 61999 891
rect 62045 845 62123 891
rect 62169 845 62247 891
rect 62293 845 62371 891
rect 62417 845 62495 891
rect 62541 845 62619 891
rect 62665 845 62743 891
rect 62789 845 62867 891
rect 62913 845 62991 891
rect 63037 845 63115 891
rect 63161 845 63239 891
rect 63285 845 63363 891
rect 63409 845 63487 891
rect 63533 845 63611 891
rect 63657 845 63735 891
rect 63781 845 63859 891
rect 63905 845 63983 891
rect 64029 845 64107 891
rect 64153 845 64231 891
rect 64277 845 64355 891
rect 64401 845 64479 891
rect 64525 845 64603 891
rect 64649 845 64727 891
rect 64773 845 64851 891
rect 64897 845 64975 891
rect 65021 845 65099 891
rect 65145 845 65223 891
rect 65269 845 65347 891
rect 65393 845 65471 891
rect 65517 845 65595 891
rect 65641 845 65719 891
rect 65765 845 65843 891
rect 65889 845 65967 891
rect 66013 845 66091 891
rect 66137 845 66215 891
rect 66261 845 66339 891
rect 66385 845 66463 891
rect 66509 845 66587 891
rect 66633 845 66711 891
rect 66757 845 66835 891
rect 66881 845 66959 891
rect 67005 845 67083 891
rect 67129 845 67207 891
rect 67253 845 67331 891
rect 67377 845 67455 891
rect 67501 845 67579 891
rect 67625 845 67703 891
rect 67749 845 67827 891
rect 67873 845 67951 891
rect 67997 845 68075 891
rect 68121 845 68199 891
rect 68245 845 68323 891
rect 68369 845 68447 891
rect 68493 845 68571 891
rect 68617 845 68695 891
rect 68741 845 68819 891
rect 68865 845 68943 891
rect 68989 845 69067 891
rect 69113 845 69191 891
rect 69237 845 69315 891
rect 69361 845 69439 891
rect 69485 845 69563 891
rect 69609 845 69687 891
rect 69733 845 69811 891
rect 69857 845 69935 891
rect 69981 845 70059 891
rect 70105 845 70183 891
rect 70229 845 70307 891
rect 70353 845 70431 891
rect 70477 845 70555 891
rect 70601 845 70679 891
rect 70725 845 70803 891
rect 70849 845 70927 891
rect 70973 845 71051 891
rect 71097 845 71175 891
rect 71221 845 71299 891
rect 71345 845 71423 891
rect 71469 845 71547 891
rect 71593 845 71671 891
rect 71717 845 71795 891
rect 71841 845 71919 891
rect 71965 845 72043 891
rect 72089 845 72167 891
rect 72213 845 72291 891
rect 72337 845 72415 891
rect 72461 845 72539 891
rect 72585 845 72663 891
rect 72709 845 72787 891
rect 72833 845 72911 891
rect 72957 845 73035 891
rect 73081 845 73159 891
rect 73205 845 73283 891
rect 73329 845 73407 891
rect 73453 845 73531 891
rect 73577 845 73655 891
rect 73701 845 73779 891
rect 73825 845 73903 891
rect 73949 845 74027 891
rect 74073 845 74151 891
rect 74197 845 74275 891
rect 74321 845 74399 891
rect 74445 845 74523 891
rect 74569 845 74647 891
rect 74693 845 74771 891
rect 74817 845 74895 891
rect 74941 845 75019 891
rect 75065 845 75143 891
rect 75189 845 75267 891
rect 75313 845 75391 891
rect 75437 845 75515 891
rect 75561 845 75639 891
rect 75685 845 75763 891
rect 75809 845 75887 891
rect 75933 845 76011 891
rect 76057 845 76135 891
rect 76181 845 76259 891
rect 76305 845 76383 891
rect 76429 845 76507 891
rect 76553 845 76631 891
rect 76677 845 76755 891
rect 76801 845 76879 891
rect 76925 845 77003 891
rect 77049 845 77127 891
rect 77173 845 77251 891
rect 77297 845 77375 891
rect 77421 845 77499 891
rect 77545 845 77623 891
rect 77669 845 77747 891
rect 77793 845 77871 891
rect 77917 845 77995 891
rect 78041 845 78119 891
rect 78165 845 78243 891
rect 78289 845 78367 891
rect 78413 845 78491 891
rect 78537 845 78615 891
rect 78661 845 78739 891
rect 78785 845 78863 891
rect 78909 845 78987 891
rect 79033 845 79111 891
rect 79157 845 79235 891
rect 79281 845 79359 891
rect 79405 845 79483 891
rect 79529 845 79607 891
rect 79653 845 79731 891
rect 79777 845 79855 891
rect 79901 845 79979 891
rect 80025 845 80103 891
rect 80149 845 80227 891
rect 80273 845 80351 891
rect 80397 845 80475 891
rect 80521 845 80599 891
rect 80645 845 80723 891
rect 80769 845 80847 891
rect 80893 845 80971 891
rect 81017 845 81095 891
rect 81141 845 81219 891
rect 81265 845 81343 891
rect 81389 845 81467 891
rect 81513 845 81591 891
rect 81637 845 81715 891
rect 81761 845 81839 891
rect 81885 845 81963 891
rect 82009 845 82087 891
rect 82133 845 82211 891
rect 82257 845 82335 891
rect 82381 845 82459 891
rect 82505 845 82583 891
rect 82629 845 82707 891
rect 82753 845 82831 891
rect 82877 845 82955 891
rect 83001 845 83079 891
rect 83125 845 83203 891
rect 83249 845 83327 891
rect 83373 845 83451 891
rect 83497 845 83575 891
rect 83621 845 83699 891
rect 83745 845 83823 891
rect 83869 845 83947 891
rect 83993 845 84071 891
rect 84117 845 84195 891
rect 84241 845 84319 891
rect 84365 845 84443 891
rect 84489 845 84567 891
rect 84613 845 84691 891
rect 84737 845 84815 891
rect 84861 845 84939 891
rect 84985 845 85063 891
rect 85109 845 85187 891
rect 85233 845 85311 891
rect 85357 845 85435 891
rect 85481 845 85559 891
rect 85605 845 85683 891
rect 85729 845 85807 891
rect 85853 845 85931 891
rect 85977 845 86090 891
rect 282 767 29090 845
rect 29142 767 29787 845
rect 29839 775 53907 845
rect 29839 767 48668 775
rect 282 721 371 767
rect 417 721 495 767
rect 541 721 619 767
rect 665 721 743 767
rect 789 721 867 767
rect 913 721 991 767
rect 1037 721 1115 767
rect 1161 721 1239 767
rect 1285 721 1363 767
rect 1409 721 1487 767
rect 1533 721 1611 767
rect 1657 721 1735 767
rect 1781 721 1859 767
rect 1905 721 1983 767
rect 2029 721 2107 767
rect 2153 721 2231 767
rect 2277 721 2355 767
rect 2401 721 2479 767
rect 2525 721 2603 767
rect 2649 721 2727 767
rect 2773 721 2851 767
rect 2897 721 2975 767
rect 3021 721 3099 767
rect 3145 721 3223 767
rect 3269 721 3347 767
rect 3393 721 3471 767
rect 3517 721 3595 767
rect 3641 721 3719 767
rect 3765 721 3843 767
rect 3889 721 3967 767
rect 4013 721 4091 767
rect 4137 721 4215 767
rect 4261 721 4339 767
rect 4385 721 4463 767
rect 4509 721 4587 767
rect 4633 721 4711 767
rect 4757 721 4835 767
rect 4881 721 4959 767
rect 5005 721 5083 767
rect 5129 721 5207 767
rect 5253 721 5331 767
rect 5377 721 5455 767
rect 5501 721 5579 767
rect 5625 721 5703 767
rect 5749 721 5827 767
rect 5873 721 5951 767
rect 5997 721 6075 767
rect 6121 721 6199 767
rect 6245 721 6323 767
rect 6369 721 6447 767
rect 6493 721 6571 767
rect 6617 721 6695 767
rect 6741 721 6819 767
rect 6865 721 6943 767
rect 6989 721 7067 767
rect 7113 721 7191 767
rect 7237 721 7315 767
rect 7361 721 7439 767
rect 7485 721 7563 767
rect 7609 721 7687 767
rect 7733 721 7811 767
rect 7857 721 7935 767
rect 7981 721 8059 767
rect 8105 721 8183 767
rect 8229 721 8307 767
rect 8353 721 8431 767
rect 8477 721 8555 767
rect 8601 721 8679 767
rect 8725 721 8803 767
rect 8849 721 8927 767
rect 8973 721 9051 767
rect 9097 721 9175 767
rect 9221 721 9299 767
rect 9345 721 9423 767
rect 9469 721 9547 767
rect 9593 721 9671 767
rect 9717 721 9795 767
rect 9841 721 9919 767
rect 9965 721 10043 767
rect 10089 721 10167 767
rect 10213 721 10291 767
rect 10337 721 10415 767
rect 10461 721 10539 767
rect 10585 721 10663 767
rect 10709 721 10787 767
rect 10833 721 10911 767
rect 10957 721 11035 767
rect 11081 721 11159 767
rect 11205 721 11283 767
rect 11329 721 11407 767
rect 11453 721 11531 767
rect 11577 721 11655 767
rect 11701 721 11779 767
rect 11825 721 11903 767
rect 11949 721 12027 767
rect 12073 721 12151 767
rect 12197 721 12275 767
rect 12321 721 12399 767
rect 12445 721 12523 767
rect 12569 721 12647 767
rect 12693 721 12771 767
rect 12817 721 12895 767
rect 12941 721 13019 767
rect 13065 721 13143 767
rect 13189 721 13267 767
rect 13313 721 13391 767
rect 13437 721 13515 767
rect 13561 721 13639 767
rect 13685 721 13763 767
rect 13809 721 13887 767
rect 13933 721 14011 767
rect 14057 721 14135 767
rect 14181 721 14259 767
rect 14305 721 14383 767
rect 14429 721 14507 767
rect 14553 721 14631 767
rect 14677 721 14755 767
rect 14801 721 14879 767
rect 14925 721 15003 767
rect 15049 721 15127 767
rect 15173 721 15251 767
rect 15297 721 15375 767
rect 15421 721 15499 767
rect 15545 721 15623 767
rect 15669 721 15747 767
rect 15793 721 15871 767
rect 15917 721 15995 767
rect 16041 721 16119 767
rect 16165 721 16243 767
rect 16289 721 16367 767
rect 16413 721 16491 767
rect 16537 721 16615 767
rect 16661 721 16739 767
rect 16785 721 16863 767
rect 16909 721 16987 767
rect 17033 721 17111 767
rect 17157 721 17235 767
rect 17281 721 17359 767
rect 17405 721 17483 767
rect 17529 721 17607 767
rect 17653 721 17731 767
rect 17777 721 17855 767
rect 17901 721 17979 767
rect 18025 721 18103 767
rect 18149 721 18227 767
rect 18273 721 18351 767
rect 18397 721 18475 767
rect 18521 721 18599 767
rect 18645 721 18723 767
rect 18769 721 18847 767
rect 18893 721 18971 767
rect 19017 721 19095 767
rect 19141 721 19219 767
rect 19265 721 19343 767
rect 19389 721 19467 767
rect 19513 721 19591 767
rect 19637 721 19715 767
rect 19761 721 19839 767
rect 19885 721 19963 767
rect 20009 721 20087 767
rect 20133 721 20211 767
rect 20257 721 20335 767
rect 20381 721 20459 767
rect 20505 721 20583 767
rect 20629 721 20707 767
rect 20753 721 20831 767
rect 20877 721 20955 767
rect 21001 721 21079 767
rect 21125 721 21203 767
rect 21249 721 21327 767
rect 21373 721 21451 767
rect 21497 721 21575 767
rect 21621 721 21699 767
rect 21745 721 21823 767
rect 21869 721 21947 767
rect 21993 721 22071 767
rect 22117 721 22195 767
rect 22241 721 22319 767
rect 22365 721 22443 767
rect 22489 721 22567 767
rect 22613 721 22691 767
rect 22737 721 22815 767
rect 22861 721 22939 767
rect 22985 721 23063 767
rect 23109 721 23187 767
rect 23233 721 23311 767
rect 23357 721 23435 767
rect 23481 721 23559 767
rect 23605 721 23683 767
rect 23729 721 23807 767
rect 23853 721 23931 767
rect 23977 721 24055 767
rect 24101 721 24179 767
rect 24225 721 24303 767
rect 24349 721 24427 767
rect 24473 721 24551 767
rect 24597 721 24675 767
rect 24721 721 24799 767
rect 24845 721 24923 767
rect 24969 721 25047 767
rect 25093 721 25171 767
rect 25217 721 25295 767
rect 25341 721 25419 767
rect 25465 721 25543 767
rect 25589 721 25667 767
rect 25713 721 25791 767
rect 25837 721 25915 767
rect 25961 721 26039 767
rect 26085 721 26163 767
rect 26209 721 26287 767
rect 26333 721 26411 767
rect 26457 721 26535 767
rect 26581 721 26659 767
rect 26705 721 26783 767
rect 26829 721 26907 767
rect 26953 721 27031 767
rect 27077 721 27155 767
rect 27201 721 27279 767
rect 27325 721 27403 767
rect 27449 721 27527 767
rect 27573 721 27651 767
rect 27697 721 27775 767
rect 27821 721 27899 767
rect 27945 721 28023 767
rect 28069 721 28147 767
rect 28193 721 28271 767
rect 28317 721 28395 767
rect 28441 721 28519 767
rect 28565 721 28643 767
rect 28689 721 28767 767
rect 28813 721 28891 767
rect 28937 721 29015 767
rect 29061 721 29090 767
rect 29185 721 29263 767
rect 29309 721 29387 767
rect 29433 721 29511 767
rect 29557 721 29635 767
rect 29681 721 29759 767
rect 29839 721 29883 767
rect 29929 721 30007 767
rect 30053 721 30131 767
rect 30177 721 30255 767
rect 30301 721 30379 767
rect 30425 721 30503 767
rect 30549 721 30627 767
rect 30673 721 30751 767
rect 30797 721 30875 767
rect 30921 721 30999 767
rect 31045 721 31123 767
rect 31169 721 31247 767
rect 31293 721 31371 767
rect 31417 721 31495 767
rect 31541 721 31619 767
rect 31665 721 31743 767
rect 31789 721 31867 767
rect 31913 721 31991 767
rect 32037 721 32115 767
rect 32161 721 32239 767
rect 32285 721 32363 767
rect 32409 721 32487 767
rect 32533 721 32611 767
rect 32657 721 32735 767
rect 32781 721 32859 767
rect 32905 721 32983 767
rect 33029 721 33107 767
rect 33153 721 33231 767
rect 33277 721 33355 767
rect 33401 721 33479 767
rect 33525 721 33603 767
rect 33649 721 33727 767
rect 33773 721 33851 767
rect 33897 721 33975 767
rect 34021 721 34099 767
rect 34145 721 34223 767
rect 34269 721 34347 767
rect 34393 721 34471 767
rect 34517 721 34595 767
rect 34641 721 34719 767
rect 34765 721 34843 767
rect 34889 721 34967 767
rect 35013 721 35091 767
rect 35137 721 35215 767
rect 35261 721 35339 767
rect 35385 721 35463 767
rect 35509 721 35587 767
rect 35633 721 35711 767
rect 35757 721 35835 767
rect 35881 721 35959 767
rect 36005 721 36083 767
rect 36129 721 36207 767
rect 36253 721 36331 767
rect 36377 721 36455 767
rect 36501 721 36579 767
rect 36625 721 36703 767
rect 36749 721 36827 767
rect 36873 721 36951 767
rect 36997 721 37075 767
rect 37121 721 37199 767
rect 37245 721 37323 767
rect 37369 721 37447 767
rect 37493 721 37571 767
rect 37617 721 37695 767
rect 37741 721 37819 767
rect 37865 721 37943 767
rect 37989 721 38067 767
rect 38113 721 38191 767
rect 38237 721 38315 767
rect 38361 721 38439 767
rect 38485 721 38563 767
rect 38609 721 38687 767
rect 38733 721 38811 767
rect 38857 721 38935 767
rect 38981 721 39059 767
rect 39105 721 39183 767
rect 39229 721 39307 767
rect 39353 721 39431 767
rect 39477 721 39555 767
rect 39601 721 39679 767
rect 39725 721 39803 767
rect 39849 721 39927 767
rect 39973 721 40051 767
rect 40097 721 40175 767
rect 40221 721 40299 767
rect 40345 721 40423 767
rect 40469 721 40547 767
rect 40593 721 40671 767
rect 40717 721 40795 767
rect 40841 721 40919 767
rect 40965 721 41043 767
rect 41089 721 41167 767
rect 41213 721 41291 767
rect 41337 721 41415 767
rect 41461 721 41539 767
rect 41585 721 41663 767
rect 41709 721 41787 767
rect 41833 721 41911 767
rect 41957 721 42035 767
rect 42081 721 42159 767
rect 42205 721 42283 767
rect 42329 721 42407 767
rect 42453 721 42531 767
rect 42577 721 42655 767
rect 42701 721 42779 767
rect 42825 721 42903 767
rect 42949 721 43027 767
rect 43073 721 43151 767
rect 43197 721 43275 767
rect 43321 721 43399 767
rect 43445 721 43523 767
rect 43569 721 43647 767
rect 43693 721 43771 767
rect 43817 721 43895 767
rect 43941 721 44019 767
rect 44065 721 44143 767
rect 44189 721 44267 767
rect 44313 721 44391 767
rect 44437 721 44515 767
rect 44561 721 44639 767
rect 44685 721 44763 767
rect 44809 721 44887 767
rect 44933 721 45011 767
rect 45057 721 45135 767
rect 45181 721 45259 767
rect 45305 721 45383 767
rect 45429 721 45507 767
rect 45553 721 45631 767
rect 45677 721 45755 767
rect 45801 721 45879 767
rect 45925 721 46003 767
rect 46049 721 46127 767
rect 46173 721 46251 767
rect 46297 721 46375 767
rect 46421 721 46499 767
rect 46545 721 46623 767
rect 46669 721 46747 767
rect 46793 721 46871 767
rect 46917 721 46995 767
rect 47041 721 47119 767
rect 47165 721 47243 767
rect 47289 721 47367 767
rect 47413 721 47491 767
rect 47537 721 47615 767
rect 47661 721 47739 767
rect 47785 721 47863 767
rect 47909 721 47987 767
rect 48033 721 48111 767
rect 48157 721 48235 767
rect 48281 721 48359 767
rect 48405 721 48483 767
rect 48529 721 48607 767
rect 48653 723 48668 767
rect 48720 767 48792 775
rect 48720 723 48731 767
rect 48653 721 48731 723
rect 48777 723 48792 767
rect 48844 767 48916 775
rect 48844 723 48855 767
rect 48777 721 48855 723
rect 48901 723 48916 767
rect 48968 767 53907 775
rect 53959 767 86090 845
rect 48968 723 48979 767
rect 48901 721 48979 723
rect 49025 721 49103 767
rect 49149 721 49227 767
rect 49273 721 49351 767
rect 49397 721 49475 767
rect 49521 721 49599 767
rect 49645 721 49723 767
rect 49769 721 49847 767
rect 49893 721 49971 767
rect 50017 721 50095 767
rect 50141 721 50219 767
rect 50265 721 50343 767
rect 50389 721 50467 767
rect 50513 721 50591 767
rect 50637 721 50715 767
rect 50761 721 50839 767
rect 50885 721 50963 767
rect 51009 721 51087 767
rect 51133 721 51211 767
rect 51257 721 51335 767
rect 51381 721 51459 767
rect 51505 721 51583 767
rect 51629 721 51707 767
rect 51753 721 51831 767
rect 51877 721 51955 767
rect 52001 721 52079 767
rect 52125 721 52203 767
rect 52249 721 52327 767
rect 52373 721 52451 767
rect 52497 721 52575 767
rect 52621 721 52699 767
rect 52745 721 52823 767
rect 52869 721 52947 767
rect 52993 721 53071 767
rect 53117 721 53195 767
rect 53241 721 53319 767
rect 53365 721 53443 767
rect 53489 721 53567 767
rect 53613 721 53691 767
rect 53737 721 53815 767
rect 53861 721 53907 767
rect 53985 721 54063 767
rect 54109 721 54187 767
rect 54233 721 54311 767
rect 54357 721 54435 767
rect 54481 721 54559 767
rect 54605 721 54683 767
rect 54729 721 54807 767
rect 54853 721 54931 767
rect 54977 721 55055 767
rect 55101 721 55179 767
rect 55225 721 55303 767
rect 55349 721 55427 767
rect 55473 721 55551 767
rect 55597 721 55675 767
rect 55721 721 55799 767
rect 55845 721 55923 767
rect 55969 721 56047 767
rect 56093 721 56171 767
rect 56217 721 56295 767
rect 56341 721 56419 767
rect 56465 721 56543 767
rect 56589 721 56667 767
rect 56713 721 56791 767
rect 56837 721 56915 767
rect 56961 721 57039 767
rect 57085 721 57163 767
rect 57209 721 57287 767
rect 57333 721 57411 767
rect 57457 721 57535 767
rect 57581 721 57659 767
rect 57705 721 57783 767
rect 57829 721 57907 767
rect 57953 721 58031 767
rect 58077 721 58155 767
rect 58201 721 58279 767
rect 58325 721 58403 767
rect 58449 721 58527 767
rect 58573 721 58651 767
rect 58697 721 58775 767
rect 58821 721 58899 767
rect 58945 721 59023 767
rect 59069 721 59147 767
rect 59193 721 59271 767
rect 59317 721 59395 767
rect 59441 721 59519 767
rect 59565 721 59643 767
rect 59689 721 59767 767
rect 59813 721 59891 767
rect 59937 721 60015 767
rect 60061 721 60139 767
rect 60185 721 60263 767
rect 60309 721 60387 767
rect 60433 721 60511 767
rect 60557 721 60635 767
rect 60681 721 60759 767
rect 60805 721 60883 767
rect 60929 721 61007 767
rect 61053 721 61131 767
rect 61177 721 61255 767
rect 61301 721 61379 767
rect 61425 721 61503 767
rect 61549 721 61627 767
rect 61673 721 61751 767
rect 61797 721 61875 767
rect 61921 721 61999 767
rect 62045 721 62123 767
rect 62169 721 62247 767
rect 62293 721 62371 767
rect 62417 721 62495 767
rect 62541 721 62619 767
rect 62665 721 62743 767
rect 62789 721 62867 767
rect 62913 721 62991 767
rect 63037 721 63115 767
rect 63161 721 63239 767
rect 63285 721 63363 767
rect 63409 721 63487 767
rect 63533 721 63611 767
rect 63657 721 63735 767
rect 63781 721 63859 767
rect 63905 721 63983 767
rect 64029 721 64107 767
rect 64153 721 64231 767
rect 64277 721 64355 767
rect 64401 721 64479 767
rect 64525 721 64603 767
rect 64649 721 64727 767
rect 64773 721 64851 767
rect 64897 721 64975 767
rect 65021 721 65099 767
rect 65145 721 65223 767
rect 65269 721 65347 767
rect 65393 721 65471 767
rect 65517 721 65595 767
rect 65641 721 65719 767
rect 65765 721 65843 767
rect 65889 721 65967 767
rect 66013 721 66091 767
rect 66137 721 66215 767
rect 66261 721 66339 767
rect 66385 721 66463 767
rect 66509 721 66587 767
rect 66633 721 66711 767
rect 66757 721 66835 767
rect 66881 721 66959 767
rect 67005 721 67083 767
rect 67129 721 67207 767
rect 67253 721 67331 767
rect 67377 721 67455 767
rect 67501 721 67579 767
rect 67625 721 67703 767
rect 67749 721 67827 767
rect 67873 721 67951 767
rect 67997 721 68075 767
rect 68121 721 68199 767
rect 68245 721 68323 767
rect 68369 721 68447 767
rect 68493 721 68571 767
rect 68617 721 68695 767
rect 68741 721 68819 767
rect 68865 721 68943 767
rect 68989 721 69067 767
rect 69113 721 69191 767
rect 69237 721 69315 767
rect 69361 721 69439 767
rect 69485 721 69563 767
rect 69609 721 69687 767
rect 69733 721 69811 767
rect 69857 721 69935 767
rect 69981 721 70059 767
rect 70105 721 70183 767
rect 70229 721 70307 767
rect 70353 721 70431 767
rect 70477 721 70555 767
rect 70601 721 70679 767
rect 70725 721 70803 767
rect 70849 721 70927 767
rect 70973 721 71051 767
rect 71097 721 71175 767
rect 71221 721 71299 767
rect 71345 721 71423 767
rect 71469 721 71547 767
rect 71593 721 71671 767
rect 71717 721 71795 767
rect 71841 721 71919 767
rect 71965 721 72043 767
rect 72089 721 72167 767
rect 72213 721 72291 767
rect 72337 721 72415 767
rect 72461 721 72539 767
rect 72585 721 72663 767
rect 72709 721 72787 767
rect 72833 721 72911 767
rect 72957 721 73035 767
rect 73081 721 73159 767
rect 73205 721 73283 767
rect 73329 721 73407 767
rect 73453 721 73531 767
rect 73577 721 73655 767
rect 73701 721 73779 767
rect 73825 721 73903 767
rect 73949 721 74027 767
rect 74073 721 74151 767
rect 74197 721 74275 767
rect 74321 721 74399 767
rect 74445 721 74523 767
rect 74569 721 74647 767
rect 74693 721 74771 767
rect 74817 721 74895 767
rect 74941 721 75019 767
rect 75065 721 75143 767
rect 75189 721 75267 767
rect 75313 721 75391 767
rect 75437 721 75515 767
rect 75561 721 75639 767
rect 75685 721 75763 767
rect 75809 721 75887 767
rect 75933 721 76011 767
rect 76057 721 76135 767
rect 76181 721 76259 767
rect 76305 721 76383 767
rect 76429 721 76507 767
rect 76553 721 76631 767
rect 76677 721 76755 767
rect 76801 721 76879 767
rect 76925 721 77003 767
rect 77049 721 77127 767
rect 77173 721 77251 767
rect 77297 721 77375 767
rect 77421 721 77499 767
rect 77545 721 77623 767
rect 77669 721 77747 767
rect 77793 721 77871 767
rect 77917 721 77995 767
rect 78041 721 78119 767
rect 78165 721 78243 767
rect 78289 721 78367 767
rect 78413 721 78491 767
rect 78537 721 78615 767
rect 78661 721 78739 767
rect 78785 721 78863 767
rect 78909 721 78987 767
rect 79033 721 79111 767
rect 79157 721 79235 767
rect 79281 721 79359 767
rect 79405 721 79483 767
rect 79529 721 79607 767
rect 79653 721 79731 767
rect 79777 721 79855 767
rect 79901 721 79979 767
rect 80025 721 80103 767
rect 80149 721 80227 767
rect 80273 721 80351 767
rect 80397 721 80475 767
rect 80521 721 80599 767
rect 80645 721 80723 767
rect 80769 721 80847 767
rect 80893 721 80971 767
rect 81017 721 81095 767
rect 81141 721 81219 767
rect 81265 721 81343 767
rect 81389 721 81467 767
rect 81513 721 81591 767
rect 81637 721 81715 767
rect 81761 721 81839 767
rect 81885 721 81963 767
rect 82009 721 82087 767
rect 82133 721 82211 767
rect 82257 721 82335 767
rect 82381 721 82459 767
rect 82505 721 82583 767
rect 82629 721 82707 767
rect 82753 721 82831 767
rect 82877 721 82955 767
rect 83001 721 83079 767
rect 83125 721 83203 767
rect 83249 721 83327 767
rect 83373 721 83451 767
rect 83497 721 83575 767
rect 83621 721 83699 767
rect 83745 721 83823 767
rect 83869 721 83947 767
rect 83993 721 84071 767
rect 84117 721 84195 767
rect 84241 721 84319 767
rect 84365 721 84443 767
rect 84489 721 84567 767
rect 84613 721 84691 767
rect 84737 721 84815 767
rect 84861 721 84939 767
rect 84985 721 85063 767
rect 85109 721 85187 767
rect 85233 721 85311 767
rect 85357 721 85435 767
rect 85481 721 85559 767
rect 85605 721 85683 767
rect 85729 721 85807 767
rect 85853 721 85931 767
rect 85977 721 86090 767
rect 282 654 29090 721
rect 29142 654 29787 721
rect 29839 654 53907 721
rect 282 651 53907 654
rect 282 643 48668 651
rect 282 597 371 643
rect 417 597 495 643
rect 541 597 619 643
rect 665 597 743 643
rect 789 597 867 643
rect 913 597 991 643
rect 1037 597 1115 643
rect 1161 597 1239 643
rect 1285 597 1363 643
rect 1409 597 1487 643
rect 1533 597 1611 643
rect 1657 597 1735 643
rect 1781 597 1859 643
rect 1905 597 1983 643
rect 2029 597 2107 643
rect 2153 597 2231 643
rect 2277 597 2355 643
rect 2401 597 2479 643
rect 2525 597 2603 643
rect 2649 597 2727 643
rect 2773 597 2851 643
rect 2897 597 2975 643
rect 3021 597 3099 643
rect 3145 597 3223 643
rect 3269 597 3347 643
rect 3393 597 3471 643
rect 3517 597 3595 643
rect 3641 597 3719 643
rect 3765 597 3843 643
rect 3889 597 3967 643
rect 4013 597 4091 643
rect 4137 597 4215 643
rect 4261 597 4339 643
rect 4385 597 4463 643
rect 4509 597 4587 643
rect 4633 597 4711 643
rect 4757 597 4835 643
rect 4881 597 4959 643
rect 5005 597 5083 643
rect 5129 597 5207 643
rect 5253 597 5331 643
rect 5377 597 5455 643
rect 5501 597 5579 643
rect 5625 597 5703 643
rect 5749 597 5827 643
rect 5873 597 5951 643
rect 5997 597 6075 643
rect 6121 597 6199 643
rect 6245 597 6323 643
rect 6369 597 6447 643
rect 6493 597 6571 643
rect 6617 597 6695 643
rect 6741 597 6819 643
rect 6865 597 6943 643
rect 6989 597 7067 643
rect 7113 597 7191 643
rect 7237 597 7315 643
rect 7361 597 7439 643
rect 7485 597 7563 643
rect 7609 597 7687 643
rect 7733 597 7811 643
rect 7857 597 7935 643
rect 7981 597 8059 643
rect 8105 597 8183 643
rect 8229 597 8307 643
rect 8353 597 8431 643
rect 8477 597 8555 643
rect 8601 597 8679 643
rect 8725 597 8803 643
rect 8849 597 8927 643
rect 8973 597 9051 643
rect 9097 597 9175 643
rect 9221 597 9299 643
rect 9345 597 9423 643
rect 9469 597 9547 643
rect 9593 597 9671 643
rect 9717 597 9795 643
rect 9841 597 9919 643
rect 9965 597 10043 643
rect 10089 597 10167 643
rect 10213 597 10291 643
rect 10337 597 10415 643
rect 10461 597 10539 643
rect 10585 597 10663 643
rect 10709 597 10787 643
rect 10833 597 10911 643
rect 10957 597 11035 643
rect 11081 597 11159 643
rect 11205 597 11283 643
rect 11329 597 11407 643
rect 11453 597 11531 643
rect 11577 597 11655 643
rect 11701 597 11779 643
rect 11825 597 11903 643
rect 11949 597 12027 643
rect 12073 597 12151 643
rect 12197 597 12275 643
rect 12321 597 12399 643
rect 12445 597 12523 643
rect 12569 597 12647 643
rect 12693 597 12771 643
rect 12817 597 12895 643
rect 12941 597 13019 643
rect 13065 597 13143 643
rect 13189 597 13267 643
rect 13313 597 13391 643
rect 13437 597 13515 643
rect 13561 597 13639 643
rect 13685 597 13763 643
rect 13809 597 13887 643
rect 13933 597 14011 643
rect 14057 597 14135 643
rect 14181 597 14259 643
rect 14305 597 14383 643
rect 14429 597 14507 643
rect 14553 597 14631 643
rect 14677 597 14755 643
rect 14801 597 14879 643
rect 14925 597 15003 643
rect 15049 597 15127 643
rect 15173 597 15251 643
rect 15297 597 15375 643
rect 15421 597 15499 643
rect 15545 597 15623 643
rect 15669 597 15747 643
rect 15793 597 15871 643
rect 15917 597 15995 643
rect 16041 597 16119 643
rect 16165 597 16243 643
rect 16289 597 16367 643
rect 16413 597 16491 643
rect 16537 597 16615 643
rect 16661 597 16739 643
rect 16785 597 16863 643
rect 16909 597 16987 643
rect 17033 597 17111 643
rect 17157 597 17235 643
rect 17281 597 17359 643
rect 17405 597 17483 643
rect 17529 597 17607 643
rect 17653 597 17731 643
rect 17777 597 17855 643
rect 17901 597 17979 643
rect 18025 597 18103 643
rect 18149 597 18227 643
rect 18273 597 18351 643
rect 18397 597 18475 643
rect 18521 597 18599 643
rect 18645 597 18723 643
rect 18769 597 18847 643
rect 18893 597 18971 643
rect 19017 597 19095 643
rect 19141 597 19219 643
rect 19265 597 19343 643
rect 19389 597 19467 643
rect 19513 597 19591 643
rect 19637 597 19715 643
rect 19761 597 19839 643
rect 19885 597 19963 643
rect 20009 597 20087 643
rect 20133 597 20211 643
rect 20257 597 20335 643
rect 20381 597 20459 643
rect 20505 597 20583 643
rect 20629 597 20707 643
rect 20753 597 20831 643
rect 20877 597 20955 643
rect 21001 597 21079 643
rect 21125 597 21203 643
rect 21249 597 21327 643
rect 21373 597 21451 643
rect 21497 597 21575 643
rect 21621 597 21699 643
rect 21745 597 21823 643
rect 21869 597 21947 643
rect 21993 597 22071 643
rect 22117 597 22195 643
rect 22241 597 22319 643
rect 22365 597 22443 643
rect 22489 597 22567 643
rect 22613 597 22691 643
rect 22737 597 22815 643
rect 22861 597 22939 643
rect 22985 597 23063 643
rect 23109 597 23187 643
rect 23233 597 23311 643
rect 23357 597 23435 643
rect 23481 597 23559 643
rect 23605 597 23683 643
rect 23729 597 23807 643
rect 23853 597 23931 643
rect 23977 597 24055 643
rect 24101 597 24179 643
rect 24225 597 24303 643
rect 24349 597 24427 643
rect 24473 597 24551 643
rect 24597 597 24675 643
rect 24721 597 24799 643
rect 24845 597 24923 643
rect 24969 597 25047 643
rect 25093 597 25171 643
rect 25217 597 25295 643
rect 25341 597 25419 643
rect 25465 597 25543 643
rect 25589 597 25667 643
rect 25713 597 25791 643
rect 25837 597 25915 643
rect 25961 597 26039 643
rect 26085 597 26163 643
rect 26209 597 26287 643
rect 26333 597 26411 643
rect 26457 597 26535 643
rect 26581 597 26659 643
rect 26705 597 26783 643
rect 26829 597 26907 643
rect 26953 597 27031 643
rect 27077 597 27155 643
rect 27201 597 27279 643
rect 27325 597 27403 643
rect 27449 597 27527 643
rect 27573 597 27651 643
rect 27697 597 27775 643
rect 27821 597 27899 643
rect 27945 597 28023 643
rect 28069 597 28147 643
rect 28193 597 28271 643
rect 28317 597 28395 643
rect 28441 597 28519 643
rect 28565 597 28643 643
rect 28689 597 28767 643
rect 28813 597 28891 643
rect 28937 597 29015 643
rect 29061 597 29139 643
rect 29185 597 29263 643
rect 29309 597 29387 643
rect 29433 597 29511 643
rect 29557 597 29635 643
rect 29681 597 29759 643
rect 29805 597 29883 643
rect 29929 597 30007 643
rect 30053 597 30131 643
rect 30177 597 30255 643
rect 30301 597 30379 643
rect 30425 597 30503 643
rect 30549 597 30627 643
rect 30673 597 30751 643
rect 30797 597 30875 643
rect 30921 597 30999 643
rect 31045 597 31123 643
rect 31169 597 31247 643
rect 31293 597 31371 643
rect 31417 597 31495 643
rect 31541 597 31619 643
rect 31665 597 31743 643
rect 31789 597 31867 643
rect 31913 597 31991 643
rect 32037 597 32115 643
rect 32161 597 32239 643
rect 32285 597 32363 643
rect 32409 597 32487 643
rect 32533 597 32611 643
rect 32657 597 32735 643
rect 32781 597 32859 643
rect 32905 597 32983 643
rect 33029 597 33107 643
rect 33153 597 33231 643
rect 33277 597 33355 643
rect 33401 597 33479 643
rect 33525 597 33603 643
rect 33649 597 33727 643
rect 33773 597 33851 643
rect 33897 597 33975 643
rect 34021 597 34099 643
rect 34145 597 34223 643
rect 34269 597 34347 643
rect 34393 597 34471 643
rect 34517 597 34595 643
rect 34641 597 34719 643
rect 34765 597 34843 643
rect 34889 597 34967 643
rect 35013 597 35091 643
rect 35137 597 35215 643
rect 35261 597 35339 643
rect 35385 597 35463 643
rect 35509 597 35587 643
rect 35633 597 35711 643
rect 35757 597 35835 643
rect 35881 597 35959 643
rect 36005 597 36083 643
rect 36129 597 36207 643
rect 36253 597 36331 643
rect 36377 597 36455 643
rect 36501 597 36579 643
rect 36625 597 36703 643
rect 36749 597 36827 643
rect 36873 597 36951 643
rect 36997 597 37075 643
rect 37121 597 37199 643
rect 37245 597 37323 643
rect 37369 597 37447 643
rect 37493 597 37571 643
rect 37617 597 37695 643
rect 37741 597 37819 643
rect 37865 597 37943 643
rect 37989 597 38067 643
rect 38113 597 38191 643
rect 38237 597 38315 643
rect 38361 597 38439 643
rect 38485 597 38563 643
rect 38609 597 38687 643
rect 38733 597 38811 643
rect 38857 597 38935 643
rect 38981 597 39059 643
rect 39105 597 39183 643
rect 39229 597 39307 643
rect 39353 597 39431 643
rect 39477 597 39555 643
rect 39601 597 39679 643
rect 39725 597 39803 643
rect 39849 597 39927 643
rect 39973 597 40051 643
rect 40097 597 40175 643
rect 40221 597 40299 643
rect 40345 597 40423 643
rect 40469 597 40547 643
rect 40593 597 40671 643
rect 40717 597 40795 643
rect 40841 597 40919 643
rect 40965 597 41043 643
rect 41089 597 41167 643
rect 41213 597 41291 643
rect 41337 597 41415 643
rect 41461 597 41539 643
rect 41585 597 41663 643
rect 41709 597 41787 643
rect 41833 597 41911 643
rect 41957 597 42035 643
rect 42081 597 42159 643
rect 42205 597 42283 643
rect 42329 597 42407 643
rect 42453 597 42531 643
rect 42577 597 42655 643
rect 42701 597 42779 643
rect 42825 597 42903 643
rect 42949 597 43027 643
rect 43073 597 43151 643
rect 43197 597 43275 643
rect 43321 597 43399 643
rect 43445 597 43523 643
rect 43569 597 43647 643
rect 43693 597 43771 643
rect 43817 597 43895 643
rect 43941 597 44019 643
rect 44065 597 44143 643
rect 44189 597 44267 643
rect 44313 597 44391 643
rect 44437 597 44515 643
rect 44561 597 44639 643
rect 44685 597 44763 643
rect 44809 597 44887 643
rect 44933 597 45011 643
rect 45057 597 45135 643
rect 45181 597 45259 643
rect 45305 597 45383 643
rect 45429 597 45507 643
rect 45553 597 45631 643
rect 45677 597 45755 643
rect 45801 597 45879 643
rect 45925 597 46003 643
rect 46049 597 46127 643
rect 46173 597 46251 643
rect 46297 597 46375 643
rect 46421 597 46499 643
rect 46545 597 46623 643
rect 46669 597 46747 643
rect 46793 597 46871 643
rect 46917 597 46995 643
rect 47041 597 47119 643
rect 47165 597 47243 643
rect 47289 597 47367 643
rect 47413 597 47491 643
rect 47537 597 47615 643
rect 47661 597 47739 643
rect 47785 597 47863 643
rect 47909 597 47987 643
rect 48033 597 48111 643
rect 48157 597 48235 643
rect 48281 597 48359 643
rect 48405 597 48483 643
rect 48529 597 48607 643
rect 48653 599 48668 643
rect 48720 643 48792 651
rect 48720 599 48731 643
rect 48653 597 48731 599
rect 48777 599 48792 643
rect 48844 643 48916 651
rect 48844 599 48855 643
rect 48777 597 48855 599
rect 48901 599 48916 643
rect 48968 643 53907 651
rect 53959 643 86090 721
rect 48968 599 48979 643
rect 48901 597 48979 599
rect 49025 597 49103 643
rect 49149 597 49227 643
rect 49273 597 49351 643
rect 49397 597 49475 643
rect 49521 597 49599 643
rect 49645 597 49723 643
rect 49769 597 49847 643
rect 49893 597 49971 643
rect 50017 597 50095 643
rect 50141 597 50219 643
rect 50265 597 50343 643
rect 50389 597 50467 643
rect 50513 597 50591 643
rect 50637 597 50715 643
rect 50761 597 50839 643
rect 50885 597 50963 643
rect 51009 597 51087 643
rect 51133 597 51211 643
rect 51257 597 51335 643
rect 51381 597 51459 643
rect 51505 597 51583 643
rect 51629 597 51707 643
rect 51753 597 51831 643
rect 51877 597 51955 643
rect 52001 597 52079 643
rect 52125 597 52203 643
rect 52249 597 52327 643
rect 52373 597 52451 643
rect 52497 597 52575 643
rect 52621 597 52699 643
rect 52745 597 52823 643
rect 52869 597 52947 643
rect 52993 597 53071 643
rect 53117 597 53195 643
rect 53241 597 53319 643
rect 53365 597 53443 643
rect 53489 597 53567 643
rect 53613 597 53691 643
rect 53737 597 53815 643
rect 53861 642 53907 643
rect 53861 597 53939 642
rect 53985 597 54063 643
rect 54109 597 54187 643
rect 54233 597 54311 643
rect 54357 597 54435 643
rect 54481 597 54559 643
rect 54605 597 54683 643
rect 54729 597 54807 643
rect 54853 597 54931 643
rect 54977 597 55055 643
rect 55101 597 55179 643
rect 55225 597 55303 643
rect 55349 597 55427 643
rect 55473 597 55551 643
rect 55597 597 55675 643
rect 55721 597 55799 643
rect 55845 597 55923 643
rect 55969 597 56047 643
rect 56093 597 56171 643
rect 56217 597 56295 643
rect 56341 597 56419 643
rect 56465 597 56543 643
rect 56589 597 56667 643
rect 56713 597 56791 643
rect 56837 597 56915 643
rect 56961 597 57039 643
rect 57085 597 57163 643
rect 57209 597 57287 643
rect 57333 597 57411 643
rect 57457 597 57535 643
rect 57581 597 57659 643
rect 57705 597 57783 643
rect 57829 597 57907 643
rect 57953 597 58031 643
rect 58077 597 58155 643
rect 58201 597 58279 643
rect 58325 597 58403 643
rect 58449 597 58527 643
rect 58573 597 58651 643
rect 58697 597 58775 643
rect 58821 597 58899 643
rect 58945 597 59023 643
rect 59069 597 59147 643
rect 59193 597 59271 643
rect 59317 597 59395 643
rect 59441 597 59519 643
rect 59565 597 59643 643
rect 59689 597 59767 643
rect 59813 597 59891 643
rect 59937 597 60015 643
rect 60061 597 60139 643
rect 60185 597 60263 643
rect 60309 597 60387 643
rect 60433 597 60511 643
rect 60557 597 60635 643
rect 60681 597 60759 643
rect 60805 597 60883 643
rect 60929 597 61007 643
rect 61053 597 61131 643
rect 61177 597 61255 643
rect 61301 597 61379 643
rect 61425 597 61503 643
rect 61549 597 61627 643
rect 61673 597 61751 643
rect 61797 597 61875 643
rect 61921 597 61999 643
rect 62045 597 62123 643
rect 62169 597 62247 643
rect 62293 597 62371 643
rect 62417 597 62495 643
rect 62541 597 62619 643
rect 62665 597 62743 643
rect 62789 597 62867 643
rect 62913 597 62991 643
rect 63037 597 63115 643
rect 63161 597 63239 643
rect 63285 597 63363 643
rect 63409 597 63487 643
rect 63533 597 63611 643
rect 63657 597 63735 643
rect 63781 597 63859 643
rect 63905 597 63983 643
rect 64029 597 64107 643
rect 64153 597 64231 643
rect 64277 597 64355 643
rect 64401 597 64479 643
rect 64525 597 64603 643
rect 64649 597 64727 643
rect 64773 597 64851 643
rect 64897 597 64975 643
rect 65021 597 65099 643
rect 65145 597 65223 643
rect 65269 597 65347 643
rect 65393 597 65471 643
rect 65517 597 65595 643
rect 65641 597 65719 643
rect 65765 597 65843 643
rect 65889 597 65967 643
rect 66013 597 66091 643
rect 66137 597 66215 643
rect 66261 597 66339 643
rect 66385 597 66463 643
rect 66509 597 66587 643
rect 66633 597 66711 643
rect 66757 597 66835 643
rect 66881 597 66959 643
rect 67005 597 67083 643
rect 67129 597 67207 643
rect 67253 597 67331 643
rect 67377 597 67455 643
rect 67501 597 67579 643
rect 67625 597 67703 643
rect 67749 597 67827 643
rect 67873 597 67951 643
rect 67997 597 68075 643
rect 68121 597 68199 643
rect 68245 597 68323 643
rect 68369 597 68447 643
rect 68493 597 68571 643
rect 68617 597 68695 643
rect 68741 597 68819 643
rect 68865 597 68943 643
rect 68989 597 69067 643
rect 69113 597 69191 643
rect 69237 597 69315 643
rect 69361 597 69439 643
rect 69485 597 69563 643
rect 69609 597 69687 643
rect 69733 597 69811 643
rect 69857 597 69935 643
rect 69981 597 70059 643
rect 70105 597 70183 643
rect 70229 597 70307 643
rect 70353 597 70431 643
rect 70477 597 70555 643
rect 70601 597 70679 643
rect 70725 597 70803 643
rect 70849 597 70927 643
rect 70973 597 71051 643
rect 71097 597 71175 643
rect 71221 597 71299 643
rect 71345 597 71423 643
rect 71469 597 71547 643
rect 71593 597 71671 643
rect 71717 597 71795 643
rect 71841 597 71919 643
rect 71965 597 72043 643
rect 72089 597 72167 643
rect 72213 597 72291 643
rect 72337 597 72415 643
rect 72461 597 72539 643
rect 72585 597 72663 643
rect 72709 597 72787 643
rect 72833 597 72911 643
rect 72957 597 73035 643
rect 73081 597 73159 643
rect 73205 597 73283 643
rect 73329 597 73407 643
rect 73453 597 73531 643
rect 73577 597 73655 643
rect 73701 597 73779 643
rect 73825 597 73903 643
rect 73949 597 74027 643
rect 74073 597 74151 643
rect 74197 597 74275 643
rect 74321 597 74399 643
rect 74445 597 74523 643
rect 74569 597 74647 643
rect 74693 597 74771 643
rect 74817 597 74895 643
rect 74941 597 75019 643
rect 75065 597 75143 643
rect 75189 597 75267 643
rect 75313 597 75391 643
rect 75437 597 75515 643
rect 75561 597 75639 643
rect 75685 597 75763 643
rect 75809 597 75887 643
rect 75933 597 76011 643
rect 76057 597 76135 643
rect 76181 597 76259 643
rect 76305 597 76383 643
rect 76429 597 76507 643
rect 76553 597 76631 643
rect 76677 597 76755 643
rect 76801 597 76879 643
rect 76925 597 77003 643
rect 77049 597 77127 643
rect 77173 597 77251 643
rect 77297 597 77375 643
rect 77421 597 77499 643
rect 77545 597 77623 643
rect 77669 597 77747 643
rect 77793 597 77871 643
rect 77917 597 77995 643
rect 78041 597 78119 643
rect 78165 597 78243 643
rect 78289 597 78367 643
rect 78413 597 78491 643
rect 78537 597 78615 643
rect 78661 597 78739 643
rect 78785 597 78863 643
rect 78909 597 78987 643
rect 79033 597 79111 643
rect 79157 597 79235 643
rect 79281 597 79359 643
rect 79405 597 79483 643
rect 79529 597 79607 643
rect 79653 597 79731 643
rect 79777 597 79855 643
rect 79901 597 79979 643
rect 80025 597 80103 643
rect 80149 597 80227 643
rect 80273 597 80351 643
rect 80397 597 80475 643
rect 80521 597 80599 643
rect 80645 597 80723 643
rect 80769 597 80847 643
rect 80893 597 80971 643
rect 81017 597 81095 643
rect 81141 597 81219 643
rect 81265 597 81343 643
rect 81389 597 81467 643
rect 81513 597 81591 643
rect 81637 597 81715 643
rect 81761 597 81839 643
rect 81885 597 81963 643
rect 82009 597 82087 643
rect 82133 597 82211 643
rect 82257 597 82335 643
rect 82381 597 82459 643
rect 82505 597 82583 643
rect 82629 597 82707 643
rect 82753 597 82831 643
rect 82877 597 82955 643
rect 83001 597 83079 643
rect 83125 597 83203 643
rect 83249 597 83327 643
rect 83373 597 83451 643
rect 83497 597 83575 643
rect 83621 597 83699 643
rect 83745 597 83823 643
rect 83869 597 83947 643
rect 83993 597 84071 643
rect 84117 597 84195 643
rect 84241 597 84319 643
rect 84365 597 84443 643
rect 84489 597 84567 643
rect 84613 597 84691 643
rect 84737 597 84815 643
rect 84861 597 84939 643
rect 84985 597 85063 643
rect 85109 597 85187 643
rect 85233 597 85311 643
rect 85357 597 85435 643
rect 85481 597 85559 643
rect 85605 597 85683 643
rect 85729 597 85807 643
rect 85853 597 85931 643
rect 85977 597 86090 643
rect 282 282 86090 597
<< via1 >>
rect 25337 44286 25389 44338
rect 25461 44286 25513 44338
rect 25585 44286 25637 44338
rect 25709 44286 25761 44338
rect 25833 44286 25885 44338
rect 25957 44286 26009 44338
rect 25337 44162 25389 44214
rect 25461 44162 25513 44214
rect 25585 44162 25637 44214
rect 25709 44162 25761 44214
rect 25833 44162 25885 44214
rect 25957 44162 26009 44214
rect 25400 34920 25452 34972
rect 25524 34920 25576 34972
rect 25648 34920 25700 34972
rect 25772 34920 25824 34972
rect 25896 34920 25948 34972
rect 27790 44201 27842 44253
rect 28001 44201 28053 44253
rect 28212 44201 28264 44253
rect 28423 44201 28475 44253
rect 28634 44201 28686 44253
rect 28845 44201 28897 44253
rect 29056 44201 29108 44253
rect 29582 44201 29634 44253
rect 29793 44250 29845 44253
rect 29793 44204 29798 44250
rect 29798 44204 29844 44250
rect 29844 44204 29845 44250
rect 29793 44201 29845 44204
rect 30005 44201 30057 44253
rect 30216 44201 30268 44253
rect 30807 44236 30859 44253
rect 31018 44236 31070 44253
rect 30807 44201 30854 44236
rect 30854 44201 30859 44236
rect 31018 44201 31058 44236
rect 31058 44201 31070 44236
rect 31229 44201 31281 44253
rect 31440 44236 31492 44253
rect 31651 44236 31703 44253
rect 31440 44201 31487 44236
rect 31487 44201 31492 44236
rect 31651 44201 31691 44236
rect 31691 44201 31703 44236
rect 31861 44201 31913 44253
rect 32072 44236 32124 44253
rect 32283 44236 32335 44253
rect 32072 44201 32119 44236
rect 32119 44201 32124 44236
rect 32283 44201 32323 44236
rect 32323 44201 32335 44236
rect 32494 44201 32546 44253
rect 30807 44027 30854 44035
rect 30854 44027 30859 44035
rect 31018 44027 31058 44035
rect 31058 44027 31070 44035
rect 30807 43983 30859 44027
rect 31018 43983 31070 44027
rect 31229 43983 31281 44035
rect 31440 44027 31487 44035
rect 31487 44027 31492 44035
rect 31651 44027 31691 44035
rect 31691 44027 31703 44035
rect 31440 43983 31492 44027
rect 31651 43983 31703 44027
rect 31861 43983 31913 44035
rect 32072 44027 32119 44035
rect 32119 44027 32124 44035
rect 32283 44027 32323 44035
rect 32323 44027 32335 44035
rect 32072 43983 32124 44027
rect 32283 43983 32335 44027
rect 32494 43983 32546 44035
rect 34290 44201 34342 44253
rect 34501 44201 34553 44253
rect 34712 44201 34764 44253
rect 34923 44201 34975 44253
rect 35443 44218 35495 44233
rect 35654 44218 35706 44233
rect 35865 44218 35917 44233
rect 36076 44218 36128 44233
rect 36287 44218 36339 44233
rect 35443 44181 35495 44218
rect 35654 44181 35706 44218
rect 35865 44181 35917 44218
rect 36076 44181 36128 44218
rect 36287 44181 36339 44218
rect 40252 44206 40304 44258
rect 40432 44206 40484 44258
rect 42710 44263 42717 44305
rect 42717 44263 42762 44305
rect 42710 44253 42762 44263
rect 42921 44253 42973 44305
rect 43132 44253 43184 44305
rect 34290 43983 34342 44035
rect 34501 43994 34553 44035
rect 34712 43994 34764 44035
rect 34923 43994 34975 44035
rect 34501 43983 34552 43994
rect 34552 43983 34553 43994
rect 34712 43983 34758 43994
rect 34758 43983 34764 43994
rect 34923 43983 34964 43994
rect 34964 43983 34975 43994
rect 30807 43766 30859 43818
rect 31018 43766 31070 43818
rect 31229 43766 31281 43818
rect 31440 43766 31492 43818
rect 31651 43766 31703 43818
rect 31861 43766 31913 43818
rect 32072 43766 32124 43818
rect 32283 43766 32335 43818
rect 32494 43766 32546 43818
rect 39053 43994 39105 44001
rect 39264 43994 39316 44001
rect 39475 43994 39527 44001
rect 42246 44192 42298 44244
rect 42458 44243 42510 44244
rect 42458 44197 42459 44243
rect 42459 44197 42510 44243
rect 43777 44253 43829 44305
rect 43988 44253 44040 44305
rect 44199 44253 44251 44305
rect 44410 44253 44462 44305
rect 42458 44192 42510 44197
rect 40252 43994 40304 44040
rect 40432 43994 40484 44040
rect 39053 43949 39102 43994
rect 39102 43949 39105 43994
rect 39264 43949 39310 43994
rect 39310 43949 39316 43994
rect 39475 43949 39518 43994
rect 39518 43949 39527 43994
rect 40252 43988 40303 43994
rect 40303 43988 40304 43994
rect 40432 43988 40463 43994
rect 40463 43988 40484 43994
rect 33050 43770 33102 43772
rect 33261 43770 33313 43772
rect 33472 43770 33524 43772
rect 33683 43770 33735 43772
rect 33894 43770 33946 43772
rect 48828 44218 48880 44233
rect 49039 44218 49091 44233
rect 49250 44218 49302 44233
rect 49461 44218 49513 44233
rect 48828 44181 48880 44218
rect 49039 44181 49053 44218
rect 49053 44181 49091 44218
rect 49250 44181 49259 44218
rect 49259 44181 49302 44218
rect 49461 44181 49465 44218
rect 49465 44181 49511 44218
rect 49511 44181 49513 44218
rect 50137 44201 50189 44253
rect 50348 44201 50400 44253
rect 50559 44201 50611 44253
rect 50770 44201 50822 44253
rect 50137 43994 50189 44035
rect 50348 43994 50400 44035
rect 50559 43994 50611 44035
rect 50770 43994 50822 44035
rect 33050 43724 33102 43770
rect 33261 43724 33313 43770
rect 33472 43724 33524 43770
rect 33683 43724 33735 43770
rect 33894 43724 33934 43770
rect 33934 43724 33946 43770
rect 35443 43724 35495 43770
rect 35654 43724 35706 43770
rect 35865 43724 35917 43770
rect 36076 43724 36128 43770
rect 36287 43724 36339 43770
rect 41010 43725 41022 43770
rect 41022 43725 41062 43770
rect 41221 43725 41228 43770
rect 41228 43725 41273 43770
rect 41432 43725 41436 43770
rect 41436 43725 41484 43770
rect 41643 43725 41644 43770
rect 41644 43725 41695 43770
rect 33050 43720 33102 43724
rect 33261 43720 33313 43724
rect 33472 43720 33524 43724
rect 33683 43720 33735 43724
rect 33894 43720 33946 43724
rect 35443 43718 35495 43724
rect 35654 43718 35706 43724
rect 35865 43718 35917 43724
rect 36076 43718 36128 43724
rect 36287 43718 36339 43724
rect 41010 43718 41062 43725
rect 41221 43718 41273 43725
rect 41432 43718 41484 43725
rect 41643 43718 41695 43725
rect 41854 43718 41906 43770
rect 42064 43718 42116 43770
rect 50137 43983 50189 43994
rect 50348 43983 50400 43994
rect 50559 43983 50611 43994
rect 50770 43983 50774 43994
rect 50774 43983 50822 43994
rect 52576 44201 52628 44253
rect 52787 44236 52839 44253
rect 52998 44236 53050 44253
rect 52787 44201 52799 44236
rect 52799 44201 52839 44236
rect 52998 44201 53003 44236
rect 53003 44201 53050 44236
rect 53209 44201 53261 44253
rect 53419 44236 53471 44253
rect 53630 44236 53682 44253
rect 53419 44201 53431 44236
rect 53431 44201 53471 44236
rect 53630 44201 53635 44236
rect 53635 44201 53682 44236
rect 53841 44201 53893 44253
rect 54052 44236 54104 44253
rect 54263 44236 54315 44253
rect 54052 44201 54064 44236
rect 54064 44201 54104 44236
rect 54263 44201 54268 44236
rect 54268 44201 54315 44236
rect 54855 44201 54907 44253
rect 55066 44201 55118 44253
rect 55278 44250 55330 44253
rect 55278 44204 55279 44250
rect 55279 44204 55325 44250
rect 55325 44204 55330 44250
rect 55278 44201 55330 44204
rect 55489 44201 55541 44253
rect 56015 44201 56067 44253
rect 56226 44201 56278 44253
rect 56437 44201 56489 44253
rect 56648 44201 56700 44253
rect 56859 44201 56911 44253
rect 57070 44201 57122 44253
rect 57281 44201 57333 44253
rect 52576 43983 52628 44035
rect 52787 44027 52799 44035
rect 52799 44027 52839 44035
rect 52998 44027 53003 44035
rect 53003 44027 53050 44035
rect 52787 43983 52839 44027
rect 52998 43983 53050 44027
rect 53209 43983 53261 44035
rect 53419 44027 53431 44035
rect 53431 44027 53471 44035
rect 53630 44027 53635 44035
rect 53635 44027 53682 44035
rect 53419 43983 53471 44027
rect 53630 43983 53682 44027
rect 53841 43983 53893 44035
rect 54052 44027 54064 44035
rect 54064 44027 54104 44035
rect 54263 44027 54268 44035
rect 54268 44027 54315 44035
rect 54052 43983 54104 44027
rect 54263 43983 54315 44027
rect 48828 43724 48880 43770
rect 49039 43724 49053 43770
rect 49053 43724 49091 43770
rect 49250 43724 49259 43770
rect 49259 43724 49302 43770
rect 49461 43724 49465 43770
rect 49465 43724 49511 43770
rect 49511 43724 49513 43770
rect 51081 43724 51083 43770
rect 51083 43724 51133 43770
rect 48828 43718 48880 43724
rect 49039 43718 49091 43724
rect 49250 43718 49302 43724
rect 49461 43718 49513 43724
rect 51081 43718 51133 43724
rect 51292 43718 51344 43770
rect 51503 43724 51552 43770
rect 51552 43724 51555 43770
rect 51714 43724 51758 43770
rect 51758 43724 51766 43770
rect 51925 43724 51964 43770
rect 51964 43724 51977 43770
rect 52576 43766 52628 43818
rect 52787 43766 52839 43818
rect 52998 43766 53050 43818
rect 53209 43766 53261 43818
rect 53419 43766 53471 43818
rect 53630 43766 53682 43818
rect 53841 43766 53893 43818
rect 54052 43766 54104 43818
rect 54263 43766 54315 43818
rect 51503 43718 51555 43724
rect 51714 43718 51766 43724
rect 51925 43718 51977 43724
rect 29582 43301 29634 43353
rect 29793 43350 29845 43353
rect 29793 43304 29798 43350
rect 29798 43304 29844 43350
rect 29844 43304 29845 43350
rect 29793 43301 29845 43304
rect 30005 43301 30057 43353
rect 30216 43301 30268 43353
rect 30854 43301 30906 43353
rect 31065 43301 31117 43353
rect 31276 43301 31328 43353
rect 31486 43350 31538 43353
rect 31697 43350 31749 43353
rect 31909 43350 31961 43353
rect 32120 43350 32172 43353
rect 32330 43350 32382 43353
rect 32541 43350 32593 43353
rect 32752 43350 32804 43353
rect 34284 43350 34336 43353
rect 34495 43350 34547 43353
rect 31486 43304 31538 43350
rect 31697 43304 31749 43350
rect 31909 43304 31961 43350
rect 32120 43304 32172 43350
rect 32330 43304 32382 43350
rect 32541 43304 32593 43350
rect 32752 43304 32804 43350
rect 34284 43304 34302 43350
rect 34302 43304 34336 43350
rect 34495 43304 34508 43350
rect 34508 43304 34547 43350
rect 31486 43301 31538 43304
rect 31697 43301 31749 43304
rect 31909 43301 31961 43304
rect 32120 43301 32172 43304
rect 32330 43301 32382 43304
rect 32541 43301 32593 43304
rect 32752 43301 32804 43304
rect 34284 43301 34336 43304
rect 34495 43301 34547 43304
rect 34707 43301 34759 43353
rect 34918 43301 34970 43353
rect 35220 43301 35272 43353
rect 35430 43301 35482 43353
rect 35641 43301 35693 43353
rect 35853 43301 35905 43353
rect 36064 43301 36116 43353
rect 36274 43301 36326 43353
rect 38330 43350 38382 43353
rect 38330 43304 38382 43350
rect 38330 43301 38382 43304
rect 38541 43301 38593 43353
rect 38752 43301 38804 43353
rect 39052 43350 39104 43353
rect 39232 43350 39284 43353
rect 39052 43304 39062 43350
rect 39062 43304 39104 43350
rect 39232 43304 39266 43350
rect 39266 43304 39284 43350
rect 39052 43301 39104 43304
rect 39232 43301 39284 43304
rect 33057 43126 33109 43129
rect 33237 43126 33289 43129
rect 33057 43080 33109 43126
rect 33237 43080 33289 43126
rect 33057 43077 33109 43080
rect 33237 43077 33289 43080
rect 33819 43126 33871 43137
rect 33999 43126 34051 43137
rect 33819 43085 33833 43126
rect 33833 43085 33871 43126
rect 33999 43085 34039 43126
rect 34039 43085 34051 43126
rect 35332 43039 35384 43051
rect 35543 43039 35595 43051
rect 35754 43039 35806 43051
rect 35965 43039 36017 43051
rect 36176 43039 36228 43051
rect 37891 43039 37943 43063
rect 38071 43039 38123 43063
rect 35332 42999 35384 43039
rect 35543 42999 35580 43039
rect 35580 42999 35595 43039
rect 35754 42999 35786 43039
rect 35786 42999 35806 43039
rect 35965 42999 35992 43039
rect 35992 42999 36017 43039
rect 36176 42999 36198 43039
rect 36198 42999 36228 43039
rect 37891 43011 37909 43039
rect 37909 43011 37943 43039
rect 38071 43011 38072 43039
rect 38072 43011 38123 43039
rect 34267 42856 34302 42891
rect 34302 42856 34319 42891
rect 34447 42856 34451 42891
rect 34451 42856 34499 42891
rect 34627 42856 34658 42891
rect 34658 42856 34679 42891
rect 34267 42839 34319 42856
rect 34447 42839 34499 42856
rect 34627 42839 34679 42856
rect 33057 42678 33109 42681
rect 33237 42678 33289 42681
rect 33057 42632 33109 42678
rect 33237 42632 33289 42678
rect 33057 42629 33109 42632
rect 33237 42629 33289 42632
rect 36678 42764 36697 42816
rect 36697 42764 36730 42816
rect 36961 42815 37013 42823
rect 37172 42815 37224 42823
rect 36961 42771 36971 42815
rect 36971 42771 37013 42815
rect 37172 42771 37206 42815
rect 37206 42771 37224 42815
rect 37384 42771 37436 42823
rect 37595 42771 37647 42823
rect 40253 43301 40305 43353
rect 40433 43301 40485 43353
rect 43790 43301 43842 43353
rect 44001 43301 44053 43353
rect 44213 43350 44265 43353
rect 44213 43304 44236 43350
rect 44236 43304 44265 43350
rect 44213 43301 44265 43304
rect 44424 43301 44476 43353
rect 44834 43350 44886 43353
rect 45045 43350 45097 43353
rect 45256 43350 45308 43353
rect 44834 43304 44858 43350
rect 44858 43304 44886 43350
rect 45045 43304 45084 43350
rect 45084 43304 45097 43350
rect 45256 43304 45264 43350
rect 45264 43304 45308 43350
rect 44834 43301 44886 43304
rect 45045 43301 45097 43304
rect 45256 43301 45308 43304
rect 48838 43301 48890 43353
rect 49048 43301 49100 43353
rect 49259 43301 49311 43353
rect 49471 43301 49523 43353
rect 49682 43301 49734 43353
rect 49892 43301 49944 43353
rect 50346 43301 50398 43353
rect 50557 43350 50609 43353
rect 50768 43350 50820 43353
rect 52316 43350 52368 43353
rect 52527 43350 52579 43353
rect 52738 43350 52790 43353
rect 52948 43350 53000 43353
rect 53159 43350 53211 43353
rect 53371 43350 53423 43353
rect 53582 43350 53634 43353
rect 50557 43304 50571 43350
rect 50571 43304 50609 43350
rect 50768 43304 50777 43350
rect 50777 43304 50820 43350
rect 52316 43304 52368 43350
rect 52527 43304 52579 43350
rect 52738 43304 52790 43350
rect 52948 43304 53000 43350
rect 53159 43304 53211 43350
rect 53371 43304 53423 43350
rect 53582 43304 53634 43350
rect 50557 43301 50609 43304
rect 50768 43301 50820 43304
rect 39775 43080 39786 43115
rect 39786 43080 39827 43115
rect 39775 43063 39827 43080
rect 39994 42848 40046 42900
rect 39994 42662 40046 42714
rect 52316 43301 52368 43304
rect 52527 43301 52579 43304
rect 52738 43301 52790 43304
rect 52948 43301 53000 43304
rect 53159 43301 53211 43304
rect 53371 43301 53423 43304
rect 53582 43301 53634 43304
rect 53792 43301 53844 43353
rect 54003 43301 54055 43353
rect 54214 43301 54266 43353
rect 54855 43301 54907 43353
rect 55066 43301 55118 43353
rect 55278 43350 55330 43353
rect 55278 43304 55279 43350
rect 55279 43304 55325 43350
rect 55325 43304 55330 43350
rect 55278 43301 55330 43304
rect 55489 43301 55541 43353
rect 41935 43063 41987 43115
rect 51073 43126 51125 43129
rect 51253 43126 51305 43129
rect 43445 42832 43497 42884
rect 51073 43080 51086 43126
rect 51086 43080 51125 43126
rect 51253 43080 51292 43126
rect 51292 43080 51305 43126
rect 48943 43039 48995 43054
rect 49154 43039 49206 43054
rect 49365 43039 49417 43054
rect 49576 43039 49628 43054
rect 49787 43039 49839 43054
rect 48943 43002 48984 43039
rect 48984 43002 48995 43039
rect 49154 43002 49190 43039
rect 49190 43002 49206 43039
rect 49365 43002 49396 43039
rect 49396 43002 49417 43039
rect 49576 43002 49602 43039
rect 49602 43002 49628 43039
rect 49787 43002 49839 43039
rect 51073 43077 51125 43080
rect 51253 43077 51305 43080
rect 44939 42856 44971 42891
rect 44971 42856 44991 42891
rect 45151 42856 45197 42891
rect 45197 42856 45203 42891
rect 48596 42895 48648 42947
rect 44939 42839 44991 42856
rect 45151 42839 45203 42856
rect 45597 42737 45604 42775
rect 45604 42737 45649 42775
rect 45597 42723 45649 42737
rect 50300 42839 50352 42891
rect 50511 42856 50513 42891
rect 50513 42856 50563 42891
rect 50511 42839 50563 42856
rect 50722 42839 50774 42891
rect 48596 42677 48648 42729
rect 51835 43080 51887 43122
rect 52015 43080 52067 43122
rect 51835 43070 51887 43080
rect 52015 43070 52067 43080
rect 35332 42545 35384 42591
rect 35543 42545 35580 42591
rect 35580 42545 35595 42591
rect 35754 42545 35786 42591
rect 35786 42545 35806 42591
rect 35965 42545 35992 42591
rect 35992 42545 36017 42591
rect 36176 42545 36198 42591
rect 36198 42545 36228 42591
rect 37891 42545 37909 42589
rect 37909 42545 37943 42589
rect 38071 42545 38072 42589
rect 38072 42545 38123 42589
rect 48943 42545 48984 42591
rect 48984 42545 48995 42591
rect 49154 42545 49190 42591
rect 49190 42545 49206 42591
rect 49365 42545 49396 42591
rect 49396 42545 49417 42591
rect 49576 42545 49602 42591
rect 49602 42545 49628 42591
rect 49787 42545 49839 42591
rect 51835 42632 51887 42659
rect 52015 42632 52067 42659
rect 51835 42607 51887 42632
rect 52015 42607 52067 42632
rect 35332 42539 35384 42545
rect 35543 42539 35595 42545
rect 35754 42539 35806 42545
rect 35965 42539 36017 42545
rect 36176 42539 36228 42545
rect 37891 42537 37943 42545
rect 38071 42537 38123 42545
rect 27790 42401 27842 42453
rect 28001 42401 28053 42453
rect 28212 42401 28264 42453
rect 28423 42401 28475 42453
rect 28634 42401 28686 42453
rect 28845 42450 28897 42453
rect 28845 42404 28856 42450
rect 28856 42404 28897 42450
rect 28845 42401 28897 42404
rect 29056 42401 29108 42453
rect 29582 42401 29634 42453
rect 29793 42450 29845 42453
rect 29793 42404 29798 42450
rect 29798 42404 29844 42450
rect 29844 42404 29845 42450
rect 29793 42401 29845 42404
rect 30005 42401 30057 42453
rect 30216 42401 30268 42453
rect 30854 42401 30906 42453
rect 31065 42401 31117 42453
rect 31276 42401 31328 42453
rect 31486 42401 31538 42453
rect 31697 42401 31749 42453
rect 31909 42401 31961 42453
rect 32120 42401 32172 42453
rect 32330 42401 32382 42453
rect 32541 42401 32593 42453
rect 32752 42401 32804 42453
rect 48943 42539 48995 42545
rect 49154 42539 49206 42545
rect 49365 42539 49417 42545
rect 49576 42539 49628 42545
rect 49787 42539 49839 42545
rect 34755 42401 34807 42453
rect 34935 42450 34987 42453
rect 34935 42404 34962 42450
rect 34962 42404 34987 42450
rect 34935 42401 34987 42404
rect 50138 42450 50190 42453
rect 50138 42404 50160 42450
rect 50160 42404 50190 42450
rect 50138 42401 50190 42404
rect 50318 42401 50370 42453
rect 35332 42309 35384 42315
rect 35543 42309 35595 42315
rect 35754 42309 35806 42315
rect 35965 42309 36017 42315
rect 36176 42309 36228 42315
rect 37891 42309 37943 42317
rect 38071 42309 38123 42317
rect 52316 42401 52368 42453
rect 52527 42401 52579 42453
rect 52738 42401 52790 42453
rect 52948 42401 53000 42453
rect 53159 42401 53211 42453
rect 53371 42401 53423 42453
rect 53582 42401 53634 42453
rect 53792 42401 53844 42453
rect 54003 42401 54055 42453
rect 54214 42401 54266 42453
rect 54855 42401 54907 42453
rect 55066 42401 55118 42453
rect 55278 42450 55330 42453
rect 55278 42404 55279 42450
rect 55279 42404 55325 42450
rect 55325 42404 55330 42450
rect 55278 42401 55330 42404
rect 55489 42401 55541 42453
rect 56015 42401 56067 42453
rect 56226 42450 56278 42453
rect 56226 42404 56267 42450
rect 56267 42404 56278 42450
rect 56226 42401 56278 42404
rect 56437 42401 56489 42453
rect 56648 42401 56700 42453
rect 56859 42401 56911 42453
rect 57070 42401 57122 42453
rect 57281 42401 57333 42453
rect 48943 42309 48995 42315
rect 49154 42309 49206 42315
rect 49365 42309 49417 42315
rect 49576 42309 49628 42315
rect 49787 42309 49839 42315
rect 33057 42222 33109 42225
rect 33237 42222 33289 42225
rect 35332 42263 35384 42309
rect 35543 42263 35580 42309
rect 35580 42263 35595 42309
rect 35754 42263 35786 42309
rect 35786 42263 35806 42309
rect 35965 42263 35992 42309
rect 35992 42263 36017 42309
rect 36176 42263 36198 42309
rect 36198 42263 36228 42309
rect 37891 42265 37909 42309
rect 37909 42265 37943 42309
rect 38071 42265 38072 42309
rect 38072 42265 38123 42309
rect 33057 42176 33109 42222
rect 33237 42176 33289 42222
rect 33057 42173 33109 42176
rect 33237 42173 33289 42176
rect 33057 41774 33109 41777
rect 33237 41774 33289 41777
rect 33057 41728 33109 41774
rect 33237 41728 33289 41774
rect 33057 41725 33109 41728
rect 33237 41725 33289 41728
rect 29582 41501 29634 41553
rect 29793 41550 29845 41553
rect 29793 41504 29798 41550
rect 29798 41504 29844 41550
rect 29844 41504 29845 41550
rect 29793 41501 29845 41504
rect 30005 41501 30057 41553
rect 30216 41501 30268 41553
rect 34267 41998 34319 42015
rect 34447 41998 34499 42015
rect 34627 41998 34679 42015
rect 34267 41963 34302 41998
rect 34302 41963 34319 41998
rect 34447 41963 34451 41998
rect 34451 41963 34499 41998
rect 34627 41963 34658 41998
rect 34658 41963 34679 41998
rect 36678 42038 36697 42090
rect 36697 42038 36730 42090
rect 48943 42263 48984 42309
rect 48984 42263 48995 42309
rect 49154 42263 49190 42309
rect 49190 42263 49206 42309
rect 49365 42263 49396 42309
rect 49396 42263 49417 42309
rect 49576 42263 49602 42309
rect 49602 42263 49628 42309
rect 49787 42263 49839 42309
rect 39994 42140 40046 42192
rect 36961 42039 36971 42083
rect 36971 42039 37013 42083
rect 37172 42039 37206 42083
rect 37206 42039 37224 42083
rect 36961 42031 37013 42039
rect 37172 42031 37224 42039
rect 37384 42031 37436 42083
rect 37595 42031 37647 42083
rect 35332 41815 35384 41855
rect 35543 41815 35580 41855
rect 35580 41815 35595 41855
rect 35754 41815 35786 41855
rect 35786 41815 35806 41855
rect 35965 41815 35992 41855
rect 35992 41815 36017 41855
rect 36176 41815 36198 41855
rect 36198 41815 36228 41855
rect 37891 41815 37909 41843
rect 37909 41815 37943 41843
rect 38071 41815 38072 41843
rect 38072 41815 38123 41843
rect 35332 41803 35384 41815
rect 35543 41803 35595 41815
rect 35754 41803 35806 41815
rect 35965 41803 36017 41815
rect 36176 41803 36228 41815
rect 33819 41728 33833 41769
rect 33833 41728 33871 41769
rect 33999 41728 34039 41769
rect 34039 41728 34051 41769
rect 37891 41791 37943 41815
rect 38071 41791 38123 41815
rect 33819 41717 33871 41728
rect 33999 41717 34051 41728
rect 30854 41501 30906 41553
rect 31065 41501 31117 41553
rect 31276 41501 31328 41553
rect 31486 41550 31538 41553
rect 31697 41550 31749 41553
rect 31909 41550 31961 41553
rect 32120 41550 32172 41553
rect 32330 41550 32382 41553
rect 32541 41550 32593 41553
rect 32752 41550 32804 41553
rect 34284 41550 34336 41553
rect 34495 41550 34547 41553
rect 31486 41504 31538 41550
rect 31697 41504 31749 41550
rect 31909 41504 31961 41550
rect 32120 41504 32172 41550
rect 32330 41504 32382 41550
rect 32541 41504 32593 41550
rect 32752 41504 32804 41550
rect 34284 41504 34302 41550
rect 34302 41504 34336 41550
rect 34495 41504 34508 41550
rect 34508 41504 34547 41550
rect 31486 41501 31538 41504
rect 31697 41501 31749 41504
rect 31909 41501 31961 41504
rect 32120 41501 32172 41504
rect 32330 41501 32382 41504
rect 32541 41501 32593 41504
rect 32752 41501 32804 41504
rect 34284 41501 34336 41504
rect 34495 41501 34547 41504
rect 34707 41501 34759 41553
rect 34918 41501 34970 41553
rect 35220 41501 35272 41553
rect 35430 41501 35482 41553
rect 35641 41501 35693 41553
rect 35853 41501 35905 41553
rect 36064 41501 36116 41553
rect 36274 41501 36326 41553
rect 38330 41550 38382 41553
rect 38330 41504 38382 41550
rect 38330 41501 38382 41504
rect 38541 41501 38593 41553
rect 38752 41501 38804 41553
rect 39052 41550 39104 41553
rect 39232 41550 39284 41553
rect 39052 41504 39062 41550
rect 39062 41504 39104 41550
rect 39232 41504 39266 41550
rect 39266 41504 39284 41550
rect 39052 41501 39104 41504
rect 39232 41501 39284 41504
rect 33057 41326 33109 41329
rect 33237 41326 33289 41329
rect 33057 41280 33109 41326
rect 33237 41280 33289 41326
rect 33057 41277 33109 41280
rect 33237 41277 33289 41280
rect 33819 41326 33871 41337
rect 33999 41326 34051 41337
rect 33819 41285 33833 41326
rect 33833 41285 33871 41326
rect 33999 41285 34039 41326
rect 34039 41285 34051 41326
rect 35332 41239 35384 41251
rect 35543 41239 35595 41251
rect 35754 41239 35806 41251
rect 35965 41239 36017 41251
rect 36176 41239 36228 41251
rect 37891 41239 37943 41263
rect 38071 41239 38123 41263
rect 35332 41199 35384 41239
rect 35543 41199 35580 41239
rect 35580 41199 35595 41239
rect 35754 41199 35786 41239
rect 35786 41199 35806 41239
rect 35965 41199 35992 41239
rect 35992 41199 36017 41239
rect 36176 41199 36198 41239
rect 36198 41199 36228 41239
rect 37891 41211 37909 41239
rect 37909 41211 37943 41239
rect 38071 41211 38072 41239
rect 38072 41211 38123 41239
rect 34267 41056 34302 41091
rect 34302 41056 34319 41091
rect 34447 41056 34451 41091
rect 34451 41056 34499 41091
rect 34627 41056 34658 41091
rect 34658 41056 34679 41091
rect 34267 41039 34319 41056
rect 34447 41039 34499 41056
rect 34627 41039 34679 41056
rect 33057 40878 33109 40881
rect 33237 40878 33289 40881
rect 33057 40832 33109 40878
rect 33237 40832 33289 40878
rect 33057 40829 33109 40832
rect 33237 40829 33289 40832
rect 36678 40964 36697 41016
rect 36697 40964 36730 41016
rect 36961 41015 37013 41023
rect 37172 41015 37224 41023
rect 36961 40971 36971 41015
rect 36971 40971 37013 41015
rect 37172 40971 37206 41015
rect 37206 40971 37224 41015
rect 37384 40971 37436 41023
rect 37595 40971 37647 41023
rect 39994 41954 40046 42006
rect 39775 41774 39827 41791
rect 39775 41739 39786 41774
rect 39786 41739 39827 41774
rect 43445 41970 43497 42022
rect 41935 41739 41987 41791
rect 45975 42079 46027 42131
rect 48596 42125 48648 42177
rect 51835 42222 51887 42247
rect 52015 42222 52067 42247
rect 51835 42195 51887 42222
rect 52015 42195 52067 42222
rect 44939 41998 44991 42015
rect 45151 41998 45203 42015
rect 44939 41963 44971 41998
rect 44971 41963 44991 41998
rect 45151 41963 45197 41998
rect 45197 41963 45203 41998
rect 48596 41907 48648 41959
rect 50300 41963 50352 42015
rect 50511 41998 50563 42015
rect 50511 41963 50513 41998
rect 50513 41963 50563 41998
rect 50722 41963 50774 42015
rect 48943 41815 48984 41852
rect 48984 41815 48995 41852
rect 49154 41815 49190 41852
rect 49190 41815 49206 41852
rect 49365 41815 49396 41852
rect 49396 41815 49417 41852
rect 49576 41815 49602 41852
rect 49602 41815 49628 41852
rect 49787 41815 49839 41852
rect 48943 41800 48995 41815
rect 49154 41800 49206 41815
rect 49365 41800 49417 41815
rect 49576 41800 49628 41815
rect 49787 41800 49839 41815
rect 51073 41774 51125 41777
rect 51253 41774 51305 41777
rect 51073 41728 51086 41774
rect 51086 41728 51125 41774
rect 51253 41728 51292 41774
rect 51292 41728 51305 41774
rect 51073 41725 51125 41728
rect 51253 41725 51305 41728
rect 51835 41774 51887 41784
rect 52015 41774 52067 41784
rect 51835 41732 51887 41774
rect 52015 41732 52067 41774
rect 40253 41501 40305 41553
rect 40433 41501 40485 41553
rect 43790 41501 43842 41553
rect 44001 41501 44053 41553
rect 44213 41550 44265 41553
rect 44213 41504 44236 41550
rect 44236 41504 44265 41550
rect 44213 41501 44265 41504
rect 44424 41501 44476 41553
rect 44834 41550 44886 41553
rect 45045 41550 45097 41553
rect 45256 41550 45308 41553
rect 44834 41504 44858 41550
rect 44858 41504 44886 41550
rect 45045 41504 45084 41550
rect 45084 41504 45097 41550
rect 45256 41504 45264 41550
rect 45264 41504 45308 41550
rect 44834 41501 44886 41504
rect 45045 41501 45097 41504
rect 45256 41501 45308 41504
rect 48838 41501 48890 41553
rect 49048 41501 49100 41553
rect 49259 41501 49311 41553
rect 49471 41501 49523 41553
rect 49682 41501 49734 41553
rect 49892 41501 49944 41553
rect 50346 41501 50398 41553
rect 50557 41550 50609 41553
rect 50768 41550 50820 41553
rect 52316 41550 52368 41553
rect 52527 41550 52579 41553
rect 52738 41550 52790 41553
rect 52948 41550 53000 41553
rect 53159 41550 53211 41553
rect 53371 41550 53423 41553
rect 53582 41550 53634 41553
rect 50557 41504 50571 41550
rect 50571 41504 50609 41550
rect 50768 41504 50777 41550
rect 50777 41504 50820 41550
rect 52316 41504 52368 41550
rect 52527 41504 52579 41550
rect 52738 41504 52790 41550
rect 52948 41504 53000 41550
rect 53159 41504 53211 41550
rect 53371 41504 53423 41550
rect 53582 41504 53634 41550
rect 50557 41501 50609 41504
rect 50768 41501 50820 41504
rect 39775 41280 39786 41315
rect 39786 41280 39827 41315
rect 39775 41263 39827 41280
rect 39994 41048 40046 41100
rect 39994 40862 40046 40914
rect 52316 41501 52368 41504
rect 52527 41501 52579 41504
rect 52738 41501 52790 41504
rect 52948 41501 53000 41504
rect 53159 41501 53211 41504
rect 53371 41501 53423 41504
rect 53582 41501 53634 41504
rect 53792 41501 53844 41553
rect 54003 41501 54055 41553
rect 54214 41501 54266 41553
rect 54855 41501 54907 41553
rect 55066 41501 55118 41553
rect 55278 41550 55330 41553
rect 55278 41504 55279 41550
rect 55279 41504 55325 41550
rect 55325 41504 55330 41550
rect 55278 41501 55330 41504
rect 55489 41501 55541 41553
rect 41935 41263 41987 41315
rect 51073 41326 51125 41329
rect 51253 41326 51305 41329
rect 43445 41032 43497 41084
rect 51073 41280 51086 41326
rect 51086 41280 51125 41326
rect 51253 41280 51292 41326
rect 51292 41280 51305 41326
rect 48943 41239 48995 41254
rect 49154 41239 49206 41254
rect 49365 41239 49417 41254
rect 49576 41239 49628 41254
rect 49787 41239 49839 41254
rect 48943 41202 48984 41239
rect 48984 41202 48995 41239
rect 49154 41202 49190 41239
rect 49190 41202 49206 41239
rect 49365 41202 49396 41239
rect 49396 41202 49417 41239
rect 49576 41202 49602 41239
rect 49602 41202 49628 41239
rect 49787 41202 49839 41239
rect 51073 41277 51125 41280
rect 51253 41277 51305 41280
rect 44939 41056 44971 41091
rect 44971 41056 44991 41091
rect 45151 41056 45197 41091
rect 45197 41056 45203 41091
rect 48596 41095 48648 41147
rect 44939 41039 44991 41056
rect 45151 41039 45203 41056
rect 46353 40923 46405 40975
rect 50300 41039 50352 41091
rect 50511 41056 50513 41091
rect 50513 41056 50563 41091
rect 50511 41039 50563 41056
rect 50722 41039 50774 41091
rect 48596 40877 48648 40929
rect 51835 41280 51887 41322
rect 52015 41280 52067 41322
rect 51835 41270 51887 41280
rect 52015 41270 52067 41280
rect 35332 40745 35384 40791
rect 35543 40745 35580 40791
rect 35580 40745 35595 40791
rect 35754 40745 35786 40791
rect 35786 40745 35806 40791
rect 35965 40745 35992 40791
rect 35992 40745 36017 40791
rect 36176 40745 36198 40791
rect 36198 40745 36228 40791
rect 37891 40745 37909 40789
rect 37909 40745 37943 40789
rect 38071 40745 38072 40789
rect 38072 40745 38123 40789
rect 48943 40745 48984 40791
rect 48984 40745 48995 40791
rect 49154 40745 49190 40791
rect 49190 40745 49206 40791
rect 49365 40745 49396 40791
rect 49396 40745 49417 40791
rect 49576 40745 49602 40791
rect 49602 40745 49628 40791
rect 49787 40745 49839 40791
rect 51835 40832 51887 40859
rect 52015 40832 52067 40859
rect 51835 40807 51887 40832
rect 52015 40807 52067 40832
rect 35332 40739 35384 40745
rect 35543 40739 35595 40745
rect 35754 40739 35806 40745
rect 35965 40739 36017 40745
rect 36176 40739 36228 40745
rect 37891 40737 37943 40745
rect 38071 40737 38123 40745
rect 27790 40601 27842 40653
rect 28001 40601 28053 40653
rect 28212 40601 28264 40653
rect 28423 40601 28475 40653
rect 28634 40601 28686 40653
rect 28845 40650 28897 40653
rect 28845 40604 28856 40650
rect 28856 40604 28897 40650
rect 28845 40601 28897 40604
rect 29056 40601 29108 40653
rect 29582 40601 29634 40653
rect 29793 40650 29845 40653
rect 29793 40604 29798 40650
rect 29798 40604 29844 40650
rect 29844 40604 29845 40650
rect 29793 40601 29845 40604
rect 30005 40601 30057 40653
rect 30216 40601 30268 40653
rect 30854 40601 30906 40653
rect 31065 40601 31117 40653
rect 31276 40601 31328 40653
rect 31486 40601 31538 40653
rect 31697 40601 31749 40653
rect 31909 40601 31961 40653
rect 32120 40601 32172 40653
rect 32330 40601 32382 40653
rect 32541 40601 32593 40653
rect 32752 40601 32804 40653
rect 48943 40739 48995 40745
rect 49154 40739 49206 40745
rect 49365 40739 49417 40745
rect 49576 40739 49628 40745
rect 49787 40739 49839 40745
rect 34755 40601 34807 40653
rect 34935 40650 34987 40653
rect 34935 40604 34962 40650
rect 34962 40604 34987 40650
rect 34935 40601 34987 40604
rect 50138 40650 50190 40653
rect 50138 40604 50160 40650
rect 50160 40604 50190 40650
rect 50138 40601 50190 40604
rect 50318 40601 50370 40653
rect 35332 40509 35384 40515
rect 35543 40509 35595 40515
rect 35754 40509 35806 40515
rect 35965 40509 36017 40515
rect 36176 40509 36228 40515
rect 37891 40509 37943 40517
rect 38071 40509 38123 40517
rect 52316 40601 52368 40653
rect 52527 40601 52579 40653
rect 52738 40601 52790 40653
rect 52948 40601 53000 40653
rect 53159 40601 53211 40653
rect 53371 40601 53423 40653
rect 53582 40601 53634 40653
rect 53792 40601 53844 40653
rect 54003 40601 54055 40653
rect 54214 40601 54266 40653
rect 54855 40601 54907 40653
rect 55066 40601 55118 40653
rect 55278 40650 55330 40653
rect 55278 40604 55279 40650
rect 55279 40604 55325 40650
rect 55325 40604 55330 40650
rect 55278 40601 55330 40604
rect 55489 40601 55541 40653
rect 56015 40601 56067 40653
rect 56226 40650 56278 40653
rect 56226 40604 56267 40650
rect 56267 40604 56278 40650
rect 56226 40601 56278 40604
rect 56437 40601 56489 40653
rect 56648 40601 56700 40653
rect 56859 40601 56911 40653
rect 57070 40601 57122 40653
rect 57281 40601 57333 40653
rect 48943 40509 48995 40515
rect 49154 40509 49206 40515
rect 49365 40509 49417 40515
rect 49576 40509 49628 40515
rect 49787 40509 49839 40515
rect 33057 40422 33109 40425
rect 33237 40422 33289 40425
rect 35332 40463 35384 40509
rect 35543 40463 35580 40509
rect 35580 40463 35595 40509
rect 35754 40463 35786 40509
rect 35786 40463 35806 40509
rect 35965 40463 35992 40509
rect 35992 40463 36017 40509
rect 36176 40463 36198 40509
rect 36198 40463 36228 40509
rect 37891 40465 37909 40509
rect 37909 40465 37943 40509
rect 38071 40465 38072 40509
rect 38072 40465 38123 40509
rect 33057 40376 33109 40422
rect 33237 40376 33289 40422
rect 33057 40373 33109 40376
rect 33237 40373 33289 40376
rect 33057 39974 33109 39977
rect 33237 39974 33289 39977
rect 33057 39928 33109 39974
rect 33237 39928 33289 39974
rect 33057 39925 33109 39928
rect 33237 39925 33289 39928
rect 29582 39701 29634 39753
rect 29793 39750 29845 39753
rect 29793 39704 29798 39750
rect 29798 39704 29844 39750
rect 29844 39704 29845 39750
rect 29793 39701 29845 39704
rect 30005 39701 30057 39753
rect 30216 39701 30268 39753
rect 34267 40198 34319 40215
rect 34447 40198 34499 40215
rect 34627 40198 34679 40215
rect 34267 40163 34302 40198
rect 34302 40163 34319 40198
rect 34447 40163 34451 40198
rect 34451 40163 34499 40198
rect 34627 40163 34658 40198
rect 34658 40163 34679 40198
rect 36678 40238 36697 40290
rect 36697 40238 36730 40290
rect 48943 40463 48984 40509
rect 48984 40463 48995 40509
rect 49154 40463 49190 40509
rect 49190 40463 49206 40509
rect 49365 40463 49396 40509
rect 49396 40463 49417 40509
rect 49576 40463 49602 40509
rect 49602 40463 49628 40509
rect 49787 40463 49839 40509
rect 39994 40340 40046 40392
rect 36961 40239 36971 40283
rect 36971 40239 37013 40283
rect 37172 40239 37206 40283
rect 37206 40239 37224 40283
rect 36961 40231 37013 40239
rect 37172 40231 37224 40239
rect 37384 40231 37436 40283
rect 37595 40231 37647 40283
rect 35332 40015 35384 40055
rect 35543 40015 35580 40055
rect 35580 40015 35595 40055
rect 35754 40015 35786 40055
rect 35786 40015 35806 40055
rect 35965 40015 35992 40055
rect 35992 40015 36017 40055
rect 36176 40015 36198 40055
rect 36198 40015 36228 40055
rect 37891 40015 37909 40043
rect 37909 40015 37943 40043
rect 38071 40015 38072 40043
rect 38072 40015 38123 40043
rect 35332 40003 35384 40015
rect 35543 40003 35595 40015
rect 35754 40003 35806 40015
rect 35965 40003 36017 40015
rect 36176 40003 36228 40015
rect 33819 39928 33833 39969
rect 33833 39928 33871 39969
rect 33999 39928 34039 39969
rect 34039 39928 34051 39969
rect 37891 39991 37943 40015
rect 38071 39991 38123 40015
rect 33819 39917 33871 39928
rect 33999 39917 34051 39928
rect 30854 39701 30906 39753
rect 31065 39701 31117 39753
rect 31276 39701 31328 39753
rect 31486 39750 31538 39753
rect 31697 39750 31749 39753
rect 31909 39750 31961 39753
rect 32120 39750 32172 39753
rect 32330 39750 32382 39753
rect 32541 39750 32593 39753
rect 32752 39750 32804 39753
rect 34284 39750 34336 39753
rect 34495 39750 34547 39753
rect 31486 39704 31538 39750
rect 31697 39704 31749 39750
rect 31909 39704 31961 39750
rect 32120 39704 32172 39750
rect 32330 39704 32382 39750
rect 32541 39704 32593 39750
rect 32752 39704 32804 39750
rect 34284 39704 34302 39750
rect 34302 39704 34336 39750
rect 34495 39704 34508 39750
rect 34508 39704 34547 39750
rect 31486 39701 31538 39704
rect 31697 39701 31749 39704
rect 31909 39701 31961 39704
rect 32120 39701 32172 39704
rect 32330 39701 32382 39704
rect 32541 39701 32593 39704
rect 32752 39701 32804 39704
rect 34284 39701 34336 39704
rect 34495 39701 34547 39704
rect 34707 39701 34759 39753
rect 34918 39701 34970 39753
rect 35220 39701 35272 39753
rect 35430 39701 35482 39753
rect 35641 39701 35693 39753
rect 35853 39701 35905 39753
rect 36064 39701 36116 39753
rect 36274 39701 36326 39753
rect 38330 39750 38382 39753
rect 38330 39704 38382 39750
rect 38330 39701 38382 39704
rect 38541 39701 38593 39753
rect 38752 39701 38804 39753
rect 39052 39750 39104 39753
rect 39232 39750 39284 39753
rect 39052 39704 39062 39750
rect 39062 39704 39104 39750
rect 39232 39704 39266 39750
rect 39266 39704 39284 39750
rect 39052 39701 39104 39704
rect 39232 39701 39284 39704
rect 33057 39526 33109 39529
rect 33237 39526 33289 39529
rect 33057 39480 33109 39526
rect 33237 39480 33289 39526
rect 33057 39477 33109 39480
rect 33237 39477 33289 39480
rect 33819 39526 33871 39537
rect 33999 39526 34051 39537
rect 33819 39485 33833 39526
rect 33833 39485 33871 39526
rect 33999 39485 34039 39526
rect 34039 39485 34051 39526
rect 35332 39439 35384 39451
rect 35543 39439 35595 39451
rect 35754 39439 35806 39451
rect 35965 39439 36017 39451
rect 36176 39439 36228 39451
rect 37891 39439 37943 39463
rect 38071 39439 38123 39463
rect 35332 39399 35384 39439
rect 35543 39399 35580 39439
rect 35580 39399 35595 39439
rect 35754 39399 35786 39439
rect 35786 39399 35806 39439
rect 35965 39399 35992 39439
rect 35992 39399 36017 39439
rect 36176 39399 36198 39439
rect 36198 39399 36228 39439
rect 37891 39411 37909 39439
rect 37909 39411 37943 39439
rect 38071 39411 38072 39439
rect 38072 39411 38123 39439
rect 34267 39256 34302 39291
rect 34302 39256 34319 39291
rect 34447 39256 34451 39291
rect 34451 39256 34499 39291
rect 34627 39256 34658 39291
rect 34658 39256 34679 39291
rect 34267 39239 34319 39256
rect 34447 39239 34499 39256
rect 34627 39239 34679 39256
rect 33057 39078 33109 39081
rect 33237 39078 33289 39081
rect 33057 39032 33109 39078
rect 33237 39032 33289 39078
rect 33057 39029 33109 39032
rect 33237 39029 33289 39032
rect 36678 39164 36697 39216
rect 36697 39164 36730 39216
rect 36961 39215 37013 39223
rect 37172 39215 37224 39223
rect 36961 39171 36971 39215
rect 36971 39171 37013 39215
rect 37172 39171 37206 39215
rect 37206 39171 37224 39215
rect 37384 39171 37436 39223
rect 37595 39171 37647 39223
rect 39994 40154 40046 40206
rect 39775 39974 39827 39991
rect 39775 39939 39786 39974
rect 39786 39939 39827 39974
rect 43445 40170 43497 40222
rect 41935 39939 41987 39991
rect 46731 40279 46783 40331
rect 48596 40325 48648 40377
rect 51835 40422 51887 40447
rect 52015 40422 52067 40447
rect 51835 40395 51887 40422
rect 52015 40395 52067 40422
rect 44939 40198 44991 40215
rect 45151 40198 45203 40215
rect 44939 40163 44971 40198
rect 44971 40163 44991 40198
rect 45151 40163 45197 40198
rect 45197 40163 45203 40198
rect 48596 40107 48648 40159
rect 50300 40163 50352 40215
rect 50511 40198 50563 40215
rect 50511 40163 50513 40198
rect 50513 40163 50563 40198
rect 50722 40163 50774 40215
rect 48943 40015 48984 40052
rect 48984 40015 48995 40052
rect 49154 40015 49190 40052
rect 49190 40015 49206 40052
rect 49365 40015 49396 40052
rect 49396 40015 49417 40052
rect 49576 40015 49602 40052
rect 49602 40015 49628 40052
rect 49787 40015 49839 40052
rect 48943 40000 48995 40015
rect 49154 40000 49206 40015
rect 49365 40000 49417 40015
rect 49576 40000 49628 40015
rect 49787 40000 49839 40015
rect 51073 39974 51125 39977
rect 51253 39974 51305 39977
rect 51073 39928 51086 39974
rect 51086 39928 51125 39974
rect 51253 39928 51292 39974
rect 51292 39928 51305 39974
rect 51073 39925 51125 39928
rect 51253 39925 51305 39928
rect 51835 39974 51887 39984
rect 52015 39974 52067 39984
rect 51835 39932 51887 39974
rect 52015 39932 52067 39974
rect 40253 39701 40305 39753
rect 40433 39701 40485 39753
rect 43790 39701 43842 39753
rect 44001 39701 44053 39753
rect 44213 39750 44265 39753
rect 44213 39704 44236 39750
rect 44236 39704 44265 39750
rect 44213 39701 44265 39704
rect 44424 39701 44476 39753
rect 44834 39750 44886 39753
rect 45045 39750 45097 39753
rect 45256 39750 45308 39753
rect 44834 39704 44858 39750
rect 44858 39704 44886 39750
rect 45045 39704 45084 39750
rect 45084 39704 45097 39750
rect 45256 39704 45264 39750
rect 45264 39704 45308 39750
rect 44834 39701 44886 39704
rect 45045 39701 45097 39704
rect 45256 39701 45308 39704
rect 48838 39701 48890 39753
rect 49048 39701 49100 39753
rect 49259 39701 49311 39753
rect 49471 39701 49523 39753
rect 49682 39701 49734 39753
rect 49892 39701 49944 39753
rect 50346 39701 50398 39753
rect 50557 39750 50609 39753
rect 50768 39750 50820 39753
rect 52316 39750 52368 39753
rect 52527 39750 52579 39753
rect 52738 39750 52790 39753
rect 52948 39750 53000 39753
rect 53159 39750 53211 39753
rect 53371 39750 53423 39753
rect 53582 39750 53634 39753
rect 50557 39704 50571 39750
rect 50571 39704 50609 39750
rect 50768 39704 50777 39750
rect 50777 39704 50820 39750
rect 52316 39704 52368 39750
rect 52527 39704 52579 39750
rect 52738 39704 52790 39750
rect 52948 39704 53000 39750
rect 53159 39704 53211 39750
rect 53371 39704 53423 39750
rect 53582 39704 53634 39750
rect 50557 39701 50609 39704
rect 50768 39701 50820 39704
rect 39775 39480 39786 39515
rect 39786 39480 39827 39515
rect 39775 39463 39827 39480
rect 39994 39248 40046 39300
rect 39994 39062 40046 39114
rect 52316 39701 52368 39704
rect 52527 39701 52579 39704
rect 52738 39701 52790 39704
rect 52948 39701 53000 39704
rect 53159 39701 53211 39704
rect 53371 39701 53423 39704
rect 53582 39701 53634 39704
rect 53792 39701 53844 39753
rect 54003 39701 54055 39753
rect 54214 39701 54266 39753
rect 54855 39701 54907 39753
rect 55066 39701 55118 39753
rect 55278 39750 55330 39753
rect 55278 39704 55279 39750
rect 55279 39704 55325 39750
rect 55325 39704 55330 39750
rect 55278 39701 55330 39704
rect 55489 39701 55541 39753
rect 41935 39463 41987 39515
rect 51073 39526 51125 39529
rect 51253 39526 51305 39529
rect 43445 39232 43497 39284
rect 51073 39480 51086 39526
rect 51086 39480 51125 39526
rect 51253 39480 51292 39526
rect 51292 39480 51305 39526
rect 48943 39439 48995 39454
rect 49154 39439 49206 39454
rect 49365 39439 49417 39454
rect 49576 39439 49628 39454
rect 49787 39439 49839 39454
rect 48943 39402 48984 39439
rect 48984 39402 48995 39439
rect 49154 39402 49190 39439
rect 49190 39402 49206 39439
rect 49365 39402 49396 39439
rect 49396 39402 49417 39439
rect 49576 39402 49602 39439
rect 49602 39402 49628 39439
rect 49787 39402 49839 39439
rect 51073 39477 51125 39480
rect 51253 39477 51305 39480
rect 44939 39256 44971 39291
rect 44971 39256 44991 39291
rect 45151 39256 45197 39291
rect 45197 39256 45203 39291
rect 48596 39295 48648 39347
rect 44939 39239 44991 39256
rect 45151 39239 45203 39256
rect 47108 39123 47160 39175
rect 50300 39239 50352 39291
rect 50511 39256 50513 39291
rect 50513 39256 50563 39291
rect 50511 39239 50563 39256
rect 50722 39239 50774 39291
rect 48596 39077 48648 39129
rect 51835 39480 51887 39522
rect 52015 39480 52067 39522
rect 51835 39470 51887 39480
rect 52015 39470 52067 39480
rect 35332 38945 35384 38991
rect 35543 38945 35580 38991
rect 35580 38945 35595 38991
rect 35754 38945 35786 38991
rect 35786 38945 35806 38991
rect 35965 38945 35992 38991
rect 35992 38945 36017 38991
rect 36176 38945 36198 38991
rect 36198 38945 36228 38991
rect 37891 38945 37909 38989
rect 37909 38945 37943 38989
rect 38071 38945 38072 38989
rect 38072 38945 38123 38989
rect 48943 38945 48984 38991
rect 48984 38945 48995 38991
rect 49154 38945 49190 38991
rect 49190 38945 49206 38991
rect 49365 38945 49396 38991
rect 49396 38945 49417 38991
rect 49576 38945 49602 38991
rect 49602 38945 49628 38991
rect 49787 38945 49839 38991
rect 51835 39032 51887 39059
rect 52015 39032 52067 39059
rect 51835 39007 51887 39032
rect 52015 39007 52067 39032
rect 35332 38939 35384 38945
rect 35543 38939 35595 38945
rect 35754 38939 35806 38945
rect 35965 38939 36017 38945
rect 36176 38939 36228 38945
rect 37891 38937 37943 38945
rect 38071 38937 38123 38945
rect 27790 38801 27842 38853
rect 28001 38801 28053 38853
rect 28212 38801 28264 38853
rect 28423 38801 28475 38853
rect 28634 38801 28686 38853
rect 28845 38850 28897 38853
rect 28845 38804 28856 38850
rect 28856 38804 28897 38850
rect 28845 38801 28897 38804
rect 29056 38801 29108 38853
rect 29582 38801 29634 38853
rect 29793 38850 29845 38853
rect 29793 38804 29798 38850
rect 29798 38804 29844 38850
rect 29844 38804 29845 38850
rect 29793 38801 29845 38804
rect 30005 38801 30057 38853
rect 30216 38801 30268 38853
rect 30854 38801 30906 38853
rect 31065 38801 31117 38853
rect 31276 38801 31328 38853
rect 31486 38801 31538 38853
rect 31697 38801 31749 38853
rect 31909 38801 31961 38853
rect 32120 38801 32172 38853
rect 32330 38801 32382 38853
rect 32541 38801 32593 38853
rect 32752 38801 32804 38853
rect 48943 38939 48995 38945
rect 49154 38939 49206 38945
rect 49365 38939 49417 38945
rect 49576 38939 49628 38945
rect 49787 38939 49839 38945
rect 34755 38801 34807 38853
rect 34935 38850 34987 38853
rect 34935 38804 34962 38850
rect 34962 38804 34987 38850
rect 34935 38801 34987 38804
rect 50138 38850 50190 38853
rect 50138 38804 50160 38850
rect 50160 38804 50190 38850
rect 50138 38801 50190 38804
rect 50318 38801 50370 38853
rect 35332 38709 35384 38715
rect 35543 38709 35595 38715
rect 35754 38709 35806 38715
rect 35965 38709 36017 38715
rect 36176 38709 36228 38715
rect 37891 38709 37943 38717
rect 38071 38709 38123 38717
rect 52316 38801 52368 38853
rect 52527 38801 52579 38853
rect 52738 38801 52790 38853
rect 52948 38801 53000 38853
rect 53159 38801 53211 38853
rect 53371 38801 53423 38853
rect 53582 38801 53634 38853
rect 53792 38801 53844 38853
rect 54003 38801 54055 38853
rect 54214 38801 54266 38853
rect 54855 38801 54907 38853
rect 55066 38801 55118 38853
rect 55278 38850 55330 38853
rect 55278 38804 55279 38850
rect 55279 38804 55325 38850
rect 55325 38804 55330 38850
rect 55278 38801 55330 38804
rect 55489 38801 55541 38853
rect 56015 38801 56067 38853
rect 56226 38850 56278 38853
rect 56226 38804 56267 38850
rect 56267 38804 56278 38850
rect 56226 38801 56278 38804
rect 56437 38801 56489 38853
rect 56648 38801 56700 38853
rect 56859 38801 56911 38853
rect 57070 38801 57122 38853
rect 57281 38801 57333 38853
rect 48943 38709 48995 38715
rect 49154 38709 49206 38715
rect 49365 38709 49417 38715
rect 49576 38709 49628 38715
rect 49787 38709 49839 38715
rect 33057 38622 33109 38625
rect 33237 38622 33289 38625
rect 35332 38663 35384 38709
rect 35543 38663 35580 38709
rect 35580 38663 35595 38709
rect 35754 38663 35786 38709
rect 35786 38663 35806 38709
rect 35965 38663 35992 38709
rect 35992 38663 36017 38709
rect 36176 38663 36198 38709
rect 36198 38663 36228 38709
rect 37891 38665 37909 38709
rect 37909 38665 37943 38709
rect 38071 38665 38072 38709
rect 38072 38665 38123 38709
rect 33057 38576 33109 38622
rect 33237 38576 33289 38622
rect 33057 38573 33109 38576
rect 33237 38573 33289 38576
rect 33057 38174 33109 38177
rect 33237 38174 33289 38177
rect 33057 38128 33109 38174
rect 33237 38128 33289 38174
rect 33057 38125 33109 38128
rect 33237 38125 33289 38128
rect 29582 37901 29634 37953
rect 29793 37950 29845 37953
rect 29793 37904 29798 37950
rect 29798 37904 29844 37950
rect 29844 37904 29845 37950
rect 29793 37901 29845 37904
rect 30005 37901 30057 37953
rect 30216 37901 30268 37953
rect 34267 38398 34319 38415
rect 34447 38398 34499 38415
rect 34627 38398 34679 38415
rect 34267 38363 34302 38398
rect 34302 38363 34319 38398
rect 34447 38363 34451 38398
rect 34451 38363 34499 38398
rect 34627 38363 34658 38398
rect 34658 38363 34679 38398
rect 36678 38438 36697 38490
rect 36697 38438 36730 38490
rect 48943 38663 48984 38709
rect 48984 38663 48995 38709
rect 49154 38663 49190 38709
rect 49190 38663 49206 38709
rect 49365 38663 49396 38709
rect 49396 38663 49417 38709
rect 49576 38663 49602 38709
rect 49602 38663 49628 38709
rect 49787 38663 49839 38709
rect 39994 38540 40046 38592
rect 36961 38439 36971 38483
rect 36971 38439 37013 38483
rect 37172 38439 37206 38483
rect 37206 38439 37224 38483
rect 36961 38431 37013 38439
rect 37172 38431 37224 38439
rect 37384 38431 37436 38483
rect 37595 38431 37647 38483
rect 35332 38215 35384 38255
rect 35543 38215 35580 38255
rect 35580 38215 35595 38255
rect 35754 38215 35786 38255
rect 35786 38215 35806 38255
rect 35965 38215 35992 38255
rect 35992 38215 36017 38255
rect 36176 38215 36198 38255
rect 36198 38215 36228 38255
rect 37891 38215 37909 38243
rect 37909 38215 37943 38243
rect 38071 38215 38072 38243
rect 38072 38215 38123 38243
rect 35332 38203 35384 38215
rect 35543 38203 35595 38215
rect 35754 38203 35806 38215
rect 35965 38203 36017 38215
rect 36176 38203 36228 38215
rect 33819 38128 33833 38169
rect 33833 38128 33871 38169
rect 33999 38128 34039 38169
rect 34039 38128 34051 38169
rect 37891 38191 37943 38215
rect 38071 38191 38123 38215
rect 33819 38117 33871 38128
rect 33999 38117 34051 38128
rect 30854 37901 30906 37953
rect 31065 37901 31117 37953
rect 31276 37901 31328 37953
rect 31486 37950 31538 37953
rect 31697 37950 31749 37953
rect 31909 37950 31961 37953
rect 32120 37950 32172 37953
rect 32330 37950 32382 37953
rect 32541 37950 32593 37953
rect 32752 37950 32804 37953
rect 34284 37950 34336 37953
rect 34495 37950 34547 37953
rect 31486 37904 31538 37950
rect 31697 37904 31749 37950
rect 31909 37904 31961 37950
rect 32120 37904 32172 37950
rect 32330 37904 32382 37950
rect 32541 37904 32593 37950
rect 32752 37904 32804 37950
rect 34284 37904 34302 37950
rect 34302 37904 34336 37950
rect 34495 37904 34508 37950
rect 34508 37904 34547 37950
rect 31486 37901 31538 37904
rect 31697 37901 31749 37904
rect 31909 37901 31961 37904
rect 32120 37901 32172 37904
rect 32330 37901 32382 37904
rect 32541 37901 32593 37904
rect 32752 37901 32804 37904
rect 34284 37901 34336 37904
rect 34495 37901 34547 37904
rect 34707 37901 34759 37953
rect 34918 37901 34970 37953
rect 35220 37901 35272 37953
rect 35430 37901 35482 37953
rect 35641 37901 35693 37953
rect 35853 37901 35905 37953
rect 36064 37901 36116 37953
rect 36274 37901 36326 37953
rect 38330 37950 38382 37953
rect 38330 37904 38382 37950
rect 38330 37901 38382 37904
rect 38541 37901 38593 37953
rect 38752 37901 38804 37953
rect 39052 37950 39104 37953
rect 39232 37950 39284 37953
rect 39052 37904 39062 37950
rect 39062 37904 39104 37950
rect 39232 37904 39266 37950
rect 39266 37904 39284 37950
rect 39052 37901 39104 37904
rect 39232 37901 39284 37904
rect 33057 37726 33109 37729
rect 33237 37726 33289 37729
rect 33057 37680 33109 37726
rect 33237 37680 33289 37726
rect 33057 37677 33109 37680
rect 33237 37677 33289 37680
rect 33819 37726 33871 37737
rect 33999 37726 34051 37737
rect 33819 37685 33833 37726
rect 33833 37685 33871 37726
rect 33999 37685 34039 37726
rect 34039 37685 34051 37726
rect 35332 37639 35384 37651
rect 35543 37639 35595 37651
rect 35754 37639 35806 37651
rect 35965 37639 36017 37651
rect 36176 37639 36228 37651
rect 37891 37639 37943 37663
rect 38071 37639 38123 37663
rect 35332 37599 35384 37639
rect 35543 37599 35580 37639
rect 35580 37599 35595 37639
rect 35754 37599 35786 37639
rect 35786 37599 35806 37639
rect 35965 37599 35992 37639
rect 35992 37599 36017 37639
rect 36176 37599 36198 37639
rect 36198 37599 36228 37639
rect 37891 37611 37909 37639
rect 37909 37611 37943 37639
rect 38071 37611 38072 37639
rect 38072 37611 38123 37639
rect 34267 37456 34302 37491
rect 34302 37456 34319 37491
rect 34447 37456 34451 37491
rect 34451 37456 34499 37491
rect 34627 37456 34658 37491
rect 34658 37456 34679 37491
rect 34267 37439 34319 37456
rect 34447 37439 34499 37456
rect 34627 37439 34679 37456
rect 33057 37278 33109 37281
rect 33237 37278 33289 37281
rect 33057 37232 33109 37278
rect 33237 37232 33289 37278
rect 33057 37229 33109 37232
rect 33237 37229 33289 37232
rect 36678 37364 36697 37416
rect 36697 37364 36730 37416
rect 36961 37415 37013 37423
rect 37172 37415 37224 37423
rect 36961 37371 36971 37415
rect 36971 37371 37013 37415
rect 37172 37371 37206 37415
rect 37206 37371 37224 37415
rect 37384 37371 37436 37423
rect 37595 37371 37647 37423
rect 39994 38354 40046 38406
rect 39775 38174 39827 38191
rect 39775 38139 39786 38174
rect 39786 38139 39827 38174
rect 43445 38370 43497 38422
rect 41935 38139 41987 38191
rect 47486 38479 47538 38531
rect 48596 38525 48648 38577
rect 51835 38622 51887 38647
rect 52015 38622 52067 38647
rect 51835 38595 51887 38622
rect 52015 38595 52067 38622
rect 44939 38398 44991 38415
rect 45151 38398 45203 38415
rect 44939 38363 44971 38398
rect 44971 38363 44991 38398
rect 45151 38363 45197 38398
rect 45197 38363 45203 38398
rect 48596 38307 48648 38359
rect 50300 38363 50352 38415
rect 50511 38398 50563 38415
rect 50511 38363 50513 38398
rect 50513 38363 50563 38398
rect 50722 38363 50774 38415
rect 48943 38215 48984 38252
rect 48984 38215 48995 38252
rect 49154 38215 49190 38252
rect 49190 38215 49206 38252
rect 49365 38215 49396 38252
rect 49396 38215 49417 38252
rect 49576 38215 49602 38252
rect 49602 38215 49628 38252
rect 49787 38215 49839 38252
rect 48943 38200 48995 38215
rect 49154 38200 49206 38215
rect 49365 38200 49417 38215
rect 49576 38200 49628 38215
rect 49787 38200 49839 38215
rect 51073 38174 51125 38177
rect 51253 38174 51305 38177
rect 51073 38128 51086 38174
rect 51086 38128 51125 38174
rect 51253 38128 51292 38174
rect 51292 38128 51305 38174
rect 51073 38125 51125 38128
rect 51253 38125 51305 38128
rect 51835 38174 51887 38184
rect 52015 38174 52067 38184
rect 51835 38132 51887 38174
rect 52015 38132 52067 38174
rect 40253 37901 40305 37953
rect 40433 37901 40485 37953
rect 43790 37901 43842 37953
rect 44001 37901 44053 37953
rect 44213 37950 44265 37953
rect 44213 37904 44236 37950
rect 44236 37904 44265 37950
rect 44213 37901 44265 37904
rect 44424 37901 44476 37953
rect 44834 37950 44886 37953
rect 45045 37950 45097 37953
rect 45256 37950 45308 37953
rect 44834 37904 44858 37950
rect 44858 37904 44886 37950
rect 45045 37904 45084 37950
rect 45084 37904 45097 37950
rect 45256 37904 45264 37950
rect 45264 37904 45308 37950
rect 44834 37901 44886 37904
rect 45045 37901 45097 37904
rect 45256 37901 45308 37904
rect 48838 37901 48890 37953
rect 49048 37901 49100 37953
rect 49259 37901 49311 37953
rect 49471 37901 49523 37953
rect 49682 37901 49734 37953
rect 49892 37901 49944 37953
rect 50346 37901 50398 37953
rect 50557 37950 50609 37953
rect 50768 37950 50820 37953
rect 52316 37950 52368 37953
rect 52527 37950 52579 37953
rect 52738 37950 52790 37953
rect 52948 37950 53000 37953
rect 53159 37950 53211 37953
rect 53371 37950 53423 37953
rect 53582 37950 53634 37953
rect 50557 37904 50571 37950
rect 50571 37904 50609 37950
rect 50768 37904 50777 37950
rect 50777 37904 50820 37950
rect 52316 37904 52368 37950
rect 52527 37904 52579 37950
rect 52738 37904 52790 37950
rect 52948 37904 53000 37950
rect 53159 37904 53211 37950
rect 53371 37904 53423 37950
rect 53582 37904 53634 37950
rect 50557 37901 50609 37904
rect 50768 37901 50820 37904
rect 39775 37680 39786 37715
rect 39786 37680 39827 37715
rect 39775 37663 39827 37680
rect 39994 37448 40046 37500
rect 39994 37262 40046 37314
rect 52316 37901 52368 37904
rect 52527 37901 52579 37904
rect 52738 37901 52790 37904
rect 52948 37901 53000 37904
rect 53159 37901 53211 37904
rect 53371 37901 53423 37904
rect 53582 37901 53634 37904
rect 53792 37901 53844 37953
rect 54003 37901 54055 37953
rect 54214 37901 54266 37953
rect 54855 37901 54907 37953
rect 55066 37901 55118 37953
rect 55278 37950 55330 37953
rect 55278 37904 55279 37950
rect 55279 37904 55325 37950
rect 55325 37904 55330 37950
rect 55278 37901 55330 37904
rect 55489 37901 55541 37953
rect 41935 37663 41987 37715
rect 51073 37726 51125 37729
rect 51253 37726 51305 37729
rect 43445 37432 43497 37484
rect 51073 37680 51086 37726
rect 51086 37680 51125 37726
rect 51253 37680 51292 37726
rect 51292 37680 51305 37726
rect 48943 37639 48995 37654
rect 49154 37639 49206 37654
rect 49365 37639 49417 37654
rect 49576 37639 49628 37654
rect 49787 37639 49839 37654
rect 48943 37602 48984 37639
rect 48984 37602 48995 37639
rect 49154 37602 49190 37639
rect 49190 37602 49206 37639
rect 49365 37602 49396 37639
rect 49396 37602 49417 37639
rect 49576 37602 49602 37639
rect 49602 37602 49628 37639
rect 49787 37602 49839 37639
rect 51073 37677 51125 37680
rect 51253 37677 51305 37680
rect 44939 37456 44971 37491
rect 44971 37456 44991 37491
rect 45151 37456 45197 37491
rect 45197 37456 45203 37491
rect 48596 37495 48648 37547
rect 44939 37439 44991 37456
rect 45151 37439 45203 37456
rect 47864 37323 47916 37375
rect 50300 37439 50352 37491
rect 50511 37456 50513 37491
rect 50513 37456 50563 37491
rect 50511 37439 50563 37456
rect 50722 37439 50774 37491
rect 48596 37277 48648 37329
rect 51835 37680 51887 37722
rect 52015 37680 52067 37722
rect 51835 37670 51887 37680
rect 52015 37670 52067 37680
rect 35332 37145 35384 37191
rect 35543 37145 35580 37191
rect 35580 37145 35595 37191
rect 35754 37145 35786 37191
rect 35786 37145 35806 37191
rect 35965 37145 35992 37191
rect 35992 37145 36017 37191
rect 36176 37145 36198 37191
rect 36198 37145 36228 37191
rect 37891 37145 37909 37189
rect 37909 37145 37943 37189
rect 38071 37145 38072 37189
rect 38072 37145 38123 37189
rect 48943 37145 48984 37191
rect 48984 37145 48995 37191
rect 49154 37145 49190 37191
rect 49190 37145 49206 37191
rect 49365 37145 49396 37191
rect 49396 37145 49417 37191
rect 49576 37145 49602 37191
rect 49602 37145 49628 37191
rect 49787 37145 49839 37191
rect 51835 37232 51887 37259
rect 52015 37232 52067 37259
rect 51835 37207 51887 37232
rect 52015 37207 52067 37232
rect 35332 37139 35384 37145
rect 35543 37139 35595 37145
rect 35754 37139 35806 37145
rect 35965 37139 36017 37145
rect 36176 37139 36228 37145
rect 37891 37137 37943 37145
rect 38071 37137 38123 37145
rect 27790 37001 27842 37053
rect 28001 37001 28053 37053
rect 28212 37001 28264 37053
rect 28423 37001 28475 37053
rect 28634 37001 28686 37053
rect 28845 37050 28897 37053
rect 28845 37004 28856 37050
rect 28856 37004 28897 37050
rect 28845 37001 28897 37004
rect 29056 37001 29108 37053
rect 29582 37001 29634 37053
rect 29793 37050 29845 37053
rect 29793 37004 29798 37050
rect 29798 37004 29844 37050
rect 29844 37004 29845 37050
rect 29793 37001 29845 37004
rect 30005 37001 30057 37053
rect 30216 37001 30268 37053
rect 30854 37001 30906 37053
rect 31065 37001 31117 37053
rect 31276 37001 31328 37053
rect 31486 37001 31538 37053
rect 31697 37001 31749 37053
rect 31909 37001 31961 37053
rect 32120 37001 32172 37053
rect 32330 37001 32382 37053
rect 32541 37001 32593 37053
rect 32752 37001 32804 37053
rect 48943 37139 48995 37145
rect 49154 37139 49206 37145
rect 49365 37139 49417 37145
rect 49576 37139 49628 37145
rect 49787 37139 49839 37145
rect 34755 37001 34807 37053
rect 34935 37050 34987 37053
rect 34935 37004 34962 37050
rect 34962 37004 34987 37050
rect 34935 37001 34987 37004
rect 50138 37050 50190 37053
rect 50138 37004 50160 37050
rect 50160 37004 50190 37050
rect 50138 37001 50190 37004
rect 50318 37001 50370 37053
rect 35332 36909 35384 36915
rect 35543 36909 35595 36915
rect 35754 36909 35806 36915
rect 35965 36909 36017 36915
rect 36176 36909 36228 36915
rect 37891 36909 37943 36917
rect 38071 36909 38123 36917
rect 52316 37001 52368 37053
rect 52527 37001 52579 37053
rect 52738 37001 52790 37053
rect 52948 37001 53000 37053
rect 53159 37001 53211 37053
rect 53371 37001 53423 37053
rect 53582 37001 53634 37053
rect 53792 37001 53844 37053
rect 54003 37001 54055 37053
rect 54214 37001 54266 37053
rect 54855 37001 54907 37053
rect 55066 37001 55118 37053
rect 55278 37050 55330 37053
rect 55278 37004 55279 37050
rect 55279 37004 55325 37050
rect 55325 37004 55330 37050
rect 55278 37001 55330 37004
rect 55489 37001 55541 37053
rect 56015 37001 56067 37053
rect 56226 37050 56278 37053
rect 56226 37004 56267 37050
rect 56267 37004 56278 37050
rect 56226 37001 56278 37004
rect 56437 37001 56489 37053
rect 56648 37001 56700 37053
rect 56859 37001 56911 37053
rect 57070 37001 57122 37053
rect 57281 37001 57333 37053
rect 48943 36909 48995 36915
rect 49154 36909 49206 36915
rect 49365 36909 49417 36915
rect 49576 36909 49628 36915
rect 49787 36909 49839 36915
rect 33057 36822 33109 36825
rect 33237 36822 33289 36825
rect 35332 36863 35384 36909
rect 35543 36863 35580 36909
rect 35580 36863 35595 36909
rect 35754 36863 35786 36909
rect 35786 36863 35806 36909
rect 35965 36863 35992 36909
rect 35992 36863 36017 36909
rect 36176 36863 36198 36909
rect 36198 36863 36228 36909
rect 37891 36865 37909 36909
rect 37909 36865 37943 36909
rect 38071 36865 38072 36909
rect 38072 36865 38123 36909
rect 33057 36776 33109 36822
rect 33237 36776 33289 36822
rect 33057 36773 33109 36776
rect 33237 36773 33289 36776
rect 33057 36374 33109 36377
rect 33237 36374 33289 36377
rect 33057 36328 33109 36374
rect 33237 36328 33289 36374
rect 33057 36325 33109 36328
rect 33237 36325 33289 36328
rect 29582 36101 29634 36153
rect 29793 36150 29845 36153
rect 29793 36104 29798 36150
rect 29798 36104 29844 36150
rect 29844 36104 29845 36150
rect 29793 36101 29845 36104
rect 30005 36101 30057 36153
rect 30216 36101 30268 36153
rect 34267 36598 34319 36615
rect 34447 36598 34499 36615
rect 34627 36598 34679 36615
rect 34267 36563 34302 36598
rect 34302 36563 34319 36598
rect 34447 36563 34451 36598
rect 34451 36563 34499 36598
rect 34627 36563 34658 36598
rect 34658 36563 34679 36598
rect 36678 36638 36697 36690
rect 36697 36638 36730 36690
rect 48943 36863 48984 36909
rect 48984 36863 48995 36909
rect 49154 36863 49190 36909
rect 49190 36863 49206 36909
rect 49365 36863 49396 36909
rect 49396 36863 49417 36909
rect 49576 36863 49602 36909
rect 49602 36863 49628 36909
rect 49787 36863 49839 36909
rect 39994 36740 40046 36792
rect 36961 36639 36971 36683
rect 36971 36639 37013 36683
rect 37172 36639 37206 36683
rect 37206 36639 37224 36683
rect 36961 36631 37013 36639
rect 37172 36631 37224 36639
rect 37384 36631 37436 36683
rect 37595 36631 37647 36683
rect 35332 36415 35384 36455
rect 35543 36415 35580 36455
rect 35580 36415 35595 36455
rect 35754 36415 35786 36455
rect 35786 36415 35806 36455
rect 35965 36415 35992 36455
rect 35992 36415 36017 36455
rect 36176 36415 36198 36455
rect 36198 36415 36228 36455
rect 37891 36415 37909 36443
rect 37909 36415 37943 36443
rect 38071 36415 38072 36443
rect 38072 36415 38123 36443
rect 35332 36403 35384 36415
rect 35543 36403 35595 36415
rect 35754 36403 35806 36415
rect 35965 36403 36017 36415
rect 36176 36403 36228 36415
rect 33819 36328 33833 36369
rect 33833 36328 33871 36369
rect 33999 36328 34039 36369
rect 34039 36328 34051 36369
rect 37891 36391 37943 36415
rect 38071 36391 38123 36415
rect 33819 36317 33871 36328
rect 33999 36317 34051 36328
rect 30854 36101 30906 36153
rect 31065 36101 31117 36153
rect 31276 36101 31328 36153
rect 31486 36150 31538 36153
rect 31697 36150 31749 36153
rect 31909 36150 31961 36153
rect 32120 36150 32172 36153
rect 32330 36150 32382 36153
rect 32541 36150 32593 36153
rect 32752 36150 32804 36153
rect 34284 36150 34336 36153
rect 34495 36150 34547 36153
rect 31486 36104 31538 36150
rect 31697 36104 31749 36150
rect 31909 36104 31961 36150
rect 32120 36104 32172 36150
rect 32330 36104 32382 36150
rect 32541 36104 32593 36150
rect 32752 36104 32804 36150
rect 34284 36104 34302 36150
rect 34302 36104 34336 36150
rect 34495 36104 34508 36150
rect 34508 36104 34547 36150
rect 31486 36101 31538 36104
rect 31697 36101 31749 36104
rect 31909 36101 31961 36104
rect 32120 36101 32172 36104
rect 32330 36101 32382 36104
rect 32541 36101 32593 36104
rect 32752 36101 32804 36104
rect 34284 36101 34336 36104
rect 34495 36101 34547 36104
rect 34707 36101 34759 36153
rect 34918 36101 34970 36153
rect 35220 36101 35272 36153
rect 35430 36101 35482 36153
rect 35641 36101 35693 36153
rect 35853 36101 35905 36153
rect 36064 36101 36116 36153
rect 36274 36101 36326 36153
rect 38330 36150 38382 36153
rect 38330 36104 38382 36150
rect 38330 36101 38382 36104
rect 38541 36101 38593 36153
rect 38752 36101 38804 36153
rect 39052 36150 39104 36153
rect 39232 36150 39284 36153
rect 39052 36104 39062 36150
rect 39062 36104 39104 36150
rect 39232 36104 39266 36150
rect 39266 36104 39284 36150
rect 39052 36101 39104 36104
rect 39232 36101 39284 36104
rect 39994 36554 40046 36606
rect 39775 36374 39827 36391
rect 39775 36339 39786 36374
rect 39786 36339 39827 36374
rect 43445 36570 43497 36622
rect 41935 36339 41987 36391
rect 48241 36679 48293 36731
rect 48596 36725 48648 36777
rect 51835 36822 51887 36847
rect 52015 36822 52067 36847
rect 51835 36795 51887 36822
rect 52015 36795 52067 36822
rect 44939 36598 44991 36615
rect 45151 36598 45203 36615
rect 44939 36563 44971 36598
rect 44971 36563 44991 36598
rect 45151 36563 45197 36598
rect 45197 36563 45203 36598
rect 48596 36507 48648 36559
rect 50300 36563 50352 36615
rect 50511 36598 50563 36615
rect 50511 36563 50513 36598
rect 50513 36563 50563 36598
rect 50722 36563 50774 36615
rect 48943 36415 48984 36452
rect 48984 36415 48995 36452
rect 49154 36415 49190 36452
rect 49190 36415 49206 36452
rect 49365 36415 49396 36452
rect 49396 36415 49417 36452
rect 49576 36415 49602 36452
rect 49602 36415 49628 36452
rect 49787 36415 49839 36452
rect 48943 36400 48995 36415
rect 49154 36400 49206 36415
rect 49365 36400 49417 36415
rect 49576 36400 49628 36415
rect 49787 36400 49839 36415
rect 51073 36374 51125 36377
rect 51253 36374 51305 36377
rect 51073 36328 51086 36374
rect 51086 36328 51125 36374
rect 51253 36328 51292 36374
rect 51292 36328 51305 36374
rect 51073 36325 51125 36328
rect 51253 36325 51305 36328
rect 51835 36374 51887 36384
rect 52015 36374 52067 36384
rect 51835 36332 51887 36374
rect 52015 36332 52067 36374
rect 40253 36101 40305 36153
rect 40433 36101 40485 36153
rect 43790 36101 43842 36153
rect 44001 36101 44053 36153
rect 44213 36150 44265 36153
rect 44213 36104 44236 36150
rect 44236 36104 44265 36150
rect 44213 36101 44265 36104
rect 44424 36101 44476 36153
rect 44834 36150 44886 36153
rect 45045 36150 45097 36153
rect 45256 36150 45308 36153
rect 44834 36104 44858 36150
rect 44858 36104 44886 36150
rect 45045 36104 45084 36150
rect 45084 36104 45097 36150
rect 45256 36104 45264 36150
rect 45264 36104 45308 36150
rect 44834 36101 44886 36104
rect 45045 36101 45097 36104
rect 45256 36101 45308 36104
rect 48838 36101 48890 36153
rect 49048 36101 49100 36153
rect 49259 36101 49311 36153
rect 49471 36101 49523 36153
rect 49682 36101 49734 36153
rect 49892 36101 49944 36153
rect 50346 36101 50398 36153
rect 50557 36150 50609 36153
rect 50768 36150 50820 36153
rect 52316 36150 52368 36153
rect 52527 36150 52579 36153
rect 52738 36150 52790 36153
rect 52948 36150 53000 36153
rect 53159 36150 53211 36153
rect 53371 36150 53423 36153
rect 53582 36150 53634 36153
rect 50557 36104 50571 36150
rect 50571 36104 50609 36150
rect 50768 36104 50777 36150
rect 50777 36104 50820 36150
rect 52316 36104 52368 36150
rect 52527 36104 52579 36150
rect 52738 36104 52790 36150
rect 52948 36104 53000 36150
rect 53159 36104 53211 36150
rect 53371 36104 53423 36150
rect 53582 36104 53634 36150
rect 50557 36101 50609 36104
rect 50768 36101 50820 36104
rect 52316 36101 52368 36104
rect 52527 36101 52579 36104
rect 52738 36101 52790 36104
rect 52948 36101 53000 36104
rect 53159 36101 53211 36104
rect 53371 36101 53423 36104
rect 53582 36101 53634 36104
rect 53792 36101 53844 36153
rect 54003 36101 54055 36153
rect 54214 36101 54266 36153
rect 54855 36101 54907 36153
rect 55066 36101 55118 36153
rect 55278 36150 55330 36153
rect 55278 36104 55279 36150
rect 55279 36104 55325 36150
rect 55325 36104 55330 36150
rect 55278 36101 55330 36104
rect 55489 36101 55541 36153
rect 27449 34886 27498 34938
rect 27498 34886 27501 34938
rect 27573 34886 27625 34938
rect 27697 34886 27744 34938
rect 27744 34886 27749 34938
rect 25400 34796 25452 34848
rect 25524 34796 25576 34848
rect 25648 34796 25700 34848
rect 25772 34796 25824 34848
rect 25896 34796 25948 34848
rect 27449 34762 27498 34814
rect 27498 34762 27501 34814
rect 27573 34762 27625 34814
rect 27697 34762 27744 34814
rect 27744 34762 27749 34814
rect 25400 34672 25452 34724
rect 25524 34672 25576 34724
rect 25648 34672 25700 34724
rect 25772 34672 25824 34724
rect 25896 34672 25948 34724
rect 27449 34638 27498 34690
rect 27498 34638 27501 34690
rect 27573 34638 27625 34690
rect 27697 34638 27744 34690
rect 27744 34638 27749 34690
rect 27449 34514 27498 34566
rect 27498 34514 27501 34566
rect 27573 34514 27625 34566
rect 27697 34514 27744 34566
rect 27744 34514 27749 34566
rect 26861 33380 26913 33432
rect 27073 33380 27125 33432
rect 26861 33163 26913 33215
rect 27073 33163 27125 33215
rect 26861 32945 26913 32997
rect 27073 32945 27125 32997
rect 26861 32727 26913 32779
rect 27073 32727 27125 32779
rect 26861 32510 26913 32562
rect 27073 32510 27125 32562
rect 26861 32292 26913 32344
rect 27073 32292 27125 32344
rect 26861 32075 26913 32127
rect 27073 32075 27125 32127
rect 26861 31857 26913 31909
rect 27073 31857 27125 31909
rect 26861 31639 26913 31691
rect 27073 31639 27125 31691
rect 26861 31422 26913 31474
rect 27073 31422 27125 31474
rect 26861 31204 26913 31256
rect 27073 31204 27125 31256
rect 26861 30986 26913 31038
rect 27073 30986 27125 31038
rect 26861 30769 26913 30821
rect 27073 30769 27125 30821
rect 26861 30551 26913 30603
rect 27073 30551 27125 30603
rect 26861 30334 26913 30386
rect 27073 30334 27125 30386
rect 26861 30116 26913 30168
rect 27073 30116 27125 30168
rect 26861 29898 26913 29950
rect 27073 29898 27125 29950
rect 26861 29681 26913 29733
rect 27073 29681 27125 29733
rect 26861 29463 26913 29515
rect 27073 29463 27125 29515
rect 26861 29245 26913 29297
rect 27073 29245 27125 29297
rect 26861 29028 26913 29080
rect 27073 29028 27125 29080
rect 26861 28810 26913 28862
rect 27073 28810 27125 28862
rect 26861 28592 26913 28644
rect 27073 28592 27125 28644
rect 26861 28375 26913 28427
rect 27073 28375 27125 28427
rect 26861 28157 26913 28209
rect 27073 28157 27125 28209
rect 26861 27940 26913 27992
rect 27073 27940 27125 27992
rect 26861 27722 26913 27774
rect 27073 27722 27125 27774
rect 26861 27504 26913 27556
rect 27073 27504 27125 27556
rect 26861 27287 26913 27339
rect 27073 27287 27125 27339
rect 26861 27069 26913 27121
rect 27073 27069 27125 27121
rect 26861 26851 26913 26903
rect 27073 26851 27125 26903
rect 26861 26634 26913 26686
rect 27073 26634 27125 26686
rect 26861 26416 26913 26468
rect 27073 26416 27125 26468
rect 26861 26198 26913 26250
rect 27073 26198 27125 26250
rect 26861 25981 26913 26033
rect 27073 25981 27125 26033
rect 26861 25763 26913 25815
rect 27073 25763 27125 25815
rect 26861 25546 26913 25598
rect 27073 25546 27125 25598
rect 26861 25328 26913 25380
rect 27073 25328 27125 25380
rect 26861 25110 26913 25162
rect 27073 25110 27125 25162
rect 26861 24893 26913 24945
rect 27073 24893 27125 24945
rect 26861 24675 26913 24727
rect 27073 24675 27125 24727
rect 26861 24457 26913 24509
rect 27073 24457 27125 24509
rect 26861 24240 26913 24292
rect 27073 24240 27125 24292
rect 26861 24022 26913 24074
rect 27073 24022 27125 24074
rect 26861 23805 26913 23857
rect 27073 23805 27125 23857
rect 26861 23587 26913 23639
rect 27073 23587 27125 23639
rect 26861 23369 26913 23421
rect 27073 23369 27125 23421
rect 26861 23152 26913 23204
rect 27073 23152 27125 23204
rect 26861 22934 26913 22986
rect 27073 22934 27125 22986
rect 26861 22716 26913 22768
rect 27073 22716 27125 22768
rect 26861 22499 26913 22551
rect 27073 22499 27125 22551
rect 26861 22281 26913 22333
rect 27073 22281 27125 22333
rect 26861 22063 26913 22115
rect 27073 22063 27125 22115
rect 26861 21846 26913 21898
rect 27073 21846 27125 21898
rect 26861 21628 26913 21680
rect 27073 21628 27125 21680
rect 26861 21411 26913 21463
rect 27073 21411 27125 21463
rect 26861 21193 26913 21245
rect 27073 21193 27125 21245
rect 26861 20975 26913 21027
rect 27073 20975 27125 21027
rect 26861 20758 26913 20810
rect 27073 20758 27125 20810
rect 26861 20540 26913 20592
rect 27073 20540 27125 20592
rect 26861 20322 26913 20374
rect 27073 20322 27125 20374
rect 26861 20105 26913 20157
rect 27073 20105 27125 20157
rect 26861 19887 26913 19939
rect 27073 19887 27125 19939
rect 26861 19670 26913 19722
rect 27073 19670 27125 19722
rect 26861 19452 26913 19504
rect 27073 19452 27125 19504
rect 26861 19234 26913 19286
rect 27073 19234 27125 19286
rect 26861 19016 26913 19068
rect 27073 19016 27125 19068
rect 26861 18799 26913 18851
rect 27073 18799 27125 18851
rect 26861 18581 26913 18633
rect 27073 18581 27125 18633
rect 26861 18364 26913 18416
rect 27073 18364 27125 18416
rect 26861 18146 26913 18198
rect 27073 18146 27125 18198
rect 26861 17928 26913 17980
rect 27073 17928 27125 17980
rect 26861 17711 26913 17763
rect 27073 17711 27125 17763
rect 26861 17493 26913 17545
rect 27073 17493 27125 17545
rect 26861 17275 26913 17327
rect 27073 17275 27125 17327
rect 26861 17058 26913 17110
rect 27073 17058 27125 17110
rect 26861 16840 26913 16892
rect 27073 16840 27125 16892
rect 26861 16623 26913 16675
rect 27073 16623 27125 16675
rect 26861 16405 26913 16457
rect 27073 16405 27125 16457
rect 26861 16187 26913 16239
rect 27073 16187 27125 16239
rect 26861 15970 26913 16022
rect 27073 15970 27125 16022
rect 26861 15752 26913 15804
rect 27073 15752 27125 15804
rect 26861 15534 26913 15586
rect 27073 15534 27125 15586
rect 26861 15317 26913 15369
rect 27073 15317 27125 15369
rect 26861 15099 26913 15151
rect 27073 15099 27125 15151
rect 26861 14881 26913 14933
rect 27073 14881 27125 14933
rect 26861 14664 26913 14716
rect 27073 14664 27125 14716
rect 26861 14446 26913 14498
rect 27073 14446 27125 14498
rect 26861 14229 26913 14281
rect 27073 14229 27125 14281
rect 26861 14011 26913 14063
rect 27073 14011 27125 14063
rect 26861 13793 26913 13845
rect 27073 13793 27125 13845
rect 26861 13576 26913 13628
rect 27073 13576 27125 13628
rect 26861 13358 26913 13410
rect 27073 13358 27125 13410
rect 26861 13140 26913 13192
rect 27073 13140 27125 13192
rect 26861 12923 26913 12975
rect 27073 12923 27125 12975
rect 26861 12705 26913 12757
rect 27073 12705 27125 12757
rect 26861 12488 26913 12540
rect 27073 12488 27125 12540
rect 26861 12270 26913 12322
rect 27073 12270 27125 12322
rect 26861 12052 26913 12104
rect 27073 12052 27125 12104
rect 26861 11835 26913 11887
rect 27073 11835 27125 11887
rect 26861 11617 26913 11669
rect 27073 11617 27125 11669
rect 26861 11399 26913 11451
rect 27073 11399 27125 11451
rect 26861 11182 26913 11234
rect 27073 11182 27125 11234
rect 26861 10964 26913 11016
rect 27073 10964 27125 11016
rect 26861 10746 26913 10798
rect 27073 10746 27125 10798
rect 26861 10529 26913 10581
rect 27073 10529 27125 10581
rect 26861 10311 26913 10363
rect 27073 10311 27125 10363
rect 26861 10094 26913 10146
rect 27073 10094 27125 10146
rect 26861 9876 26913 9928
rect 27073 9876 27125 9928
rect 26861 9658 26913 9710
rect 27073 9658 27125 9710
rect 26861 9441 26913 9493
rect 27073 9441 27125 9493
rect 26861 9223 26913 9275
rect 27073 9223 27125 9275
rect 26861 9005 26913 9057
rect 27073 9005 27125 9057
rect 26861 8788 26913 8840
rect 27073 8788 27125 8840
rect 26861 8570 26913 8622
rect 27073 8570 27125 8622
rect 26861 8352 26913 8404
rect 27073 8352 27125 8404
rect 26861 8135 26913 8187
rect 27073 8135 27125 8187
rect 26861 7917 26913 7969
rect 27073 7917 27125 7969
rect 26861 7700 26913 7752
rect 27073 7700 27125 7752
rect 26861 7482 26913 7534
rect 27073 7482 27125 7534
rect 26861 7264 26913 7316
rect 27073 7264 27125 7316
rect 26861 7047 26913 7099
rect 27073 7047 27125 7099
rect 26861 6829 26913 6881
rect 27073 6829 27125 6881
rect 26861 6611 26913 6663
rect 27073 6611 27125 6663
rect 26861 6394 26913 6446
rect 27073 6394 27125 6446
rect 26861 6176 26913 6228
rect 27073 6176 27125 6228
rect 26861 5959 26913 6011
rect 27073 5959 27125 6011
rect 26861 5741 26913 5793
rect 27073 5741 27125 5793
rect 26861 5523 26913 5575
rect 27073 5523 27125 5575
rect 26861 5306 26913 5358
rect 27073 5306 27125 5358
rect 26861 4535 26913 4587
rect 27073 4535 27125 4587
rect 26861 4318 26913 4370
rect 27073 4318 27125 4370
rect 26861 4100 26913 4152
rect 27073 4100 27125 4152
rect 26861 3882 26913 3934
rect 27073 3882 27125 3934
rect 26861 3665 26913 3717
rect 27073 3665 27125 3717
rect 27476 33380 27498 33432
rect 27498 33380 27528 33432
rect 27688 33380 27740 33432
rect 27476 33163 27498 33215
rect 27498 33163 27528 33215
rect 27688 33163 27740 33215
rect 27476 32945 27498 32997
rect 27498 32945 27528 32997
rect 27688 32945 27740 32997
rect 27476 32727 27498 32779
rect 27498 32727 27528 32779
rect 27688 32727 27740 32779
rect 27476 32510 27498 32562
rect 27498 32510 27528 32562
rect 27688 32510 27740 32562
rect 27476 32292 27498 32344
rect 27498 32292 27528 32344
rect 27688 32292 27740 32344
rect 27476 32075 27498 32127
rect 27498 32075 27528 32127
rect 27688 32075 27740 32127
rect 27476 31857 27498 31909
rect 27498 31857 27528 31909
rect 27688 31857 27740 31909
rect 27476 31639 27498 31691
rect 27498 31639 27528 31691
rect 27688 31639 27740 31691
rect 27476 31422 27498 31474
rect 27498 31422 27528 31474
rect 27688 31422 27740 31474
rect 27476 31204 27498 31256
rect 27498 31204 27528 31256
rect 27688 31204 27740 31256
rect 27476 30986 27498 31038
rect 27498 30986 27528 31038
rect 27688 30986 27740 31038
rect 27476 30769 27498 30821
rect 27498 30769 27528 30821
rect 27688 30769 27740 30821
rect 27476 30551 27498 30603
rect 27498 30551 27528 30603
rect 27688 30551 27740 30603
rect 27476 30334 27498 30386
rect 27498 30334 27528 30386
rect 27688 30334 27740 30386
rect 27476 30116 27498 30168
rect 27498 30116 27528 30168
rect 27688 30116 27740 30168
rect 27476 29898 27498 29950
rect 27498 29898 27528 29950
rect 27688 29898 27740 29950
rect 27476 29681 27498 29733
rect 27498 29681 27528 29733
rect 27688 29681 27740 29733
rect 27476 29463 27498 29515
rect 27498 29463 27528 29515
rect 27688 29463 27740 29515
rect 27476 29245 27498 29297
rect 27498 29245 27528 29297
rect 27688 29245 27740 29297
rect 27476 29028 27498 29080
rect 27498 29028 27528 29080
rect 27688 29028 27740 29080
rect 27476 28810 27498 28862
rect 27498 28810 27528 28862
rect 27688 28810 27740 28862
rect 27476 28592 27498 28644
rect 27498 28592 27528 28644
rect 27688 28592 27740 28644
rect 27476 28375 27498 28427
rect 27498 28375 27528 28427
rect 27688 28375 27740 28427
rect 27476 28157 27498 28209
rect 27498 28157 27528 28209
rect 27688 28157 27740 28209
rect 27476 27940 27498 27992
rect 27498 27940 27528 27992
rect 27688 27940 27740 27992
rect 27476 27722 27498 27774
rect 27498 27722 27528 27774
rect 27688 27722 27740 27774
rect 27476 27504 27498 27556
rect 27498 27504 27528 27556
rect 27688 27504 27740 27556
rect 27476 27287 27498 27339
rect 27498 27287 27528 27339
rect 27688 27287 27740 27339
rect 27476 27069 27498 27121
rect 27498 27069 27528 27121
rect 27688 27069 27740 27121
rect 27476 26851 27498 26903
rect 27498 26851 27528 26903
rect 27688 26851 27740 26903
rect 27476 26634 27498 26686
rect 27498 26634 27528 26686
rect 27688 26634 27740 26686
rect 27476 26416 27498 26468
rect 27498 26416 27528 26468
rect 27688 26416 27740 26468
rect 27476 26198 27498 26250
rect 27498 26198 27528 26250
rect 27688 26198 27740 26250
rect 27476 25981 27498 26033
rect 27498 25981 27528 26033
rect 27688 25981 27740 26033
rect 27476 25763 27498 25815
rect 27498 25763 27528 25815
rect 27688 25763 27740 25815
rect 27476 25546 27498 25598
rect 27498 25546 27528 25598
rect 27688 25546 27740 25598
rect 27476 25328 27498 25380
rect 27498 25328 27528 25380
rect 27688 25328 27740 25380
rect 27476 25110 27498 25162
rect 27498 25110 27528 25162
rect 27688 25110 27740 25162
rect 27476 24893 27498 24945
rect 27498 24893 27528 24945
rect 27688 24893 27740 24945
rect 27476 24675 27498 24727
rect 27498 24675 27528 24727
rect 27688 24675 27740 24727
rect 27476 24457 27498 24509
rect 27498 24457 27528 24509
rect 27688 24457 27740 24509
rect 27476 24240 27498 24292
rect 27498 24240 27528 24292
rect 27688 24240 27740 24292
rect 27476 24022 27498 24074
rect 27498 24022 27528 24074
rect 27688 24022 27740 24074
rect 27476 23805 27498 23857
rect 27498 23805 27528 23857
rect 27688 23805 27740 23857
rect 27476 23587 27498 23639
rect 27498 23587 27528 23639
rect 27688 23587 27740 23639
rect 27476 23369 27498 23421
rect 27498 23369 27528 23421
rect 27688 23369 27740 23421
rect 27476 23152 27498 23204
rect 27498 23152 27528 23204
rect 27688 23152 27740 23204
rect 27476 22934 27498 22986
rect 27498 22934 27528 22986
rect 27688 22934 27740 22986
rect 27476 22716 27498 22768
rect 27498 22716 27528 22768
rect 27688 22716 27740 22768
rect 27476 22499 27498 22551
rect 27498 22499 27528 22551
rect 27688 22499 27740 22551
rect 27476 22281 27498 22333
rect 27498 22281 27528 22333
rect 27688 22281 27740 22333
rect 27476 22063 27498 22115
rect 27498 22063 27528 22115
rect 27688 22063 27740 22115
rect 27476 21846 27498 21898
rect 27498 21846 27528 21898
rect 27688 21846 27740 21898
rect 27476 21628 27498 21680
rect 27498 21628 27528 21680
rect 27688 21628 27740 21680
rect 27476 21411 27498 21463
rect 27498 21411 27528 21463
rect 27688 21411 27740 21463
rect 27476 21193 27498 21245
rect 27498 21193 27528 21245
rect 27688 21193 27740 21245
rect 27476 20975 27498 21027
rect 27498 20975 27528 21027
rect 27688 20975 27740 21027
rect 27476 20758 27498 20810
rect 27498 20758 27528 20810
rect 27688 20758 27740 20810
rect 27476 20540 27498 20592
rect 27498 20540 27528 20592
rect 27688 20540 27740 20592
rect 27476 20322 27498 20374
rect 27498 20322 27528 20374
rect 27688 20322 27740 20374
rect 27476 20105 27498 20157
rect 27498 20105 27528 20157
rect 27688 20105 27740 20157
rect 27476 19887 27498 19939
rect 27498 19887 27528 19939
rect 27688 19887 27740 19939
rect 27476 19670 27498 19722
rect 27498 19670 27528 19722
rect 27688 19670 27740 19722
rect 27476 19452 27498 19504
rect 27498 19452 27528 19504
rect 27688 19452 27740 19504
rect 27476 19234 27498 19286
rect 27498 19234 27528 19286
rect 27688 19234 27740 19286
rect 27476 19016 27498 19068
rect 27498 19016 27528 19068
rect 27688 19016 27740 19068
rect 27476 18799 27498 18851
rect 27498 18799 27528 18851
rect 27688 18799 27740 18851
rect 27476 18581 27498 18633
rect 27498 18581 27528 18633
rect 27688 18581 27740 18633
rect 27476 18364 27498 18416
rect 27498 18364 27528 18416
rect 27688 18364 27740 18416
rect 27476 18146 27498 18198
rect 27498 18146 27528 18198
rect 27688 18146 27740 18198
rect 27476 17928 27498 17980
rect 27498 17928 27528 17980
rect 27688 17928 27740 17980
rect 27476 17711 27498 17763
rect 27498 17711 27528 17763
rect 27688 17711 27740 17763
rect 27476 17493 27498 17545
rect 27498 17493 27528 17545
rect 27688 17493 27740 17545
rect 27476 17275 27498 17327
rect 27498 17275 27528 17327
rect 27688 17275 27740 17327
rect 27476 17058 27498 17110
rect 27498 17058 27528 17110
rect 27688 17058 27740 17110
rect 27476 16840 27498 16892
rect 27498 16840 27528 16892
rect 27688 16840 27740 16892
rect 27476 16623 27498 16675
rect 27498 16623 27528 16675
rect 27688 16623 27740 16675
rect 27476 16405 27498 16457
rect 27498 16405 27528 16457
rect 27688 16405 27740 16457
rect 27476 16187 27498 16239
rect 27498 16187 27528 16239
rect 27688 16187 27740 16239
rect 27476 15970 27498 16022
rect 27498 15970 27528 16022
rect 27688 15970 27740 16022
rect 27476 15752 27498 15804
rect 27498 15752 27528 15804
rect 27688 15752 27740 15804
rect 27476 15534 27498 15586
rect 27498 15534 27528 15586
rect 27688 15534 27740 15586
rect 27476 15317 27498 15369
rect 27498 15317 27528 15369
rect 27688 15317 27740 15369
rect 27476 15099 27498 15151
rect 27498 15099 27528 15151
rect 27688 15099 27740 15151
rect 27476 14881 27498 14933
rect 27498 14881 27528 14933
rect 27688 14881 27740 14933
rect 27476 14664 27498 14716
rect 27498 14664 27528 14716
rect 27688 14664 27740 14716
rect 27476 14446 27498 14498
rect 27498 14446 27528 14498
rect 27688 14446 27740 14498
rect 27476 14229 27498 14281
rect 27498 14229 27528 14281
rect 27688 14229 27740 14281
rect 27476 14011 27498 14063
rect 27498 14011 27528 14063
rect 27688 14011 27740 14063
rect 27476 13793 27498 13845
rect 27498 13793 27528 13845
rect 27688 13793 27740 13845
rect 27476 13576 27498 13628
rect 27498 13576 27528 13628
rect 27688 13576 27740 13628
rect 27476 13358 27498 13410
rect 27498 13358 27528 13410
rect 27688 13358 27740 13410
rect 27476 13140 27498 13192
rect 27498 13140 27528 13192
rect 27688 13140 27740 13192
rect 27476 12923 27498 12975
rect 27498 12923 27528 12975
rect 27688 12923 27740 12975
rect 27476 12705 27498 12757
rect 27498 12705 27528 12757
rect 27688 12705 27740 12757
rect 27476 12488 27498 12540
rect 27498 12488 27528 12540
rect 27688 12488 27740 12540
rect 27476 12270 27498 12322
rect 27498 12270 27528 12322
rect 27688 12270 27740 12322
rect 27476 12052 27498 12104
rect 27498 12052 27528 12104
rect 27688 12052 27740 12104
rect 27476 11835 27498 11887
rect 27498 11835 27528 11887
rect 27688 11835 27740 11887
rect 27476 11617 27498 11669
rect 27498 11617 27528 11669
rect 27688 11617 27740 11669
rect 27476 11399 27498 11451
rect 27498 11399 27528 11451
rect 27688 11399 27740 11451
rect 27476 11182 27498 11234
rect 27498 11182 27528 11234
rect 27688 11182 27740 11234
rect 27476 10964 27498 11016
rect 27498 10964 27528 11016
rect 27688 10964 27740 11016
rect 27476 10746 27498 10798
rect 27498 10746 27528 10798
rect 27688 10746 27740 10798
rect 27476 10529 27498 10581
rect 27498 10529 27528 10581
rect 27688 10529 27740 10581
rect 27476 10311 27498 10363
rect 27498 10311 27528 10363
rect 27688 10311 27740 10363
rect 27476 10094 27498 10146
rect 27498 10094 27528 10146
rect 27688 10094 27740 10146
rect 27476 9876 27498 9928
rect 27498 9876 27528 9928
rect 27688 9876 27740 9928
rect 27476 9658 27498 9710
rect 27498 9658 27528 9710
rect 27688 9658 27740 9710
rect 27476 9441 27498 9493
rect 27498 9441 27528 9493
rect 27688 9441 27740 9493
rect 27476 9223 27498 9275
rect 27498 9223 27528 9275
rect 27688 9223 27740 9275
rect 27476 9005 27498 9057
rect 27498 9005 27528 9057
rect 27688 9005 27740 9057
rect 27476 8788 27498 8840
rect 27498 8788 27528 8840
rect 27688 8788 27740 8840
rect 27476 8570 27498 8622
rect 27498 8570 27528 8622
rect 27688 8570 27740 8622
rect 27476 8352 27498 8404
rect 27498 8352 27528 8404
rect 27688 8352 27740 8404
rect 27476 8135 27498 8187
rect 27498 8135 27528 8187
rect 27688 8135 27740 8187
rect 27476 7917 27498 7969
rect 27498 7917 27528 7969
rect 27688 7917 27740 7969
rect 27476 7700 27498 7752
rect 27498 7700 27528 7752
rect 27688 7700 27740 7752
rect 27476 7482 27498 7534
rect 27498 7482 27528 7534
rect 27688 7482 27740 7534
rect 27476 7264 27498 7316
rect 27498 7264 27528 7316
rect 27688 7264 27740 7316
rect 27476 7047 27498 7099
rect 27498 7047 27528 7099
rect 27688 7047 27740 7099
rect 27476 6829 27498 6881
rect 27498 6829 27528 6881
rect 27688 6829 27740 6881
rect 27476 6611 27498 6663
rect 27498 6611 27528 6663
rect 27688 6611 27740 6663
rect 27476 6394 27498 6446
rect 27498 6394 27528 6446
rect 27688 6394 27740 6446
rect 27476 6176 27498 6228
rect 27498 6176 27528 6228
rect 27688 6176 27740 6228
rect 27476 5959 27498 6011
rect 27498 5959 27528 6011
rect 27688 5959 27740 6011
rect 27476 5741 27498 5793
rect 27498 5741 27528 5793
rect 27688 5741 27740 5793
rect 27476 5523 27498 5575
rect 27498 5523 27528 5575
rect 27688 5523 27740 5575
rect 27476 5306 27498 5358
rect 27498 5306 27528 5358
rect 27688 5306 27740 5358
rect 27476 4535 27498 4587
rect 27498 4535 27528 4587
rect 27688 4535 27740 4587
rect 27476 4318 27498 4370
rect 27498 4318 27528 4370
rect 27688 4318 27740 4370
rect 27476 4100 27498 4152
rect 27498 4100 27528 4152
rect 27688 4100 27740 4152
rect 27476 3882 27498 3934
rect 27498 3882 27528 3934
rect 27688 3882 27740 3934
rect 27476 3665 27498 3717
rect 27498 3665 27528 3717
rect 27688 3665 27740 3717
rect 2574 1637 2730 1689
rect 12639 1637 12795 1689
rect 13089 1637 13245 1689
rect 23439 1637 23595 1689
rect 49908 6297 50064 6349
rect 51654 5147 51810 5199
rect 40623 3230 40779 3282
rect 58814 44286 58866 44338
rect 58938 44286 58990 44338
rect 59062 44286 59114 44338
rect 59186 44286 59238 44338
rect 59310 44286 59362 44338
rect 59434 44286 59486 44338
rect 58814 44162 58866 44214
rect 58938 44162 58990 44214
rect 59062 44162 59114 44214
rect 59186 44162 59238 44214
rect 59310 44162 59362 44214
rect 59434 44162 59486 44214
rect 60575 35338 60627 35494
rect 57998 33380 58050 33432
rect 58210 33380 58262 33432
rect 57998 33163 58050 33215
rect 58210 33163 58262 33215
rect 57998 32945 58050 32997
rect 58210 32945 58262 32997
rect 57998 32727 58050 32779
rect 58210 32727 58262 32779
rect 57998 32510 58050 32562
rect 58210 32510 58262 32562
rect 57998 32292 58050 32344
rect 58210 32292 58262 32344
rect 57998 32075 58050 32127
rect 58210 32075 58262 32127
rect 57998 31857 58050 31909
rect 58210 31857 58262 31909
rect 57998 31639 58050 31691
rect 58210 31639 58262 31691
rect 57998 31422 58050 31474
rect 58210 31422 58262 31474
rect 57998 31204 58050 31256
rect 58210 31204 58262 31256
rect 57998 30986 58050 31038
rect 58210 30986 58262 31038
rect 57998 30769 58050 30821
rect 58210 30769 58262 30821
rect 57998 30551 58050 30603
rect 58210 30551 58262 30603
rect 57998 30334 58050 30386
rect 58210 30334 58262 30386
rect 57998 30116 58050 30168
rect 58210 30116 58262 30168
rect 57998 29898 58050 29950
rect 58210 29898 58262 29950
rect 57998 29681 58050 29733
rect 58210 29681 58262 29733
rect 57998 29463 58050 29515
rect 58210 29463 58262 29515
rect 57998 29245 58050 29297
rect 58210 29245 58262 29297
rect 57998 29028 58050 29080
rect 58210 29028 58262 29080
rect 57998 28810 58050 28862
rect 58210 28810 58262 28862
rect 57998 28592 58050 28644
rect 58210 28592 58262 28644
rect 57998 28375 58050 28427
rect 58210 28375 58262 28427
rect 57998 28157 58050 28209
rect 58210 28157 58262 28209
rect 57998 27940 58050 27992
rect 58210 27940 58262 27992
rect 57998 27722 58050 27774
rect 58210 27722 58262 27774
rect 57998 27504 58050 27556
rect 58210 27504 58262 27556
rect 57998 27287 58050 27339
rect 58210 27287 58262 27339
rect 57998 27069 58050 27121
rect 58210 27069 58262 27121
rect 57998 26851 58050 26903
rect 58210 26851 58262 26903
rect 57998 26634 58050 26686
rect 58210 26634 58262 26686
rect 57998 26416 58050 26468
rect 58210 26416 58262 26468
rect 57998 26198 58050 26250
rect 58210 26198 58262 26250
rect 57998 25981 58050 26033
rect 58210 25981 58262 26033
rect 57998 25763 58050 25815
rect 58210 25763 58262 25815
rect 57998 25546 58050 25598
rect 58210 25546 58262 25598
rect 57998 25328 58050 25380
rect 58210 25328 58262 25380
rect 57998 25110 58050 25162
rect 58210 25110 58262 25162
rect 57998 24893 58050 24945
rect 58210 24893 58262 24945
rect 57998 24675 58050 24727
rect 58210 24675 58262 24727
rect 57998 24457 58050 24509
rect 58210 24457 58262 24509
rect 57998 24240 58050 24292
rect 58210 24240 58262 24292
rect 57998 24022 58050 24074
rect 58210 24022 58262 24074
rect 57998 23805 58050 23857
rect 58210 23805 58262 23857
rect 57998 23587 58050 23639
rect 58210 23587 58262 23639
rect 57998 23369 58050 23421
rect 58210 23369 58262 23421
rect 57998 23152 58050 23204
rect 58210 23152 58262 23204
rect 57998 22934 58050 22986
rect 58210 22934 58262 22986
rect 57998 22716 58050 22768
rect 58210 22716 58262 22768
rect 57998 22499 58050 22551
rect 58210 22499 58262 22551
rect 57998 22281 58050 22333
rect 58210 22281 58262 22333
rect 57998 22063 58050 22115
rect 58210 22063 58262 22115
rect 57998 21846 58050 21898
rect 58210 21846 58262 21898
rect 57998 21628 58050 21680
rect 58210 21628 58262 21680
rect 57998 21411 58050 21463
rect 58210 21411 58262 21463
rect 57998 21193 58050 21245
rect 58210 21193 58262 21245
rect 57998 20975 58050 21027
rect 58210 20975 58262 21027
rect 57998 20758 58050 20810
rect 58210 20758 58262 20810
rect 57998 20540 58050 20592
rect 58210 20540 58262 20592
rect 57998 20322 58050 20374
rect 58210 20322 58262 20374
rect 57998 20105 58050 20157
rect 58210 20105 58262 20157
rect 57998 19887 58050 19939
rect 58210 19887 58262 19939
rect 57998 19670 58050 19722
rect 58210 19670 58262 19722
rect 57998 19452 58050 19504
rect 58210 19452 58262 19504
rect 57998 19234 58050 19286
rect 58210 19234 58262 19286
rect 57998 19016 58050 19068
rect 58210 19016 58262 19068
rect 57998 18799 58050 18851
rect 58210 18799 58262 18851
rect 57998 18581 58050 18633
rect 58210 18581 58262 18633
rect 57998 18364 58050 18416
rect 58210 18364 58262 18416
rect 57998 18146 58050 18198
rect 58210 18146 58262 18198
rect 57998 17928 58050 17980
rect 58210 17928 58262 17980
rect 57998 17711 58050 17763
rect 58210 17711 58262 17763
rect 57998 17493 58050 17545
rect 58210 17493 58262 17545
rect 57998 17275 58050 17327
rect 58210 17275 58262 17327
rect 57998 17058 58050 17110
rect 58210 17058 58262 17110
rect 57998 16840 58050 16892
rect 58210 16840 58262 16892
rect 57998 16623 58050 16675
rect 58210 16623 58262 16675
rect 57998 16405 58050 16457
rect 58210 16405 58262 16457
rect 57998 16187 58050 16239
rect 58210 16187 58262 16239
rect 57998 15970 58050 16022
rect 58210 15970 58262 16022
rect 57998 15752 58050 15804
rect 58210 15752 58262 15804
rect 57998 15534 58050 15586
rect 58210 15534 58262 15586
rect 57998 15317 58050 15369
rect 58210 15317 58262 15369
rect 57998 15099 58050 15151
rect 58210 15099 58262 15151
rect 57998 14881 58050 14933
rect 58210 14881 58262 14933
rect 57998 14664 58050 14716
rect 58210 14664 58262 14716
rect 57998 14446 58050 14498
rect 58210 14446 58262 14498
rect 57998 14229 58050 14281
rect 58210 14229 58262 14281
rect 57998 14011 58050 14063
rect 58210 14011 58262 14063
rect 57998 13793 58050 13845
rect 58210 13793 58262 13845
rect 57998 13576 58050 13628
rect 58210 13576 58262 13628
rect 57998 13358 58050 13410
rect 58210 13358 58262 13410
rect 57998 13140 58050 13192
rect 58210 13140 58262 13192
rect 57998 12923 58050 12975
rect 58210 12923 58262 12975
rect 57998 12705 58050 12757
rect 58210 12705 58262 12757
rect 57998 12488 58050 12540
rect 58210 12488 58262 12540
rect 57998 12270 58050 12322
rect 58210 12270 58262 12322
rect 57998 12052 58050 12104
rect 58210 12052 58262 12104
rect 57998 11835 58050 11887
rect 58210 11835 58262 11887
rect 57998 11617 58050 11669
rect 58210 11617 58262 11669
rect 57998 11399 58050 11451
rect 58210 11399 58262 11451
rect 57998 11182 58050 11234
rect 58210 11182 58262 11234
rect 57998 10964 58050 11016
rect 58210 10964 58262 11016
rect 57998 10746 58050 10798
rect 58210 10746 58262 10798
rect 57998 10529 58050 10581
rect 58210 10529 58262 10581
rect 57998 10311 58050 10363
rect 58210 10311 58262 10363
rect 57998 10094 58050 10146
rect 58210 10094 58262 10146
rect 57998 9876 58050 9928
rect 58210 9876 58262 9928
rect 57998 9658 58050 9710
rect 58210 9658 58262 9710
rect 57998 9441 58050 9493
rect 58210 9441 58262 9493
rect 57998 9223 58050 9275
rect 58210 9223 58262 9275
rect 57998 9005 58050 9057
rect 58210 9005 58262 9057
rect 57998 8788 58050 8840
rect 58210 8788 58262 8840
rect 57998 8570 58050 8622
rect 58210 8570 58262 8622
rect 57998 8352 58050 8404
rect 58210 8352 58262 8404
rect 57998 8135 58050 8187
rect 58210 8135 58262 8187
rect 57998 7917 58050 7969
rect 58210 7917 58262 7969
rect 57998 7700 58050 7752
rect 58210 7700 58262 7752
rect 57998 7482 58050 7534
rect 58210 7482 58262 7534
rect 57998 7264 58050 7316
rect 58210 7264 58262 7316
rect 57998 7047 58050 7099
rect 58210 7047 58262 7099
rect 57998 6829 58050 6881
rect 58210 6829 58262 6881
rect 57998 6611 58050 6663
rect 58210 6611 58262 6663
rect 57998 6394 58050 6446
rect 58210 6394 58262 6446
rect 57998 6176 58050 6228
rect 58210 6176 58262 6228
rect 57998 5959 58050 6011
rect 58210 5959 58262 6011
rect 57998 5741 58050 5793
rect 58210 5741 58262 5793
rect 57998 5523 58050 5575
rect 58210 5523 58262 5575
rect 57998 5306 58050 5358
rect 58210 5306 58262 5358
rect 57383 4535 57435 4587
rect 57595 4535 57626 4587
rect 57626 4535 57647 4587
rect 57383 4318 57435 4370
rect 57595 4318 57626 4370
rect 57626 4318 57647 4370
rect 57383 4100 57435 4152
rect 57595 4100 57626 4152
rect 57626 4100 57647 4152
rect 57383 3882 57435 3934
rect 57595 3882 57626 3934
rect 57626 3882 57647 3934
rect 57383 3665 57435 3717
rect 57595 3665 57626 3717
rect 57626 3665 57647 3717
rect 57998 4535 58050 4587
rect 58210 4535 58262 4587
rect 57998 4318 58050 4370
rect 58210 4318 58262 4370
rect 57998 4100 58050 4152
rect 58210 4100 58262 4152
rect 57998 3882 58050 3934
rect 58210 3882 58262 3934
rect 57998 3665 58050 3717
rect 58210 3665 58262 3717
rect 62150 1637 62306 1689
rect 72215 1637 72371 1689
rect 72665 1637 72821 1689
rect 82730 1637 82886 1689
rect 48668 971 48720 1023
rect 48792 971 48844 1023
rect 48916 971 48968 1023
rect 53907 969 53939 1006
rect 53939 969 53959 1006
rect 29090 891 29142 914
rect 29787 891 29839 914
rect 29090 845 29139 891
rect 29139 845 29142 891
rect 29787 845 29805 891
rect 29805 845 29839 891
rect 48668 847 48720 899
rect 48792 847 48844 899
rect 48916 847 48968 899
rect 53907 891 53959 969
rect 53907 845 53939 891
rect 53939 845 53959 891
rect 29090 767 29142 845
rect 29787 767 29839 845
rect 29090 721 29139 767
rect 29139 721 29142 767
rect 29787 721 29805 767
rect 29805 721 29839 767
rect 48668 723 48720 775
rect 48792 723 48844 775
rect 48916 723 48968 775
rect 53907 767 53959 845
rect 53907 721 53939 767
rect 53939 721 53959 767
rect 29090 654 29142 721
rect 29787 654 29839 721
rect 48668 599 48720 651
rect 48792 599 48844 651
rect 48916 599 48968 651
rect 53907 643 53959 721
rect 53907 642 53939 643
rect 53939 642 53959 643
<< metal2 >>
rect 282 45968 86090 46294
rect 706 44776 85666 45776
rect 706 403 1706 44776
rect 25313 44338 26039 44375
rect 25313 44314 25337 44338
rect 25389 44314 25461 44338
rect 25513 44314 25585 44338
rect 25637 44314 25709 44338
rect 25761 44314 25833 44338
rect 25885 44314 25957 44338
rect 26009 44314 26039 44338
rect 25313 44258 25335 44314
rect 25391 44258 25459 44314
rect 25515 44258 25583 44314
rect 25639 44258 25707 44314
rect 25763 44258 25831 44314
rect 25887 44258 25955 44314
rect 26011 44258 26039 44314
rect 25313 44214 26039 44258
rect 25313 44190 25337 44214
rect 25389 44190 25461 44214
rect 25513 44190 25585 44214
rect 25637 44190 25709 44214
rect 25761 44190 25833 44214
rect 25885 44190 25957 44214
rect 26009 44190 26039 44214
rect 25313 44134 25335 44190
rect 25391 44134 25459 44190
rect 25515 44134 25583 44190
rect 25639 44134 25707 44190
rect 25763 44134 25831 44190
rect 25887 44134 25955 44190
rect 26011 44134 26039 44190
rect 25313 34972 26039 44134
rect 25313 34920 25400 34972
rect 25452 34920 25524 34972
rect 25576 34920 25648 34972
rect 25700 34920 25772 34972
rect 25824 34920 25896 34972
rect 25948 34920 26039 34972
rect 25313 34877 26039 34920
rect 25313 34821 25398 34877
rect 25454 34821 25522 34877
rect 25578 34821 25646 34877
rect 25702 34821 25770 34877
rect 25826 34821 25894 34877
rect 25950 34821 26039 34877
rect 25313 34796 25400 34821
rect 25452 34796 25524 34821
rect 25576 34796 25648 34821
rect 25700 34796 25772 34821
rect 25824 34796 25896 34821
rect 25948 34796 26039 34821
rect 25313 34753 26039 34796
rect 25313 34697 25398 34753
rect 25454 34697 25522 34753
rect 25578 34697 25646 34753
rect 25702 34697 25770 34753
rect 25826 34697 25894 34753
rect 25950 34697 26039 34753
rect 25313 34672 25400 34697
rect 25452 34672 25524 34697
rect 25576 34672 25648 34697
rect 25700 34672 25772 34697
rect 25824 34672 25896 34697
rect 25948 34672 26039 34697
rect 25313 34629 26039 34672
rect 25313 34573 25398 34629
rect 25454 34573 25522 34629
rect 25578 34573 25646 34629
rect 25702 34573 25770 34629
rect 25826 34573 25894 34629
rect 25950 34573 26039 34629
rect 25313 31248 26039 34573
rect 25313 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31192 26039 31248
rect 25313 31124 26039 31192
rect 25313 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 26039 31124
rect 25313 31000 26039 31068
rect 25313 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30944 26039 31000
rect 25313 30793 26039 30944
rect 25313 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30737 26039 30793
rect 25313 30669 26039 30737
rect 25313 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 26039 30669
rect 25313 30545 26039 30613
rect 25313 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30489 26039 30545
rect 25313 28282 26039 30489
rect 25313 28226 25404 28282
rect 25460 28226 25528 28282
rect 25584 28226 25652 28282
rect 25708 28226 25776 28282
rect 25832 28226 25900 28282
rect 25956 28226 26039 28282
rect 25313 28158 26039 28226
rect 25313 28102 25404 28158
rect 25460 28102 25528 28158
rect 25584 28102 25652 28158
rect 25708 28102 25776 28158
rect 25832 28102 25900 28158
rect 25956 28102 26039 28158
rect 25313 28034 26039 28102
rect 25313 27978 25404 28034
rect 25460 27978 25528 28034
rect 25584 27978 25652 28034
rect 25708 27978 25776 28034
rect 25832 27978 25900 28034
rect 25956 27978 26039 28034
rect 25313 27910 26039 27978
rect 25313 27854 25404 27910
rect 25460 27854 25528 27910
rect 25584 27854 25652 27910
rect 25708 27854 25776 27910
rect 25832 27854 25900 27910
rect 25956 27854 26039 27910
rect 25313 27786 26039 27854
rect 25313 27730 25404 27786
rect 25460 27730 25528 27786
rect 25584 27730 25652 27786
rect 25708 27730 25776 27786
rect 25832 27730 25900 27786
rect 25956 27730 26039 27786
rect 25313 27662 26039 27730
rect 25313 27606 25404 27662
rect 25460 27606 25528 27662
rect 25584 27606 25652 27662
rect 25708 27606 25776 27662
rect 25832 27606 25900 27662
rect 25956 27606 26039 27662
rect 25313 27538 26039 27606
rect 25313 27482 25404 27538
rect 25460 27482 25528 27538
rect 25584 27482 25652 27538
rect 25708 27482 25776 27538
rect 25832 27482 25900 27538
rect 25956 27482 26039 27538
rect 25313 27414 26039 27482
rect 25313 27358 25404 27414
rect 25460 27358 25528 27414
rect 25584 27358 25652 27414
rect 25708 27358 25776 27414
rect 25832 27358 25900 27414
rect 25956 27358 26039 27414
rect 25313 27290 26039 27358
rect 25313 27234 25404 27290
rect 25460 27234 25528 27290
rect 25584 27234 25652 27290
rect 25708 27234 25776 27290
rect 25832 27234 25900 27290
rect 25956 27234 26039 27290
rect 25313 27166 26039 27234
rect 25313 27110 25404 27166
rect 25460 27110 25528 27166
rect 25584 27110 25652 27166
rect 25708 27110 25776 27166
rect 25832 27110 25900 27166
rect 25956 27110 26039 27166
rect 25313 27042 26039 27110
rect 25313 26986 25404 27042
rect 25460 26986 25528 27042
rect 25584 26986 25652 27042
rect 25708 26986 25776 27042
rect 25832 26986 25900 27042
rect 25956 26986 26039 27042
rect 25313 26918 26039 26986
rect 25313 26862 25404 26918
rect 25460 26862 25528 26918
rect 25584 26862 25652 26918
rect 25708 26862 25776 26918
rect 25832 26862 25900 26918
rect 25956 26862 26039 26918
rect 25313 26794 26039 26862
rect 25313 26738 25404 26794
rect 25460 26738 25528 26794
rect 25584 26738 25652 26794
rect 25708 26738 25776 26794
rect 25832 26738 25900 26794
rect 25956 26738 26039 26794
rect 25313 26670 26039 26738
rect 25313 26614 25404 26670
rect 25460 26614 25528 26670
rect 25584 26614 25652 26670
rect 25708 26614 25776 26670
rect 25832 26614 25900 26670
rect 25956 26614 26039 26670
rect 25313 26546 26039 26614
rect 25313 26490 25404 26546
rect 25460 26490 25528 26546
rect 25584 26490 25652 26546
rect 25708 26490 25776 26546
rect 25832 26490 25900 26546
rect 25956 26490 26039 26546
rect 25313 26433 26039 26490
rect 26823 43417 27163 44776
rect 29486 44328 30364 44776
rect 26823 43361 26838 43417
rect 26894 43361 26962 43417
rect 27018 43361 27086 43417
rect 27142 43361 27163 43417
rect 26823 43293 27163 43361
rect 26823 43237 26838 43293
rect 26894 43237 26962 43293
rect 27018 43237 27086 43293
rect 27142 43237 27163 43293
rect 26823 36218 27163 43237
rect 26823 36162 26838 36218
rect 26894 36162 26962 36218
rect 27018 36162 27086 36218
rect 27142 36162 27163 36218
rect 26823 36094 27163 36162
rect 26823 36038 26838 36094
rect 26894 36038 26962 36094
rect 27018 36038 27086 36094
rect 27142 36038 27163 36094
rect 26823 34011 27163 36038
rect 26823 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27163 34011
rect 26823 33793 27163 33955
rect 26823 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27163 33793
rect 26823 33576 27163 33737
rect 26823 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27163 33576
rect 26823 33432 27163 33520
rect 26823 33380 26861 33432
rect 26913 33380 27073 33432
rect 27125 33380 27163 33432
rect 26823 33358 27163 33380
rect 26823 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27163 33358
rect 26823 33215 27163 33302
rect 26823 33163 26861 33215
rect 26913 33163 27073 33215
rect 27125 33163 27163 33215
rect 26823 33140 27163 33163
rect 26823 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27163 33140
rect 26823 32997 27163 33084
rect 26823 32945 26861 32997
rect 26913 32945 27073 32997
rect 27125 32945 27163 32997
rect 26823 32922 27163 32945
rect 26823 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27163 32922
rect 26823 32779 27163 32866
rect 26823 32727 26861 32779
rect 26913 32727 27073 32779
rect 27125 32727 27163 32779
rect 26823 32705 27163 32727
rect 26823 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27163 32705
rect 26823 32562 27163 32649
rect 26823 32510 26861 32562
rect 26913 32510 27073 32562
rect 27125 32510 27163 32562
rect 26823 32487 27163 32510
rect 26823 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27163 32487
rect 26823 32344 27163 32431
rect 26823 32292 26861 32344
rect 26913 32292 27073 32344
rect 27125 32292 27163 32344
rect 26823 32127 27163 32292
rect 26823 32088 26861 32127
rect 26913 32088 27073 32127
rect 27125 32088 27163 32127
rect 26823 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 27163 32088
rect 26823 31909 27163 32032
rect 26823 31870 26861 31909
rect 26913 31870 27073 31909
rect 27125 31870 27163 31909
rect 26823 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 27163 31870
rect 26823 31691 27163 31814
rect 26823 31652 26861 31691
rect 26913 31652 27073 31691
rect 27125 31652 27163 31691
rect 26823 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 27163 31652
rect 26823 31474 27163 31596
rect 26823 31422 26861 31474
rect 26913 31422 27073 31474
rect 27125 31422 27163 31474
rect 26823 31256 27163 31422
rect 26823 31204 26861 31256
rect 26913 31204 27073 31256
rect 27125 31204 27163 31256
rect 26823 31038 27163 31204
rect 26823 30986 26861 31038
rect 26913 30986 27073 31038
rect 27125 30986 27163 31038
rect 26823 30821 27163 30986
rect 26823 30769 26861 30821
rect 26913 30769 27073 30821
rect 27125 30769 27163 30821
rect 26823 30603 27163 30769
rect 26823 30551 26861 30603
rect 26913 30551 27073 30603
rect 27125 30551 27163 30603
rect 26823 30386 27163 30551
rect 26823 30334 26861 30386
rect 26913 30334 27073 30386
rect 27125 30334 27163 30386
rect 26823 30168 27163 30334
rect 26823 30116 26861 30168
rect 26913 30116 27073 30168
rect 27125 30116 27163 30168
rect 26823 29968 27163 30116
rect 26823 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 27163 29968
rect 26823 29898 26861 29912
rect 26913 29898 27073 29912
rect 27125 29898 27163 29912
rect 26823 29750 27163 29898
rect 26823 29694 26859 29750
rect 26915 29694 27071 29750
rect 27127 29694 27163 29750
rect 26823 29681 26861 29694
rect 26913 29681 27073 29694
rect 27125 29681 27163 29694
rect 26823 29533 27163 29681
rect 26823 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 27163 29533
rect 26823 29463 26861 29477
rect 26913 29463 27073 29477
rect 27125 29463 27163 29477
rect 26823 29315 27163 29463
rect 26823 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 27163 29315
rect 26823 29245 26861 29259
rect 26913 29245 27073 29259
rect 27125 29245 27163 29259
rect 26823 29098 27163 29245
rect 26823 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 27163 29098
rect 26823 29028 26861 29042
rect 26913 29028 27073 29042
rect 27125 29028 27163 29042
rect 26823 28880 27163 29028
rect 26823 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 27163 28880
rect 26823 28810 26861 28824
rect 26913 28810 27073 28824
rect 27125 28810 27163 28824
rect 26823 28662 27163 28810
rect 26823 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 27163 28662
rect 26823 28592 26861 28606
rect 26913 28592 27073 28606
rect 27125 28592 27163 28606
rect 26823 28444 27163 28592
rect 26823 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 27163 28444
rect 26823 28375 26861 28388
rect 26913 28375 27073 28388
rect 27125 28375 27163 28388
rect 26823 28227 27163 28375
rect 26823 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 27163 28227
rect 26823 28157 26861 28171
rect 26913 28157 27073 28171
rect 27125 28157 27163 28171
rect 26823 28009 27163 28157
rect 26823 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 27163 28009
rect 26823 27940 26861 27953
rect 26913 27940 27073 27953
rect 27125 27940 27163 27953
rect 26823 27792 27163 27940
rect 26823 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 27163 27792
rect 26823 27722 26861 27736
rect 26913 27722 27073 27736
rect 27125 27722 27163 27736
rect 26823 27574 27163 27722
rect 26823 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 27163 27574
rect 26823 27504 26861 27518
rect 26913 27504 27073 27518
rect 27125 27504 27163 27518
rect 26823 27339 27163 27504
rect 26823 27287 26861 27339
rect 26913 27287 27073 27339
rect 27125 27287 27163 27339
rect 26823 27121 27163 27287
rect 26823 27069 26861 27121
rect 26913 27069 27073 27121
rect 27125 27069 27163 27121
rect 26823 26903 27163 27069
rect 26823 26851 26861 26903
rect 26913 26851 27073 26903
rect 27125 26851 27163 26903
rect 26823 26686 27163 26851
rect 26823 26634 26861 26686
rect 26913 26634 27073 26686
rect 27125 26634 27163 26686
rect 26823 26468 27163 26634
rect 26823 26416 26861 26468
rect 26913 26416 27073 26468
rect 27125 26416 27163 26468
rect 26435 26286 26643 26321
rect 26435 26126 26450 26286
rect 26610 26126 26643 26286
rect 26077 25967 26285 26002
rect 26077 25807 26092 25967
rect 26252 25807 26285 25967
rect 25741 25647 25949 25676
rect 25741 25487 25756 25647
rect 25916 25487 25949 25647
rect 25406 25328 25614 25357
rect 25406 25168 25421 25328
rect 25581 25168 25614 25328
rect 25066 24637 25274 24666
rect 25066 24477 25081 24637
rect 25241 24477 25274 24637
rect 24729 24316 24937 24345
rect 24729 24156 24744 24316
rect 24904 24156 24937 24316
rect 24401 23995 24609 24024
rect 24401 23835 24416 23995
rect 24576 23835 24609 23995
rect 24042 23673 24250 23702
rect 24042 23513 24057 23673
rect 24217 23513 24250 23673
rect 24042 17317 24250 23513
rect 24401 17656 24609 23835
rect 24729 17977 24937 24156
rect 25066 18350 25274 24477
rect 25406 18684 25614 25168
rect 25741 19027 25949 25487
rect 26077 19347 26285 25807
rect 26435 19692 26643 26126
rect 26435 19532 26465 19692
rect 26625 19532 26643 19692
rect 26435 19502 26643 19532
rect 26823 26250 27163 26416
rect 26823 26198 26861 26250
rect 26913 26198 27073 26250
rect 27125 26198 27163 26250
rect 26823 26033 27163 26198
rect 26823 25981 26861 26033
rect 26913 25981 27073 26033
rect 27125 25981 27163 26033
rect 26823 25815 27163 25981
rect 26823 25763 26861 25815
rect 26913 25763 27073 25815
rect 27125 25763 27163 25815
rect 26823 25598 27163 25763
rect 26823 25546 26861 25598
rect 26913 25546 27073 25598
rect 27125 25546 27163 25598
rect 26823 25380 27163 25546
rect 26823 25328 26861 25380
rect 26913 25328 27073 25380
rect 27125 25328 27163 25380
rect 26823 25162 27163 25328
rect 26823 25110 26861 25162
rect 26913 25110 27073 25162
rect 27125 25110 27163 25162
rect 26823 24945 27163 25110
rect 26823 24893 26861 24945
rect 26913 24893 27073 24945
rect 27125 24893 27163 24945
rect 26823 24727 27163 24893
rect 26823 24675 26861 24727
rect 26913 24675 27073 24727
rect 27125 24675 27163 24727
rect 26823 24509 27163 24675
rect 26823 24457 26861 24509
rect 26913 24457 27073 24509
rect 27125 24457 27163 24509
rect 26823 24292 27163 24457
rect 26823 24240 26861 24292
rect 26913 24240 27073 24292
rect 27125 24240 27163 24292
rect 26823 24227 27163 24240
rect 26823 24171 26858 24227
rect 27122 24171 27163 24227
rect 26823 24085 27163 24171
rect 26823 24029 26858 24085
rect 27122 24074 27163 24085
rect 26823 24022 26861 24029
rect 26913 24022 27073 24029
rect 27125 24022 27163 24074
rect 26823 23943 27163 24022
rect 26823 23887 26858 23943
rect 27122 23887 27163 23943
rect 26823 23857 27163 23887
rect 26823 23805 26861 23857
rect 26913 23805 27073 23857
rect 27125 23805 27163 23857
rect 26823 23801 27163 23805
rect 26823 23745 26858 23801
rect 27122 23745 27163 23801
rect 26823 23659 27163 23745
rect 26823 23603 26858 23659
rect 27122 23639 27163 23659
rect 26823 23587 26861 23603
rect 26913 23587 27073 23603
rect 27125 23587 27163 23639
rect 26823 23517 27163 23587
rect 26823 23461 26858 23517
rect 27122 23461 27163 23517
rect 26823 23421 27163 23461
rect 26823 23375 26861 23421
rect 26913 23375 27073 23421
rect 26823 23319 26858 23375
rect 27125 23369 27163 23421
rect 27122 23319 27163 23369
rect 26823 23233 27163 23319
rect 26823 23177 26858 23233
rect 27122 23204 27163 23233
rect 26823 23152 26861 23177
rect 26913 23152 27073 23177
rect 27125 23152 27163 23204
rect 26823 23091 27163 23152
rect 26823 23035 26858 23091
rect 27122 23035 27163 23091
rect 26823 22986 27163 23035
rect 26823 22934 26861 22986
rect 26913 22934 27073 22986
rect 27125 22934 27163 22986
rect 26823 22768 27163 22934
rect 26823 22716 26861 22768
rect 26913 22716 27073 22768
rect 27125 22716 27163 22768
rect 26823 22551 27163 22716
rect 26823 22499 26861 22551
rect 26913 22499 27073 22551
rect 27125 22499 27163 22551
rect 26823 22333 27163 22499
rect 26823 22281 26861 22333
rect 26913 22281 27073 22333
rect 27125 22281 27163 22333
rect 26823 22115 27163 22281
rect 26823 22063 26861 22115
rect 26913 22063 27073 22115
rect 27125 22063 27163 22115
rect 26823 21898 27163 22063
rect 26823 21846 26861 21898
rect 26913 21846 27073 21898
rect 27125 21846 27163 21898
rect 26823 21680 27163 21846
rect 26823 21628 26861 21680
rect 26913 21628 27073 21680
rect 27125 21628 27163 21680
rect 26823 21463 27163 21628
rect 26823 21411 26861 21463
rect 26913 21411 27073 21463
rect 27125 21411 27163 21463
rect 26823 21245 27163 21411
rect 26823 21193 26861 21245
rect 26913 21193 27073 21245
rect 27125 21193 27163 21245
rect 26823 21027 27163 21193
rect 26823 20975 26861 21027
rect 26913 20975 27073 21027
rect 27125 20975 27163 21027
rect 26823 20810 27163 20975
rect 26823 20758 26861 20810
rect 26913 20758 27073 20810
rect 27125 20758 27163 20810
rect 26823 20592 27163 20758
rect 26823 20540 26861 20592
rect 26913 20570 27073 20592
rect 26913 20540 26924 20570
rect 27125 20540 27163 20592
rect 26823 20410 26924 20540
rect 27084 20410 27163 20540
rect 26823 20374 27163 20410
rect 26823 20322 26861 20374
rect 26913 20322 27073 20374
rect 27125 20322 27163 20374
rect 26823 20226 27163 20322
rect 26823 20157 26924 20226
rect 27084 20157 27163 20226
rect 26823 20105 26861 20157
rect 26913 20105 26924 20157
rect 27125 20105 27163 20157
rect 26823 20066 26924 20105
rect 27084 20066 27163 20105
rect 26823 19939 27163 20066
rect 26823 19887 26861 19939
rect 26913 19887 27073 19939
rect 27125 19887 27163 19939
rect 26823 19722 27163 19887
rect 26823 19670 26861 19722
rect 26913 19670 27073 19722
rect 27125 19670 27163 19722
rect 26823 19504 27163 19670
rect 26077 19187 26107 19347
rect 26267 19187 26285 19347
rect 26077 19162 26285 19187
rect 26823 19452 26861 19504
rect 26913 19452 27073 19504
rect 27125 19452 27163 19504
rect 26823 19286 27163 19452
rect 26823 19234 26861 19286
rect 26913 19234 27073 19286
rect 27125 19234 27163 19286
rect 25741 18867 25771 19027
rect 25931 18867 25949 19027
rect 25741 18822 25949 18867
rect 26823 19068 27163 19234
rect 26823 19016 26861 19068
rect 26913 19016 27073 19068
rect 27125 19016 27163 19068
rect 26823 18851 27163 19016
rect 25406 18524 25434 18684
rect 25594 18524 25614 18684
rect 25406 18482 25614 18524
rect 26823 18799 26861 18851
rect 26913 18799 27073 18851
rect 27125 18799 27163 18851
rect 26823 18633 27163 18799
rect 26823 18581 26861 18633
rect 26913 18581 27073 18633
rect 27125 18581 27163 18633
rect 25066 18190 25094 18350
rect 25254 18190 25274 18350
rect 25066 18142 25274 18190
rect 26823 18416 27163 18581
rect 26823 18364 26861 18416
rect 26913 18364 27073 18416
rect 27125 18364 27163 18416
rect 26823 18198 27163 18364
rect 26823 18146 26861 18198
rect 26913 18146 27073 18198
rect 27125 18146 27163 18198
rect 24729 17817 24757 17977
rect 24917 17817 24937 17977
rect 24729 17803 24937 17817
rect 26823 17980 27163 18146
rect 26823 17928 26861 17980
rect 26913 17928 27073 17980
rect 27125 17928 27163 17980
rect 24401 17496 24429 17656
rect 24589 17496 24609 17656
rect 24401 17462 24609 17496
rect 26823 17763 27163 17928
rect 26823 17711 26861 17763
rect 26913 17711 27073 17763
rect 27125 17711 27163 17763
rect 26823 17545 27163 17711
rect 26823 17493 26861 17545
rect 26913 17493 27073 17545
rect 27125 17493 27163 17545
rect 24042 17157 24069 17317
rect 24229 17157 24250 17317
rect 24042 17122 24250 17157
rect 26823 17327 27163 17493
rect 26823 17275 26861 17327
rect 26913 17275 27073 17327
rect 27125 17275 27163 17327
rect 26823 17110 27163 17275
rect 26823 17058 26861 17110
rect 26913 17058 27073 17110
rect 27125 17058 27163 17110
rect 26823 16892 27163 17058
rect 26823 16840 26861 16892
rect 26913 16840 27073 16892
rect 27125 16840 27163 16892
rect 26823 16675 27163 16840
rect 26823 16623 26861 16675
rect 26913 16623 27073 16675
rect 27125 16623 27163 16675
rect 26823 16457 27163 16623
rect 26823 16405 26861 16457
rect 26913 16405 27073 16457
rect 27125 16405 27163 16457
rect 26823 16239 27163 16405
rect 26823 16187 26861 16239
rect 26913 16187 27073 16239
rect 27125 16187 27163 16239
rect 26823 16022 27163 16187
rect 26823 15970 26861 16022
rect 26913 15970 27073 16022
rect 27125 15970 27163 16022
rect 26823 15804 27163 15970
rect 26823 15752 26861 15804
rect 26913 15752 27073 15804
rect 27125 15752 27163 15804
rect 26823 15586 27163 15752
rect 26823 15534 26861 15586
rect 26913 15534 27073 15586
rect 27125 15534 27163 15586
rect 26823 15369 27163 15534
rect 26823 15317 26861 15369
rect 26913 15317 27073 15369
rect 27125 15317 27163 15369
rect 26823 15151 27163 15317
rect 26823 15099 26861 15151
rect 26913 15099 27073 15151
rect 27125 15099 27163 15151
rect 26823 14933 27163 15099
rect 26823 14881 26861 14933
rect 26913 14881 27073 14933
rect 27125 14881 27163 14933
rect 26823 14716 27163 14881
rect 26823 14664 26861 14716
rect 26913 14664 27073 14716
rect 27125 14664 27163 14716
rect 26823 14498 27163 14664
rect 26823 14446 26861 14498
rect 26913 14446 27073 14498
rect 27125 14446 27163 14498
rect 26823 14281 27163 14446
rect 26823 14229 26861 14281
rect 26913 14229 27073 14281
rect 27125 14229 27163 14281
rect 26823 14119 27163 14229
rect 26823 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27163 14119
rect 26823 14011 26861 14063
rect 26913 14011 27073 14063
rect 27125 14011 27163 14063
rect 26823 13902 27163 14011
rect 26823 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27163 13902
rect 26823 13845 27163 13846
rect 26823 13793 26861 13845
rect 26913 13793 27073 13845
rect 27125 13793 27163 13845
rect 26823 13684 27163 13793
rect 26823 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27163 13684
rect 26823 13576 26861 13628
rect 26913 13576 27073 13628
rect 27125 13576 27163 13628
rect 26823 13467 27163 13576
rect 26823 13411 26859 13467
rect 26915 13411 27071 13467
rect 27127 13411 27163 13467
rect 26823 13410 27163 13411
rect 26823 13358 26861 13410
rect 26913 13358 27073 13410
rect 27125 13358 27163 13410
rect 26823 13249 27163 13358
rect 26823 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27163 13249
rect 26823 13192 27163 13193
rect 26823 13140 26861 13192
rect 26913 13140 27073 13192
rect 27125 13140 27163 13192
rect 26823 13031 27163 13140
rect 26823 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27163 13031
rect 26823 12923 26861 12975
rect 26913 12923 27073 12975
rect 27125 12923 27163 12975
rect 26823 12813 27163 12923
rect 26823 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 27163 12813
rect 26823 12705 26861 12757
rect 26913 12705 27073 12757
rect 27125 12705 27163 12757
rect 26823 12596 27163 12705
rect 26823 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12540 27163 12596
rect 26823 12488 26861 12540
rect 26913 12488 27073 12540
rect 27125 12488 27163 12540
rect 26823 12378 27163 12488
rect 26823 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 27163 12378
rect 26823 12270 26861 12322
rect 26913 12270 27073 12322
rect 27125 12270 27163 12322
rect 26823 12161 27163 12270
rect 26823 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 27163 12161
rect 26823 12104 27163 12105
rect 26823 12052 26861 12104
rect 26913 12052 27073 12104
rect 27125 12052 27163 12104
rect 26823 11887 27163 12052
rect 26823 11835 26861 11887
rect 26913 11835 27073 11887
rect 27125 11835 27163 11887
rect 26823 11669 27163 11835
rect 26823 11617 26861 11669
rect 26913 11617 27073 11669
rect 27125 11617 27163 11669
rect 26823 11451 27163 11617
rect 26823 11399 26861 11451
rect 26913 11399 27073 11451
rect 27125 11399 27163 11451
rect 26823 11234 27163 11399
rect 26823 11182 26861 11234
rect 26913 11182 27073 11234
rect 27125 11182 27163 11234
rect 26823 11016 27163 11182
rect 26823 10964 26861 11016
rect 26913 10964 27073 11016
rect 27125 10964 27163 11016
rect 26823 10798 27163 10964
rect 26823 10746 26861 10798
rect 26913 10746 27073 10798
rect 27125 10746 27163 10798
rect 26823 10581 27163 10746
rect 26823 10529 26861 10581
rect 26913 10529 27073 10581
rect 27125 10529 27163 10581
rect 26823 10363 27163 10529
rect 26823 10311 26861 10363
rect 26913 10311 27073 10363
rect 27125 10311 27163 10363
rect 26823 10146 27163 10311
rect 26823 10094 26861 10146
rect 26913 10094 27073 10146
rect 27125 10094 27163 10146
rect 26823 9928 27163 10094
rect 26823 9876 26861 9928
rect 26913 9876 27073 9928
rect 27125 9876 27163 9928
rect 26823 9710 27163 9876
rect 26823 9658 26861 9710
rect 26913 9658 27073 9710
rect 27125 9658 27163 9710
rect 26823 9493 27163 9658
rect 26823 9441 26861 9493
rect 26913 9441 27073 9493
rect 27125 9441 27163 9493
rect 26823 9407 27163 9441
rect 26823 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 27163 9407
rect 26823 9275 27163 9351
rect 26823 9223 26861 9275
rect 26913 9223 27073 9275
rect 27125 9223 27163 9275
rect 26823 9190 27163 9223
rect 26823 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 27163 9190
rect 26823 9057 27163 9134
rect 26823 9005 26861 9057
rect 26913 9005 27073 9057
rect 27125 9005 27163 9057
rect 26823 8972 27163 9005
rect 26823 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 27163 8972
rect 26823 8840 27163 8916
rect 26823 8788 26861 8840
rect 26913 8788 27073 8840
rect 27125 8788 27163 8840
rect 26823 8754 27163 8788
rect 26823 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 27163 8754
rect 26823 8622 27163 8698
rect 26823 8570 26861 8622
rect 26913 8570 27073 8622
rect 27125 8570 27163 8622
rect 26823 8536 27163 8570
rect 26823 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 27163 8536
rect 26823 8404 27163 8480
rect 26823 8352 26861 8404
rect 26913 8352 27073 8404
rect 27125 8352 27163 8404
rect 26823 8319 27163 8352
rect 26823 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 27163 8319
rect 26823 8187 27163 8263
rect 26823 8135 26861 8187
rect 26913 8135 27073 8187
rect 27125 8135 27163 8187
rect 26823 7969 27163 8135
rect 26823 7917 26861 7969
rect 26913 7917 27073 7969
rect 27125 7917 27163 7969
rect 26823 7752 27163 7917
rect 26823 7700 26861 7752
rect 26913 7700 27073 7752
rect 27125 7700 27163 7752
rect 26823 7534 27163 7700
rect 26823 7482 26861 7534
rect 26913 7482 27073 7534
rect 27125 7482 27163 7534
rect 26823 7316 27163 7482
rect 26823 7264 26861 7316
rect 26913 7264 27073 7316
rect 27125 7264 27163 7316
rect 26823 7099 27163 7264
rect 26823 7047 26861 7099
rect 26913 7047 27073 7099
rect 27125 7047 27163 7099
rect 26823 6881 27163 7047
rect 26823 6829 26861 6881
rect 26913 6829 27073 6881
rect 27125 6829 27163 6881
rect 26823 6663 27163 6829
rect 26823 6611 26861 6663
rect 26913 6611 27073 6663
rect 27125 6611 27163 6663
rect 26823 6446 27163 6611
rect 26823 6394 26861 6446
rect 26913 6394 27073 6446
rect 27125 6394 27163 6446
rect 26823 6228 27163 6394
rect 26823 6176 26861 6228
rect 26913 6176 27073 6228
rect 27125 6176 27163 6228
rect 26823 6011 27163 6176
rect 26823 5959 26861 6011
rect 26913 5959 27073 6011
rect 27125 5959 27163 6011
rect 26823 5793 27163 5959
rect 26823 5741 26861 5793
rect 26913 5741 27073 5793
rect 27125 5741 27163 5793
rect 26823 5575 27163 5741
rect 26823 5539 26861 5575
rect 26913 5539 27073 5575
rect 27125 5539 27163 5575
rect 26823 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27163 5539
rect 26823 5358 27163 5483
rect 26823 5321 26861 5358
rect 26913 5321 27073 5358
rect 27125 5321 27163 5358
rect 26823 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27163 5321
rect 26823 5226 27163 5265
rect 27387 44255 29146 44294
rect 27387 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 29146 44255
rect 27387 44160 29146 44199
rect 29485 44253 30365 44328
rect 29485 44201 29582 44253
rect 29634 44201 29793 44253
rect 29845 44201 30005 44253
rect 30057 44201 30216 44253
rect 30268 44201 30365 44253
rect 27387 42494 27828 44160
rect 29485 43355 30365 44201
rect 29485 43299 29580 43355
rect 29636 43299 29791 43355
rect 29847 43299 30003 43355
rect 30059 43299 30214 43355
rect 30270 43299 30365 43355
rect 30769 44253 32888 44776
rect 30769 44201 30807 44253
rect 30859 44201 31018 44253
rect 31070 44201 31229 44253
rect 31281 44201 31440 44253
rect 31492 44201 31651 44253
rect 31703 44201 31861 44253
rect 31913 44201 32072 44253
rect 32124 44201 32283 44253
rect 32335 44201 32494 44253
rect 32546 44201 32888 44253
rect 30769 44035 32888 44201
rect 30769 43983 30807 44035
rect 30859 43983 31018 44035
rect 31070 43983 31229 44035
rect 31281 43983 31440 44035
rect 31492 43983 31651 44035
rect 31703 43983 31861 44035
rect 31913 43983 32072 44035
rect 32124 43983 32283 44035
rect 32335 43983 32494 44035
rect 32546 43983 32888 44035
rect 30769 43818 32888 43983
rect 30769 43766 30807 43818
rect 30859 43766 31018 43818
rect 31070 43766 31229 43818
rect 31281 43766 31440 43818
rect 31492 43766 31651 43818
rect 31703 43766 31861 43818
rect 31913 43766 32072 43818
rect 32124 43766 32283 43818
rect 32335 43766 32494 43818
rect 32546 43766 32888 43818
rect 34227 44255 35024 44328
rect 34227 44199 34288 44255
rect 34344 44199 34499 44255
rect 34555 44199 34710 44255
rect 34766 44199 34921 44255
rect 34977 44199 35024 44255
rect 34227 44035 35024 44199
rect 34227 43983 34290 44035
rect 34342 43983 34501 44035
rect 34553 43983 34712 44035
rect 34764 43983 34923 44035
rect 34975 43983 35024 44035
rect 30769 43478 32888 43766
rect 33011 43774 33984 43813
rect 33011 43718 33048 43774
rect 33104 43718 33259 43774
rect 33315 43718 33470 43774
rect 33526 43718 33681 43774
rect 33737 43718 33892 43774
rect 33948 43718 33984 43774
rect 33011 43680 33984 43718
rect 34227 43478 35024 43983
rect 35128 44233 36415 44776
rect 35128 44181 35443 44233
rect 35495 44181 35654 44233
rect 35706 44181 35865 44233
rect 35917 44181 36076 44233
rect 36128 44181 36287 44233
rect 36339 44181 36415 44233
rect 35128 43770 36415 44181
rect 35128 43718 35443 43770
rect 35495 43718 35654 43770
rect 35706 43718 35865 43770
rect 35917 43718 36076 43770
rect 36128 43718 36287 43770
rect 36339 43718 36415 43770
rect 30769 43355 32889 43478
rect 30769 43340 30852 43355
rect 27387 42455 29146 42494
rect 27387 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 29146 42455
rect 27387 42360 29146 42399
rect 29485 42453 30365 43299
rect 29485 42401 29582 42453
rect 29634 42401 29793 42453
rect 29845 42401 30005 42453
rect 30057 42401 30216 42453
rect 30268 42401 30365 42453
rect 27387 40694 27828 42360
rect 29485 41555 30365 42401
rect 29485 41499 29580 41555
rect 29636 41499 29791 41555
rect 29847 41499 30003 41555
rect 30059 41499 30214 41555
rect 30270 41499 30365 41555
rect 27387 40655 29146 40694
rect 27387 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 29146 40655
rect 27387 40560 29146 40599
rect 29485 40653 30365 41499
rect 29485 40601 29582 40653
rect 29634 40601 29793 40653
rect 29845 40601 30005 40653
rect 30057 40601 30216 40653
rect 30268 40601 30365 40653
rect 27387 38894 27828 40560
rect 29485 39755 30365 40601
rect 29485 39699 29580 39755
rect 29636 39699 29791 39755
rect 29847 39699 30003 39755
rect 30059 39699 30214 39755
rect 30270 39699 30365 39755
rect 27387 38855 29146 38894
rect 27387 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 29146 38855
rect 27387 38760 29146 38799
rect 29485 38853 30365 39699
rect 29485 38801 29582 38853
rect 29634 38801 29793 38853
rect 29845 38801 30005 38853
rect 30057 38801 30216 38853
rect 30268 38801 30365 38853
rect 27387 37094 27828 38760
rect 29485 37955 30365 38801
rect 29485 37899 29580 37955
rect 29636 37899 29791 37955
rect 29847 37899 30003 37955
rect 30059 37899 30214 37955
rect 30270 37899 30365 37955
rect 27387 37055 29146 37094
rect 27387 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 29146 37055
rect 27387 36960 29146 36999
rect 29485 37053 30365 37899
rect 29485 37001 29582 37053
rect 29634 37001 29793 37053
rect 29845 37001 30005 37053
rect 30057 37001 30216 37053
rect 30268 37001 30365 37053
rect 27387 34940 27828 36960
rect 29485 36155 30365 37001
rect 29485 36099 29580 36155
rect 29636 36099 29791 36155
rect 29847 36099 30003 36155
rect 30059 36099 30214 36155
rect 30270 36099 30365 36155
rect 29485 36027 30365 36099
rect 30770 43299 30852 43340
rect 30908 43299 31063 43355
rect 31119 43299 31274 43355
rect 31330 43299 31484 43355
rect 31540 43299 31695 43355
rect 31751 43299 31907 43355
rect 31963 43299 32118 43355
rect 32174 43299 32328 43355
rect 32384 43299 32539 43355
rect 32595 43299 32750 43355
rect 32806 43299 32889 43355
rect 34227 43353 35025 43478
rect 34227 43340 34284 43353
rect 30770 42453 32889 43299
rect 34228 43301 34284 43340
rect 34336 43301 34495 43353
rect 34547 43301 34707 43353
rect 34759 43301 34918 43353
rect 34970 43301 35025 43353
rect 35128 43355 36415 43718
rect 35128 43340 35218 43355
rect 33019 43129 33327 43170
rect 33019 43077 33057 43129
rect 33109 43077 33237 43129
rect 33289 43077 33327 43129
rect 33019 42922 33327 43077
rect 33019 42866 33055 42922
rect 33111 42866 33235 42922
rect 33291 42866 33327 42922
rect 33019 42681 33327 42866
rect 33731 43137 34090 43178
rect 33731 43085 33819 43137
rect 33871 43085 33999 43137
rect 34051 43085 34090 43137
rect 33731 42915 34090 43085
rect 33731 42859 33817 42915
rect 33873 42859 33997 42915
rect 34053 42859 34090 42915
rect 33731 42786 34090 42859
rect 34228 42891 35025 43301
rect 34228 42839 34267 42891
rect 34319 42839 34447 42891
rect 34499 42839 34627 42891
rect 34679 42839 35025 42891
rect 33019 42629 33057 42681
rect 33109 42629 33237 42681
rect 33289 42629 33327 42681
rect 33019 42589 33327 42629
rect 30770 42401 30854 42453
rect 30906 42401 31065 42453
rect 31117 42401 31276 42453
rect 31328 42401 31486 42453
rect 31538 42401 31697 42453
rect 31749 42401 31909 42453
rect 31961 42401 32120 42453
rect 32172 42401 32330 42453
rect 32382 42401 32541 42453
rect 32593 42401 32752 42453
rect 32804 42401 32889 42453
rect 30770 41555 32889 42401
rect 34228 42455 35025 42839
rect 34228 42399 34282 42455
rect 34338 42399 34493 42455
rect 34549 42399 34705 42455
rect 34761 42453 34916 42455
rect 34972 42453 35025 42455
rect 34807 42401 34916 42453
rect 34987 42401 35025 42453
rect 34761 42399 34916 42401
rect 34972 42399 35025 42401
rect 33019 42225 33327 42265
rect 33019 42173 33057 42225
rect 33109 42173 33237 42225
rect 33289 42173 33327 42225
rect 33019 41988 33327 42173
rect 33019 41932 33055 41988
rect 33111 41932 33235 41988
rect 33291 41932 33327 41988
rect 33019 41777 33327 41932
rect 33019 41725 33057 41777
rect 33109 41725 33237 41777
rect 33289 41725 33327 41777
rect 33019 41684 33327 41725
rect 33731 41995 34090 42068
rect 33731 41939 33817 41995
rect 33873 41939 33997 41995
rect 34053 41939 34090 41995
rect 33731 41769 34090 41939
rect 33731 41717 33819 41769
rect 33871 41717 33999 41769
rect 34051 41717 34090 41769
rect 33731 41676 34090 41717
rect 34228 42015 35025 42399
rect 34228 41963 34267 42015
rect 34319 41963 34447 42015
rect 34499 41963 34627 42015
rect 34679 41963 35025 42015
rect 30770 41499 30852 41555
rect 30908 41499 31063 41555
rect 31119 41499 31274 41555
rect 31330 41499 31484 41555
rect 31540 41499 31695 41555
rect 31751 41499 31907 41555
rect 31963 41499 32118 41555
rect 32174 41499 32328 41555
rect 32384 41499 32539 41555
rect 32595 41499 32750 41555
rect 32806 41499 32889 41555
rect 30770 40653 32889 41499
rect 34228 41553 35025 41963
rect 34228 41501 34284 41553
rect 34336 41501 34495 41553
rect 34547 41501 34707 41553
rect 34759 41501 34918 41553
rect 34970 41501 35025 41553
rect 33019 41329 33327 41370
rect 33019 41277 33057 41329
rect 33109 41277 33237 41329
rect 33289 41277 33327 41329
rect 33019 41122 33327 41277
rect 33019 41066 33055 41122
rect 33111 41066 33235 41122
rect 33291 41066 33327 41122
rect 33019 40881 33327 41066
rect 33731 41337 34090 41378
rect 33731 41285 33819 41337
rect 33871 41285 33999 41337
rect 34051 41285 34090 41337
rect 33731 41115 34090 41285
rect 33731 41059 33817 41115
rect 33873 41059 33997 41115
rect 34053 41059 34090 41115
rect 33731 40986 34090 41059
rect 34228 41091 35025 41501
rect 34228 41039 34267 41091
rect 34319 41039 34447 41091
rect 34499 41039 34627 41091
rect 34679 41039 35025 41091
rect 33019 40829 33057 40881
rect 33109 40829 33237 40881
rect 33289 40829 33327 40881
rect 33019 40789 33327 40829
rect 30770 40601 30854 40653
rect 30906 40601 31065 40653
rect 31117 40601 31276 40653
rect 31328 40601 31486 40653
rect 31538 40601 31697 40653
rect 31749 40601 31909 40653
rect 31961 40601 32120 40653
rect 32172 40601 32330 40653
rect 32382 40601 32541 40653
rect 32593 40601 32752 40653
rect 32804 40601 32889 40653
rect 30770 39755 32889 40601
rect 34228 40655 35025 41039
rect 34228 40599 34282 40655
rect 34338 40599 34493 40655
rect 34549 40599 34705 40655
rect 34761 40653 34916 40655
rect 34972 40653 35025 40655
rect 34807 40601 34916 40653
rect 34987 40601 35025 40653
rect 34761 40599 34916 40601
rect 34972 40599 35025 40601
rect 33019 40425 33327 40465
rect 33019 40373 33057 40425
rect 33109 40373 33237 40425
rect 33289 40373 33327 40425
rect 33019 40188 33327 40373
rect 33019 40132 33055 40188
rect 33111 40132 33235 40188
rect 33291 40132 33327 40188
rect 33019 39977 33327 40132
rect 33019 39925 33057 39977
rect 33109 39925 33237 39977
rect 33289 39925 33327 39977
rect 33019 39884 33327 39925
rect 33731 40195 34090 40268
rect 33731 40139 33817 40195
rect 33873 40139 33997 40195
rect 34053 40139 34090 40195
rect 33731 39969 34090 40139
rect 33731 39917 33819 39969
rect 33871 39917 33999 39969
rect 34051 39917 34090 39969
rect 33731 39876 34090 39917
rect 34228 40215 35025 40599
rect 34228 40163 34267 40215
rect 34319 40163 34447 40215
rect 34499 40163 34627 40215
rect 34679 40163 35025 40215
rect 30770 39699 30852 39755
rect 30908 39699 31063 39755
rect 31119 39699 31274 39755
rect 31330 39699 31484 39755
rect 31540 39699 31695 39755
rect 31751 39699 31907 39755
rect 31963 39699 32118 39755
rect 32174 39699 32328 39755
rect 32384 39699 32539 39755
rect 32595 39699 32750 39755
rect 32806 39699 32889 39755
rect 30770 38853 32889 39699
rect 34228 39753 35025 40163
rect 34228 39701 34284 39753
rect 34336 39701 34495 39753
rect 34547 39701 34707 39753
rect 34759 39701 34918 39753
rect 34970 39701 35025 39753
rect 33019 39529 33327 39570
rect 33019 39477 33057 39529
rect 33109 39477 33237 39529
rect 33289 39477 33327 39529
rect 33019 39322 33327 39477
rect 33019 39266 33055 39322
rect 33111 39266 33235 39322
rect 33291 39266 33327 39322
rect 33019 39081 33327 39266
rect 33731 39537 34090 39578
rect 33731 39485 33819 39537
rect 33871 39485 33999 39537
rect 34051 39485 34090 39537
rect 33731 39315 34090 39485
rect 33731 39259 33817 39315
rect 33873 39259 33997 39315
rect 34053 39259 34090 39315
rect 33731 39186 34090 39259
rect 34228 39291 35025 39701
rect 34228 39239 34267 39291
rect 34319 39239 34447 39291
rect 34499 39239 34627 39291
rect 34679 39239 35025 39291
rect 33019 39029 33057 39081
rect 33109 39029 33237 39081
rect 33289 39029 33327 39081
rect 33019 38989 33327 39029
rect 30770 38801 30854 38853
rect 30906 38801 31065 38853
rect 31117 38801 31276 38853
rect 31328 38801 31486 38853
rect 31538 38801 31697 38853
rect 31749 38801 31909 38853
rect 31961 38801 32120 38853
rect 32172 38801 32330 38853
rect 32382 38801 32541 38853
rect 32593 38801 32752 38853
rect 32804 38801 32889 38853
rect 30770 37955 32889 38801
rect 34228 38855 35025 39239
rect 34228 38799 34282 38855
rect 34338 38799 34493 38855
rect 34549 38799 34705 38855
rect 34761 38853 34916 38855
rect 34972 38853 35025 38855
rect 34807 38801 34916 38853
rect 34987 38801 35025 38853
rect 34761 38799 34916 38801
rect 34972 38799 35025 38801
rect 33019 38625 33327 38665
rect 33019 38573 33057 38625
rect 33109 38573 33237 38625
rect 33289 38573 33327 38625
rect 33019 38388 33327 38573
rect 33019 38332 33055 38388
rect 33111 38332 33235 38388
rect 33291 38332 33327 38388
rect 33019 38177 33327 38332
rect 33019 38125 33057 38177
rect 33109 38125 33237 38177
rect 33289 38125 33327 38177
rect 33019 38084 33327 38125
rect 33731 38395 34090 38468
rect 33731 38339 33817 38395
rect 33873 38339 33997 38395
rect 34053 38339 34090 38395
rect 33731 38169 34090 38339
rect 33731 38117 33819 38169
rect 33871 38117 33999 38169
rect 34051 38117 34090 38169
rect 33731 38076 34090 38117
rect 34228 38415 35025 38799
rect 34228 38363 34267 38415
rect 34319 38363 34447 38415
rect 34499 38363 34627 38415
rect 34679 38363 35025 38415
rect 30770 37899 30852 37955
rect 30908 37899 31063 37955
rect 31119 37899 31274 37955
rect 31330 37899 31484 37955
rect 31540 37899 31695 37955
rect 31751 37899 31907 37955
rect 31963 37899 32118 37955
rect 32174 37899 32328 37955
rect 32384 37899 32539 37955
rect 32595 37899 32750 37955
rect 32806 37899 32889 37955
rect 30770 37053 32889 37899
rect 34228 37953 35025 38363
rect 34228 37901 34284 37953
rect 34336 37901 34495 37953
rect 34547 37901 34707 37953
rect 34759 37901 34918 37953
rect 34970 37901 35025 37953
rect 33019 37729 33327 37770
rect 33019 37677 33057 37729
rect 33109 37677 33237 37729
rect 33289 37677 33327 37729
rect 33019 37522 33327 37677
rect 33019 37466 33055 37522
rect 33111 37466 33235 37522
rect 33291 37466 33327 37522
rect 33019 37281 33327 37466
rect 33731 37737 34090 37778
rect 33731 37685 33819 37737
rect 33871 37685 33999 37737
rect 34051 37685 34090 37737
rect 33731 37515 34090 37685
rect 33731 37459 33817 37515
rect 33873 37459 33997 37515
rect 34053 37459 34090 37515
rect 33731 37386 34090 37459
rect 34228 37491 35025 37901
rect 34228 37439 34267 37491
rect 34319 37439 34447 37491
rect 34499 37439 34627 37491
rect 34679 37439 35025 37491
rect 33019 37229 33057 37281
rect 33109 37229 33237 37281
rect 33289 37229 33327 37281
rect 33019 37189 33327 37229
rect 30770 37001 30854 37053
rect 30906 37001 31065 37053
rect 31117 37001 31276 37053
rect 31328 37001 31486 37053
rect 31538 37001 31697 37053
rect 31749 37001 31909 37053
rect 31961 37001 32120 37053
rect 32172 37001 32330 37053
rect 32382 37001 32541 37053
rect 32593 37001 32752 37053
rect 32804 37001 32889 37053
rect 30770 36155 32889 37001
rect 34228 37055 35025 37439
rect 34228 36999 34282 37055
rect 34338 36999 34493 37055
rect 34549 36999 34705 37055
rect 34761 37053 34916 37055
rect 34972 37053 35025 37055
rect 34807 37001 34916 37053
rect 34987 37001 35025 37053
rect 34761 36999 34916 37001
rect 34972 36999 35025 37001
rect 33019 36825 33327 36865
rect 33019 36773 33057 36825
rect 33109 36773 33237 36825
rect 33289 36773 33327 36825
rect 33019 36588 33327 36773
rect 33019 36532 33055 36588
rect 33111 36532 33235 36588
rect 33291 36532 33327 36588
rect 33019 36377 33327 36532
rect 33019 36325 33057 36377
rect 33109 36325 33237 36377
rect 33289 36325 33327 36377
rect 33019 36284 33327 36325
rect 33731 36595 34090 36668
rect 33731 36539 33817 36595
rect 33873 36539 33997 36595
rect 34053 36539 34090 36595
rect 33731 36369 34090 36539
rect 33731 36317 33819 36369
rect 33871 36317 33999 36369
rect 34051 36317 34090 36369
rect 33731 36276 34090 36317
rect 34228 36615 35025 36999
rect 34228 36563 34267 36615
rect 34319 36563 34447 36615
rect 34499 36563 34627 36615
rect 34679 36563 35025 36615
rect 30770 36099 30852 36155
rect 30908 36099 31063 36155
rect 31119 36099 31274 36155
rect 31330 36099 31484 36155
rect 31540 36099 31695 36155
rect 31751 36099 31907 36155
rect 31963 36099 32118 36155
rect 32174 36099 32328 36155
rect 32384 36099 32539 36155
rect 32595 36099 32750 36155
rect 32806 36099 32889 36155
rect 30770 35976 32889 36099
rect 34228 36153 35025 36563
rect 34228 36101 34284 36153
rect 34336 36101 34495 36153
rect 34547 36101 34707 36153
rect 34759 36101 34918 36153
rect 34970 36101 35025 36153
rect 34228 35976 35025 36101
rect 35131 43299 35218 43340
rect 35274 43299 35428 43355
rect 35484 43299 35639 43355
rect 35695 43299 35851 43355
rect 35907 43299 36062 43355
rect 36118 43299 36272 43355
rect 36328 43299 36415 43355
rect 36863 43772 37743 43811
rect 36863 43716 36899 43772
rect 36955 43716 37110 43772
rect 37166 43716 37321 43772
rect 37377 43716 37532 43772
rect 37588 43716 37743 43772
rect 36863 43478 37743 43716
rect 38268 43478 38863 44328
rect 38953 44001 39618 44776
rect 38953 43949 39053 44001
rect 39105 43949 39264 44001
rect 39316 43949 39475 44001
rect 39527 43949 39618 44001
rect 38953 43478 39618 43949
rect 40214 44258 40523 44328
rect 42671 44305 43222 44346
rect 40214 44255 40252 44258
rect 40304 44255 40432 44258
rect 40484 44255 40523 44258
rect 40214 44199 40250 44255
rect 40306 44199 40430 44255
rect 40486 44199 40523 44255
rect 40214 44040 40523 44199
rect 42208 44244 42548 44285
rect 42208 44192 42246 44244
rect 42298 44192 42458 44244
rect 42510 44192 42548 44244
rect 42208 44151 42548 44192
rect 42671 44253 42710 44305
rect 42762 44253 42921 44305
rect 42973 44253 43132 44305
rect 43184 44253 43222 44305
rect 40214 43988 40252 44040
rect 40304 43988 40432 44040
rect 40484 43988 40523 44040
rect 40214 43478 40523 43988
rect 40971 43772 42155 43811
rect 40971 43716 41008 43772
rect 41064 43716 41219 43772
rect 41275 43716 41430 43772
rect 41486 43716 41641 43772
rect 41697 43716 41852 43772
rect 41908 43716 42062 43772
rect 42118 43716 42155 43772
rect 40971 43677 42155 43716
rect 42671 43765 43222 44253
rect 42671 43709 42708 43765
rect 42764 43709 42919 43765
rect 42975 43709 43130 43765
rect 43186 43709 43222 43765
rect 42671 43491 43222 43709
rect 43703 44305 44564 44346
rect 43703 44253 43777 44305
rect 43829 44253 43988 44305
rect 44040 44253 44199 44305
rect 44251 44253 44410 44305
rect 44462 44253 44564 44305
rect 40717 43478 41316 43491
rect 36863 43340 37744 43478
rect 38268 43353 38864 43478
rect 38268 43340 38330 43353
rect 35131 43051 36415 43299
rect 35131 42999 35332 43051
rect 35384 42999 35543 43051
rect 35595 42999 35754 43051
rect 35806 42999 35965 43051
rect 36017 42999 36176 43051
rect 36228 42999 36415 43051
rect 35131 42591 36415 42999
rect 36640 42963 36768 43002
rect 36640 42907 36676 42963
rect 36732 42940 36768 42963
rect 36732 42907 36769 42940
rect 36640 42816 36769 42907
rect 36640 42764 36678 42816
rect 36730 42764 36769 42816
rect 36640 42723 36769 42764
rect 36864 42823 37744 43340
rect 38269 43301 38330 43340
rect 38382 43301 38541 43353
rect 38593 43301 38752 43353
rect 38804 43301 38864 43353
rect 38953 43355 39619 43478
rect 38953 43340 39050 43355
rect 36864 42771 36961 42823
rect 37013 42771 37172 42823
rect 37224 42771 37384 42823
rect 37436 42771 37595 42823
rect 37647 42771 37744 42823
rect 35131 42539 35332 42591
rect 35384 42539 35543 42591
rect 35595 42539 35754 42591
rect 35806 42539 35965 42591
rect 36017 42539 36176 42591
rect 36228 42539 36415 42591
rect 35131 42315 36415 42539
rect 35131 42263 35332 42315
rect 35384 42263 35543 42315
rect 35595 42263 35754 42315
rect 35806 42263 35965 42315
rect 36017 42263 36176 42315
rect 36228 42263 36415 42315
rect 35131 41855 36415 42263
rect 35131 41803 35332 41855
rect 35384 41803 35543 41855
rect 35595 41803 35754 41855
rect 35806 41803 35965 41855
rect 36017 41803 36176 41855
rect 36228 41803 36415 41855
rect 36640 42090 36769 42131
rect 36640 42038 36678 42090
rect 36730 42038 36769 42090
rect 36640 41947 36769 42038
rect 36640 41891 36676 41947
rect 36732 41914 36769 41947
rect 36864 42083 37744 42771
rect 37852 43063 38161 43104
rect 37852 43011 37891 43063
rect 37943 43011 38071 43063
rect 38123 43011 38161 43063
rect 37852 42732 38161 43011
rect 37852 42676 37889 42732
rect 37945 42676 38069 42732
rect 38125 42676 38161 42732
rect 37852 42589 38161 42676
rect 37852 42537 37891 42589
rect 37943 42537 38071 42589
rect 38123 42537 38161 42589
rect 37852 42496 38161 42537
rect 38269 42455 38864 43301
rect 38269 42399 38328 42455
rect 38384 42399 38539 42455
rect 38595 42399 38750 42455
rect 38806 42399 38864 42455
rect 36864 42031 36961 42083
rect 37013 42031 37172 42083
rect 37224 42031 37384 42083
rect 37436 42031 37595 42083
rect 37647 42031 37744 42083
rect 36732 41891 36768 41914
rect 36640 41852 36768 41891
rect 35131 41555 36415 41803
rect 35131 41499 35218 41555
rect 35274 41499 35428 41555
rect 35484 41499 35639 41555
rect 35695 41499 35851 41555
rect 35907 41499 36062 41555
rect 36118 41499 36272 41555
rect 36328 41499 36415 41555
rect 35131 41251 36415 41499
rect 35131 41199 35332 41251
rect 35384 41199 35543 41251
rect 35595 41199 35754 41251
rect 35806 41199 35965 41251
rect 36017 41199 36176 41251
rect 36228 41199 36415 41251
rect 35131 40791 36415 41199
rect 36640 41163 36768 41202
rect 36640 41107 36676 41163
rect 36732 41140 36768 41163
rect 36732 41107 36769 41140
rect 36640 41016 36769 41107
rect 36640 40964 36678 41016
rect 36730 40964 36769 41016
rect 36640 40923 36769 40964
rect 36864 41023 37744 42031
rect 37852 42317 38161 42358
rect 37852 42265 37891 42317
rect 37943 42265 38071 42317
rect 38123 42265 38161 42317
rect 37852 42178 38161 42265
rect 37852 42122 37889 42178
rect 37945 42122 38069 42178
rect 38125 42122 38161 42178
rect 37852 41843 38161 42122
rect 37852 41791 37891 41843
rect 37943 41791 38071 41843
rect 38123 41791 38161 41843
rect 37852 41750 38161 41791
rect 38269 41553 38864 42399
rect 38269 41501 38330 41553
rect 38382 41501 38541 41553
rect 38593 41501 38752 41553
rect 38804 41501 38864 41553
rect 36864 40971 36961 41023
rect 37013 40971 37172 41023
rect 37224 40971 37384 41023
rect 37436 40971 37595 41023
rect 37647 40971 37744 41023
rect 35131 40739 35332 40791
rect 35384 40739 35543 40791
rect 35595 40739 35754 40791
rect 35806 40739 35965 40791
rect 36017 40739 36176 40791
rect 36228 40739 36415 40791
rect 35131 40515 36415 40739
rect 35131 40463 35332 40515
rect 35384 40463 35543 40515
rect 35595 40463 35754 40515
rect 35806 40463 35965 40515
rect 36017 40463 36176 40515
rect 36228 40463 36415 40515
rect 35131 40055 36415 40463
rect 35131 40003 35332 40055
rect 35384 40003 35543 40055
rect 35595 40003 35754 40055
rect 35806 40003 35965 40055
rect 36017 40003 36176 40055
rect 36228 40003 36415 40055
rect 36640 40290 36769 40331
rect 36640 40238 36678 40290
rect 36730 40238 36769 40290
rect 36640 40147 36769 40238
rect 36640 40091 36676 40147
rect 36732 40114 36769 40147
rect 36864 40283 37744 40971
rect 37852 41263 38161 41304
rect 37852 41211 37891 41263
rect 37943 41211 38071 41263
rect 38123 41211 38161 41263
rect 37852 40932 38161 41211
rect 37852 40876 37889 40932
rect 37945 40876 38069 40932
rect 38125 40876 38161 40932
rect 37852 40789 38161 40876
rect 37852 40737 37891 40789
rect 37943 40737 38071 40789
rect 38123 40737 38161 40789
rect 37852 40696 38161 40737
rect 38269 40655 38864 41501
rect 38269 40599 38328 40655
rect 38384 40599 38539 40655
rect 38595 40599 38750 40655
rect 38806 40599 38864 40655
rect 36864 40231 36961 40283
rect 37013 40231 37172 40283
rect 37224 40231 37384 40283
rect 37436 40231 37595 40283
rect 37647 40231 37744 40283
rect 36732 40091 36768 40114
rect 36640 40052 36768 40091
rect 35131 39755 36415 40003
rect 35131 39699 35218 39755
rect 35274 39699 35428 39755
rect 35484 39699 35639 39755
rect 35695 39699 35851 39755
rect 35907 39699 36062 39755
rect 36118 39699 36272 39755
rect 36328 39699 36415 39755
rect 35131 39451 36415 39699
rect 35131 39399 35332 39451
rect 35384 39399 35543 39451
rect 35595 39399 35754 39451
rect 35806 39399 35965 39451
rect 36017 39399 36176 39451
rect 36228 39399 36415 39451
rect 35131 38991 36415 39399
rect 36640 39363 36768 39402
rect 36640 39307 36676 39363
rect 36732 39340 36768 39363
rect 36732 39307 36769 39340
rect 36640 39216 36769 39307
rect 36640 39164 36678 39216
rect 36730 39164 36769 39216
rect 36640 39123 36769 39164
rect 36864 39223 37744 40231
rect 37852 40517 38161 40558
rect 37852 40465 37891 40517
rect 37943 40465 38071 40517
rect 38123 40465 38161 40517
rect 37852 40378 38161 40465
rect 37852 40322 37889 40378
rect 37945 40322 38069 40378
rect 38125 40322 38161 40378
rect 37852 40043 38161 40322
rect 37852 39991 37891 40043
rect 37943 39991 38071 40043
rect 38123 39991 38161 40043
rect 37852 39950 38161 39991
rect 38269 39753 38864 40599
rect 38269 39701 38330 39753
rect 38382 39701 38541 39753
rect 38593 39701 38752 39753
rect 38804 39701 38864 39753
rect 36864 39171 36961 39223
rect 37013 39171 37172 39223
rect 37224 39171 37384 39223
rect 37436 39171 37595 39223
rect 37647 39171 37744 39223
rect 35131 38939 35332 38991
rect 35384 38939 35543 38991
rect 35595 38939 35754 38991
rect 35806 38939 35965 38991
rect 36017 38939 36176 38991
rect 36228 38939 36415 38991
rect 35131 38715 36415 38939
rect 35131 38663 35332 38715
rect 35384 38663 35543 38715
rect 35595 38663 35754 38715
rect 35806 38663 35965 38715
rect 36017 38663 36176 38715
rect 36228 38663 36415 38715
rect 35131 38255 36415 38663
rect 35131 38203 35332 38255
rect 35384 38203 35543 38255
rect 35595 38203 35754 38255
rect 35806 38203 35965 38255
rect 36017 38203 36176 38255
rect 36228 38203 36415 38255
rect 36640 38490 36769 38531
rect 36640 38438 36678 38490
rect 36730 38438 36769 38490
rect 36640 38347 36769 38438
rect 36640 38291 36676 38347
rect 36732 38314 36769 38347
rect 36864 38483 37744 39171
rect 37852 39463 38161 39504
rect 37852 39411 37891 39463
rect 37943 39411 38071 39463
rect 38123 39411 38161 39463
rect 37852 39132 38161 39411
rect 37852 39076 37889 39132
rect 37945 39076 38069 39132
rect 38125 39076 38161 39132
rect 37852 38989 38161 39076
rect 37852 38937 37891 38989
rect 37943 38937 38071 38989
rect 38123 38937 38161 38989
rect 37852 38896 38161 38937
rect 38269 38855 38864 39701
rect 38269 38799 38328 38855
rect 38384 38799 38539 38855
rect 38595 38799 38750 38855
rect 38806 38799 38864 38855
rect 36864 38431 36961 38483
rect 37013 38431 37172 38483
rect 37224 38431 37384 38483
rect 37436 38431 37595 38483
rect 37647 38431 37744 38483
rect 36732 38291 36768 38314
rect 36640 38252 36768 38291
rect 35131 37955 36415 38203
rect 35131 37899 35218 37955
rect 35274 37899 35428 37955
rect 35484 37899 35639 37955
rect 35695 37899 35851 37955
rect 35907 37899 36062 37955
rect 36118 37899 36272 37955
rect 36328 37899 36415 37955
rect 35131 37651 36415 37899
rect 35131 37599 35332 37651
rect 35384 37599 35543 37651
rect 35595 37599 35754 37651
rect 35806 37599 35965 37651
rect 36017 37599 36176 37651
rect 36228 37599 36415 37651
rect 35131 37191 36415 37599
rect 36640 37563 36768 37602
rect 36640 37507 36676 37563
rect 36732 37540 36768 37563
rect 36732 37507 36769 37540
rect 36640 37416 36769 37507
rect 36640 37364 36678 37416
rect 36730 37364 36769 37416
rect 36640 37323 36769 37364
rect 36864 37423 37744 38431
rect 37852 38717 38161 38758
rect 37852 38665 37891 38717
rect 37943 38665 38071 38717
rect 38123 38665 38161 38717
rect 37852 38578 38161 38665
rect 37852 38522 37889 38578
rect 37945 38522 38069 38578
rect 38125 38522 38161 38578
rect 37852 38243 38161 38522
rect 37852 38191 37891 38243
rect 37943 38191 38071 38243
rect 38123 38191 38161 38243
rect 37852 38150 38161 38191
rect 38269 37953 38864 38799
rect 38269 37901 38330 37953
rect 38382 37901 38541 37953
rect 38593 37901 38752 37953
rect 38804 37901 38864 37953
rect 36864 37371 36961 37423
rect 37013 37371 37172 37423
rect 37224 37371 37384 37423
rect 37436 37371 37595 37423
rect 37647 37371 37744 37423
rect 35131 37139 35332 37191
rect 35384 37139 35543 37191
rect 35595 37139 35754 37191
rect 35806 37139 35965 37191
rect 36017 37139 36176 37191
rect 36228 37139 36415 37191
rect 35131 36915 36415 37139
rect 35131 36863 35332 36915
rect 35384 36863 35543 36915
rect 35595 36863 35754 36915
rect 35806 36863 35965 36915
rect 36017 36863 36176 36915
rect 36228 36863 36415 36915
rect 35131 36455 36415 36863
rect 35131 36403 35332 36455
rect 35384 36403 35543 36455
rect 35595 36403 35754 36455
rect 35806 36403 35965 36455
rect 36017 36403 36176 36455
rect 36228 36403 36415 36455
rect 36640 36690 36769 36731
rect 36640 36638 36678 36690
rect 36730 36638 36769 36690
rect 36864 36683 37744 37371
rect 37852 37663 38161 37704
rect 37852 37611 37891 37663
rect 37943 37611 38071 37663
rect 38123 37611 38161 37663
rect 37852 37332 38161 37611
rect 37852 37276 37889 37332
rect 37945 37276 38069 37332
rect 38125 37276 38161 37332
rect 37852 37189 38161 37276
rect 37852 37137 37891 37189
rect 37943 37137 38071 37189
rect 38123 37137 38161 37189
rect 37852 37096 38161 37137
rect 38269 37055 38864 37901
rect 38269 36999 38328 37055
rect 38384 36999 38539 37055
rect 38595 36999 38750 37055
rect 38806 36999 38864 37055
rect 36864 36650 36961 36683
rect 36640 36547 36769 36638
rect 36640 36491 36676 36547
rect 36732 36514 36769 36547
rect 36863 36631 36961 36650
rect 37013 36631 37172 36683
rect 37224 36631 37384 36683
rect 37436 36631 37595 36683
rect 37647 36631 37744 36683
rect 36732 36491 36768 36514
rect 36640 36452 36768 36491
rect 35131 36155 36415 36403
rect 35131 36099 35218 36155
rect 35274 36099 35428 36155
rect 35484 36099 35639 36155
rect 35695 36099 35851 36155
rect 35907 36099 36062 36155
rect 36118 36099 36272 36155
rect 36328 36099 36415 36155
rect 35131 35976 36415 36099
rect 36863 35976 37744 36631
rect 37852 36917 38161 36958
rect 37852 36865 37891 36917
rect 37943 36865 38071 36917
rect 38123 36865 38161 36917
rect 37852 36778 38161 36865
rect 37852 36722 37889 36778
rect 37945 36722 38069 36778
rect 38125 36722 38161 36778
rect 37852 36443 38161 36722
rect 37852 36391 37891 36443
rect 37943 36391 38071 36443
rect 38123 36391 38161 36443
rect 37852 36350 38161 36391
rect 38269 36153 38864 36999
rect 38269 36101 38330 36153
rect 38382 36101 38541 36153
rect 38593 36101 38752 36153
rect 38804 36101 38864 36153
rect 38269 35976 38864 36101
rect 38967 43299 39050 43340
rect 39106 43299 39230 43355
rect 39286 43299 39619 43355
rect 40214 43353 40524 43478
rect 40214 43340 40253 43353
rect 38967 41555 39619 43299
rect 40215 43301 40253 43340
rect 40305 43301 40433 43353
rect 40485 43301 40524 43353
rect 39736 43115 39865 43156
rect 39736 43063 39775 43115
rect 39827 43063 39865 43115
rect 39736 42732 39865 43063
rect 39736 42676 39773 42732
rect 39829 42676 39865 42732
rect 39736 42637 39865 42676
rect 39956 42963 40084 43002
rect 39956 42907 39992 42963
rect 40048 42941 40084 42963
rect 40048 42907 40085 42941
rect 39956 42900 40085 42907
rect 39956 42848 39994 42900
rect 40046 42848 40085 42900
rect 39956 42714 40085 42848
rect 39956 42662 39994 42714
rect 40046 42662 40085 42714
rect 39956 42621 40085 42662
rect 40215 42455 40524 43301
rect 40717 43355 41317 43478
rect 40717 43299 40777 43355
rect 40833 43299 40988 43355
rect 41044 43299 41199 43355
rect 41255 43299 41317 43355
rect 40717 43226 41317 43299
rect 40215 42399 40251 42455
rect 40307 42399 40431 42455
rect 40487 42399 40524 42455
rect 39736 42178 39865 42217
rect 39736 42122 39773 42178
rect 39829 42122 39865 42178
rect 39736 41791 39865 42122
rect 39956 42192 40085 42233
rect 39956 42140 39994 42192
rect 40046 42140 40085 42192
rect 39956 42006 40085 42140
rect 39956 41954 39994 42006
rect 40046 41954 40085 42006
rect 39956 41947 40085 41954
rect 39956 41891 39992 41947
rect 40048 41913 40085 41947
rect 40048 41891 40084 41913
rect 39956 41852 40084 41891
rect 39736 41739 39775 41791
rect 39827 41739 39865 41791
rect 39736 41698 39865 41739
rect 38967 41499 39050 41555
rect 39106 41499 39230 41555
rect 39286 41499 39619 41555
rect 38967 39755 39619 41499
rect 40215 41553 40524 42399
rect 40215 41501 40253 41553
rect 40305 41501 40433 41553
rect 40485 41501 40524 41553
rect 39736 41315 39865 41356
rect 39736 41263 39775 41315
rect 39827 41263 39865 41315
rect 39736 40932 39865 41263
rect 39736 40876 39773 40932
rect 39829 40876 39865 40932
rect 39736 40837 39865 40876
rect 39956 41163 40084 41202
rect 39956 41107 39992 41163
rect 40048 41141 40084 41163
rect 40048 41107 40085 41141
rect 39956 41100 40085 41107
rect 39956 41048 39994 41100
rect 40046 41048 40085 41100
rect 39956 40914 40085 41048
rect 39956 40862 39994 40914
rect 40046 40862 40085 40914
rect 39956 40821 40085 40862
rect 40215 40655 40524 41501
rect 40215 40599 40251 40655
rect 40307 40599 40431 40655
rect 40487 40599 40524 40655
rect 39736 40378 39865 40417
rect 39736 40322 39773 40378
rect 39829 40322 39865 40378
rect 39736 39991 39865 40322
rect 39956 40392 40085 40433
rect 39956 40340 39994 40392
rect 40046 40340 40085 40392
rect 39956 40206 40085 40340
rect 39956 40154 39994 40206
rect 40046 40154 40085 40206
rect 39956 40147 40085 40154
rect 39956 40091 39992 40147
rect 40048 40113 40085 40147
rect 40048 40091 40084 40113
rect 39956 40052 40084 40091
rect 39736 39939 39775 39991
rect 39827 39939 39865 39991
rect 39736 39898 39865 39939
rect 38967 39699 39050 39755
rect 39106 39699 39230 39755
rect 39286 39699 39619 39755
rect 38967 37955 39619 39699
rect 40215 39753 40524 40599
rect 40215 39701 40253 39753
rect 40305 39701 40433 39753
rect 40485 39701 40524 39753
rect 39736 39515 39865 39556
rect 39736 39463 39775 39515
rect 39827 39463 39865 39515
rect 39736 39132 39865 39463
rect 39736 39076 39773 39132
rect 39829 39076 39865 39132
rect 39736 39037 39865 39076
rect 39956 39363 40084 39402
rect 39956 39307 39992 39363
rect 40048 39341 40084 39363
rect 40048 39307 40085 39341
rect 39956 39300 40085 39307
rect 39956 39248 39994 39300
rect 40046 39248 40085 39300
rect 39956 39114 40085 39248
rect 39956 39062 39994 39114
rect 40046 39062 40085 39114
rect 39956 39021 40085 39062
rect 40215 38855 40524 39701
rect 40215 38799 40251 38855
rect 40307 38799 40431 38855
rect 40487 38799 40524 38855
rect 39736 38578 39865 38617
rect 39736 38522 39773 38578
rect 39829 38522 39865 38578
rect 39736 38191 39865 38522
rect 39956 38592 40085 38633
rect 39956 38540 39994 38592
rect 40046 38540 40085 38592
rect 39956 38406 40085 38540
rect 39956 38354 39994 38406
rect 40046 38354 40085 38406
rect 39956 38347 40085 38354
rect 39956 38291 39992 38347
rect 40048 38313 40085 38347
rect 40048 38291 40084 38313
rect 39956 38252 40084 38291
rect 39736 38139 39775 38191
rect 39827 38139 39865 38191
rect 39736 38098 39865 38139
rect 38967 37899 39050 37955
rect 39106 37899 39230 37955
rect 39286 37899 39619 37955
rect 38967 36155 39619 37899
rect 40215 37953 40524 38799
rect 40215 37901 40253 37953
rect 40305 37901 40433 37953
rect 40485 37901 40524 37953
rect 39736 37715 39865 37756
rect 39736 37663 39775 37715
rect 39827 37663 39865 37715
rect 39736 37332 39865 37663
rect 39736 37276 39773 37332
rect 39829 37276 39865 37332
rect 39736 37237 39865 37276
rect 39956 37563 40084 37602
rect 39956 37507 39992 37563
rect 40048 37541 40084 37563
rect 40048 37507 40085 37541
rect 39956 37500 40085 37507
rect 39956 37448 39994 37500
rect 40046 37448 40085 37500
rect 39956 37314 40085 37448
rect 39956 37262 39994 37314
rect 40046 37262 40085 37314
rect 39956 37221 40085 37262
rect 40215 37055 40524 37901
rect 40215 36999 40251 37055
rect 40307 36999 40431 37055
rect 40487 36999 40524 37055
rect 39736 36778 39865 36817
rect 39736 36722 39773 36778
rect 39829 36722 39865 36778
rect 39736 36391 39865 36722
rect 39956 36792 40085 36833
rect 39956 36740 39994 36792
rect 40046 36740 40085 36792
rect 39956 36606 40085 36740
rect 39956 36554 39994 36606
rect 40046 36554 40085 36606
rect 39956 36547 40085 36554
rect 39956 36491 39992 36547
rect 40048 36513 40085 36547
rect 40048 36491 40084 36513
rect 39956 36452 40084 36491
rect 39736 36339 39775 36391
rect 39827 36339 39865 36391
rect 39736 36298 39865 36339
rect 38967 36099 39050 36155
rect 39106 36099 39230 36155
rect 39286 36099 39619 36155
rect 38967 35976 39619 36099
rect 40215 36153 40524 36999
rect 40215 36101 40253 36153
rect 40305 36101 40433 36153
rect 40485 36101 40524 36153
rect 40215 35976 40524 36101
rect 40718 35976 40939 43226
rect 41095 35976 41317 43226
rect 41473 43250 43583 43491
rect 43703 43353 44564 44253
rect 48789 44233 49990 44776
rect 48789 44181 48828 44233
rect 48880 44181 49039 44233
rect 49091 44181 49250 44233
rect 49302 44181 49461 44233
rect 49513 44181 49990 44233
rect 48789 43770 49990 44181
rect 48789 43718 48828 43770
rect 48880 43718 49039 43770
rect 49091 43718 49250 43770
rect 49302 43718 49461 43770
rect 49513 43718 49990 43770
rect 43703 43340 43790 43353
rect 41473 36096 41695 43250
rect 41851 43115 42072 43250
rect 41851 43063 41935 43115
rect 41987 43063 42072 43115
rect 41851 41791 42072 43063
rect 41851 41739 41935 41791
rect 41987 41739 42072 41791
rect 41851 41315 42072 41739
rect 41851 41263 41935 41315
rect 41987 41263 42072 41315
rect 41851 39991 42072 41263
rect 41851 39939 41935 39991
rect 41987 39939 42072 39991
rect 41851 39515 42072 39939
rect 41851 39463 41935 39515
rect 41987 39463 42072 39515
rect 41851 38191 42072 39463
rect 41851 38139 41935 38191
rect 41987 38139 42072 38191
rect 41851 37715 42072 38139
rect 41851 37663 41935 37715
rect 41987 37663 42072 37715
rect 41851 36391 42072 37663
rect 41851 36339 41935 36391
rect 41987 36339 42072 36391
rect 41851 36096 42072 36339
rect 42229 36096 42450 43250
rect 36863 35881 37743 35976
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 36863 35786 37743 35825
rect 41472 35963 41695 36096
rect 41472 35809 41694 35963
rect 38596 35532 41102 35761
rect 41359 35532 41694 35809
rect 38596 35516 38817 35532
rect 27387 34884 27447 34940
rect 27503 34884 27571 34940
rect 27627 34884 27695 34940
rect 27751 34884 27828 34940
rect 27387 34816 27828 34884
rect 27387 34760 27447 34816
rect 27503 34760 27571 34816
rect 27627 34760 27695 34816
rect 27751 34760 27828 34816
rect 27387 34692 27828 34760
rect 27387 34636 27447 34692
rect 27503 34636 27571 34692
rect 27627 34636 27695 34692
rect 27751 34636 27828 34692
rect 27387 34568 27828 34636
rect 27387 34512 27447 34568
rect 27503 34512 27571 34568
rect 27627 34512 27695 34568
rect 27751 34512 27828 34568
rect 27387 33432 27828 34512
rect 27387 33380 27476 33432
rect 27528 33380 27688 33432
rect 27740 33380 27828 33432
rect 27387 33215 27828 33380
rect 31615 35287 38817 35516
rect 41850 35425 42072 36096
rect 31615 33349 31836 35287
rect 39077 35197 41102 35425
rect 41482 35197 42072 35425
rect 42228 35963 42450 36096
rect 42606 36085 42828 43250
rect 42984 36096 43205 43250
rect 42603 35963 42828 36085
rect 39077 35171 39298 35197
rect 31970 34943 39298 35171
rect 42228 35090 42449 35963
rect 31970 33349 32192 34943
rect 39755 34861 41102 35090
rect 41482 34861 42449 35090
rect 39755 34675 39977 34861
rect 42603 34754 42825 35963
rect 38301 34491 39977 34675
rect 37201 34446 39977 34491
rect 40106 34526 41102 34754
rect 41482 34526 42825 34754
rect 37201 34263 38523 34446
rect 40106 34312 40328 34526
rect 42983 34419 43205 36096
rect 43362 42884 43583 43250
rect 43362 42832 43445 42884
rect 43497 42832 43583 42884
rect 43362 42022 43583 42832
rect 43362 41970 43445 42022
rect 43497 41970 43583 42022
rect 43362 41084 43583 41970
rect 43362 41032 43445 41084
rect 43497 41032 43583 41084
rect 43362 40222 43583 41032
rect 43362 40170 43445 40222
rect 43497 40170 43583 40222
rect 43362 39284 43583 40170
rect 43362 39232 43445 39284
rect 43497 39232 43583 39284
rect 43362 38422 43583 39232
rect 43362 38370 43445 38422
rect 43497 38370 43583 38422
rect 43362 37484 43583 38370
rect 43362 37432 43445 37484
rect 43497 37432 43583 37484
rect 43362 36622 43583 37432
rect 43362 36570 43445 36622
rect 43497 36570 43583 36622
rect 43362 36085 43583 36570
rect 37201 33360 37423 34263
rect 38642 34156 40328 34312
rect 37557 34084 40328 34156
rect 40458 34190 41102 34419
rect 41482 34190 43205 34419
rect 43359 35963 43583 36085
rect 43704 43301 43790 43340
rect 43842 43301 44001 43353
rect 44053 43301 44213 43353
rect 44265 43301 44424 43353
rect 44476 43340 44564 43353
rect 44758 43355 45384 43478
rect 44476 43301 44563 43340
rect 43704 42455 44563 43301
rect 43704 42399 43788 42455
rect 43844 42399 43999 42455
rect 44055 42399 44211 42455
rect 44267 42399 44422 42455
rect 44478 42399 44563 42455
rect 43704 41553 44563 42399
rect 43704 41501 43790 41553
rect 43842 41501 44001 41553
rect 44053 41501 44213 41553
rect 44265 41501 44424 41553
rect 44476 41501 44563 41553
rect 43704 40655 44563 41501
rect 43704 40599 43788 40655
rect 43844 40599 43999 40655
rect 44055 40599 44211 40655
rect 44267 40599 44422 40655
rect 44478 40599 44563 40655
rect 43704 39753 44563 40599
rect 43704 39701 43790 39753
rect 43842 39701 44001 39753
rect 44053 39701 44213 39753
rect 44265 39701 44424 39753
rect 44476 39701 44563 39753
rect 43704 38855 44563 39701
rect 43704 38799 43788 38855
rect 43844 38799 43999 38855
rect 44055 38799 44211 38855
rect 44267 38799 44422 38855
rect 44478 38799 44563 38855
rect 43704 37953 44563 38799
rect 43704 37901 43790 37953
rect 43842 37901 44001 37953
rect 44053 37901 44213 37953
rect 44265 37901 44424 37953
rect 44476 37901 44563 37953
rect 43704 37055 44563 37901
rect 43704 36999 43788 37055
rect 43844 36999 43999 37055
rect 44055 36999 44211 37055
rect 44267 36999 44422 37055
rect 44478 36999 44563 37055
rect 43704 36153 44563 36999
rect 43704 36101 43790 36153
rect 43842 36101 44001 36153
rect 44053 36101 44213 36153
rect 44265 36101 44424 36153
rect 44476 36101 44563 36153
rect 43704 35976 44563 36101
rect 44758 43299 44832 43355
rect 44888 43299 45043 43355
rect 45099 43299 45254 43355
rect 45310 43299 45384 43355
rect 44758 42891 45384 43299
rect 44758 42839 44939 42891
rect 44991 42839 45151 42891
rect 45203 42839 45384 42891
rect 44758 42015 45384 42839
rect 44758 41963 44939 42015
rect 44991 41963 45151 42015
rect 45203 41963 45384 42015
rect 44758 41555 45384 41963
rect 44758 41499 44832 41555
rect 44888 41499 45043 41555
rect 45099 41499 45254 41555
rect 45310 41499 45384 41555
rect 44758 41091 45384 41499
rect 44758 41039 44939 41091
rect 44991 41039 45151 41091
rect 45203 41039 45384 41091
rect 44758 40215 45384 41039
rect 44758 40163 44939 40215
rect 44991 40163 45151 40215
rect 45203 40163 45384 40215
rect 44758 39755 45384 40163
rect 44758 39699 44832 39755
rect 44888 39699 45043 39755
rect 45099 39699 45254 39755
rect 45310 39699 45384 39755
rect 44758 39291 45384 39699
rect 44758 39239 44939 39291
rect 44991 39239 45151 39291
rect 45203 39239 45384 39291
rect 44758 38415 45384 39239
rect 44758 38363 44939 38415
rect 44991 38363 45151 38415
rect 45203 38363 45384 38415
rect 44758 37955 45384 38363
rect 44758 37899 44832 37955
rect 44888 37899 45043 37955
rect 45099 37899 45254 37955
rect 45310 37899 45384 37955
rect 44758 37491 45384 37899
rect 44758 37439 44939 37491
rect 44991 37439 45151 37491
rect 45203 37439 45384 37491
rect 44758 36615 45384 37439
rect 44758 36563 44939 36615
rect 44991 36563 45151 36615
rect 45203 36563 45384 36615
rect 44758 36155 45384 36563
rect 44758 36099 44832 36155
rect 44888 36099 45043 36155
rect 45099 36099 45254 36155
rect 45310 36099 45384 36155
rect 44758 35976 45384 36099
rect 45514 42775 45735 43491
rect 45514 42723 45597 42775
rect 45649 42723 45735 42775
rect 45514 36096 45735 42723
rect 37557 33927 38863 34084
rect 40458 33977 40679 34190
rect 43359 34083 43580 35963
rect 45513 35842 45735 36096
rect 37557 33349 37778 33927
rect 38993 33748 40679 33977
rect 40809 33855 41102 34083
rect 41482 33855 43580 34083
rect 44646 35614 45735 35842
rect 45891 42131 46113 43491
rect 45891 42079 45975 42131
rect 46027 42079 46113 42131
rect 45891 35963 46113 42079
rect 46269 40975 46491 43491
rect 46269 40923 46353 40975
rect 46405 40923 46491 40975
rect 46269 36096 46491 40923
rect 46268 35963 46491 36096
rect 46647 40331 46868 43491
rect 46647 40279 46731 40331
rect 46783 40279 46868 40331
rect 46647 36085 46868 40279
rect 38993 33360 39215 33748
rect 40809 33625 41031 33855
rect 39349 33397 41031 33625
rect 44646 33576 44867 35614
rect 45891 35507 46112 35963
rect 44997 35278 46112 35507
rect 46268 35681 46490 35963
rect 46268 35453 46501 35681
rect 44997 33576 45219 35278
rect 46279 33576 46501 35453
rect 46646 35346 46868 36085
rect 47025 39175 47246 43491
rect 47025 39123 47108 39175
rect 47160 39123 47246 39175
rect 47025 36085 47246 39123
rect 47402 38531 47624 43491
rect 47402 38479 47486 38531
rect 47538 38479 47624 38531
rect 47025 35963 47248 36085
rect 46631 35117 46868 35346
rect 46631 33564 46852 35117
rect 47026 34836 47248 35963
rect 47402 35963 47624 38479
rect 47780 37375 48002 43491
rect 47780 37323 47864 37375
rect 47916 37323 48002 37375
rect 47780 36096 48002 37323
rect 48158 36731 48379 43491
rect 48789 43478 49990 43718
rect 50098 44255 50913 44346
rect 50098 44199 50135 44255
rect 50191 44199 50346 44255
rect 50402 44199 50557 44255
rect 50613 44199 50768 44255
rect 50824 44199 50913 44255
rect 50098 44035 50913 44199
rect 50098 43983 50137 44035
rect 50189 43983 50348 44035
rect 50400 43983 50559 44035
rect 50611 43983 50770 44035
rect 50822 43983 50913 44035
rect 48789 43355 49991 43478
rect 48789 43340 48836 43355
rect 48790 43299 48836 43340
rect 48892 43299 49046 43355
rect 49102 43299 49257 43355
rect 49313 43299 49469 43355
rect 49525 43299 49680 43355
rect 49736 43299 49890 43355
rect 49946 43299 49991 43355
rect 50098 43353 50913 43983
rect 52226 44253 54354 44776
rect 52226 44201 52576 44253
rect 52628 44201 52787 44253
rect 52839 44201 52998 44253
rect 53050 44201 53209 44253
rect 53261 44201 53419 44253
rect 53471 44201 53630 44253
rect 53682 44201 53841 44253
rect 53893 44201 54052 44253
rect 54104 44201 54263 44253
rect 54315 44201 54354 44253
rect 52226 44035 54354 44201
rect 52226 43983 52576 44035
rect 52628 43983 52787 44035
rect 52839 43983 52998 44035
rect 53050 43983 53209 44035
rect 53261 43983 53419 44035
rect 53471 43983 53630 44035
rect 53682 43983 53841 44035
rect 53893 43983 54052 44035
rect 54104 43983 54263 44035
rect 54315 43983 54354 44035
rect 52226 43818 54354 43983
rect 51042 43772 52015 43811
rect 51042 43716 51079 43772
rect 51135 43716 51290 43772
rect 51346 43716 51501 43772
rect 51557 43716 51712 43772
rect 51768 43716 51923 43772
rect 51979 43716 52015 43772
rect 51042 43678 52015 43716
rect 52226 43766 52576 43818
rect 52628 43766 52787 43818
rect 52839 43766 52998 43818
rect 53050 43766 53209 43818
rect 53261 43766 53419 43818
rect 53471 43766 53630 43818
rect 53682 43766 53841 43818
rect 53893 43766 54052 43818
rect 54104 43766 54263 43818
rect 54315 43766 54354 43818
rect 50098 43340 50346 43353
rect 48790 43054 49991 43299
rect 48790 43002 48943 43054
rect 48995 43002 49154 43054
rect 49206 43002 49365 43054
rect 49417 43002 49576 43054
rect 49628 43002 49787 43054
rect 49839 43002 49991 43054
rect 48557 42949 48687 42988
rect 48557 42893 48594 42949
rect 48650 42893 48687 42949
rect 48557 42731 48687 42893
rect 48557 42675 48594 42731
rect 48650 42675 48687 42731
rect 48557 42637 48687 42675
rect 48790 42591 49991 43002
rect 48790 42539 48943 42591
rect 48995 42539 49154 42591
rect 49206 42539 49365 42591
rect 49417 42539 49576 42591
rect 49628 42539 49787 42591
rect 49839 42539 49991 42591
rect 48790 42315 49991 42539
rect 48790 42263 48943 42315
rect 48995 42263 49154 42315
rect 49206 42263 49365 42315
rect 49417 42263 49576 42315
rect 49628 42263 49787 42315
rect 49839 42263 49991 42315
rect 48557 42179 48687 42217
rect 48557 42123 48594 42179
rect 48650 42123 48687 42179
rect 48557 41961 48687 42123
rect 48557 41905 48594 41961
rect 48650 41905 48687 41961
rect 48557 41866 48687 41905
rect 48790 41852 49991 42263
rect 48790 41800 48943 41852
rect 48995 41800 49154 41852
rect 49206 41800 49365 41852
rect 49417 41800 49576 41852
rect 49628 41800 49787 41852
rect 49839 41800 49991 41852
rect 48790 41555 49991 41800
rect 48790 41499 48836 41555
rect 48892 41499 49046 41555
rect 49102 41499 49257 41555
rect 49313 41499 49469 41555
rect 49525 41499 49680 41555
rect 49736 41499 49890 41555
rect 49946 41499 49991 41555
rect 48790 41254 49991 41499
rect 48790 41202 48943 41254
rect 48995 41202 49154 41254
rect 49206 41202 49365 41254
rect 49417 41202 49576 41254
rect 49628 41202 49787 41254
rect 49839 41202 49991 41254
rect 48557 41149 48687 41188
rect 48557 41093 48594 41149
rect 48650 41093 48687 41149
rect 48557 40931 48687 41093
rect 48557 40875 48594 40931
rect 48650 40875 48687 40931
rect 48557 40837 48687 40875
rect 48790 40791 49991 41202
rect 48790 40739 48943 40791
rect 48995 40739 49154 40791
rect 49206 40739 49365 40791
rect 49417 40739 49576 40791
rect 49628 40739 49787 40791
rect 49839 40739 49991 40791
rect 48790 40515 49991 40739
rect 48790 40463 48943 40515
rect 48995 40463 49154 40515
rect 49206 40463 49365 40515
rect 49417 40463 49576 40515
rect 49628 40463 49787 40515
rect 49839 40463 49991 40515
rect 48557 40379 48687 40417
rect 48557 40323 48594 40379
rect 48650 40323 48687 40379
rect 48557 40161 48687 40323
rect 48557 40105 48594 40161
rect 48650 40105 48687 40161
rect 48557 40066 48687 40105
rect 48790 40052 49991 40463
rect 48790 40000 48943 40052
rect 48995 40000 49154 40052
rect 49206 40000 49365 40052
rect 49417 40000 49576 40052
rect 49628 40000 49787 40052
rect 49839 40000 49991 40052
rect 48790 39755 49991 40000
rect 48790 39699 48836 39755
rect 48892 39699 49046 39755
rect 49102 39699 49257 39755
rect 49313 39699 49469 39755
rect 49525 39699 49680 39755
rect 49736 39699 49890 39755
rect 49946 39699 49991 39755
rect 48790 39454 49991 39699
rect 48790 39402 48943 39454
rect 48995 39402 49154 39454
rect 49206 39402 49365 39454
rect 49417 39402 49576 39454
rect 49628 39402 49787 39454
rect 49839 39402 49991 39454
rect 48557 39349 48687 39388
rect 48557 39293 48594 39349
rect 48650 39293 48687 39349
rect 48557 39131 48687 39293
rect 48557 39075 48594 39131
rect 48650 39075 48687 39131
rect 48557 39037 48687 39075
rect 48790 38991 49991 39402
rect 48790 38939 48943 38991
rect 48995 38939 49154 38991
rect 49206 38939 49365 38991
rect 49417 38939 49576 38991
rect 49628 38939 49787 38991
rect 49839 38939 49991 38991
rect 48790 38715 49991 38939
rect 48790 38663 48943 38715
rect 48995 38663 49154 38715
rect 49206 38663 49365 38715
rect 49417 38663 49576 38715
rect 49628 38663 49787 38715
rect 49839 38663 49991 38715
rect 48557 38579 48687 38617
rect 48557 38523 48594 38579
rect 48650 38523 48687 38579
rect 48557 38361 48687 38523
rect 48557 38305 48594 38361
rect 48650 38305 48687 38361
rect 48557 38266 48687 38305
rect 48790 38252 49991 38663
rect 48790 38200 48943 38252
rect 48995 38200 49154 38252
rect 49206 38200 49365 38252
rect 49417 38200 49576 38252
rect 49628 38200 49787 38252
rect 49839 38200 49991 38252
rect 48790 37955 49991 38200
rect 48790 37899 48836 37955
rect 48892 37899 49046 37955
rect 49102 37899 49257 37955
rect 49313 37899 49469 37955
rect 49525 37899 49680 37955
rect 49736 37899 49890 37955
rect 49946 37899 49991 37955
rect 48790 37654 49991 37899
rect 48790 37602 48943 37654
rect 48995 37602 49154 37654
rect 49206 37602 49365 37654
rect 49417 37602 49576 37654
rect 49628 37602 49787 37654
rect 49839 37602 49991 37654
rect 48557 37549 48687 37588
rect 48557 37493 48594 37549
rect 48650 37493 48687 37549
rect 48557 37331 48687 37493
rect 48557 37275 48594 37331
rect 48650 37275 48687 37331
rect 48557 37237 48687 37275
rect 48790 37191 49991 37602
rect 48790 37139 48943 37191
rect 48995 37139 49154 37191
rect 49206 37139 49365 37191
rect 49417 37139 49576 37191
rect 49628 37139 49787 37191
rect 49839 37139 49991 37191
rect 48790 36915 49991 37139
rect 48790 36863 48943 36915
rect 48995 36863 49154 36915
rect 49206 36863 49365 36915
rect 49417 36863 49576 36915
rect 49628 36863 49787 36915
rect 49839 36863 49991 36915
rect 48158 36679 48241 36731
rect 48293 36679 48379 36731
rect 48158 36096 48379 36679
rect 48557 36779 48687 36817
rect 48557 36723 48594 36779
rect 48650 36723 48687 36779
rect 48557 36561 48687 36723
rect 48557 36505 48594 36561
rect 48650 36505 48687 36561
rect 48557 36466 48687 36505
rect 47779 35963 48002 36096
rect 47402 35171 47623 35963
rect 47779 35507 48001 35963
rect 48157 35842 48379 36096
rect 48790 36452 49991 36863
rect 48790 36400 48943 36452
rect 48995 36400 49154 36452
rect 49206 36400 49365 36452
rect 49417 36400 49576 36452
rect 49628 36400 49787 36452
rect 49839 36400 49991 36452
rect 48790 36155 49991 36400
rect 48790 36099 48836 36155
rect 48892 36099 49046 36155
rect 49102 36099 49257 36155
rect 49313 36099 49469 36155
rect 49525 36099 49680 36155
rect 49736 36099 49890 36155
rect 49946 36099 49991 36155
rect 48790 35976 49991 36099
rect 50099 43301 50346 43340
rect 50398 43301 50557 43353
rect 50609 43301 50768 43353
rect 50820 43301 50913 43353
rect 52226 43478 54354 43766
rect 54758 44253 55638 44776
rect 54758 44201 54855 44253
rect 54907 44201 55066 44253
rect 55118 44201 55278 44253
rect 55330 44201 55489 44253
rect 55541 44201 55638 44253
rect 52226 43355 54355 43478
rect 52226 43340 52314 43355
rect 50099 42891 50913 43301
rect 52227 43299 52314 43340
rect 52370 43299 52525 43355
rect 52581 43299 52736 43355
rect 52792 43299 52946 43355
rect 53002 43299 53157 43355
rect 53213 43299 53369 43355
rect 53425 43299 53580 43355
rect 53636 43299 53790 43355
rect 53846 43299 54001 43355
rect 54057 43299 54212 43355
rect 54268 43299 54355 43355
rect 50099 42839 50300 42891
rect 50352 42839 50511 42891
rect 50563 42839 50722 42891
rect 50774 42839 50913 42891
rect 50099 42455 50913 42839
rect 51034 43129 51344 43170
rect 51034 43077 51073 43129
rect 51125 43077 51253 43129
rect 51305 43077 51344 43129
rect 51034 42915 51344 43077
rect 51034 42859 51071 42915
rect 51127 42859 51251 42915
rect 51307 42859 51344 42915
rect 51034 42786 51344 42859
rect 51796 43122 52106 43163
rect 51796 43070 51835 43122
rect 51887 43070 52015 43122
rect 52067 43070 52106 43122
rect 51796 42915 52106 43070
rect 51796 42859 51833 42915
rect 51889 42859 52013 42915
rect 52069 42859 52106 42915
rect 51796 42659 52106 42859
rect 51796 42607 51835 42659
rect 51887 42607 52015 42659
rect 52067 42607 52106 42659
rect 51796 42567 52106 42607
rect 50099 42453 50161 42455
rect 50217 42453 50372 42455
rect 50099 42401 50138 42453
rect 50217 42401 50318 42453
rect 50370 42401 50372 42453
rect 50099 42399 50161 42401
rect 50217 42399 50372 42401
rect 50428 42399 50584 42455
rect 50640 42399 50795 42455
rect 50851 42399 50913 42455
rect 50099 42015 50913 42399
rect 52227 42453 54355 43299
rect 52227 42401 52316 42453
rect 52368 42401 52527 42453
rect 52579 42401 52738 42453
rect 52790 42401 52948 42453
rect 53000 42401 53159 42453
rect 53211 42401 53371 42453
rect 53423 42401 53582 42453
rect 53634 42401 53792 42453
rect 53844 42401 54003 42453
rect 54055 42401 54214 42453
rect 54266 42401 54355 42453
rect 51796 42247 52106 42287
rect 51796 42195 51835 42247
rect 51887 42195 52015 42247
rect 52067 42195 52106 42247
rect 50099 41963 50300 42015
rect 50352 41963 50511 42015
rect 50563 41963 50722 42015
rect 50774 41963 50913 42015
rect 50099 41553 50913 41963
rect 51034 41995 51344 42068
rect 51034 41939 51071 41995
rect 51127 41939 51251 41995
rect 51307 41939 51344 41995
rect 51034 41777 51344 41939
rect 51034 41725 51073 41777
rect 51125 41725 51253 41777
rect 51305 41725 51344 41777
rect 51034 41684 51344 41725
rect 51796 41995 52106 42195
rect 51796 41939 51833 41995
rect 51889 41939 52013 41995
rect 52069 41939 52106 41995
rect 51796 41784 52106 41939
rect 51796 41732 51835 41784
rect 51887 41732 52015 41784
rect 52067 41732 52106 41784
rect 51796 41691 52106 41732
rect 50099 41501 50346 41553
rect 50398 41501 50557 41553
rect 50609 41501 50768 41553
rect 50820 41501 50913 41553
rect 50099 41091 50913 41501
rect 52227 41555 54355 42401
rect 52227 41499 52314 41555
rect 52370 41499 52525 41555
rect 52581 41499 52736 41555
rect 52792 41499 52946 41555
rect 53002 41499 53157 41555
rect 53213 41499 53369 41555
rect 53425 41499 53580 41555
rect 53636 41499 53790 41555
rect 53846 41499 54001 41555
rect 54057 41499 54212 41555
rect 54268 41499 54355 41555
rect 50099 41039 50300 41091
rect 50352 41039 50511 41091
rect 50563 41039 50722 41091
rect 50774 41039 50913 41091
rect 50099 40655 50913 41039
rect 51034 41329 51344 41370
rect 51034 41277 51073 41329
rect 51125 41277 51253 41329
rect 51305 41277 51344 41329
rect 51034 41115 51344 41277
rect 51034 41059 51071 41115
rect 51127 41059 51251 41115
rect 51307 41059 51344 41115
rect 51034 40986 51344 41059
rect 51796 41322 52106 41363
rect 51796 41270 51835 41322
rect 51887 41270 52015 41322
rect 52067 41270 52106 41322
rect 51796 41115 52106 41270
rect 51796 41059 51833 41115
rect 51889 41059 52013 41115
rect 52069 41059 52106 41115
rect 51796 40859 52106 41059
rect 51796 40807 51835 40859
rect 51887 40807 52015 40859
rect 52067 40807 52106 40859
rect 51796 40767 52106 40807
rect 50099 40653 50161 40655
rect 50217 40653 50372 40655
rect 50099 40601 50138 40653
rect 50217 40601 50318 40653
rect 50370 40601 50372 40653
rect 50099 40599 50161 40601
rect 50217 40599 50372 40601
rect 50428 40599 50584 40655
rect 50640 40599 50795 40655
rect 50851 40599 50913 40655
rect 50099 40215 50913 40599
rect 52227 40653 54355 41499
rect 52227 40601 52316 40653
rect 52368 40601 52527 40653
rect 52579 40601 52738 40653
rect 52790 40601 52948 40653
rect 53000 40601 53159 40653
rect 53211 40601 53371 40653
rect 53423 40601 53582 40653
rect 53634 40601 53792 40653
rect 53844 40601 54003 40653
rect 54055 40601 54214 40653
rect 54266 40601 54355 40653
rect 51796 40447 52106 40487
rect 51796 40395 51835 40447
rect 51887 40395 52015 40447
rect 52067 40395 52106 40447
rect 50099 40163 50300 40215
rect 50352 40163 50511 40215
rect 50563 40163 50722 40215
rect 50774 40163 50913 40215
rect 50099 39753 50913 40163
rect 51034 40195 51344 40268
rect 51034 40139 51071 40195
rect 51127 40139 51251 40195
rect 51307 40139 51344 40195
rect 51034 39977 51344 40139
rect 51034 39925 51073 39977
rect 51125 39925 51253 39977
rect 51305 39925 51344 39977
rect 51034 39884 51344 39925
rect 51796 40195 52106 40395
rect 51796 40139 51833 40195
rect 51889 40139 52013 40195
rect 52069 40139 52106 40195
rect 51796 39984 52106 40139
rect 51796 39932 51835 39984
rect 51887 39932 52015 39984
rect 52067 39932 52106 39984
rect 51796 39891 52106 39932
rect 50099 39701 50346 39753
rect 50398 39701 50557 39753
rect 50609 39701 50768 39753
rect 50820 39701 50913 39753
rect 50099 39291 50913 39701
rect 52227 39755 54355 40601
rect 52227 39699 52314 39755
rect 52370 39699 52525 39755
rect 52581 39699 52736 39755
rect 52792 39699 52946 39755
rect 53002 39699 53157 39755
rect 53213 39699 53369 39755
rect 53425 39699 53580 39755
rect 53636 39699 53790 39755
rect 53846 39699 54001 39755
rect 54057 39699 54212 39755
rect 54268 39699 54355 39755
rect 50099 39239 50300 39291
rect 50352 39239 50511 39291
rect 50563 39239 50722 39291
rect 50774 39239 50913 39291
rect 50099 38855 50913 39239
rect 51034 39529 51344 39570
rect 51034 39477 51073 39529
rect 51125 39477 51253 39529
rect 51305 39477 51344 39529
rect 51034 39315 51344 39477
rect 51034 39259 51071 39315
rect 51127 39259 51251 39315
rect 51307 39259 51344 39315
rect 51034 39186 51344 39259
rect 51796 39522 52106 39563
rect 51796 39470 51835 39522
rect 51887 39470 52015 39522
rect 52067 39470 52106 39522
rect 51796 39315 52106 39470
rect 51796 39259 51833 39315
rect 51889 39259 52013 39315
rect 52069 39259 52106 39315
rect 51796 39059 52106 39259
rect 51796 39007 51835 39059
rect 51887 39007 52015 39059
rect 52067 39007 52106 39059
rect 51796 38967 52106 39007
rect 50099 38853 50161 38855
rect 50217 38853 50372 38855
rect 50099 38801 50138 38853
rect 50217 38801 50318 38853
rect 50370 38801 50372 38853
rect 50099 38799 50161 38801
rect 50217 38799 50372 38801
rect 50428 38799 50584 38855
rect 50640 38799 50795 38855
rect 50851 38799 50913 38855
rect 50099 38415 50913 38799
rect 52227 38853 54355 39699
rect 52227 38801 52316 38853
rect 52368 38801 52527 38853
rect 52579 38801 52738 38853
rect 52790 38801 52948 38853
rect 53000 38801 53159 38853
rect 53211 38801 53371 38853
rect 53423 38801 53582 38853
rect 53634 38801 53792 38853
rect 53844 38801 54003 38853
rect 54055 38801 54214 38853
rect 54266 38801 54355 38853
rect 51796 38647 52106 38687
rect 51796 38595 51835 38647
rect 51887 38595 52015 38647
rect 52067 38595 52106 38647
rect 50099 38363 50300 38415
rect 50352 38363 50511 38415
rect 50563 38363 50722 38415
rect 50774 38363 50913 38415
rect 50099 37953 50913 38363
rect 51034 38395 51344 38468
rect 51034 38339 51071 38395
rect 51127 38339 51251 38395
rect 51307 38339 51344 38395
rect 51034 38177 51344 38339
rect 51034 38125 51073 38177
rect 51125 38125 51253 38177
rect 51305 38125 51344 38177
rect 51034 38084 51344 38125
rect 51796 38395 52106 38595
rect 51796 38339 51833 38395
rect 51889 38339 52013 38395
rect 52069 38339 52106 38395
rect 51796 38184 52106 38339
rect 51796 38132 51835 38184
rect 51887 38132 52015 38184
rect 52067 38132 52106 38184
rect 51796 38091 52106 38132
rect 50099 37901 50346 37953
rect 50398 37901 50557 37953
rect 50609 37901 50768 37953
rect 50820 37901 50913 37953
rect 50099 37491 50913 37901
rect 52227 37955 54355 38801
rect 52227 37899 52314 37955
rect 52370 37899 52525 37955
rect 52581 37899 52736 37955
rect 52792 37899 52946 37955
rect 53002 37899 53157 37955
rect 53213 37899 53369 37955
rect 53425 37899 53580 37955
rect 53636 37899 53790 37955
rect 53846 37899 54001 37955
rect 54057 37899 54212 37955
rect 54268 37899 54355 37955
rect 50099 37439 50300 37491
rect 50352 37439 50511 37491
rect 50563 37439 50722 37491
rect 50774 37439 50913 37491
rect 50099 37055 50913 37439
rect 51034 37729 51344 37770
rect 51034 37677 51073 37729
rect 51125 37677 51253 37729
rect 51305 37677 51344 37729
rect 51034 37515 51344 37677
rect 51034 37459 51071 37515
rect 51127 37459 51251 37515
rect 51307 37459 51344 37515
rect 51034 37386 51344 37459
rect 51796 37722 52106 37763
rect 51796 37670 51835 37722
rect 51887 37670 52015 37722
rect 52067 37670 52106 37722
rect 51796 37515 52106 37670
rect 51796 37459 51833 37515
rect 51889 37459 52013 37515
rect 52069 37459 52106 37515
rect 51796 37259 52106 37459
rect 51796 37207 51835 37259
rect 51887 37207 52015 37259
rect 52067 37207 52106 37259
rect 51796 37167 52106 37207
rect 50099 37053 50161 37055
rect 50217 37053 50372 37055
rect 50099 37001 50138 37053
rect 50217 37001 50318 37053
rect 50370 37001 50372 37053
rect 50099 36999 50161 37001
rect 50217 36999 50372 37001
rect 50428 36999 50584 37055
rect 50640 36999 50795 37055
rect 50851 36999 50913 37055
rect 50099 36615 50913 36999
rect 52227 37053 54355 37899
rect 52227 37001 52316 37053
rect 52368 37001 52527 37053
rect 52579 37001 52738 37053
rect 52790 37001 52948 37053
rect 53000 37001 53159 37053
rect 53211 37001 53371 37053
rect 53423 37001 53582 37053
rect 53634 37001 53792 37053
rect 53844 37001 54003 37053
rect 54055 37001 54214 37053
rect 54266 37001 54355 37053
rect 51796 36847 52106 36887
rect 51796 36795 51835 36847
rect 51887 36795 52015 36847
rect 52067 36795 52106 36847
rect 50099 36563 50300 36615
rect 50352 36563 50511 36615
rect 50563 36563 50722 36615
rect 50774 36563 50913 36615
rect 50099 36153 50913 36563
rect 51034 36595 51344 36668
rect 51034 36539 51071 36595
rect 51127 36539 51251 36595
rect 51307 36539 51344 36595
rect 51034 36377 51344 36539
rect 51034 36325 51073 36377
rect 51125 36325 51253 36377
rect 51305 36325 51344 36377
rect 51034 36284 51344 36325
rect 51796 36595 52106 36795
rect 51796 36539 51833 36595
rect 51889 36539 52013 36595
rect 52069 36539 52106 36595
rect 51796 36384 52106 36539
rect 51796 36332 51835 36384
rect 51887 36332 52015 36384
rect 52067 36332 52106 36384
rect 51796 36291 52106 36332
rect 50099 36101 50346 36153
rect 50398 36101 50557 36153
rect 50609 36101 50768 36153
rect 50820 36101 50913 36153
rect 50099 35976 50913 36101
rect 52227 36155 54355 37001
rect 52227 36099 52314 36155
rect 52370 36099 52525 36155
rect 52581 36099 52736 36155
rect 52792 36099 52946 36155
rect 53002 36099 53157 36155
rect 53213 36099 53369 36155
rect 53425 36099 53580 36155
rect 53636 36099 53790 36155
rect 53846 36099 54001 36155
rect 54057 36099 54212 36155
rect 54268 36099 54355 36155
rect 52227 35976 54355 36099
rect 54758 43355 55638 44201
rect 55977 44255 57736 44294
rect 55977 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 57736 44255
rect 55977 44160 57736 44199
rect 54758 43299 54853 43355
rect 54909 43299 55064 43355
rect 55120 43299 55276 43355
rect 55332 43299 55487 43355
rect 55543 43299 55638 43355
rect 54758 42453 55638 43299
rect 57295 42494 57736 44160
rect 54758 42401 54855 42453
rect 54907 42401 55066 42453
rect 55118 42401 55278 42453
rect 55330 42401 55489 42453
rect 55541 42401 55638 42453
rect 54758 41555 55638 42401
rect 55977 42455 57736 42494
rect 55977 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 57736 42455
rect 55977 42360 57736 42399
rect 54758 41499 54853 41555
rect 54909 41499 55064 41555
rect 55120 41499 55276 41555
rect 55332 41499 55487 41555
rect 55543 41499 55638 41555
rect 54758 40653 55638 41499
rect 57295 40694 57736 42360
rect 54758 40601 54855 40653
rect 54907 40601 55066 40653
rect 55118 40601 55278 40653
rect 55330 40601 55489 40653
rect 55541 40601 55638 40653
rect 54758 39755 55638 40601
rect 55977 40655 57736 40694
rect 55977 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 57736 40655
rect 55977 40560 57736 40599
rect 54758 39699 54853 39755
rect 54909 39699 55064 39755
rect 55120 39699 55276 39755
rect 55332 39699 55487 39755
rect 55543 39699 55638 39755
rect 54758 38853 55638 39699
rect 57295 38894 57736 40560
rect 54758 38801 54855 38853
rect 54907 38801 55066 38853
rect 55118 38801 55278 38853
rect 55330 38801 55489 38853
rect 55541 38801 55638 38853
rect 54758 37955 55638 38801
rect 55977 38855 57736 38894
rect 55977 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 57736 38855
rect 55977 38760 57736 38799
rect 54758 37899 54853 37955
rect 54909 37899 55064 37955
rect 55120 37899 55276 37955
rect 55332 37899 55487 37955
rect 55543 37899 55638 37955
rect 54758 37053 55638 37899
rect 57295 37094 57736 38760
rect 54758 37001 54855 37053
rect 54907 37001 55066 37053
rect 55118 37001 55278 37053
rect 55330 37001 55489 37053
rect 55541 37001 55638 37053
rect 54758 36155 55638 37001
rect 55977 37055 57736 37094
rect 55977 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 57736 37055
rect 55977 36960 57736 36999
rect 54758 36099 54853 36155
rect 54909 36099 55064 36155
rect 55120 36099 55276 36155
rect 55332 36099 55487 36155
rect 55543 36099 55638 36155
rect 54758 36027 55638 36099
rect 48157 35614 50120 35842
rect 47779 35278 49769 35507
rect 47402 34943 48486 35171
rect 47026 34607 48135 34836
rect 47913 33564 48135 34607
rect 48265 33576 48486 34943
rect 49547 33576 49769 35278
rect 49898 33576 50120 35614
rect 27387 33163 27476 33215
rect 27528 33163 27688 33215
rect 27740 33163 27828 33215
rect 27387 33141 27828 33163
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 27828 33141
rect 27387 32997 27828 33085
rect 27387 32945 27476 32997
rect 27528 32945 27688 32997
rect 27740 32945 27828 32997
rect 27387 32923 27828 32945
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 27828 32923
rect 27387 32779 27828 32867
rect 27387 32727 27476 32779
rect 27528 32727 27688 32779
rect 27740 32727 27828 32779
rect 27387 32705 27828 32727
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 27828 32705
rect 27387 32562 27828 32649
rect 27387 32510 27476 32562
rect 27528 32510 27688 32562
rect 27740 32510 27828 32562
rect 27387 32487 27828 32510
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 27828 32487
rect 27387 32344 27828 32431
rect 27387 32292 27476 32344
rect 27528 32292 27688 32344
rect 27740 32292 27828 32344
rect 27387 32127 27828 32292
rect 27387 32075 27476 32127
rect 27528 32075 27688 32127
rect 27740 32075 27828 32127
rect 27387 31909 27828 32075
rect 27387 31857 27476 31909
rect 27528 31857 27688 31909
rect 27740 31857 27828 31909
rect 27387 31691 27828 31857
rect 27387 31639 27476 31691
rect 27528 31639 27688 31691
rect 27740 31639 27828 31691
rect 27387 31474 27828 31639
rect 27387 31422 27476 31474
rect 27528 31422 27688 31474
rect 27740 31422 27828 31474
rect 27387 31256 27828 31422
rect 27387 31252 27476 31256
rect 27528 31252 27688 31256
rect 27740 31252 27828 31256
rect 27387 31196 27474 31252
rect 27530 31196 27686 31252
rect 27742 31196 27828 31252
rect 27387 31038 27828 31196
rect 27387 31034 27476 31038
rect 27528 31034 27688 31038
rect 27740 31034 27828 31038
rect 27387 30978 27474 31034
rect 27530 30978 27686 31034
rect 27742 30978 27828 31034
rect 27387 30821 27828 30978
rect 27387 30816 27476 30821
rect 27528 30816 27688 30821
rect 27740 30816 27828 30821
rect 27387 30760 27474 30816
rect 27530 30760 27686 30816
rect 27742 30760 27828 30816
rect 27387 30603 27828 30760
rect 27387 30598 27476 30603
rect 27528 30598 27688 30603
rect 27740 30598 27828 30603
rect 27387 30542 27474 30598
rect 27530 30542 27686 30598
rect 27742 30542 27828 30598
rect 27387 30386 27828 30542
rect 27387 30334 27476 30386
rect 27528 30334 27688 30386
rect 27740 30334 27828 30386
rect 27387 30168 27828 30334
rect 27387 30116 27476 30168
rect 27528 30116 27688 30168
rect 27740 30116 27828 30168
rect 27387 29950 27828 30116
rect 27387 29898 27476 29950
rect 27528 29898 27688 29950
rect 27740 29898 27828 29950
rect 27387 29733 27828 29898
rect 27387 29681 27476 29733
rect 27528 29681 27688 29733
rect 27740 29681 27828 29733
rect 27387 29515 27828 29681
rect 27387 29463 27476 29515
rect 27528 29463 27688 29515
rect 27740 29463 27828 29515
rect 27387 29297 27828 29463
rect 27387 29245 27476 29297
rect 27528 29245 27688 29297
rect 27740 29245 27828 29297
rect 27387 29080 27828 29245
rect 27387 29028 27476 29080
rect 27528 29028 27688 29080
rect 27740 29028 27828 29080
rect 27387 28862 27828 29028
rect 27387 28810 27476 28862
rect 27528 28810 27688 28862
rect 27740 28810 27828 28862
rect 27387 28644 27828 28810
rect 27387 28592 27476 28644
rect 27528 28592 27688 28644
rect 27740 28592 27828 28644
rect 27387 28427 27828 28592
rect 27387 28375 27476 28427
rect 27528 28375 27688 28427
rect 27740 28375 27828 28427
rect 27387 28209 27828 28375
rect 27387 28157 27476 28209
rect 27528 28157 27688 28209
rect 27740 28157 27828 28209
rect 27387 27992 27828 28157
rect 27387 27940 27476 27992
rect 27528 27940 27688 27992
rect 27740 27940 27828 27992
rect 27387 27774 27828 27940
rect 27387 27722 27476 27774
rect 27528 27722 27688 27774
rect 27740 27722 27828 27774
rect 27387 27556 27828 27722
rect 27387 27504 27476 27556
rect 27528 27504 27688 27556
rect 27740 27504 27828 27556
rect 27387 27339 27828 27504
rect 27387 27287 27476 27339
rect 27528 27287 27688 27339
rect 27740 27287 27828 27339
rect 27387 27121 27828 27287
rect 27387 27069 27476 27121
rect 27528 27069 27688 27121
rect 27740 27069 27828 27121
rect 27387 26903 27828 27069
rect 27387 26851 27476 26903
rect 27528 26851 27688 26903
rect 27740 26851 27828 26903
rect 27387 26799 27828 26851
rect 27387 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 27387 26686 27828 26743
rect 27387 26634 27476 26686
rect 27528 26634 27688 26686
rect 27740 26634 27828 26686
rect 27387 26581 27828 26634
rect 27387 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 27387 26468 27828 26525
rect 27387 26416 27476 26468
rect 27528 26416 27688 26468
rect 27740 26416 27828 26468
rect 27387 26250 27828 26416
rect 27387 26198 27476 26250
rect 27528 26198 27688 26250
rect 27740 26198 27828 26250
rect 27387 26033 27828 26198
rect 27387 25981 27476 26033
rect 27528 25981 27688 26033
rect 27740 25981 27828 26033
rect 27387 25815 27828 25981
rect 27387 25763 27476 25815
rect 27528 25763 27688 25815
rect 27740 25763 27828 25815
rect 27387 25598 27828 25763
rect 27387 25546 27476 25598
rect 27528 25546 27688 25598
rect 27740 25546 27828 25598
rect 27387 25380 27828 25546
rect 27387 25328 27476 25380
rect 27528 25328 27688 25380
rect 27740 25328 27828 25380
rect 27387 25162 27828 25328
rect 27387 25110 27476 25162
rect 27528 25110 27688 25162
rect 27740 25110 27828 25162
rect 27387 25028 27828 25110
rect 27387 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 27828 25028
rect 27387 24945 27828 24972
rect 27387 24893 27476 24945
rect 27528 24893 27688 24945
rect 27740 24893 27828 24945
rect 27387 24810 27828 24893
rect 27387 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 27828 24810
rect 27387 24727 27828 24754
rect 27387 24675 27476 24727
rect 27528 24675 27688 24727
rect 27740 24675 27828 24727
rect 27387 24509 27828 24675
rect 27387 24457 27476 24509
rect 27528 24457 27688 24509
rect 27740 24457 27828 24509
rect 27387 24292 27828 24457
rect 27387 24240 27476 24292
rect 27528 24240 27688 24292
rect 27740 24240 27828 24292
rect 27387 24074 27828 24240
rect 27387 24022 27476 24074
rect 27528 24022 27688 24074
rect 27740 24022 27828 24074
rect 27387 23857 27828 24022
rect 27387 23805 27476 23857
rect 27528 23805 27688 23857
rect 27740 23805 27828 23857
rect 27387 23639 27828 23805
rect 27387 23587 27476 23639
rect 27528 23587 27688 23639
rect 27740 23587 27828 23639
rect 27387 23421 27828 23587
rect 27387 23369 27476 23421
rect 27528 23369 27688 23421
rect 27740 23369 27828 23421
rect 27387 23204 27828 23369
rect 27387 23152 27476 23204
rect 27528 23152 27688 23204
rect 27740 23152 27828 23204
rect 27387 22986 27828 23152
rect 27387 22936 27476 22986
rect 27528 22936 27688 22986
rect 27387 22048 27475 22936
rect 27740 22934 27828 22986
rect 27739 22768 27828 22934
rect 27740 22716 27828 22768
rect 27739 22551 27828 22716
rect 27740 22499 27828 22551
rect 27739 22333 27828 22499
rect 27740 22281 27828 22333
rect 27739 22115 27828 22281
rect 27740 22063 27828 22115
rect 27739 22048 27828 22063
rect 27387 21898 27828 22048
rect 27387 21846 27476 21898
rect 27528 21846 27688 21898
rect 27740 21846 27828 21898
rect 27387 21680 27828 21846
rect 27387 21628 27476 21680
rect 27528 21628 27688 21680
rect 27740 21628 27828 21680
rect 27387 21463 27828 21628
rect 27387 21411 27476 21463
rect 27528 21411 27688 21463
rect 27740 21411 27828 21463
rect 27387 21245 27828 21411
rect 27387 21193 27476 21245
rect 27528 21193 27688 21245
rect 27740 21193 27828 21245
rect 27387 21027 27828 21193
rect 27387 20975 27476 21027
rect 27528 20975 27688 21027
rect 27740 20975 27828 21027
rect 27387 20810 27828 20975
rect 27387 20758 27476 20810
rect 27528 20758 27688 20810
rect 27740 20758 27828 20810
rect 27387 20592 27828 20758
rect 27387 20540 27476 20592
rect 27528 20540 27688 20592
rect 27740 20540 27828 20592
rect 27387 20374 27828 20540
rect 27387 20322 27476 20374
rect 27528 20322 27688 20374
rect 27740 20322 27828 20374
rect 27387 20157 27828 20322
rect 27387 20105 27476 20157
rect 27528 20105 27688 20157
rect 27740 20105 27828 20157
rect 27387 19939 27828 20105
rect 27387 19887 27476 19939
rect 27528 19887 27688 19939
rect 27740 19887 27828 19939
rect 27387 19722 27828 19887
rect 27387 19670 27476 19722
rect 27528 19670 27688 19722
rect 27740 19670 27828 19722
rect 27387 19504 27828 19670
rect 27387 19452 27476 19504
rect 27528 19452 27688 19504
rect 27740 19452 27828 19504
rect 27387 19286 27828 19452
rect 27387 19234 27476 19286
rect 27528 19234 27688 19286
rect 27740 19234 27828 19286
rect 27387 19068 27828 19234
rect 27387 19016 27476 19068
rect 27528 19016 27688 19068
rect 27740 19016 27828 19068
rect 27387 18851 27828 19016
rect 27387 18799 27476 18851
rect 27528 18799 27688 18851
rect 27740 18799 27828 18851
rect 27387 18633 27828 18799
rect 27387 18581 27476 18633
rect 27528 18581 27688 18633
rect 27740 18581 27828 18633
rect 27387 18416 27828 18581
rect 27387 18364 27476 18416
rect 27528 18364 27688 18416
rect 27740 18364 27828 18416
rect 27387 18198 27828 18364
rect 27387 18146 27476 18198
rect 27528 18146 27688 18198
rect 27740 18146 27828 18198
rect 27387 17980 27828 18146
rect 27387 17928 27476 17980
rect 27528 17928 27688 17980
rect 27740 17928 27828 17980
rect 27387 17763 27828 17928
rect 27387 17711 27476 17763
rect 27528 17711 27688 17763
rect 27740 17711 27828 17763
rect 27387 17545 27828 17711
rect 27387 17493 27476 17545
rect 27528 17493 27688 17545
rect 27740 17493 27828 17545
rect 27387 17327 27828 17493
rect 27387 17275 27476 17327
rect 27528 17275 27688 17327
rect 27740 17275 27828 17327
rect 27387 17110 27828 17275
rect 27387 17058 27476 17110
rect 27528 17058 27688 17110
rect 27740 17058 27828 17110
rect 27387 16892 27828 17058
rect 27387 16840 27476 16892
rect 27528 16840 27688 16892
rect 27740 16840 27828 16892
rect 27387 16675 27828 16840
rect 27387 16623 27476 16675
rect 27528 16623 27688 16675
rect 27740 16623 27828 16675
rect 27387 16470 27828 16623
rect 27387 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 27387 16405 27476 16414
rect 27528 16405 27688 16414
rect 27740 16405 27828 16414
rect 27387 16253 27828 16405
rect 27387 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 27387 16187 27476 16197
rect 27528 16187 27688 16197
rect 27740 16187 27828 16197
rect 27387 16035 27828 16187
rect 27387 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 27387 15970 27476 15979
rect 27528 15970 27688 15979
rect 27740 15970 27828 15979
rect 27387 15818 27828 15970
rect 27387 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 27387 15752 27476 15762
rect 27528 15752 27688 15762
rect 27740 15752 27828 15762
rect 27387 15600 27828 15752
rect 27387 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 27387 15534 27476 15544
rect 27528 15534 27688 15544
rect 27740 15534 27828 15544
rect 27387 15382 27828 15534
rect 27387 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 27387 15317 27476 15326
rect 27528 15317 27688 15326
rect 27740 15317 27828 15326
rect 27387 15164 27828 15317
rect 27387 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 27387 15099 27476 15108
rect 27528 15099 27688 15108
rect 27740 15099 27828 15108
rect 27387 14947 27828 15099
rect 27387 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14891 27828 14947
rect 27387 14881 27476 14891
rect 27528 14881 27688 14891
rect 27740 14881 27828 14891
rect 27387 14729 27828 14881
rect 27387 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 27828 14729
rect 27387 14664 27476 14673
rect 27528 14664 27688 14673
rect 27740 14664 27828 14673
rect 27387 14512 27828 14664
rect 27387 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14456 27828 14512
rect 27387 14446 27476 14456
rect 27528 14446 27688 14456
rect 27740 14446 27828 14456
rect 27387 14281 27828 14446
rect 27387 14231 27476 14281
rect 27528 14231 27688 14281
rect 27740 14231 27828 14281
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 27828 14231
rect 27387 14063 27828 14175
rect 27387 14014 27476 14063
rect 27528 14014 27688 14063
rect 27740 14014 27828 14063
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 27828 14014
rect 27387 13845 27828 13958
rect 27387 13796 27476 13845
rect 27528 13796 27688 13845
rect 27740 13796 27828 13845
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13740 27828 13796
rect 27387 13628 27828 13740
rect 27387 13578 27476 13628
rect 27528 13578 27688 13628
rect 27740 13578 27828 13628
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 27828 13578
rect 27387 13410 27828 13522
rect 27387 13361 27476 13410
rect 27528 13361 27688 13410
rect 27740 13361 27828 13410
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 27828 13361
rect 27387 13192 27828 13305
rect 27387 13140 27476 13192
rect 27528 13140 27688 13192
rect 27740 13140 27828 13192
rect 27387 12975 27828 13140
rect 27387 12923 27476 12975
rect 27528 12923 27688 12975
rect 27740 12923 27828 12975
rect 27387 12757 27828 12923
rect 27387 12705 27476 12757
rect 27528 12705 27688 12757
rect 27740 12705 27828 12757
rect 27387 12540 27828 12705
rect 27387 12488 27476 12540
rect 27528 12488 27688 12540
rect 27740 12488 27828 12540
rect 27387 12322 27828 12488
rect 27387 12270 27476 12322
rect 27528 12270 27688 12322
rect 27740 12270 27828 12322
rect 27387 12104 27828 12270
rect 27387 12052 27476 12104
rect 27528 12052 27688 12104
rect 27740 12052 27828 12104
rect 27387 11887 27828 12052
rect 27387 11835 27476 11887
rect 27528 11835 27688 11887
rect 27740 11835 27828 11887
rect 27387 11669 27828 11835
rect 27387 11617 27476 11669
rect 27528 11617 27688 11669
rect 27740 11617 27828 11669
rect 27387 11451 27828 11617
rect 27387 11406 27476 11451
rect 27528 11406 27688 11451
rect 27740 11406 27828 11451
rect 27387 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 27387 11234 27828 11350
rect 27387 11189 27476 11234
rect 27528 11189 27688 11234
rect 27740 11189 27828 11234
rect 27387 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 27387 11016 27828 11133
rect 27387 10971 27476 11016
rect 27528 10971 27688 11016
rect 27740 10971 27828 11016
rect 27387 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 27387 10798 27828 10915
rect 27387 10753 27476 10798
rect 27528 10753 27688 10798
rect 27740 10753 27828 10798
rect 27387 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 27387 10581 27828 10697
rect 27387 10535 27476 10581
rect 27528 10535 27688 10581
rect 27740 10535 27828 10581
rect 27387 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 27387 10363 27828 10479
rect 27387 10318 27476 10363
rect 27528 10318 27688 10363
rect 27740 10318 27828 10363
rect 27387 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 27387 10146 27828 10262
rect 27387 10094 27476 10146
rect 27528 10094 27688 10146
rect 27740 10094 27828 10146
rect 27387 9928 27828 10094
rect 57295 33141 57736 36960
rect 57295 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 57295 32923 57736 33085
rect 57295 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 57295 32705 57736 32867
rect 57295 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 57295 32487 57736 32649
rect 57295 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 57295 31252 57736 32431
rect 57295 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31196 57736 31252
rect 57295 31034 57736 31196
rect 57295 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30978 57736 31034
rect 57295 30816 57736 30978
rect 57295 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30760 57736 30816
rect 57295 30598 57736 30760
rect 57295 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30542 57736 30598
rect 57295 26799 57736 30542
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 57736 26799
rect 57295 26581 57736 26743
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 57736 26581
rect 57295 22923 57736 26525
rect 57295 22035 57363 22923
rect 57627 22035 57736 22923
rect 57295 16678 57736 22035
rect 57295 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 57736 16678
rect 57295 16461 57736 16622
rect 57295 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 57736 16461
rect 57295 16243 57736 16405
rect 57295 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 57736 16243
rect 57295 16026 57736 16187
rect 57295 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 57736 16026
rect 57295 15808 57736 15970
rect 57295 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 57736 15808
rect 57295 15590 57736 15752
rect 57295 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 57736 15590
rect 57295 15372 57736 15534
rect 57295 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 57736 15372
rect 57295 15155 57736 15316
rect 57295 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 57736 15155
rect 57295 14937 57736 15099
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 57736 14937
rect 57295 14720 57736 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 57736 14720
rect 57295 11406 57736 14664
rect 57295 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 57736 11406
rect 57295 11189 57736 11350
rect 57295 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 57736 11189
rect 57295 10971 57736 11133
rect 57295 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 57736 10971
rect 57295 10753 57736 10915
rect 57295 10697 57381 10753
rect 57437 10697 57593 10753
rect 57649 10697 57736 10753
rect 57295 10535 57736 10697
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 57736 10535
rect 57295 10318 57736 10479
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 57736 10318
rect 27387 9876 27476 9928
rect 27528 9876 27688 9928
rect 27740 9876 27828 9928
rect 27387 9710 27828 9876
rect 51756 9971 51832 9981
rect 51756 9811 51766 9971
rect 51822 9811 51832 9971
rect 51756 9801 51832 9811
rect 27387 9658 27476 9710
rect 27528 9658 27688 9710
rect 27740 9658 27828 9710
rect 27387 9493 27828 9658
rect 27387 9441 27476 9493
rect 27528 9441 27688 9493
rect 27740 9441 27828 9493
rect 27387 9275 27828 9441
rect 27387 9223 27476 9275
rect 27528 9223 27688 9275
rect 27740 9223 27828 9275
rect 27387 9057 27828 9223
rect 27387 9005 27476 9057
rect 27528 9005 27688 9057
rect 27740 9005 27828 9057
rect 27387 8840 27828 9005
rect 49887 8953 50067 8963
rect 49887 8897 49897 8953
rect 50057 8897 50067 8953
rect 49887 8887 50067 8897
rect 27387 8788 27476 8840
rect 27528 8788 27688 8840
rect 27740 8788 27828 8840
rect 27387 8622 27828 8788
rect 27387 8570 27476 8622
rect 27528 8570 27688 8622
rect 27740 8570 27828 8622
rect 27387 8404 27828 8570
rect 27387 8352 27476 8404
rect 27528 8352 27688 8404
rect 27740 8352 27828 8404
rect 27387 8187 27828 8352
rect 27387 8135 27476 8187
rect 27528 8135 27688 8187
rect 27740 8135 27828 8187
rect 27387 7969 27828 8135
rect 27387 7917 27476 7969
rect 27528 7917 27688 7969
rect 27740 7917 27828 7969
rect 27387 7752 27828 7917
rect 27387 7700 27476 7752
rect 27528 7700 27688 7752
rect 27740 7700 27828 7752
rect 27387 7535 27828 7700
rect 27387 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 27387 7317 27828 7479
rect 27387 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 27387 7099 27828 7261
rect 27387 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 27387 6881 27828 7043
rect 27387 6829 27476 6881
rect 27528 6829 27688 6881
rect 27740 6829 27828 6881
rect 27387 6663 27828 6829
rect 27387 6611 27476 6663
rect 27528 6611 27688 6663
rect 27740 6611 27828 6663
rect 27387 6446 27828 6611
rect 27387 6394 27476 6446
rect 27528 6394 27688 6446
rect 27740 6394 27828 6446
rect 27387 6228 27828 6394
rect 28237 6836 28999 6874
rect 28237 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 28999 6836
rect 28237 6618 28999 6780
rect 28237 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 28999 6618
rect 28237 6400 28999 6562
rect 28237 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 28999 6400
rect 49958 6361 50014 8887
rect 28237 6306 28999 6344
rect 49896 6349 50076 6361
rect 49896 6297 49908 6349
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6176 27476 6228
rect 27528 6176 27688 6228
rect 27740 6176 27828 6228
rect 27387 6120 27828 6176
rect 27387 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 27828 6120
rect 27387 6011 27828 6064
rect 27387 5959 27476 6011
rect 27528 5959 27688 6011
rect 27740 5959 27828 6011
rect 27387 5902 27828 5959
rect 27387 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 27828 5902
rect 27387 5793 27828 5846
rect 27387 5741 27476 5793
rect 27528 5741 27688 5793
rect 27740 5741 27828 5793
rect 27387 5575 27828 5741
rect 27387 5523 27476 5575
rect 27528 5523 27688 5575
rect 27740 5523 27828 5575
rect 27387 5358 27828 5523
rect 27387 5306 27476 5358
rect 27528 5306 27688 5358
rect 27740 5306 27828 5358
rect 1864 5024 2509 5135
rect 11727 5073 11783 5140
rect 1864 0 2088 5024
rect 3263 5001 3357 5062
rect 11617 5017 11783 5073
rect 3263 4880 3604 5001
rect 2539 1689 2763 1701
rect 2539 1637 2574 1689
rect 2730 1637 2763 1689
rect 2539 0 2763 1637
rect 3380 0 3604 4880
rect 11617 1700 11673 5017
rect 12575 4740 12631 5185
rect 12290 4684 12631 4740
rect 13253 4740 13309 5185
rect 14101 5073 14157 5140
rect 23375 5134 23953 5135
rect 14101 5017 14267 5073
rect 13253 4684 13594 4740
rect 12290 1700 12346 4684
rect 11533 0 11757 1700
rect 12206 0 12430 1700
rect 12604 1689 12828 1701
rect 12604 1637 12639 1689
rect 12795 1637 12828 1689
rect 12604 0 12828 1637
rect 13054 1689 13278 1701
rect 13538 1700 13594 4684
rect 14211 1700 14267 5017
rect 22527 5001 22621 5062
rect 23375 5024 24019 5134
rect 22345 4880 22621 5001
rect 22345 1701 22439 4880
rect 13054 1637 13089 1689
rect 13245 1637 13278 1689
rect 13054 0 13278 1637
rect 13454 0 13678 1700
rect 14127 0 14351 1700
rect 22279 0 22503 1701
rect 23404 1689 23628 1701
rect 23404 1637 23439 1689
rect 23595 1637 23628 1689
rect 23404 0 23628 1637
rect 23795 0 24019 5024
rect 26823 4587 27163 4628
rect 26823 4535 26861 4587
rect 26913 4535 27073 4587
rect 27125 4535 27163 4587
rect 26823 4528 27163 4535
rect 26823 4472 26859 4528
rect 26915 4472 27071 4528
rect 27127 4472 27163 4528
rect 26823 4370 27163 4472
rect 26823 4318 26861 4370
rect 26913 4318 27073 4370
rect 27125 4318 27163 4370
rect 26823 4310 27163 4318
rect 26823 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 27163 4310
rect 26823 4152 27163 4254
rect 26823 4100 26861 4152
rect 26913 4100 27073 4152
rect 27125 4100 27163 4152
rect 26823 3934 27163 4100
rect 26823 3882 26861 3934
rect 26913 3882 27073 3934
rect 27125 3882 27163 3934
rect 26823 3717 27163 3882
rect 26823 3665 26861 3717
rect 26913 3665 27073 3717
rect 27125 3665 27163 3717
rect 26823 3624 27163 3665
rect 27387 4587 27828 5306
rect 27387 4535 27476 4587
rect 27528 4535 27688 4587
rect 27740 4535 27828 4587
rect 27387 4370 27828 4535
rect 27387 4318 27476 4370
rect 27528 4318 27688 4370
rect 27740 4318 27828 4370
rect 27387 4152 27828 4318
rect 27387 4100 27476 4152
rect 27528 4100 27688 4152
rect 27740 4100 27828 4152
rect 27387 3934 27828 4100
rect 27387 3882 27476 3934
rect 27528 3882 27688 3934
rect 27740 3882 27828 3934
rect 27387 3837 27828 3882
rect 27387 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 27828 3837
rect 27387 3717 27828 3781
rect 27387 3665 27476 3717
rect 27528 3665 27688 3717
rect 27740 3665 27828 3717
rect 27387 3619 27828 3665
rect 27387 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 27828 3619
rect 27387 3524 27828 3563
rect 28764 3837 28894 3876
rect 28764 3781 28801 3837
rect 28857 3781 28894 3837
rect 28764 3619 28894 3781
rect 28764 3563 28801 3619
rect 28857 3563 28894 3619
rect 28764 3525 28894 3563
rect 27936 2730 28070 3418
rect 27936 0 28160 2730
rect 29006 2433 29135 3418
rect 29247 2944 29377 3418
rect 29247 2720 29929 2944
rect 29006 914 29230 2433
rect 29006 654 29090 914
rect 29142 654 29230 914
rect 29006 0 29230 654
rect 29705 914 29929 2720
rect 29705 654 29787 914
rect 29839 654 29929 914
rect 29705 0 29929 654
rect 30859 0 31083 6229
rect 32552 0 32776 6229
rect 34243 0 34467 6229
rect 51766 5211 51822 9801
rect 57295 8934 57736 10262
rect 57295 8878 57386 8934
rect 57442 8878 57510 8934
rect 57566 8878 57634 8934
rect 57690 8878 57736 8934
rect 57295 8810 57736 8878
rect 57295 8754 57386 8810
rect 57442 8754 57510 8810
rect 57566 8754 57634 8810
rect 57690 8754 57736 8810
rect 57295 8686 57736 8754
rect 57295 8630 57386 8686
rect 57442 8630 57510 8686
rect 57566 8630 57634 8686
rect 57690 8630 57736 8686
rect 57295 8562 57736 8630
rect 57295 8506 57386 8562
rect 57442 8506 57510 8562
rect 57566 8506 57634 8562
rect 57690 8506 57736 8562
rect 57295 8438 57736 8506
rect 57295 8382 57386 8438
rect 57442 8382 57510 8438
rect 57566 8382 57634 8438
rect 57690 8382 57736 8438
rect 57295 8314 57736 8382
rect 57295 8258 57386 8314
rect 57442 8258 57510 8314
rect 57566 8258 57634 8314
rect 57690 8258 57736 8314
rect 57295 8190 57736 8258
rect 57295 8134 57386 8190
rect 57442 8134 57510 8190
rect 57566 8134 57634 8190
rect 57690 8134 57736 8190
rect 57295 8066 57736 8134
rect 57295 8010 57386 8066
rect 57442 8010 57510 8066
rect 57566 8010 57634 8066
rect 57690 8010 57736 8066
rect 57295 7942 57736 8010
rect 57295 7886 57386 7942
rect 57442 7886 57510 7942
rect 57566 7886 57634 7942
rect 57690 7886 57736 7942
rect 57295 7818 57736 7886
rect 57295 7762 57386 7818
rect 57442 7762 57510 7818
rect 57566 7762 57634 7818
rect 57690 7762 57736 7818
rect 57295 7694 57736 7762
rect 57295 7638 57386 7694
rect 57442 7638 57510 7694
rect 57566 7638 57634 7694
rect 57690 7638 57736 7694
rect 57295 7570 57736 7638
rect 57295 7514 57386 7570
rect 57442 7514 57510 7570
rect 57566 7514 57634 7570
rect 57690 7514 57736 7570
rect 57295 7446 57736 7514
rect 57295 7390 57386 7446
rect 57442 7390 57510 7446
rect 57566 7390 57634 7446
rect 57690 7390 57736 7446
rect 57295 7322 57736 7390
rect 57295 7266 57386 7322
rect 57442 7266 57510 7322
rect 57566 7266 57634 7322
rect 57690 7266 57736 7322
rect 57295 7198 57736 7266
rect 57295 7142 57386 7198
rect 57442 7142 57510 7198
rect 57566 7142 57634 7198
rect 57690 7142 57736 7198
rect 56124 6836 56886 6874
rect 56124 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 56886 6836
rect 56124 6618 56886 6780
rect 56124 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 56886 6618
rect 56124 6400 56886 6562
rect 56124 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 56886 6400
rect 56124 6306 56886 6344
rect 51642 5199 51822 5211
rect 51642 5147 51654 5199
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 6120 57736 7142
rect 57295 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 57736 6120
rect 57295 5902 57736 6064
rect 57295 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 57736 5902
rect 40588 3282 40812 3294
rect 40588 3230 40623 3282
rect 40779 3230 40812 3282
rect 40588 0 40812 3230
rect 43790 3044 43970 3054
rect 43790 2988 43800 3044
rect 43960 2988 43970 3044
rect 43790 2978 43970 2988
rect 48644 2822 48997 3873
rect 48644 2766 48671 2822
rect 48727 2766 48795 2822
rect 48851 2766 48919 2822
rect 48975 2766 48997 2822
rect 48644 2698 48997 2766
rect 48644 2642 48671 2698
rect 48727 2642 48795 2698
rect 48851 2642 48919 2698
rect 48975 2642 48997 2698
rect 48644 2574 48997 2642
rect 48644 2518 48671 2574
rect 48727 2518 48795 2574
rect 48851 2518 48919 2574
rect 48975 2518 48997 2574
rect 48644 1023 48997 2518
rect 48644 971 48668 1023
rect 48720 971 48792 1023
rect 48844 971 48916 1023
rect 48968 971 48997 1023
rect 48644 899 48997 971
rect 48644 847 48668 899
rect 48720 847 48792 899
rect 48844 847 48916 899
rect 48968 847 48997 899
rect 48644 775 48997 847
rect 48644 723 48668 775
rect 48720 723 48792 775
rect 48844 723 48916 775
rect 48968 723 48997 775
rect 48644 651 48997 723
rect 48644 599 48668 651
rect 48720 599 48792 651
rect 48844 599 48916 651
rect 48968 599 48997 651
rect 48644 0 48997 599
rect 49145 2143 49498 4618
rect 57295 4587 57736 5846
rect 57295 4535 57383 4587
rect 57435 4535 57595 4587
rect 57647 4535 57736 4587
rect 49145 2087 49161 2143
rect 49217 2087 49285 2143
rect 49341 2087 49409 2143
rect 49465 2087 49498 2143
rect 49145 2019 49498 2087
rect 49145 1963 49161 2019
rect 49217 1963 49285 2019
rect 49341 1963 49409 2019
rect 49465 1963 49498 2019
rect 49145 1895 49498 1963
rect 49145 1839 49161 1895
rect 49217 1839 49285 1895
rect 49341 1839 49409 1895
rect 49465 1839 49498 1895
rect 49145 0 49498 1839
rect 50342 0 50566 4382
rect 57295 4370 57736 4535
rect 57295 4318 57383 4370
rect 57435 4318 57595 4370
rect 57647 4318 57736 4370
rect 57295 4152 57736 4318
rect 57295 4100 57383 4152
rect 57435 4100 57595 4152
rect 57647 4100 57736 4152
rect 57295 3934 57736 4100
rect 57295 3882 57383 3934
rect 57435 3882 57595 3934
rect 57647 3882 57736 3934
rect 57295 3837 57736 3882
rect 57295 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 57736 3837
rect 57295 3717 57736 3781
rect 57295 3665 57383 3717
rect 57435 3665 57595 3717
rect 57647 3665 57736 3717
rect 57295 3619 57736 3665
rect 57295 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 57736 3619
rect 57295 3524 57736 3563
rect 57909 34011 58351 44776
rect 57909 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 58351 34011
rect 57909 33793 58351 33955
rect 57909 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 58351 33793
rect 57909 33576 58351 33737
rect 57909 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 58351 33576
rect 57909 33432 58351 33520
rect 57909 33380 57998 33432
rect 58050 33380 58210 33432
rect 58262 33380 58351 33432
rect 57909 33358 58351 33380
rect 57909 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 58351 33358
rect 57909 33215 58351 33302
rect 57909 33163 57998 33215
rect 58050 33163 58210 33215
rect 58262 33163 58351 33215
rect 57909 33140 58351 33163
rect 57909 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 58351 33140
rect 57909 32997 58351 33084
rect 57909 32945 57998 32997
rect 58050 32945 58210 32997
rect 58262 32945 58351 32997
rect 57909 32922 58351 32945
rect 57909 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 58351 32922
rect 57909 32779 58351 32866
rect 57909 32727 57998 32779
rect 58050 32727 58210 32779
rect 58262 32727 58351 32779
rect 57909 32705 58351 32727
rect 57909 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 58351 32705
rect 57909 32562 58351 32649
rect 57909 32510 57998 32562
rect 58050 32510 58210 32562
rect 58262 32510 58351 32562
rect 57909 32487 58351 32510
rect 57909 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 58351 32487
rect 57909 32344 58351 32431
rect 57909 32292 57998 32344
rect 58050 32292 58210 32344
rect 58262 32292 58351 32344
rect 57909 32127 58351 32292
rect 57909 32088 57998 32127
rect 58050 32088 58210 32127
rect 58262 32088 58351 32127
rect 57909 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 57909 31909 58351 32032
rect 57909 31870 57998 31909
rect 58050 31870 58210 31909
rect 58262 31870 58351 31909
rect 57909 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 57909 31691 58351 31814
rect 57909 31652 57998 31691
rect 58050 31652 58210 31691
rect 58262 31652 58351 31691
rect 57909 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 57909 31474 58351 31596
rect 57909 31422 57998 31474
rect 58050 31422 58210 31474
rect 58262 31422 58351 31474
rect 57909 31256 58351 31422
rect 57909 31204 57998 31256
rect 58050 31204 58210 31256
rect 58262 31204 58351 31256
rect 57909 31038 58351 31204
rect 57909 30986 57998 31038
rect 58050 30986 58210 31038
rect 58262 30986 58351 31038
rect 57909 30821 58351 30986
rect 57909 30769 57998 30821
rect 58050 30769 58210 30821
rect 58262 30769 58351 30821
rect 57909 30603 58351 30769
rect 57909 30551 57998 30603
rect 58050 30551 58210 30603
rect 58262 30551 58351 30603
rect 57909 30386 58351 30551
rect 57909 30334 57998 30386
rect 58050 30334 58210 30386
rect 58262 30334 58351 30386
rect 57909 30168 58351 30334
rect 57909 30116 57998 30168
rect 58050 30116 58210 30168
rect 58262 30116 58351 30168
rect 57909 29968 58351 30116
rect 57909 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 57909 29898 57998 29912
rect 58050 29898 58210 29912
rect 58262 29898 58351 29912
rect 57909 29750 58351 29898
rect 57909 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29694 58351 29750
rect 57909 29681 57998 29694
rect 58050 29681 58210 29694
rect 58262 29681 58351 29694
rect 57909 29533 58351 29681
rect 57909 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 58351 29533
rect 57909 29463 57998 29477
rect 58050 29463 58210 29477
rect 58262 29463 58351 29477
rect 57909 29315 58351 29463
rect 57909 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 57909 29245 57998 29259
rect 58050 29245 58210 29259
rect 58262 29245 58351 29259
rect 57909 29098 58351 29245
rect 57909 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 57909 29028 57998 29042
rect 58050 29028 58210 29042
rect 58262 29028 58351 29042
rect 57909 28880 58351 29028
rect 57909 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 57909 28810 57998 28824
rect 58050 28810 58210 28824
rect 58262 28810 58351 28824
rect 57909 28662 58351 28810
rect 57909 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 57909 28592 57998 28606
rect 58050 28592 58210 28606
rect 58262 28592 58351 28606
rect 57909 28444 58351 28592
rect 57909 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 57909 28375 57998 28388
rect 58050 28375 58210 28388
rect 58262 28375 58351 28388
rect 57909 28227 58351 28375
rect 57909 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 57909 28157 57998 28171
rect 58050 28157 58210 28171
rect 58262 28157 58351 28171
rect 57909 28009 58351 28157
rect 57909 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 57909 27940 57998 27953
rect 58050 27940 58210 27953
rect 58262 27940 58351 27953
rect 57909 27792 58351 27940
rect 57909 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 57909 27722 57998 27736
rect 58050 27722 58210 27736
rect 58262 27722 58351 27736
rect 57909 27574 58351 27722
rect 57909 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 57909 27504 57998 27518
rect 58050 27504 58210 27518
rect 58262 27504 58351 27518
rect 57909 27339 58351 27504
rect 57909 27287 57998 27339
rect 58050 27287 58210 27339
rect 58262 27287 58351 27339
rect 57909 27121 58351 27287
rect 57909 27069 57998 27121
rect 58050 27069 58210 27121
rect 58262 27069 58351 27121
rect 57909 26903 58351 27069
rect 57909 26851 57998 26903
rect 58050 26851 58210 26903
rect 58262 26851 58351 26903
rect 57909 26686 58351 26851
rect 57909 26634 57998 26686
rect 58050 26634 58210 26686
rect 58262 26634 58351 26686
rect 57909 26468 58351 26634
rect 57909 26416 57998 26468
rect 58050 26416 58210 26468
rect 58262 26416 58351 26468
rect 58791 44338 59517 44384
rect 58791 44314 58814 44338
rect 58866 44314 58938 44338
rect 58990 44314 59062 44338
rect 59114 44314 59186 44338
rect 59238 44314 59310 44338
rect 59362 44314 59434 44338
rect 59486 44314 59517 44338
rect 58791 44258 58812 44314
rect 58868 44258 58936 44314
rect 58992 44258 59060 44314
rect 59116 44258 59184 44314
rect 59240 44258 59308 44314
rect 59364 44258 59432 44314
rect 59488 44258 59517 44314
rect 58791 44214 59517 44258
rect 58791 44190 58814 44214
rect 58866 44190 58938 44214
rect 58990 44190 59062 44214
rect 59114 44190 59186 44214
rect 59238 44190 59310 44214
rect 59362 44190 59434 44214
rect 59486 44190 59517 44214
rect 58791 44134 58812 44190
rect 58868 44134 58936 44190
rect 58992 44134 59060 44190
rect 59116 44134 59184 44190
rect 59240 44134 59308 44190
rect 59364 44134 59432 44190
rect 59488 44134 59517 44190
rect 58791 31298 59517 44134
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 84368 35316 84493 35943
rect 58791 31242 58873 31298
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59517 31298
rect 58791 31174 59517 31242
rect 58791 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59517 31174
rect 58791 31050 59517 31118
rect 58791 30994 58873 31050
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59517 31050
rect 58791 30853 59517 30994
rect 58791 30797 58873 30853
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59517 30853
rect 58791 30729 59517 30797
rect 58791 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59517 30729
rect 58791 30605 59517 30673
rect 58791 30549 58873 30605
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59517 30605
rect 58791 28272 59517 30549
rect 58791 28216 58859 28272
rect 58915 28216 58983 28272
rect 59039 28216 59107 28272
rect 59163 28216 59231 28272
rect 59287 28216 59355 28272
rect 59411 28216 59517 28272
rect 58791 28148 59517 28216
rect 58791 28092 58859 28148
rect 58915 28092 58983 28148
rect 59039 28092 59107 28148
rect 59163 28092 59231 28148
rect 59287 28092 59355 28148
rect 59411 28092 59517 28148
rect 58791 28024 59517 28092
rect 58791 27968 58859 28024
rect 58915 27968 58983 28024
rect 59039 27968 59107 28024
rect 59163 27968 59231 28024
rect 59287 27968 59355 28024
rect 59411 27968 59517 28024
rect 58791 27900 59517 27968
rect 58791 27844 58859 27900
rect 58915 27844 58983 27900
rect 59039 27844 59107 27900
rect 59163 27844 59231 27900
rect 59287 27844 59355 27900
rect 59411 27844 59517 27900
rect 58791 27776 59517 27844
rect 58791 27720 58859 27776
rect 58915 27720 58983 27776
rect 59039 27720 59107 27776
rect 59163 27720 59231 27776
rect 59287 27720 59355 27776
rect 59411 27720 59517 27776
rect 58791 27652 59517 27720
rect 58791 27596 58859 27652
rect 58915 27596 58983 27652
rect 59039 27596 59107 27652
rect 59163 27596 59231 27652
rect 59287 27596 59355 27652
rect 59411 27596 59517 27652
rect 58791 27528 59517 27596
rect 58791 27472 58859 27528
rect 58915 27472 58983 27528
rect 59039 27472 59107 27528
rect 59163 27472 59231 27528
rect 59287 27472 59355 27528
rect 59411 27472 59517 27528
rect 58791 27404 59517 27472
rect 58791 27348 58859 27404
rect 58915 27348 58983 27404
rect 59039 27348 59107 27404
rect 59163 27348 59231 27404
rect 59287 27348 59355 27404
rect 59411 27348 59517 27404
rect 58791 27280 59517 27348
rect 58791 27224 58859 27280
rect 58915 27224 58983 27280
rect 59039 27224 59107 27280
rect 59163 27224 59231 27280
rect 59287 27224 59355 27280
rect 59411 27224 59517 27280
rect 58791 27156 59517 27224
rect 58791 27100 58859 27156
rect 58915 27100 58983 27156
rect 59039 27100 59107 27156
rect 59163 27100 59231 27156
rect 59287 27100 59355 27156
rect 59411 27100 59517 27156
rect 58791 27032 59517 27100
rect 58791 26976 58859 27032
rect 58915 26976 58983 27032
rect 59039 26976 59107 27032
rect 59163 26976 59231 27032
rect 59287 26976 59355 27032
rect 59411 26976 59517 27032
rect 58791 26908 59517 26976
rect 58791 26852 58859 26908
rect 58915 26852 58983 26908
rect 59039 26852 59107 26908
rect 59163 26852 59231 26908
rect 59287 26852 59355 26908
rect 59411 26852 59517 26908
rect 58791 26784 59517 26852
rect 58791 26728 58859 26784
rect 58915 26728 58983 26784
rect 59039 26728 59107 26784
rect 59163 26728 59231 26784
rect 59287 26728 59355 26784
rect 59411 26728 59517 26784
rect 58791 26660 59517 26728
rect 58791 26604 58859 26660
rect 58915 26604 58983 26660
rect 59039 26604 59107 26660
rect 59163 26604 59231 26660
rect 59287 26604 59355 26660
rect 59411 26604 59517 26660
rect 58791 26536 59517 26604
rect 58791 26480 58859 26536
rect 58915 26480 58983 26536
rect 59039 26480 59107 26536
rect 59163 26480 59231 26536
rect 59287 26480 59355 26536
rect 59411 26480 59517 26536
rect 58791 26433 59517 26480
rect 57909 26250 58351 26416
rect 57909 26198 57998 26250
rect 58050 26198 58210 26250
rect 58262 26198 58351 26250
rect 57909 26033 58351 26198
rect 57909 25981 57998 26033
rect 58050 25981 58210 26033
rect 58262 25981 58351 26033
rect 57909 25815 58351 25981
rect 57909 25763 57998 25815
rect 58050 25763 58210 25815
rect 58262 25763 58351 25815
rect 57909 25598 58351 25763
rect 57909 25546 57998 25598
rect 58050 25546 58210 25598
rect 58262 25546 58351 25598
rect 57909 25380 58351 25546
rect 57909 25328 57998 25380
rect 58050 25328 58210 25380
rect 58262 25328 58351 25380
rect 57909 25162 58351 25328
rect 57909 25110 57998 25162
rect 58050 25110 58210 25162
rect 58262 25110 58351 25162
rect 57909 24945 58351 25110
rect 57909 24893 57998 24945
rect 58050 24893 58210 24945
rect 58262 24893 58351 24945
rect 57909 24727 58351 24893
rect 57909 24675 57998 24727
rect 58050 24675 58210 24727
rect 58262 24675 58351 24727
rect 57909 24509 58351 24675
rect 57909 24457 57998 24509
rect 58050 24457 58210 24509
rect 58262 24457 58351 24509
rect 57909 24292 58351 24457
rect 57909 24240 57998 24292
rect 58050 24240 58210 24292
rect 58262 24240 58351 24292
rect 57909 24075 58351 24240
rect 57909 23187 57994 24075
rect 58258 24074 58351 24075
rect 58262 24022 58351 24074
rect 58258 23857 58351 24022
rect 58262 23805 58351 23857
rect 58258 23639 58351 23805
rect 58262 23587 58351 23639
rect 58258 23421 58351 23587
rect 58262 23369 58351 23421
rect 58258 23204 58351 23369
rect 57909 23152 57998 23187
rect 58050 23152 58210 23187
rect 58262 23152 58351 23204
rect 57909 22986 58351 23152
rect 57909 22934 57998 22986
rect 58050 22934 58210 22986
rect 58262 22934 58351 22986
rect 57909 22768 58351 22934
rect 57909 22716 57998 22768
rect 58050 22716 58210 22768
rect 58262 22716 58351 22768
rect 57909 22551 58351 22716
rect 57909 22499 57998 22551
rect 58050 22499 58210 22551
rect 58262 22499 58351 22551
rect 57909 22333 58351 22499
rect 57909 22281 57998 22333
rect 58050 22281 58210 22333
rect 58262 22281 58351 22333
rect 57909 22115 58351 22281
rect 57909 22063 57998 22115
rect 58050 22063 58210 22115
rect 58262 22063 58351 22115
rect 57909 21898 58351 22063
rect 57909 21846 57998 21898
rect 58050 21846 58210 21898
rect 58262 21846 58351 21898
rect 57909 21680 58351 21846
rect 57909 21628 57998 21680
rect 58050 21628 58210 21680
rect 58262 21628 58351 21680
rect 57909 21463 58351 21628
rect 57909 21411 57998 21463
rect 58050 21411 58210 21463
rect 58262 21411 58351 21463
rect 57909 21245 58351 21411
rect 57909 21193 57998 21245
rect 58050 21193 58210 21245
rect 58262 21193 58351 21245
rect 57909 21027 58351 21193
rect 57909 20975 57998 21027
rect 58050 20975 58210 21027
rect 58262 20975 58351 21027
rect 57909 20810 58351 20975
rect 57909 20758 57998 20810
rect 58050 20758 58210 20810
rect 58262 20758 58351 20810
rect 57909 20592 58351 20758
rect 57909 20540 57998 20592
rect 58050 20570 58210 20592
rect 58208 20540 58210 20570
rect 58262 20540 58351 20592
rect 57909 20410 58048 20540
rect 58208 20410 58351 20540
rect 57909 20374 58351 20410
rect 57909 20322 57998 20374
rect 58050 20322 58210 20374
rect 58262 20322 58351 20374
rect 57909 20226 58351 20322
rect 57909 20157 58048 20226
rect 58208 20157 58351 20226
rect 57909 20105 57998 20157
rect 58208 20105 58210 20157
rect 58262 20105 58351 20157
rect 57909 20066 58048 20105
rect 58208 20066 58351 20105
rect 57909 19939 58351 20066
rect 57909 19887 57998 19939
rect 58050 19887 58210 19939
rect 58262 19887 58351 19939
rect 57909 19722 58351 19887
rect 57909 19670 57998 19722
rect 58050 19670 58210 19722
rect 58262 19670 58351 19722
rect 57909 19504 58351 19670
rect 57909 19452 57998 19504
rect 58050 19452 58210 19504
rect 58262 19452 58351 19504
rect 57909 19286 58351 19452
rect 57909 19234 57998 19286
rect 58050 19234 58210 19286
rect 58262 19234 58351 19286
rect 57909 19068 58351 19234
rect 57909 19016 57998 19068
rect 58050 19016 58210 19068
rect 58262 19016 58351 19068
rect 57909 18851 58351 19016
rect 57909 18799 57998 18851
rect 58050 18799 58210 18851
rect 58262 18799 58351 18851
rect 57909 18633 58351 18799
rect 57909 18581 57998 18633
rect 58050 18581 58210 18633
rect 58262 18581 58351 18633
rect 57909 18416 58351 18581
rect 57909 18364 57998 18416
rect 58050 18364 58210 18416
rect 58262 18364 58351 18416
rect 57909 18198 58351 18364
rect 57909 18146 57998 18198
rect 58050 18146 58210 18198
rect 58262 18146 58351 18198
rect 57909 17980 58351 18146
rect 57909 17928 57998 17980
rect 58050 17928 58210 17980
rect 58262 17928 58351 17980
rect 57909 17763 58351 17928
rect 57909 17711 57998 17763
rect 58050 17711 58210 17763
rect 58262 17711 58351 17763
rect 57909 17545 58351 17711
rect 57909 17493 57998 17545
rect 58050 17493 58210 17545
rect 58262 17493 58351 17545
rect 57909 17327 58351 17493
rect 57909 17275 57998 17327
rect 58050 17275 58210 17327
rect 58262 17275 58351 17327
rect 57909 17110 58351 17275
rect 57909 17058 57998 17110
rect 58050 17058 58210 17110
rect 58262 17058 58351 17110
rect 57909 16892 58351 17058
rect 57909 16840 57998 16892
rect 58050 16840 58210 16892
rect 58262 16840 58351 16892
rect 57909 16675 58351 16840
rect 57909 16623 57998 16675
rect 58050 16623 58210 16675
rect 58262 16623 58351 16675
rect 57909 16457 58351 16623
rect 57909 16405 57998 16457
rect 58050 16405 58210 16457
rect 58262 16405 58351 16457
rect 57909 16239 58351 16405
rect 57909 16187 57998 16239
rect 58050 16187 58210 16239
rect 58262 16187 58351 16239
rect 57909 16022 58351 16187
rect 57909 15970 57998 16022
rect 58050 15970 58210 16022
rect 58262 15970 58351 16022
rect 57909 15804 58351 15970
rect 57909 15752 57998 15804
rect 58050 15752 58210 15804
rect 58262 15752 58351 15804
rect 57909 15586 58351 15752
rect 57909 15534 57998 15586
rect 58050 15534 58210 15586
rect 58262 15534 58351 15586
rect 57909 15369 58351 15534
rect 57909 15317 57998 15369
rect 58050 15317 58210 15369
rect 58262 15317 58351 15369
rect 57909 15151 58351 15317
rect 57909 15099 57998 15151
rect 58050 15099 58210 15151
rect 58262 15099 58351 15151
rect 57909 14933 58351 15099
rect 57909 14881 57998 14933
rect 58050 14881 58210 14933
rect 58262 14881 58351 14933
rect 57909 14716 58351 14881
rect 57909 14664 57998 14716
rect 58050 14664 58210 14716
rect 58262 14664 58351 14716
rect 57909 14498 58351 14664
rect 57909 14446 57998 14498
rect 58050 14446 58210 14498
rect 58262 14446 58351 14498
rect 57909 14281 58351 14446
rect 57909 14229 57998 14281
rect 58050 14229 58210 14281
rect 58262 14229 58351 14281
rect 57909 14063 58351 14229
rect 57909 14011 57998 14063
rect 58050 14011 58210 14063
rect 58262 14011 58351 14063
rect 57909 13845 58351 14011
rect 57909 13793 57998 13845
rect 58050 13793 58210 13845
rect 58262 13793 58351 13845
rect 57909 13790 58351 13793
rect 57909 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 58351 13790
rect 57909 13628 58351 13734
rect 57909 13576 57998 13628
rect 58050 13576 58210 13628
rect 58262 13576 58351 13628
rect 57909 13573 58351 13576
rect 57909 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 58351 13573
rect 57909 13410 58351 13517
rect 57909 13358 57998 13410
rect 58050 13358 58210 13410
rect 58262 13358 58351 13410
rect 57909 13355 58351 13358
rect 57909 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58351 13355
rect 57909 13192 58351 13299
rect 57909 13140 57998 13192
rect 58050 13140 58210 13192
rect 58262 13140 58351 13192
rect 57909 13138 58351 13140
rect 57909 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58351 13138
rect 57909 12975 58351 13082
rect 57909 12923 57998 12975
rect 58050 12923 58210 12975
rect 58262 12923 58351 12975
rect 57909 12920 58351 12923
rect 57909 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58351 12920
rect 57909 12757 58351 12864
rect 57909 12705 57998 12757
rect 58050 12705 58210 12757
rect 58262 12705 58351 12757
rect 57909 12702 58351 12705
rect 57909 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 58351 12702
rect 57909 12540 58351 12646
rect 57909 12488 57998 12540
rect 58050 12488 58210 12540
rect 58262 12488 58351 12540
rect 57909 12484 58351 12488
rect 57909 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 58351 12484
rect 57909 12322 58351 12428
rect 57909 12270 57998 12322
rect 58050 12270 58210 12322
rect 58262 12270 58351 12322
rect 57909 12267 58351 12270
rect 57909 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 58351 12267
rect 57909 12104 58351 12211
rect 57909 12052 57998 12104
rect 58050 12052 58210 12104
rect 58262 12052 58351 12104
rect 57909 12049 58351 12052
rect 57909 11993 57996 12049
rect 58052 11993 58208 12049
rect 58264 11993 58351 12049
rect 57909 11887 58351 11993
rect 57909 11835 57998 11887
rect 58050 11835 58210 11887
rect 58262 11835 58351 11887
rect 57909 11832 58351 11835
rect 57909 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 57909 11669 58351 11776
rect 57909 11617 57998 11669
rect 58050 11617 58210 11669
rect 58262 11617 58351 11669
rect 57909 11451 58351 11617
rect 57909 11399 57998 11451
rect 58050 11399 58210 11451
rect 58262 11399 58351 11451
rect 57909 11234 58351 11399
rect 57909 11182 57998 11234
rect 58050 11182 58210 11234
rect 58262 11182 58351 11234
rect 57909 11016 58351 11182
rect 57909 10964 57998 11016
rect 58050 10964 58210 11016
rect 58262 10964 58351 11016
rect 57909 10798 58351 10964
rect 57909 10746 57998 10798
rect 58050 10746 58210 10798
rect 58262 10746 58351 10798
rect 57909 10581 58351 10746
rect 57909 10529 57998 10581
rect 58050 10529 58210 10581
rect 58262 10529 58351 10581
rect 57909 10363 58351 10529
rect 57909 10311 57998 10363
rect 58050 10311 58210 10363
rect 58262 10311 58351 10363
rect 57909 10146 58351 10311
rect 57909 10094 57998 10146
rect 58050 10094 58210 10146
rect 58262 10094 58351 10146
rect 57909 9928 58351 10094
rect 57909 9876 57998 9928
rect 58050 9876 58210 9928
rect 58262 9876 58351 9928
rect 57909 9710 58351 9876
rect 57909 9658 57998 9710
rect 58050 9658 58210 9710
rect 58262 9658 58351 9710
rect 57909 9493 58351 9658
rect 57909 9441 57998 9493
rect 58050 9441 58210 9493
rect 58262 9441 58351 9493
rect 57909 9407 58351 9441
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 58351 9407
rect 57909 9275 58351 9351
rect 57909 9223 57998 9275
rect 58050 9223 58210 9275
rect 58262 9223 58351 9275
rect 57909 9190 58351 9223
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 58351 9190
rect 57909 9057 58351 9134
rect 57909 9005 57998 9057
rect 58050 9005 58210 9057
rect 58262 9005 58351 9057
rect 57909 8972 58351 9005
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 58351 8972
rect 57909 8840 58351 8916
rect 57909 8788 57998 8840
rect 58050 8788 58210 8840
rect 58262 8788 58351 8840
rect 57909 8754 58351 8788
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 58351 8754
rect 57909 8622 58351 8698
rect 57909 8570 57998 8622
rect 58050 8570 58210 8622
rect 58262 8570 58351 8622
rect 57909 8536 58351 8570
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 58351 8536
rect 57909 8404 58351 8480
rect 57909 8352 57998 8404
rect 58050 8352 58210 8404
rect 58262 8352 58351 8404
rect 57909 8319 58351 8352
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 58351 8319
rect 57909 8187 58351 8263
rect 57909 8135 57998 8187
rect 58050 8135 58210 8187
rect 58262 8135 58351 8187
rect 57909 7969 58351 8135
rect 57909 7917 57998 7969
rect 58050 7917 58210 7969
rect 58262 7917 58351 7969
rect 57909 7752 58351 7917
rect 57909 7700 57998 7752
rect 58050 7700 58210 7752
rect 58262 7700 58351 7752
rect 57909 7534 58351 7700
rect 57909 7482 57998 7534
rect 58050 7482 58210 7534
rect 58262 7482 58351 7534
rect 57909 7316 58351 7482
rect 57909 7264 57998 7316
rect 58050 7264 58210 7316
rect 58262 7264 58351 7316
rect 57909 7099 58351 7264
rect 57909 7047 57998 7099
rect 58050 7047 58210 7099
rect 58262 7047 58351 7099
rect 57909 6881 58351 7047
rect 57909 6829 57998 6881
rect 58050 6829 58210 6881
rect 58262 6829 58351 6881
rect 57909 6663 58351 6829
rect 57909 6611 57998 6663
rect 58050 6611 58210 6663
rect 58262 6611 58351 6663
rect 57909 6446 58351 6611
rect 57909 6394 57998 6446
rect 58050 6394 58210 6446
rect 58262 6394 58351 6446
rect 57909 6228 58351 6394
rect 57909 6176 57998 6228
rect 58050 6176 58210 6228
rect 58262 6176 58351 6228
rect 57909 6011 58351 6176
rect 57909 5959 57998 6011
rect 58050 5959 58210 6011
rect 58262 5959 58351 6011
rect 57909 5793 58351 5959
rect 57909 5741 57998 5793
rect 58050 5741 58210 5793
rect 58262 5741 58351 5793
rect 57909 5575 58351 5741
rect 57909 5539 57998 5575
rect 58050 5539 58210 5575
rect 58262 5539 58351 5575
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 58351 5539
rect 57909 5358 58351 5483
rect 57909 5321 57998 5358
rect 58050 5321 58210 5358
rect 58262 5321 58351 5358
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 58351 5321
rect 57909 4587 58351 5265
rect 57909 4535 57998 4587
rect 58050 4535 58210 4587
rect 58262 4535 58351 4587
rect 57909 4528 58351 4535
rect 57909 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4472 58351 4528
rect 57909 4370 58351 4472
rect 57909 4318 57998 4370
rect 58050 4318 58210 4370
rect 58262 4318 58351 4370
rect 57909 4310 58351 4318
rect 57909 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 58351 4310
rect 57909 4152 58351 4254
rect 57909 4100 57998 4152
rect 58050 4100 58210 4152
rect 58262 4100 58351 4152
rect 57909 3934 58351 4100
rect 57909 3882 57998 3934
rect 58050 3882 58210 3934
rect 58262 3882 58351 3934
rect 57909 3717 58351 3882
rect 57909 3665 57998 3717
rect 58050 3665 58210 3717
rect 58262 3665 58351 3717
rect 57909 3524 58351 3665
rect 61447 5024 62085 5135
rect 71303 5073 71359 5140
rect 53772 3218 55669 3418
rect 53772 1006 53996 3218
rect 55781 2983 55911 3418
rect 53772 642 53907 1006
rect 53959 642 53996 1006
rect 53772 0 53996 642
rect 54417 2783 55911 2983
rect 54417 0 54641 2783
rect 56023 2567 56152 3418
rect 55164 2367 56152 2567
rect 55164 0 55388 2367
rect 56265 0 56489 3418
rect 61447 0 61671 5024
rect 62839 5001 62933 5062
rect 71193 5017 71359 5073
rect 62839 4880 63115 5001
rect 63021 1701 63115 4880
rect 71193 1701 71249 5017
rect 72151 4740 72207 5185
rect 71866 4684 72207 4740
rect 72829 4740 72885 5185
rect 73677 5073 73733 5140
rect 73677 5017 73843 5073
rect 72829 4684 73170 4740
rect 71866 1701 71922 4684
rect 73114 1701 73170 4684
rect 73787 1701 73843 5017
rect 82103 5001 82197 5062
rect 82951 5024 83596 5135
rect 81921 4880 82197 5001
rect 81921 1701 82015 4880
rect 62115 1689 62339 1701
rect 62115 1637 62150 1689
rect 62306 1637 62339 1689
rect 62115 0 62339 1637
rect 62958 0 63182 1701
rect 71109 0 71333 1701
rect 71782 0 72006 1701
rect 72180 1689 72404 1701
rect 72180 1637 72215 1689
rect 72371 1637 72404 1689
rect 72180 0 72404 1637
rect 72630 1689 72854 1701
rect 72630 1637 72665 1689
rect 72821 1637 72854 1689
rect 72630 0 72854 1637
rect 73030 0 73254 1701
rect 73703 0 73927 1701
rect 81855 0 82079 1701
rect 82695 1689 82919 1701
rect 82695 1637 82730 1689
rect 82886 1637 82919 1689
rect 82695 0 82919 1637
rect 83372 0 83596 5024
<< via2 >>
rect 25335 44286 25337 44314
rect 25337 44286 25389 44314
rect 25389 44286 25391 44314
rect 25335 44258 25391 44286
rect 25459 44286 25461 44314
rect 25461 44286 25513 44314
rect 25513 44286 25515 44314
rect 25459 44258 25515 44286
rect 25583 44286 25585 44314
rect 25585 44286 25637 44314
rect 25637 44286 25639 44314
rect 25583 44258 25639 44286
rect 25707 44286 25709 44314
rect 25709 44286 25761 44314
rect 25761 44286 25763 44314
rect 25707 44258 25763 44286
rect 25831 44286 25833 44314
rect 25833 44286 25885 44314
rect 25885 44286 25887 44314
rect 25831 44258 25887 44286
rect 25955 44286 25957 44314
rect 25957 44286 26009 44314
rect 26009 44286 26011 44314
rect 25955 44258 26011 44286
rect 25335 44162 25337 44190
rect 25337 44162 25389 44190
rect 25389 44162 25391 44190
rect 25335 44134 25391 44162
rect 25459 44162 25461 44190
rect 25461 44162 25513 44190
rect 25513 44162 25515 44190
rect 25459 44134 25515 44162
rect 25583 44162 25585 44190
rect 25585 44162 25637 44190
rect 25637 44162 25639 44190
rect 25583 44134 25639 44162
rect 25707 44162 25709 44190
rect 25709 44162 25761 44190
rect 25761 44162 25763 44190
rect 25707 44134 25763 44162
rect 25831 44162 25833 44190
rect 25833 44162 25885 44190
rect 25885 44162 25887 44190
rect 25831 44134 25887 44162
rect 25955 44162 25957 44190
rect 25957 44162 26009 44190
rect 26009 44162 26011 44190
rect 25955 44134 26011 44162
rect 25398 34848 25454 34877
rect 25398 34821 25400 34848
rect 25400 34821 25452 34848
rect 25452 34821 25454 34848
rect 25522 34848 25578 34877
rect 25522 34821 25524 34848
rect 25524 34821 25576 34848
rect 25576 34821 25578 34848
rect 25646 34848 25702 34877
rect 25646 34821 25648 34848
rect 25648 34821 25700 34848
rect 25700 34821 25702 34848
rect 25770 34848 25826 34877
rect 25770 34821 25772 34848
rect 25772 34821 25824 34848
rect 25824 34821 25826 34848
rect 25894 34848 25950 34877
rect 25894 34821 25896 34848
rect 25896 34821 25948 34848
rect 25948 34821 25950 34848
rect 25398 34724 25454 34753
rect 25398 34697 25400 34724
rect 25400 34697 25452 34724
rect 25452 34697 25454 34724
rect 25522 34724 25578 34753
rect 25522 34697 25524 34724
rect 25524 34697 25576 34724
rect 25576 34697 25578 34724
rect 25646 34724 25702 34753
rect 25646 34697 25648 34724
rect 25648 34697 25700 34724
rect 25700 34697 25702 34724
rect 25770 34724 25826 34753
rect 25770 34697 25772 34724
rect 25772 34697 25824 34724
rect 25824 34697 25826 34724
rect 25894 34724 25950 34753
rect 25894 34697 25896 34724
rect 25896 34697 25948 34724
rect 25948 34697 25950 34724
rect 25398 34573 25454 34629
rect 25522 34573 25578 34629
rect 25646 34573 25702 34629
rect 25770 34573 25826 34629
rect 25894 34573 25950 34629
rect 25398 31192 25454 31248
rect 25522 31192 25578 31248
rect 25646 31192 25702 31248
rect 25770 31192 25826 31248
rect 25894 31192 25950 31248
rect 25398 31068 25454 31124
rect 25522 31068 25578 31124
rect 25646 31068 25702 31124
rect 25770 31068 25826 31124
rect 25894 31068 25950 31124
rect 25398 30944 25454 31000
rect 25522 30944 25578 31000
rect 25646 30944 25702 31000
rect 25770 30944 25826 31000
rect 25894 30944 25950 31000
rect 25398 30737 25454 30793
rect 25522 30737 25578 30793
rect 25646 30737 25702 30793
rect 25770 30737 25826 30793
rect 25894 30737 25950 30793
rect 25398 30613 25454 30669
rect 25522 30613 25578 30669
rect 25646 30613 25702 30669
rect 25770 30613 25826 30669
rect 25894 30613 25950 30669
rect 25398 30489 25454 30545
rect 25522 30489 25578 30545
rect 25646 30489 25702 30545
rect 25770 30489 25826 30545
rect 25894 30489 25950 30545
rect 25404 28226 25460 28282
rect 25528 28226 25584 28282
rect 25652 28226 25708 28282
rect 25776 28226 25832 28282
rect 25900 28226 25956 28282
rect 25404 28102 25460 28158
rect 25528 28102 25584 28158
rect 25652 28102 25708 28158
rect 25776 28102 25832 28158
rect 25900 28102 25956 28158
rect 25404 27978 25460 28034
rect 25528 27978 25584 28034
rect 25652 27978 25708 28034
rect 25776 27978 25832 28034
rect 25900 27978 25956 28034
rect 25404 27854 25460 27910
rect 25528 27854 25584 27910
rect 25652 27854 25708 27910
rect 25776 27854 25832 27910
rect 25900 27854 25956 27910
rect 25404 27730 25460 27786
rect 25528 27730 25584 27786
rect 25652 27730 25708 27786
rect 25776 27730 25832 27786
rect 25900 27730 25956 27786
rect 25404 27606 25460 27662
rect 25528 27606 25584 27662
rect 25652 27606 25708 27662
rect 25776 27606 25832 27662
rect 25900 27606 25956 27662
rect 25404 27482 25460 27538
rect 25528 27482 25584 27538
rect 25652 27482 25708 27538
rect 25776 27482 25832 27538
rect 25900 27482 25956 27538
rect 25404 27358 25460 27414
rect 25528 27358 25584 27414
rect 25652 27358 25708 27414
rect 25776 27358 25832 27414
rect 25900 27358 25956 27414
rect 25404 27234 25460 27290
rect 25528 27234 25584 27290
rect 25652 27234 25708 27290
rect 25776 27234 25832 27290
rect 25900 27234 25956 27290
rect 25404 27110 25460 27166
rect 25528 27110 25584 27166
rect 25652 27110 25708 27166
rect 25776 27110 25832 27166
rect 25900 27110 25956 27166
rect 25404 26986 25460 27042
rect 25528 26986 25584 27042
rect 25652 26986 25708 27042
rect 25776 26986 25832 27042
rect 25900 26986 25956 27042
rect 25404 26862 25460 26918
rect 25528 26862 25584 26918
rect 25652 26862 25708 26918
rect 25776 26862 25832 26918
rect 25900 26862 25956 26918
rect 25404 26738 25460 26794
rect 25528 26738 25584 26794
rect 25652 26738 25708 26794
rect 25776 26738 25832 26794
rect 25900 26738 25956 26794
rect 25404 26614 25460 26670
rect 25528 26614 25584 26670
rect 25652 26614 25708 26670
rect 25776 26614 25832 26670
rect 25900 26614 25956 26670
rect 25404 26490 25460 26546
rect 25528 26490 25584 26546
rect 25652 26490 25708 26546
rect 25776 26490 25832 26546
rect 25900 26490 25956 26546
rect 26838 43361 26894 43417
rect 26962 43361 27018 43417
rect 27086 43361 27142 43417
rect 26838 43237 26894 43293
rect 26962 43237 27018 43293
rect 27086 43237 27142 43293
rect 26838 36162 26894 36218
rect 26962 36162 27018 36218
rect 27086 36162 27142 36218
rect 26838 36038 26894 36094
rect 26962 36038 27018 36094
rect 27086 36038 27142 36094
rect 26859 33955 26915 34011
rect 27071 33955 27127 34011
rect 26859 33737 26915 33793
rect 27071 33737 27127 33793
rect 26859 33520 26915 33576
rect 27071 33520 27127 33576
rect 26859 33302 26915 33358
rect 27071 33302 27127 33358
rect 26859 33084 26915 33140
rect 27071 33084 27127 33140
rect 26859 32866 26915 32922
rect 27071 32866 27127 32922
rect 26859 32649 26915 32705
rect 27071 32649 27127 32705
rect 26859 32431 26915 32487
rect 27071 32431 27127 32487
rect 26859 32075 26861 32088
rect 26861 32075 26913 32088
rect 26913 32075 26915 32088
rect 26859 32032 26915 32075
rect 27071 32075 27073 32088
rect 27073 32075 27125 32088
rect 27125 32075 27127 32088
rect 27071 32032 27127 32075
rect 26859 31857 26861 31870
rect 26861 31857 26913 31870
rect 26913 31857 26915 31870
rect 26859 31814 26915 31857
rect 27071 31857 27073 31870
rect 27073 31857 27125 31870
rect 27125 31857 27127 31870
rect 27071 31814 27127 31857
rect 26859 31639 26861 31652
rect 26861 31639 26913 31652
rect 26913 31639 26915 31652
rect 26859 31596 26915 31639
rect 27071 31639 27073 31652
rect 27073 31639 27125 31652
rect 27125 31639 27127 31652
rect 27071 31596 27127 31639
rect 26859 29950 26915 29968
rect 26859 29912 26861 29950
rect 26861 29912 26913 29950
rect 26913 29912 26915 29950
rect 27071 29950 27127 29968
rect 27071 29912 27073 29950
rect 27073 29912 27125 29950
rect 27125 29912 27127 29950
rect 26859 29733 26915 29750
rect 26859 29694 26861 29733
rect 26861 29694 26913 29733
rect 26913 29694 26915 29733
rect 27071 29733 27127 29750
rect 27071 29694 27073 29733
rect 27073 29694 27125 29733
rect 27125 29694 27127 29733
rect 26859 29515 26915 29533
rect 26859 29477 26861 29515
rect 26861 29477 26913 29515
rect 26913 29477 26915 29515
rect 27071 29515 27127 29533
rect 27071 29477 27073 29515
rect 27073 29477 27125 29515
rect 27125 29477 27127 29515
rect 26859 29297 26915 29315
rect 26859 29259 26861 29297
rect 26861 29259 26913 29297
rect 26913 29259 26915 29297
rect 27071 29297 27127 29315
rect 27071 29259 27073 29297
rect 27073 29259 27125 29297
rect 27125 29259 27127 29297
rect 26859 29080 26915 29098
rect 26859 29042 26861 29080
rect 26861 29042 26913 29080
rect 26913 29042 26915 29080
rect 27071 29080 27127 29098
rect 27071 29042 27073 29080
rect 27073 29042 27125 29080
rect 27125 29042 27127 29080
rect 26859 28862 26915 28880
rect 26859 28824 26861 28862
rect 26861 28824 26913 28862
rect 26913 28824 26915 28862
rect 27071 28862 27127 28880
rect 27071 28824 27073 28862
rect 27073 28824 27125 28862
rect 27125 28824 27127 28862
rect 26859 28644 26915 28662
rect 26859 28606 26861 28644
rect 26861 28606 26913 28644
rect 26913 28606 26915 28644
rect 27071 28644 27127 28662
rect 27071 28606 27073 28644
rect 27073 28606 27125 28644
rect 27125 28606 27127 28644
rect 26859 28427 26915 28444
rect 26859 28388 26861 28427
rect 26861 28388 26913 28427
rect 26913 28388 26915 28427
rect 27071 28427 27127 28444
rect 27071 28388 27073 28427
rect 27073 28388 27125 28427
rect 27125 28388 27127 28427
rect 26859 28209 26915 28227
rect 26859 28171 26861 28209
rect 26861 28171 26913 28209
rect 26913 28171 26915 28209
rect 27071 28209 27127 28227
rect 27071 28171 27073 28209
rect 27073 28171 27125 28209
rect 27125 28171 27127 28209
rect 26859 27992 26915 28009
rect 26859 27953 26861 27992
rect 26861 27953 26913 27992
rect 26913 27953 26915 27992
rect 27071 27992 27127 28009
rect 27071 27953 27073 27992
rect 27073 27953 27125 27992
rect 27125 27953 27127 27992
rect 26859 27774 26915 27792
rect 26859 27736 26861 27774
rect 26861 27736 26913 27774
rect 26913 27736 26915 27774
rect 27071 27774 27127 27792
rect 27071 27736 27073 27774
rect 27073 27736 27125 27774
rect 27125 27736 27127 27774
rect 26859 27556 26915 27574
rect 26859 27518 26861 27556
rect 26861 27518 26913 27556
rect 26913 27518 26915 27556
rect 27071 27556 27127 27574
rect 27071 27518 27073 27556
rect 27073 27518 27125 27556
rect 27125 27518 27127 27556
rect 26450 26126 26610 26286
rect 26092 25807 26252 25967
rect 25756 25487 25916 25647
rect 25421 25168 25581 25328
rect 25081 24477 25241 24637
rect 24744 24156 24904 24316
rect 24416 23835 24576 23995
rect 24057 23513 24217 23673
rect 26465 19532 26625 19692
rect 26858 24171 27122 24227
rect 26858 24074 27122 24085
rect 26858 24029 26861 24074
rect 26861 24029 26913 24074
rect 26913 24029 27073 24074
rect 27073 24029 27122 24074
rect 26858 23887 27122 23943
rect 26858 23745 27122 23801
rect 26858 23639 27122 23659
rect 26858 23603 26861 23639
rect 26861 23603 26913 23639
rect 26913 23603 27073 23639
rect 27073 23603 27122 23639
rect 26858 23461 27122 23517
rect 26858 23369 26861 23375
rect 26861 23369 26913 23375
rect 26913 23369 27073 23375
rect 27073 23369 27122 23375
rect 26858 23319 27122 23369
rect 26858 23204 27122 23233
rect 26858 23177 26861 23204
rect 26861 23177 26913 23204
rect 26913 23177 27073 23204
rect 27073 23177 27122 23204
rect 26858 23035 27122 23091
rect 26924 20540 27073 20570
rect 27073 20540 27084 20570
rect 26924 20410 27084 20540
rect 26924 20157 27084 20226
rect 26924 20105 27073 20157
rect 27073 20105 27084 20157
rect 26924 20066 27084 20105
rect 26107 19187 26267 19347
rect 25771 18867 25931 19027
rect 25434 18524 25594 18684
rect 25094 18190 25254 18350
rect 24757 17817 24917 17977
rect 24429 17496 24589 17656
rect 24069 17157 24229 17317
rect 26859 14063 26915 14119
rect 27071 14063 27127 14119
rect 26859 13846 26915 13902
rect 27071 13846 27127 13902
rect 26859 13628 26915 13684
rect 27071 13628 27127 13684
rect 26859 13411 26915 13467
rect 27071 13411 27127 13467
rect 26859 13193 26915 13249
rect 27071 13193 27127 13249
rect 26859 12975 26915 13031
rect 27071 12975 27127 13031
rect 26859 12757 26915 12813
rect 27071 12757 27127 12813
rect 26859 12540 26915 12596
rect 27071 12540 27127 12596
rect 26859 12322 26915 12378
rect 27071 12322 27127 12378
rect 26859 12105 26915 12161
rect 27071 12105 27127 12161
rect 26859 9351 26915 9407
rect 27071 9351 27127 9407
rect 26859 9134 26915 9190
rect 27071 9134 27127 9190
rect 26859 8916 26915 8972
rect 27071 8916 27127 8972
rect 26859 8698 26915 8754
rect 27071 8698 27127 8754
rect 26859 8480 26915 8536
rect 27071 8480 27127 8536
rect 26859 8263 26915 8319
rect 27071 8263 27127 8319
rect 26859 5523 26861 5539
rect 26861 5523 26913 5539
rect 26913 5523 26915 5539
rect 26859 5483 26915 5523
rect 27071 5523 27073 5539
rect 27073 5523 27125 5539
rect 27125 5523 27127 5539
rect 27071 5483 27127 5523
rect 26859 5306 26861 5321
rect 26861 5306 26913 5321
rect 26913 5306 26915 5321
rect 26859 5265 26915 5306
rect 27071 5306 27073 5321
rect 27073 5306 27125 5321
rect 27125 5306 27127 5321
rect 27071 5265 27127 5306
rect 27788 44253 27844 44255
rect 27788 44201 27790 44253
rect 27790 44201 27842 44253
rect 27842 44201 27844 44253
rect 27788 44199 27844 44201
rect 27999 44253 28055 44255
rect 27999 44201 28001 44253
rect 28001 44201 28053 44253
rect 28053 44201 28055 44253
rect 27999 44199 28055 44201
rect 28210 44253 28266 44255
rect 28210 44201 28212 44253
rect 28212 44201 28264 44253
rect 28264 44201 28266 44253
rect 28210 44199 28266 44201
rect 28421 44253 28477 44255
rect 28421 44201 28423 44253
rect 28423 44201 28475 44253
rect 28475 44201 28477 44253
rect 28421 44199 28477 44201
rect 28632 44253 28688 44255
rect 28632 44201 28634 44253
rect 28634 44201 28686 44253
rect 28686 44201 28688 44253
rect 28632 44199 28688 44201
rect 28843 44253 28899 44255
rect 28843 44201 28845 44253
rect 28845 44201 28897 44253
rect 28897 44201 28899 44253
rect 28843 44199 28899 44201
rect 29054 44253 29110 44255
rect 29054 44201 29056 44253
rect 29056 44201 29108 44253
rect 29108 44201 29110 44253
rect 29054 44199 29110 44201
rect 29580 43353 29636 43355
rect 29580 43301 29582 43353
rect 29582 43301 29634 43353
rect 29634 43301 29636 43353
rect 29580 43299 29636 43301
rect 29791 43353 29847 43355
rect 29791 43301 29793 43353
rect 29793 43301 29845 43353
rect 29845 43301 29847 43353
rect 29791 43299 29847 43301
rect 30003 43353 30059 43355
rect 30003 43301 30005 43353
rect 30005 43301 30057 43353
rect 30057 43301 30059 43353
rect 30003 43299 30059 43301
rect 30214 43353 30270 43355
rect 30214 43301 30216 43353
rect 30216 43301 30268 43353
rect 30268 43301 30270 43353
rect 30214 43299 30270 43301
rect 34288 44253 34344 44255
rect 34288 44201 34290 44253
rect 34290 44201 34342 44253
rect 34342 44201 34344 44253
rect 34288 44199 34344 44201
rect 34499 44253 34555 44255
rect 34499 44201 34501 44253
rect 34501 44201 34553 44253
rect 34553 44201 34555 44253
rect 34499 44199 34555 44201
rect 34710 44253 34766 44255
rect 34710 44201 34712 44253
rect 34712 44201 34764 44253
rect 34764 44201 34766 44253
rect 34710 44199 34766 44201
rect 34921 44253 34977 44255
rect 34921 44201 34923 44253
rect 34923 44201 34975 44253
rect 34975 44201 34977 44253
rect 34921 44199 34977 44201
rect 33048 43772 33104 43774
rect 33048 43720 33050 43772
rect 33050 43720 33102 43772
rect 33102 43720 33104 43772
rect 33048 43718 33104 43720
rect 33259 43772 33315 43774
rect 33259 43720 33261 43772
rect 33261 43720 33313 43772
rect 33313 43720 33315 43772
rect 33259 43718 33315 43720
rect 33470 43772 33526 43774
rect 33470 43720 33472 43772
rect 33472 43720 33524 43772
rect 33524 43720 33526 43772
rect 33470 43718 33526 43720
rect 33681 43772 33737 43774
rect 33681 43720 33683 43772
rect 33683 43720 33735 43772
rect 33735 43720 33737 43772
rect 33681 43718 33737 43720
rect 33892 43772 33948 43774
rect 33892 43720 33894 43772
rect 33894 43720 33946 43772
rect 33946 43720 33948 43772
rect 33892 43718 33948 43720
rect 30852 43353 30908 43355
rect 27788 42453 27844 42455
rect 27788 42401 27790 42453
rect 27790 42401 27842 42453
rect 27842 42401 27844 42453
rect 27788 42399 27844 42401
rect 27999 42453 28055 42455
rect 27999 42401 28001 42453
rect 28001 42401 28053 42453
rect 28053 42401 28055 42453
rect 27999 42399 28055 42401
rect 28210 42453 28266 42455
rect 28210 42401 28212 42453
rect 28212 42401 28264 42453
rect 28264 42401 28266 42453
rect 28210 42399 28266 42401
rect 28421 42453 28477 42455
rect 28421 42401 28423 42453
rect 28423 42401 28475 42453
rect 28475 42401 28477 42453
rect 28421 42399 28477 42401
rect 28632 42453 28688 42455
rect 28632 42401 28634 42453
rect 28634 42401 28686 42453
rect 28686 42401 28688 42453
rect 28632 42399 28688 42401
rect 28843 42453 28899 42455
rect 28843 42401 28845 42453
rect 28845 42401 28897 42453
rect 28897 42401 28899 42453
rect 28843 42399 28899 42401
rect 29054 42453 29110 42455
rect 29054 42401 29056 42453
rect 29056 42401 29108 42453
rect 29108 42401 29110 42453
rect 29054 42399 29110 42401
rect 29580 41553 29636 41555
rect 29580 41501 29582 41553
rect 29582 41501 29634 41553
rect 29634 41501 29636 41553
rect 29580 41499 29636 41501
rect 29791 41553 29847 41555
rect 29791 41501 29793 41553
rect 29793 41501 29845 41553
rect 29845 41501 29847 41553
rect 29791 41499 29847 41501
rect 30003 41553 30059 41555
rect 30003 41501 30005 41553
rect 30005 41501 30057 41553
rect 30057 41501 30059 41553
rect 30003 41499 30059 41501
rect 30214 41553 30270 41555
rect 30214 41501 30216 41553
rect 30216 41501 30268 41553
rect 30268 41501 30270 41553
rect 30214 41499 30270 41501
rect 27788 40653 27844 40655
rect 27788 40601 27790 40653
rect 27790 40601 27842 40653
rect 27842 40601 27844 40653
rect 27788 40599 27844 40601
rect 27999 40653 28055 40655
rect 27999 40601 28001 40653
rect 28001 40601 28053 40653
rect 28053 40601 28055 40653
rect 27999 40599 28055 40601
rect 28210 40653 28266 40655
rect 28210 40601 28212 40653
rect 28212 40601 28264 40653
rect 28264 40601 28266 40653
rect 28210 40599 28266 40601
rect 28421 40653 28477 40655
rect 28421 40601 28423 40653
rect 28423 40601 28475 40653
rect 28475 40601 28477 40653
rect 28421 40599 28477 40601
rect 28632 40653 28688 40655
rect 28632 40601 28634 40653
rect 28634 40601 28686 40653
rect 28686 40601 28688 40653
rect 28632 40599 28688 40601
rect 28843 40653 28899 40655
rect 28843 40601 28845 40653
rect 28845 40601 28897 40653
rect 28897 40601 28899 40653
rect 28843 40599 28899 40601
rect 29054 40653 29110 40655
rect 29054 40601 29056 40653
rect 29056 40601 29108 40653
rect 29108 40601 29110 40653
rect 29054 40599 29110 40601
rect 29580 39753 29636 39755
rect 29580 39701 29582 39753
rect 29582 39701 29634 39753
rect 29634 39701 29636 39753
rect 29580 39699 29636 39701
rect 29791 39753 29847 39755
rect 29791 39701 29793 39753
rect 29793 39701 29845 39753
rect 29845 39701 29847 39753
rect 29791 39699 29847 39701
rect 30003 39753 30059 39755
rect 30003 39701 30005 39753
rect 30005 39701 30057 39753
rect 30057 39701 30059 39753
rect 30003 39699 30059 39701
rect 30214 39753 30270 39755
rect 30214 39701 30216 39753
rect 30216 39701 30268 39753
rect 30268 39701 30270 39753
rect 30214 39699 30270 39701
rect 27788 38853 27844 38855
rect 27788 38801 27790 38853
rect 27790 38801 27842 38853
rect 27842 38801 27844 38853
rect 27788 38799 27844 38801
rect 27999 38853 28055 38855
rect 27999 38801 28001 38853
rect 28001 38801 28053 38853
rect 28053 38801 28055 38853
rect 27999 38799 28055 38801
rect 28210 38853 28266 38855
rect 28210 38801 28212 38853
rect 28212 38801 28264 38853
rect 28264 38801 28266 38853
rect 28210 38799 28266 38801
rect 28421 38853 28477 38855
rect 28421 38801 28423 38853
rect 28423 38801 28475 38853
rect 28475 38801 28477 38853
rect 28421 38799 28477 38801
rect 28632 38853 28688 38855
rect 28632 38801 28634 38853
rect 28634 38801 28686 38853
rect 28686 38801 28688 38853
rect 28632 38799 28688 38801
rect 28843 38853 28899 38855
rect 28843 38801 28845 38853
rect 28845 38801 28897 38853
rect 28897 38801 28899 38853
rect 28843 38799 28899 38801
rect 29054 38853 29110 38855
rect 29054 38801 29056 38853
rect 29056 38801 29108 38853
rect 29108 38801 29110 38853
rect 29054 38799 29110 38801
rect 29580 37953 29636 37955
rect 29580 37901 29582 37953
rect 29582 37901 29634 37953
rect 29634 37901 29636 37953
rect 29580 37899 29636 37901
rect 29791 37953 29847 37955
rect 29791 37901 29793 37953
rect 29793 37901 29845 37953
rect 29845 37901 29847 37953
rect 29791 37899 29847 37901
rect 30003 37953 30059 37955
rect 30003 37901 30005 37953
rect 30005 37901 30057 37953
rect 30057 37901 30059 37953
rect 30003 37899 30059 37901
rect 30214 37953 30270 37955
rect 30214 37901 30216 37953
rect 30216 37901 30268 37953
rect 30268 37901 30270 37953
rect 30214 37899 30270 37901
rect 27788 37053 27844 37055
rect 27788 37001 27790 37053
rect 27790 37001 27842 37053
rect 27842 37001 27844 37053
rect 27788 36999 27844 37001
rect 27999 37053 28055 37055
rect 27999 37001 28001 37053
rect 28001 37001 28053 37053
rect 28053 37001 28055 37053
rect 27999 36999 28055 37001
rect 28210 37053 28266 37055
rect 28210 37001 28212 37053
rect 28212 37001 28264 37053
rect 28264 37001 28266 37053
rect 28210 36999 28266 37001
rect 28421 37053 28477 37055
rect 28421 37001 28423 37053
rect 28423 37001 28475 37053
rect 28475 37001 28477 37053
rect 28421 36999 28477 37001
rect 28632 37053 28688 37055
rect 28632 37001 28634 37053
rect 28634 37001 28686 37053
rect 28686 37001 28688 37053
rect 28632 36999 28688 37001
rect 28843 37053 28899 37055
rect 28843 37001 28845 37053
rect 28845 37001 28897 37053
rect 28897 37001 28899 37053
rect 28843 36999 28899 37001
rect 29054 37053 29110 37055
rect 29054 37001 29056 37053
rect 29056 37001 29108 37053
rect 29108 37001 29110 37053
rect 29054 36999 29110 37001
rect 29580 36153 29636 36155
rect 29580 36101 29582 36153
rect 29582 36101 29634 36153
rect 29634 36101 29636 36153
rect 29580 36099 29636 36101
rect 29791 36153 29847 36155
rect 29791 36101 29793 36153
rect 29793 36101 29845 36153
rect 29845 36101 29847 36153
rect 29791 36099 29847 36101
rect 30003 36153 30059 36155
rect 30003 36101 30005 36153
rect 30005 36101 30057 36153
rect 30057 36101 30059 36153
rect 30003 36099 30059 36101
rect 30214 36153 30270 36155
rect 30214 36101 30216 36153
rect 30216 36101 30268 36153
rect 30268 36101 30270 36153
rect 30214 36099 30270 36101
rect 30852 43301 30854 43353
rect 30854 43301 30906 43353
rect 30906 43301 30908 43353
rect 30852 43299 30908 43301
rect 31063 43353 31119 43355
rect 31063 43301 31065 43353
rect 31065 43301 31117 43353
rect 31117 43301 31119 43353
rect 31063 43299 31119 43301
rect 31274 43353 31330 43355
rect 31274 43301 31276 43353
rect 31276 43301 31328 43353
rect 31328 43301 31330 43353
rect 31274 43299 31330 43301
rect 31484 43353 31540 43355
rect 31484 43301 31486 43353
rect 31486 43301 31538 43353
rect 31538 43301 31540 43353
rect 31484 43299 31540 43301
rect 31695 43353 31751 43355
rect 31695 43301 31697 43353
rect 31697 43301 31749 43353
rect 31749 43301 31751 43353
rect 31695 43299 31751 43301
rect 31907 43353 31963 43355
rect 31907 43301 31909 43353
rect 31909 43301 31961 43353
rect 31961 43301 31963 43353
rect 31907 43299 31963 43301
rect 32118 43353 32174 43355
rect 32118 43301 32120 43353
rect 32120 43301 32172 43353
rect 32172 43301 32174 43353
rect 32118 43299 32174 43301
rect 32328 43353 32384 43355
rect 32328 43301 32330 43353
rect 32330 43301 32382 43353
rect 32382 43301 32384 43353
rect 32328 43299 32384 43301
rect 32539 43353 32595 43355
rect 32539 43301 32541 43353
rect 32541 43301 32593 43353
rect 32593 43301 32595 43353
rect 32539 43299 32595 43301
rect 32750 43353 32806 43355
rect 32750 43301 32752 43353
rect 32752 43301 32804 43353
rect 32804 43301 32806 43353
rect 32750 43299 32806 43301
rect 35218 43353 35274 43355
rect 33055 42866 33111 42922
rect 33235 42866 33291 42922
rect 33817 42859 33873 42915
rect 33997 42859 34053 42915
rect 34282 42399 34338 42455
rect 34493 42399 34549 42455
rect 34705 42453 34761 42455
rect 34916 42453 34972 42455
rect 34705 42401 34755 42453
rect 34755 42401 34761 42453
rect 34916 42401 34935 42453
rect 34935 42401 34972 42453
rect 34705 42399 34761 42401
rect 34916 42399 34972 42401
rect 33055 41932 33111 41988
rect 33235 41932 33291 41988
rect 33817 41939 33873 41995
rect 33997 41939 34053 41995
rect 30852 41553 30908 41555
rect 30852 41501 30854 41553
rect 30854 41501 30906 41553
rect 30906 41501 30908 41553
rect 30852 41499 30908 41501
rect 31063 41553 31119 41555
rect 31063 41501 31065 41553
rect 31065 41501 31117 41553
rect 31117 41501 31119 41553
rect 31063 41499 31119 41501
rect 31274 41553 31330 41555
rect 31274 41501 31276 41553
rect 31276 41501 31328 41553
rect 31328 41501 31330 41553
rect 31274 41499 31330 41501
rect 31484 41553 31540 41555
rect 31484 41501 31486 41553
rect 31486 41501 31538 41553
rect 31538 41501 31540 41553
rect 31484 41499 31540 41501
rect 31695 41553 31751 41555
rect 31695 41501 31697 41553
rect 31697 41501 31749 41553
rect 31749 41501 31751 41553
rect 31695 41499 31751 41501
rect 31907 41553 31963 41555
rect 31907 41501 31909 41553
rect 31909 41501 31961 41553
rect 31961 41501 31963 41553
rect 31907 41499 31963 41501
rect 32118 41553 32174 41555
rect 32118 41501 32120 41553
rect 32120 41501 32172 41553
rect 32172 41501 32174 41553
rect 32118 41499 32174 41501
rect 32328 41553 32384 41555
rect 32328 41501 32330 41553
rect 32330 41501 32382 41553
rect 32382 41501 32384 41553
rect 32328 41499 32384 41501
rect 32539 41553 32595 41555
rect 32539 41501 32541 41553
rect 32541 41501 32593 41553
rect 32593 41501 32595 41553
rect 32539 41499 32595 41501
rect 32750 41553 32806 41555
rect 32750 41501 32752 41553
rect 32752 41501 32804 41553
rect 32804 41501 32806 41553
rect 32750 41499 32806 41501
rect 33055 41066 33111 41122
rect 33235 41066 33291 41122
rect 33817 41059 33873 41115
rect 33997 41059 34053 41115
rect 34282 40599 34338 40655
rect 34493 40599 34549 40655
rect 34705 40653 34761 40655
rect 34916 40653 34972 40655
rect 34705 40601 34755 40653
rect 34755 40601 34761 40653
rect 34916 40601 34935 40653
rect 34935 40601 34972 40653
rect 34705 40599 34761 40601
rect 34916 40599 34972 40601
rect 33055 40132 33111 40188
rect 33235 40132 33291 40188
rect 33817 40139 33873 40195
rect 33997 40139 34053 40195
rect 30852 39753 30908 39755
rect 30852 39701 30854 39753
rect 30854 39701 30906 39753
rect 30906 39701 30908 39753
rect 30852 39699 30908 39701
rect 31063 39753 31119 39755
rect 31063 39701 31065 39753
rect 31065 39701 31117 39753
rect 31117 39701 31119 39753
rect 31063 39699 31119 39701
rect 31274 39753 31330 39755
rect 31274 39701 31276 39753
rect 31276 39701 31328 39753
rect 31328 39701 31330 39753
rect 31274 39699 31330 39701
rect 31484 39753 31540 39755
rect 31484 39701 31486 39753
rect 31486 39701 31538 39753
rect 31538 39701 31540 39753
rect 31484 39699 31540 39701
rect 31695 39753 31751 39755
rect 31695 39701 31697 39753
rect 31697 39701 31749 39753
rect 31749 39701 31751 39753
rect 31695 39699 31751 39701
rect 31907 39753 31963 39755
rect 31907 39701 31909 39753
rect 31909 39701 31961 39753
rect 31961 39701 31963 39753
rect 31907 39699 31963 39701
rect 32118 39753 32174 39755
rect 32118 39701 32120 39753
rect 32120 39701 32172 39753
rect 32172 39701 32174 39753
rect 32118 39699 32174 39701
rect 32328 39753 32384 39755
rect 32328 39701 32330 39753
rect 32330 39701 32382 39753
rect 32382 39701 32384 39753
rect 32328 39699 32384 39701
rect 32539 39753 32595 39755
rect 32539 39701 32541 39753
rect 32541 39701 32593 39753
rect 32593 39701 32595 39753
rect 32539 39699 32595 39701
rect 32750 39753 32806 39755
rect 32750 39701 32752 39753
rect 32752 39701 32804 39753
rect 32804 39701 32806 39753
rect 32750 39699 32806 39701
rect 33055 39266 33111 39322
rect 33235 39266 33291 39322
rect 33817 39259 33873 39315
rect 33997 39259 34053 39315
rect 34282 38799 34338 38855
rect 34493 38799 34549 38855
rect 34705 38853 34761 38855
rect 34916 38853 34972 38855
rect 34705 38801 34755 38853
rect 34755 38801 34761 38853
rect 34916 38801 34935 38853
rect 34935 38801 34972 38853
rect 34705 38799 34761 38801
rect 34916 38799 34972 38801
rect 33055 38332 33111 38388
rect 33235 38332 33291 38388
rect 33817 38339 33873 38395
rect 33997 38339 34053 38395
rect 30852 37953 30908 37955
rect 30852 37901 30854 37953
rect 30854 37901 30906 37953
rect 30906 37901 30908 37953
rect 30852 37899 30908 37901
rect 31063 37953 31119 37955
rect 31063 37901 31065 37953
rect 31065 37901 31117 37953
rect 31117 37901 31119 37953
rect 31063 37899 31119 37901
rect 31274 37953 31330 37955
rect 31274 37901 31276 37953
rect 31276 37901 31328 37953
rect 31328 37901 31330 37953
rect 31274 37899 31330 37901
rect 31484 37953 31540 37955
rect 31484 37901 31486 37953
rect 31486 37901 31538 37953
rect 31538 37901 31540 37953
rect 31484 37899 31540 37901
rect 31695 37953 31751 37955
rect 31695 37901 31697 37953
rect 31697 37901 31749 37953
rect 31749 37901 31751 37953
rect 31695 37899 31751 37901
rect 31907 37953 31963 37955
rect 31907 37901 31909 37953
rect 31909 37901 31961 37953
rect 31961 37901 31963 37953
rect 31907 37899 31963 37901
rect 32118 37953 32174 37955
rect 32118 37901 32120 37953
rect 32120 37901 32172 37953
rect 32172 37901 32174 37953
rect 32118 37899 32174 37901
rect 32328 37953 32384 37955
rect 32328 37901 32330 37953
rect 32330 37901 32382 37953
rect 32382 37901 32384 37953
rect 32328 37899 32384 37901
rect 32539 37953 32595 37955
rect 32539 37901 32541 37953
rect 32541 37901 32593 37953
rect 32593 37901 32595 37953
rect 32539 37899 32595 37901
rect 32750 37953 32806 37955
rect 32750 37901 32752 37953
rect 32752 37901 32804 37953
rect 32804 37901 32806 37953
rect 32750 37899 32806 37901
rect 33055 37466 33111 37522
rect 33235 37466 33291 37522
rect 33817 37459 33873 37515
rect 33997 37459 34053 37515
rect 34282 36999 34338 37055
rect 34493 36999 34549 37055
rect 34705 37053 34761 37055
rect 34916 37053 34972 37055
rect 34705 37001 34755 37053
rect 34755 37001 34761 37053
rect 34916 37001 34935 37053
rect 34935 37001 34972 37053
rect 34705 36999 34761 37001
rect 34916 36999 34972 37001
rect 33055 36532 33111 36588
rect 33235 36532 33291 36588
rect 33817 36539 33873 36595
rect 33997 36539 34053 36595
rect 30852 36153 30908 36155
rect 30852 36101 30854 36153
rect 30854 36101 30906 36153
rect 30906 36101 30908 36153
rect 30852 36099 30908 36101
rect 31063 36153 31119 36155
rect 31063 36101 31065 36153
rect 31065 36101 31117 36153
rect 31117 36101 31119 36153
rect 31063 36099 31119 36101
rect 31274 36153 31330 36155
rect 31274 36101 31276 36153
rect 31276 36101 31328 36153
rect 31328 36101 31330 36153
rect 31274 36099 31330 36101
rect 31484 36153 31540 36155
rect 31484 36101 31486 36153
rect 31486 36101 31538 36153
rect 31538 36101 31540 36153
rect 31484 36099 31540 36101
rect 31695 36153 31751 36155
rect 31695 36101 31697 36153
rect 31697 36101 31749 36153
rect 31749 36101 31751 36153
rect 31695 36099 31751 36101
rect 31907 36153 31963 36155
rect 31907 36101 31909 36153
rect 31909 36101 31961 36153
rect 31961 36101 31963 36153
rect 31907 36099 31963 36101
rect 32118 36153 32174 36155
rect 32118 36101 32120 36153
rect 32120 36101 32172 36153
rect 32172 36101 32174 36153
rect 32118 36099 32174 36101
rect 32328 36153 32384 36155
rect 32328 36101 32330 36153
rect 32330 36101 32382 36153
rect 32382 36101 32384 36153
rect 32328 36099 32384 36101
rect 32539 36153 32595 36155
rect 32539 36101 32541 36153
rect 32541 36101 32593 36153
rect 32593 36101 32595 36153
rect 32539 36099 32595 36101
rect 32750 36153 32806 36155
rect 32750 36101 32752 36153
rect 32752 36101 32804 36153
rect 32804 36101 32806 36153
rect 32750 36099 32806 36101
rect 35218 43301 35220 43353
rect 35220 43301 35272 43353
rect 35272 43301 35274 43353
rect 35218 43299 35274 43301
rect 35428 43353 35484 43355
rect 35428 43301 35430 43353
rect 35430 43301 35482 43353
rect 35482 43301 35484 43353
rect 35428 43299 35484 43301
rect 35639 43353 35695 43355
rect 35639 43301 35641 43353
rect 35641 43301 35693 43353
rect 35693 43301 35695 43353
rect 35639 43299 35695 43301
rect 35851 43353 35907 43355
rect 35851 43301 35853 43353
rect 35853 43301 35905 43353
rect 35905 43301 35907 43353
rect 35851 43299 35907 43301
rect 36062 43353 36118 43355
rect 36062 43301 36064 43353
rect 36064 43301 36116 43353
rect 36116 43301 36118 43353
rect 36062 43299 36118 43301
rect 36272 43353 36328 43355
rect 36272 43301 36274 43353
rect 36274 43301 36326 43353
rect 36326 43301 36328 43353
rect 36272 43299 36328 43301
rect 36899 43716 36955 43772
rect 37110 43716 37166 43772
rect 37321 43716 37377 43772
rect 37532 43716 37588 43772
rect 40250 44206 40252 44255
rect 40252 44206 40304 44255
rect 40304 44206 40306 44255
rect 40250 44199 40306 44206
rect 40430 44206 40432 44255
rect 40432 44206 40484 44255
rect 40484 44206 40486 44255
rect 40430 44199 40486 44206
rect 41008 43770 41064 43772
rect 41008 43718 41010 43770
rect 41010 43718 41062 43770
rect 41062 43718 41064 43770
rect 41008 43716 41064 43718
rect 41219 43770 41275 43772
rect 41219 43718 41221 43770
rect 41221 43718 41273 43770
rect 41273 43718 41275 43770
rect 41219 43716 41275 43718
rect 41430 43770 41486 43772
rect 41430 43718 41432 43770
rect 41432 43718 41484 43770
rect 41484 43718 41486 43770
rect 41430 43716 41486 43718
rect 41641 43770 41697 43772
rect 41641 43718 41643 43770
rect 41643 43718 41695 43770
rect 41695 43718 41697 43770
rect 41641 43716 41697 43718
rect 41852 43770 41908 43772
rect 41852 43718 41854 43770
rect 41854 43718 41906 43770
rect 41906 43718 41908 43770
rect 41852 43716 41908 43718
rect 42062 43770 42118 43772
rect 42062 43718 42064 43770
rect 42064 43718 42116 43770
rect 42116 43718 42118 43770
rect 42062 43716 42118 43718
rect 42708 43709 42764 43765
rect 42919 43709 42975 43765
rect 43130 43709 43186 43765
rect 36676 42907 36732 42963
rect 39050 43353 39106 43355
rect 36676 41891 36732 41947
rect 37889 42676 37945 42732
rect 38069 42676 38125 42732
rect 38328 42399 38384 42455
rect 38539 42399 38595 42455
rect 38750 42399 38806 42455
rect 35218 41553 35274 41555
rect 35218 41501 35220 41553
rect 35220 41501 35272 41553
rect 35272 41501 35274 41553
rect 35218 41499 35274 41501
rect 35428 41553 35484 41555
rect 35428 41501 35430 41553
rect 35430 41501 35482 41553
rect 35482 41501 35484 41553
rect 35428 41499 35484 41501
rect 35639 41553 35695 41555
rect 35639 41501 35641 41553
rect 35641 41501 35693 41553
rect 35693 41501 35695 41553
rect 35639 41499 35695 41501
rect 35851 41553 35907 41555
rect 35851 41501 35853 41553
rect 35853 41501 35905 41553
rect 35905 41501 35907 41553
rect 35851 41499 35907 41501
rect 36062 41553 36118 41555
rect 36062 41501 36064 41553
rect 36064 41501 36116 41553
rect 36116 41501 36118 41553
rect 36062 41499 36118 41501
rect 36272 41553 36328 41555
rect 36272 41501 36274 41553
rect 36274 41501 36326 41553
rect 36326 41501 36328 41553
rect 36272 41499 36328 41501
rect 36676 41107 36732 41163
rect 37889 42122 37945 42178
rect 38069 42122 38125 42178
rect 36676 40091 36732 40147
rect 37889 40876 37945 40932
rect 38069 40876 38125 40932
rect 38328 40599 38384 40655
rect 38539 40599 38595 40655
rect 38750 40599 38806 40655
rect 35218 39753 35274 39755
rect 35218 39701 35220 39753
rect 35220 39701 35272 39753
rect 35272 39701 35274 39753
rect 35218 39699 35274 39701
rect 35428 39753 35484 39755
rect 35428 39701 35430 39753
rect 35430 39701 35482 39753
rect 35482 39701 35484 39753
rect 35428 39699 35484 39701
rect 35639 39753 35695 39755
rect 35639 39701 35641 39753
rect 35641 39701 35693 39753
rect 35693 39701 35695 39753
rect 35639 39699 35695 39701
rect 35851 39753 35907 39755
rect 35851 39701 35853 39753
rect 35853 39701 35905 39753
rect 35905 39701 35907 39753
rect 35851 39699 35907 39701
rect 36062 39753 36118 39755
rect 36062 39701 36064 39753
rect 36064 39701 36116 39753
rect 36116 39701 36118 39753
rect 36062 39699 36118 39701
rect 36272 39753 36328 39755
rect 36272 39701 36274 39753
rect 36274 39701 36326 39753
rect 36326 39701 36328 39753
rect 36272 39699 36328 39701
rect 36676 39307 36732 39363
rect 37889 40322 37945 40378
rect 38069 40322 38125 40378
rect 36676 38291 36732 38347
rect 37889 39076 37945 39132
rect 38069 39076 38125 39132
rect 38328 38799 38384 38855
rect 38539 38799 38595 38855
rect 38750 38799 38806 38855
rect 35218 37953 35274 37955
rect 35218 37901 35220 37953
rect 35220 37901 35272 37953
rect 35272 37901 35274 37953
rect 35218 37899 35274 37901
rect 35428 37953 35484 37955
rect 35428 37901 35430 37953
rect 35430 37901 35482 37953
rect 35482 37901 35484 37953
rect 35428 37899 35484 37901
rect 35639 37953 35695 37955
rect 35639 37901 35641 37953
rect 35641 37901 35693 37953
rect 35693 37901 35695 37953
rect 35639 37899 35695 37901
rect 35851 37953 35907 37955
rect 35851 37901 35853 37953
rect 35853 37901 35905 37953
rect 35905 37901 35907 37953
rect 35851 37899 35907 37901
rect 36062 37953 36118 37955
rect 36062 37901 36064 37953
rect 36064 37901 36116 37953
rect 36116 37901 36118 37953
rect 36062 37899 36118 37901
rect 36272 37953 36328 37955
rect 36272 37901 36274 37953
rect 36274 37901 36326 37953
rect 36326 37901 36328 37953
rect 36272 37899 36328 37901
rect 36676 37507 36732 37563
rect 37889 38522 37945 38578
rect 38069 38522 38125 38578
rect 37889 37276 37945 37332
rect 38069 37276 38125 37332
rect 38328 36999 38384 37055
rect 38539 36999 38595 37055
rect 38750 36999 38806 37055
rect 36676 36491 36732 36547
rect 35218 36153 35274 36155
rect 35218 36101 35220 36153
rect 35220 36101 35272 36153
rect 35272 36101 35274 36153
rect 35218 36099 35274 36101
rect 35428 36153 35484 36155
rect 35428 36101 35430 36153
rect 35430 36101 35482 36153
rect 35482 36101 35484 36153
rect 35428 36099 35484 36101
rect 35639 36153 35695 36155
rect 35639 36101 35641 36153
rect 35641 36101 35693 36153
rect 35693 36101 35695 36153
rect 35639 36099 35695 36101
rect 35851 36153 35907 36155
rect 35851 36101 35853 36153
rect 35853 36101 35905 36153
rect 35905 36101 35907 36153
rect 35851 36099 35907 36101
rect 36062 36153 36118 36155
rect 36062 36101 36064 36153
rect 36064 36101 36116 36153
rect 36116 36101 36118 36153
rect 36062 36099 36118 36101
rect 36272 36153 36328 36155
rect 36272 36101 36274 36153
rect 36274 36101 36326 36153
rect 36326 36101 36328 36153
rect 36272 36099 36328 36101
rect 37889 36722 37945 36778
rect 38069 36722 38125 36778
rect 39050 43301 39052 43353
rect 39052 43301 39104 43353
rect 39104 43301 39106 43353
rect 39050 43299 39106 43301
rect 39230 43353 39286 43355
rect 39230 43301 39232 43353
rect 39232 43301 39284 43353
rect 39284 43301 39286 43353
rect 39230 43299 39286 43301
rect 39773 42676 39829 42732
rect 39992 42907 40048 42963
rect 40777 43299 40833 43355
rect 40988 43299 41044 43355
rect 41199 43299 41255 43355
rect 40251 42399 40307 42455
rect 40431 42399 40487 42455
rect 39773 42122 39829 42178
rect 39992 41891 40048 41947
rect 39050 41553 39106 41555
rect 39050 41501 39052 41553
rect 39052 41501 39104 41553
rect 39104 41501 39106 41553
rect 39050 41499 39106 41501
rect 39230 41553 39286 41555
rect 39230 41501 39232 41553
rect 39232 41501 39284 41553
rect 39284 41501 39286 41553
rect 39230 41499 39286 41501
rect 39773 40876 39829 40932
rect 39992 41107 40048 41163
rect 40251 40599 40307 40655
rect 40431 40599 40487 40655
rect 39773 40322 39829 40378
rect 39992 40091 40048 40147
rect 39050 39753 39106 39755
rect 39050 39701 39052 39753
rect 39052 39701 39104 39753
rect 39104 39701 39106 39753
rect 39050 39699 39106 39701
rect 39230 39753 39286 39755
rect 39230 39701 39232 39753
rect 39232 39701 39284 39753
rect 39284 39701 39286 39753
rect 39230 39699 39286 39701
rect 39773 39076 39829 39132
rect 39992 39307 40048 39363
rect 40251 38799 40307 38855
rect 40431 38799 40487 38855
rect 39773 38522 39829 38578
rect 39992 38291 40048 38347
rect 39050 37953 39106 37955
rect 39050 37901 39052 37953
rect 39052 37901 39104 37953
rect 39104 37901 39106 37953
rect 39050 37899 39106 37901
rect 39230 37953 39286 37955
rect 39230 37901 39232 37953
rect 39232 37901 39284 37953
rect 39284 37901 39286 37953
rect 39230 37899 39286 37901
rect 39773 37276 39829 37332
rect 39992 37507 40048 37563
rect 40251 36999 40307 37055
rect 40431 36999 40487 37055
rect 39773 36722 39829 36778
rect 39992 36491 40048 36547
rect 39050 36153 39106 36155
rect 39050 36101 39052 36153
rect 39052 36101 39104 36153
rect 39104 36101 39106 36153
rect 39050 36099 39106 36101
rect 39230 36153 39286 36155
rect 39230 36101 39232 36153
rect 39232 36101 39284 36153
rect 39284 36101 39286 36153
rect 39230 36099 39286 36101
rect 36958 35825 37014 35881
rect 37169 35825 37225 35881
rect 37381 35825 37437 35881
rect 37592 35825 37648 35881
rect 27447 34938 27503 34940
rect 27447 34886 27449 34938
rect 27449 34886 27501 34938
rect 27501 34886 27503 34938
rect 27447 34884 27503 34886
rect 27571 34938 27627 34940
rect 27571 34886 27573 34938
rect 27573 34886 27625 34938
rect 27625 34886 27627 34938
rect 27571 34884 27627 34886
rect 27695 34938 27751 34940
rect 27695 34886 27697 34938
rect 27697 34886 27749 34938
rect 27749 34886 27751 34938
rect 27695 34884 27751 34886
rect 27447 34814 27503 34816
rect 27447 34762 27449 34814
rect 27449 34762 27501 34814
rect 27501 34762 27503 34814
rect 27447 34760 27503 34762
rect 27571 34814 27627 34816
rect 27571 34762 27573 34814
rect 27573 34762 27625 34814
rect 27625 34762 27627 34814
rect 27571 34760 27627 34762
rect 27695 34814 27751 34816
rect 27695 34762 27697 34814
rect 27697 34762 27749 34814
rect 27749 34762 27751 34814
rect 27695 34760 27751 34762
rect 27447 34690 27503 34692
rect 27447 34638 27449 34690
rect 27449 34638 27501 34690
rect 27501 34638 27503 34690
rect 27447 34636 27503 34638
rect 27571 34690 27627 34692
rect 27571 34638 27573 34690
rect 27573 34638 27625 34690
rect 27625 34638 27627 34690
rect 27571 34636 27627 34638
rect 27695 34690 27751 34692
rect 27695 34638 27697 34690
rect 27697 34638 27749 34690
rect 27749 34638 27751 34690
rect 27695 34636 27751 34638
rect 27447 34566 27503 34568
rect 27447 34514 27449 34566
rect 27449 34514 27501 34566
rect 27501 34514 27503 34566
rect 27447 34512 27503 34514
rect 27571 34566 27627 34568
rect 27571 34514 27573 34566
rect 27573 34514 27625 34566
rect 27625 34514 27627 34566
rect 27571 34512 27627 34514
rect 27695 34566 27751 34568
rect 27695 34514 27697 34566
rect 27697 34514 27749 34566
rect 27749 34514 27751 34566
rect 27695 34512 27751 34514
rect 43788 42399 43844 42455
rect 43999 42399 44055 42455
rect 44211 42399 44267 42455
rect 44422 42399 44478 42455
rect 43788 40599 43844 40655
rect 43999 40599 44055 40655
rect 44211 40599 44267 40655
rect 44422 40599 44478 40655
rect 43788 38799 43844 38855
rect 43999 38799 44055 38855
rect 44211 38799 44267 38855
rect 44422 38799 44478 38855
rect 43788 36999 43844 37055
rect 43999 36999 44055 37055
rect 44211 36999 44267 37055
rect 44422 36999 44478 37055
rect 44832 43353 44888 43355
rect 44832 43301 44834 43353
rect 44834 43301 44886 43353
rect 44886 43301 44888 43353
rect 44832 43299 44888 43301
rect 45043 43353 45099 43355
rect 45043 43301 45045 43353
rect 45045 43301 45097 43353
rect 45097 43301 45099 43353
rect 45043 43299 45099 43301
rect 45254 43353 45310 43355
rect 45254 43301 45256 43353
rect 45256 43301 45308 43353
rect 45308 43301 45310 43353
rect 45254 43299 45310 43301
rect 44832 41553 44888 41555
rect 44832 41501 44834 41553
rect 44834 41501 44886 41553
rect 44886 41501 44888 41553
rect 44832 41499 44888 41501
rect 45043 41553 45099 41555
rect 45043 41501 45045 41553
rect 45045 41501 45097 41553
rect 45097 41501 45099 41553
rect 45043 41499 45099 41501
rect 45254 41553 45310 41555
rect 45254 41501 45256 41553
rect 45256 41501 45308 41553
rect 45308 41501 45310 41553
rect 45254 41499 45310 41501
rect 44832 39753 44888 39755
rect 44832 39701 44834 39753
rect 44834 39701 44886 39753
rect 44886 39701 44888 39753
rect 44832 39699 44888 39701
rect 45043 39753 45099 39755
rect 45043 39701 45045 39753
rect 45045 39701 45097 39753
rect 45097 39701 45099 39753
rect 45043 39699 45099 39701
rect 45254 39753 45310 39755
rect 45254 39701 45256 39753
rect 45256 39701 45308 39753
rect 45308 39701 45310 39753
rect 45254 39699 45310 39701
rect 44832 37953 44888 37955
rect 44832 37901 44834 37953
rect 44834 37901 44886 37953
rect 44886 37901 44888 37953
rect 44832 37899 44888 37901
rect 45043 37953 45099 37955
rect 45043 37901 45045 37953
rect 45045 37901 45097 37953
rect 45097 37901 45099 37953
rect 45043 37899 45099 37901
rect 45254 37953 45310 37955
rect 45254 37901 45256 37953
rect 45256 37901 45308 37953
rect 45308 37901 45310 37953
rect 45254 37899 45310 37901
rect 44832 36153 44888 36155
rect 44832 36101 44834 36153
rect 44834 36101 44886 36153
rect 44886 36101 44888 36153
rect 44832 36099 44888 36101
rect 45043 36153 45099 36155
rect 45043 36101 45045 36153
rect 45045 36101 45097 36153
rect 45097 36101 45099 36153
rect 45043 36099 45099 36101
rect 45254 36153 45310 36155
rect 45254 36101 45256 36153
rect 45256 36101 45308 36153
rect 45308 36101 45310 36153
rect 45254 36099 45310 36101
rect 50135 44253 50191 44255
rect 50135 44201 50137 44253
rect 50137 44201 50189 44253
rect 50189 44201 50191 44253
rect 50135 44199 50191 44201
rect 50346 44253 50402 44255
rect 50346 44201 50348 44253
rect 50348 44201 50400 44253
rect 50400 44201 50402 44253
rect 50346 44199 50402 44201
rect 50557 44253 50613 44255
rect 50557 44201 50559 44253
rect 50559 44201 50611 44253
rect 50611 44201 50613 44253
rect 50557 44199 50613 44201
rect 50768 44253 50824 44255
rect 50768 44201 50770 44253
rect 50770 44201 50822 44253
rect 50822 44201 50824 44253
rect 50768 44199 50824 44201
rect 48836 43353 48892 43355
rect 48836 43301 48838 43353
rect 48838 43301 48890 43353
rect 48890 43301 48892 43353
rect 48836 43299 48892 43301
rect 49046 43353 49102 43355
rect 49046 43301 49048 43353
rect 49048 43301 49100 43353
rect 49100 43301 49102 43353
rect 49046 43299 49102 43301
rect 49257 43353 49313 43355
rect 49257 43301 49259 43353
rect 49259 43301 49311 43353
rect 49311 43301 49313 43353
rect 49257 43299 49313 43301
rect 49469 43353 49525 43355
rect 49469 43301 49471 43353
rect 49471 43301 49523 43353
rect 49523 43301 49525 43353
rect 49469 43299 49525 43301
rect 49680 43353 49736 43355
rect 49680 43301 49682 43353
rect 49682 43301 49734 43353
rect 49734 43301 49736 43353
rect 49680 43299 49736 43301
rect 49890 43353 49946 43355
rect 49890 43301 49892 43353
rect 49892 43301 49944 43353
rect 49944 43301 49946 43353
rect 49890 43299 49946 43301
rect 51079 43770 51135 43772
rect 51079 43718 51081 43770
rect 51081 43718 51133 43770
rect 51133 43718 51135 43770
rect 51079 43716 51135 43718
rect 51290 43770 51346 43772
rect 51290 43718 51292 43770
rect 51292 43718 51344 43770
rect 51344 43718 51346 43770
rect 51290 43716 51346 43718
rect 51501 43770 51557 43772
rect 51501 43718 51503 43770
rect 51503 43718 51555 43770
rect 51555 43718 51557 43770
rect 51501 43716 51557 43718
rect 51712 43770 51768 43772
rect 51712 43718 51714 43770
rect 51714 43718 51766 43770
rect 51766 43718 51768 43770
rect 51712 43716 51768 43718
rect 51923 43770 51979 43772
rect 51923 43718 51925 43770
rect 51925 43718 51977 43770
rect 51977 43718 51979 43770
rect 51923 43716 51979 43718
rect 48594 42947 48650 42949
rect 48594 42895 48596 42947
rect 48596 42895 48648 42947
rect 48648 42895 48650 42947
rect 48594 42893 48650 42895
rect 48594 42729 48650 42731
rect 48594 42677 48596 42729
rect 48596 42677 48648 42729
rect 48648 42677 48650 42729
rect 48594 42675 48650 42677
rect 48594 42177 48650 42179
rect 48594 42125 48596 42177
rect 48596 42125 48648 42177
rect 48648 42125 48650 42177
rect 48594 42123 48650 42125
rect 48594 41959 48650 41961
rect 48594 41907 48596 41959
rect 48596 41907 48648 41959
rect 48648 41907 48650 41959
rect 48594 41905 48650 41907
rect 48836 41553 48892 41555
rect 48836 41501 48838 41553
rect 48838 41501 48890 41553
rect 48890 41501 48892 41553
rect 48836 41499 48892 41501
rect 49046 41553 49102 41555
rect 49046 41501 49048 41553
rect 49048 41501 49100 41553
rect 49100 41501 49102 41553
rect 49046 41499 49102 41501
rect 49257 41553 49313 41555
rect 49257 41501 49259 41553
rect 49259 41501 49311 41553
rect 49311 41501 49313 41553
rect 49257 41499 49313 41501
rect 49469 41553 49525 41555
rect 49469 41501 49471 41553
rect 49471 41501 49523 41553
rect 49523 41501 49525 41553
rect 49469 41499 49525 41501
rect 49680 41553 49736 41555
rect 49680 41501 49682 41553
rect 49682 41501 49734 41553
rect 49734 41501 49736 41553
rect 49680 41499 49736 41501
rect 49890 41553 49946 41555
rect 49890 41501 49892 41553
rect 49892 41501 49944 41553
rect 49944 41501 49946 41553
rect 49890 41499 49946 41501
rect 48594 41147 48650 41149
rect 48594 41095 48596 41147
rect 48596 41095 48648 41147
rect 48648 41095 48650 41147
rect 48594 41093 48650 41095
rect 48594 40929 48650 40931
rect 48594 40877 48596 40929
rect 48596 40877 48648 40929
rect 48648 40877 48650 40929
rect 48594 40875 48650 40877
rect 48594 40377 48650 40379
rect 48594 40325 48596 40377
rect 48596 40325 48648 40377
rect 48648 40325 48650 40377
rect 48594 40323 48650 40325
rect 48594 40159 48650 40161
rect 48594 40107 48596 40159
rect 48596 40107 48648 40159
rect 48648 40107 48650 40159
rect 48594 40105 48650 40107
rect 48836 39753 48892 39755
rect 48836 39701 48838 39753
rect 48838 39701 48890 39753
rect 48890 39701 48892 39753
rect 48836 39699 48892 39701
rect 49046 39753 49102 39755
rect 49046 39701 49048 39753
rect 49048 39701 49100 39753
rect 49100 39701 49102 39753
rect 49046 39699 49102 39701
rect 49257 39753 49313 39755
rect 49257 39701 49259 39753
rect 49259 39701 49311 39753
rect 49311 39701 49313 39753
rect 49257 39699 49313 39701
rect 49469 39753 49525 39755
rect 49469 39701 49471 39753
rect 49471 39701 49523 39753
rect 49523 39701 49525 39753
rect 49469 39699 49525 39701
rect 49680 39753 49736 39755
rect 49680 39701 49682 39753
rect 49682 39701 49734 39753
rect 49734 39701 49736 39753
rect 49680 39699 49736 39701
rect 49890 39753 49946 39755
rect 49890 39701 49892 39753
rect 49892 39701 49944 39753
rect 49944 39701 49946 39753
rect 49890 39699 49946 39701
rect 48594 39347 48650 39349
rect 48594 39295 48596 39347
rect 48596 39295 48648 39347
rect 48648 39295 48650 39347
rect 48594 39293 48650 39295
rect 48594 39129 48650 39131
rect 48594 39077 48596 39129
rect 48596 39077 48648 39129
rect 48648 39077 48650 39129
rect 48594 39075 48650 39077
rect 48594 38577 48650 38579
rect 48594 38525 48596 38577
rect 48596 38525 48648 38577
rect 48648 38525 48650 38577
rect 48594 38523 48650 38525
rect 48594 38359 48650 38361
rect 48594 38307 48596 38359
rect 48596 38307 48648 38359
rect 48648 38307 48650 38359
rect 48594 38305 48650 38307
rect 48836 37953 48892 37955
rect 48836 37901 48838 37953
rect 48838 37901 48890 37953
rect 48890 37901 48892 37953
rect 48836 37899 48892 37901
rect 49046 37953 49102 37955
rect 49046 37901 49048 37953
rect 49048 37901 49100 37953
rect 49100 37901 49102 37953
rect 49046 37899 49102 37901
rect 49257 37953 49313 37955
rect 49257 37901 49259 37953
rect 49259 37901 49311 37953
rect 49311 37901 49313 37953
rect 49257 37899 49313 37901
rect 49469 37953 49525 37955
rect 49469 37901 49471 37953
rect 49471 37901 49523 37953
rect 49523 37901 49525 37953
rect 49469 37899 49525 37901
rect 49680 37953 49736 37955
rect 49680 37901 49682 37953
rect 49682 37901 49734 37953
rect 49734 37901 49736 37953
rect 49680 37899 49736 37901
rect 49890 37953 49946 37955
rect 49890 37901 49892 37953
rect 49892 37901 49944 37953
rect 49944 37901 49946 37953
rect 49890 37899 49946 37901
rect 48594 37547 48650 37549
rect 48594 37495 48596 37547
rect 48596 37495 48648 37547
rect 48648 37495 48650 37547
rect 48594 37493 48650 37495
rect 48594 37329 48650 37331
rect 48594 37277 48596 37329
rect 48596 37277 48648 37329
rect 48648 37277 48650 37329
rect 48594 37275 48650 37277
rect 48594 36777 48650 36779
rect 48594 36725 48596 36777
rect 48596 36725 48648 36777
rect 48648 36725 48650 36777
rect 48594 36723 48650 36725
rect 48594 36559 48650 36561
rect 48594 36507 48596 36559
rect 48596 36507 48648 36559
rect 48648 36507 48650 36559
rect 48594 36505 48650 36507
rect 48836 36153 48892 36155
rect 48836 36101 48838 36153
rect 48838 36101 48890 36153
rect 48890 36101 48892 36153
rect 48836 36099 48892 36101
rect 49046 36153 49102 36155
rect 49046 36101 49048 36153
rect 49048 36101 49100 36153
rect 49100 36101 49102 36153
rect 49046 36099 49102 36101
rect 49257 36153 49313 36155
rect 49257 36101 49259 36153
rect 49259 36101 49311 36153
rect 49311 36101 49313 36153
rect 49257 36099 49313 36101
rect 49469 36153 49525 36155
rect 49469 36101 49471 36153
rect 49471 36101 49523 36153
rect 49523 36101 49525 36153
rect 49469 36099 49525 36101
rect 49680 36153 49736 36155
rect 49680 36101 49682 36153
rect 49682 36101 49734 36153
rect 49734 36101 49736 36153
rect 49680 36099 49736 36101
rect 49890 36153 49946 36155
rect 49890 36101 49892 36153
rect 49892 36101 49944 36153
rect 49944 36101 49946 36153
rect 49890 36099 49946 36101
rect 52314 43353 52370 43355
rect 52314 43301 52316 43353
rect 52316 43301 52368 43353
rect 52368 43301 52370 43353
rect 52314 43299 52370 43301
rect 52525 43353 52581 43355
rect 52525 43301 52527 43353
rect 52527 43301 52579 43353
rect 52579 43301 52581 43353
rect 52525 43299 52581 43301
rect 52736 43353 52792 43355
rect 52736 43301 52738 43353
rect 52738 43301 52790 43353
rect 52790 43301 52792 43353
rect 52736 43299 52792 43301
rect 52946 43353 53002 43355
rect 52946 43301 52948 43353
rect 52948 43301 53000 43353
rect 53000 43301 53002 43353
rect 52946 43299 53002 43301
rect 53157 43353 53213 43355
rect 53157 43301 53159 43353
rect 53159 43301 53211 43353
rect 53211 43301 53213 43353
rect 53157 43299 53213 43301
rect 53369 43353 53425 43355
rect 53369 43301 53371 43353
rect 53371 43301 53423 43353
rect 53423 43301 53425 43353
rect 53369 43299 53425 43301
rect 53580 43353 53636 43355
rect 53580 43301 53582 43353
rect 53582 43301 53634 43353
rect 53634 43301 53636 43353
rect 53580 43299 53636 43301
rect 53790 43353 53846 43355
rect 53790 43301 53792 43353
rect 53792 43301 53844 43353
rect 53844 43301 53846 43353
rect 53790 43299 53846 43301
rect 54001 43353 54057 43355
rect 54001 43301 54003 43353
rect 54003 43301 54055 43353
rect 54055 43301 54057 43353
rect 54001 43299 54057 43301
rect 54212 43353 54268 43355
rect 54212 43301 54214 43353
rect 54214 43301 54266 43353
rect 54266 43301 54268 43353
rect 54212 43299 54268 43301
rect 51071 42859 51127 42915
rect 51251 42859 51307 42915
rect 51833 42859 51889 42915
rect 52013 42859 52069 42915
rect 50161 42453 50217 42455
rect 50161 42401 50190 42453
rect 50190 42401 50217 42453
rect 50161 42399 50217 42401
rect 50372 42399 50428 42455
rect 50584 42399 50640 42455
rect 50795 42399 50851 42455
rect 51071 41939 51127 41995
rect 51251 41939 51307 41995
rect 51833 41939 51889 41995
rect 52013 41939 52069 41995
rect 52314 41553 52370 41555
rect 52314 41501 52316 41553
rect 52316 41501 52368 41553
rect 52368 41501 52370 41553
rect 52314 41499 52370 41501
rect 52525 41553 52581 41555
rect 52525 41501 52527 41553
rect 52527 41501 52579 41553
rect 52579 41501 52581 41553
rect 52525 41499 52581 41501
rect 52736 41553 52792 41555
rect 52736 41501 52738 41553
rect 52738 41501 52790 41553
rect 52790 41501 52792 41553
rect 52736 41499 52792 41501
rect 52946 41553 53002 41555
rect 52946 41501 52948 41553
rect 52948 41501 53000 41553
rect 53000 41501 53002 41553
rect 52946 41499 53002 41501
rect 53157 41553 53213 41555
rect 53157 41501 53159 41553
rect 53159 41501 53211 41553
rect 53211 41501 53213 41553
rect 53157 41499 53213 41501
rect 53369 41553 53425 41555
rect 53369 41501 53371 41553
rect 53371 41501 53423 41553
rect 53423 41501 53425 41553
rect 53369 41499 53425 41501
rect 53580 41553 53636 41555
rect 53580 41501 53582 41553
rect 53582 41501 53634 41553
rect 53634 41501 53636 41553
rect 53580 41499 53636 41501
rect 53790 41553 53846 41555
rect 53790 41501 53792 41553
rect 53792 41501 53844 41553
rect 53844 41501 53846 41553
rect 53790 41499 53846 41501
rect 54001 41553 54057 41555
rect 54001 41501 54003 41553
rect 54003 41501 54055 41553
rect 54055 41501 54057 41553
rect 54001 41499 54057 41501
rect 54212 41553 54268 41555
rect 54212 41501 54214 41553
rect 54214 41501 54266 41553
rect 54266 41501 54268 41553
rect 54212 41499 54268 41501
rect 51071 41059 51127 41115
rect 51251 41059 51307 41115
rect 51833 41059 51889 41115
rect 52013 41059 52069 41115
rect 50161 40653 50217 40655
rect 50161 40601 50190 40653
rect 50190 40601 50217 40653
rect 50161 40599 50217 40601
rect 50372 40599 50428 40655
rect 50584 40599 50640 40655
rect 50795 40599 50851 40655
rect 51071 40139 51127 40195
rect 51251 40139 51307 40195
rect 51833 40139 51889 40195
rect 52013 40139 52069 40195
rect 52314 39753 52370 39755
rect 52314 39701 52316 39753
rect 52316 39701 52368 39753
rect 52368 39701 52370 39753
rect 52314 39699 52370 39701
rect 52525 39753 52581 39755
rect 52525 39701 52527 39753
rect 52527 39701 52579 39753
rect 52579 39701 52581 39753
rect 52525 39699 52581 39701
rect 52736 39753 52792 39755
rect 52736 39701 52738 39753
rect 52738 39701 52790 39753
rect 52790 39701 52792 39753
rect 52736 39699 52792 39701
rect 52946 39753 53002 39755
rect 52946 39701 52948 39753
rect 52948 39701 53000 39753
rect 53000 39701 53002 39753
rect 52946 39699 53002 39701
rect 53157 39753 53213 39755
rect 53157 39701 53159 39753
rect 53159 39701 53211 39753
rect 53211 39701 53213 39753
rect 53157 39699 53213 39701
rect 53369 39753 53425 39755
rect 53369 39701 53371 39753
rect 53371 39701 53423 39753
rect 53423 39701 53425 39753
rect 53369 39699 53425 39701
rect 53580 39753 53636 39755
rect 53580 39701 53582 39753
rect 53582 39701 53634 39753
rect 53634 39701 53636 39753
rect 53580 39699 53636 39701
rect 53790 39753 53846 39755
rect 53790 39701 53792 39753
rect 53792 39701 53844 39753
rect 53844 39701 53846 39753
rect 53790 39699 53846 39701
rect 54001 39753 54057 39755
rect 54001 39701 54003 39753
rect 54003 39701 54055 39753
rect 54055 39701 54057 39753
rect 54001 39699 54057 39701
rect 54212 39753 54268 39755
rect 54212 39701 54214 39753
rect 54214 39701 54266 39753
rect 54266 39701 54268 39753
rect 54212 39699 54268 39701
rect 51071 39259 51127 39315
rect 51251 39259 51307 39315
rect 51833 39259 51889 39315
rect 52013 39259 52069 39315
rect 50161 38853 50217 38855
rect 50161 38801 50190 38853
rect 50190 38801 50217 38853
rect 50161 38799 50217 38801
rect 50372 38799 50428 38855
rect 50584 38799 50640 38855
rect 50795 38799 50851 38855
rect 51071 38339 51127 38395
rect 51251 38339 51307 38395
rect 51833 38339 51889 38395
rect 52013 38339 52069 38395
rect 52314 37953 52370 37955
rect 52314 37901 52316 37953
rect 52316 37901 52368 37953
rect 52368 37901 52370 37953
rect 52314 37899 52370 37901
rect 52525 37953 52581 37955
rect 52525 37901 52527 37953
rect 52527 37901 52579 37953
rect 52579 37901 52581 37953
rect 52525 37899 52581 37901
rect 52736 37953 52792 37955
rect 52736 37901 52738 37953
rect 52738 37901 52790 37953
rect 52790 37901 52792 37953
rect 52736 37899 52792 37901
rect 52946 37953 53002 37955
rect 52946 37901 52948 37953
rect 52948 37901 53000 37953
rect 53000 37901 53002 37953
rect 52946 37899 53002 37901
rect 53157 37953 53213 37955
rect 53157 37901 53159 37953
rect 53159 37901 53211 37953
rect 53211 37901 53213 37953
rect 53157 37899 53213 37901
rect 53369 37953 53425 37955
rect 53369 37901 53371 37953
rect 53371 37901 53423 37953
rect 53423 37901 53425 37953
rect 53369 37899 53425 37901
rect 53580 37953 53636 37955
rect 53580 37901 53582 37953
rect 53582 37901 53634 37953
rect 53634 37901 53636 37953
rect 53580 37899 53636 37901
rect 53790 37953 53846 37955
rect 53790 37901 53792 37953
rect 53792 37901 53844 37953
rect 53844 37901 53846 37953
rect 53790 37899 53846 37901
rect 54001 37953 54057 37955
rect 54001 37901 54003 37953
rect 54003 37901 54055 37953
rect 54055 37901 54057 37953
rect 54001 37899 54057 37901
rect 54212 37953 54268 37955
rect 54212 37901 54214 37953
rect 54214 37901 54266 37953
rect 54266 37901 54268 37953
rect 54212 37899 54268 37901
rect 51071 37459 51127 37515
rect 51251 37459 51307 37515
rect 51833 37459 51889 37515
rect 52013 37459 52069 37515
rect 50161 37053 50217 37055
rect 50161 37001 50190 37053
rect 50190 37001 50217 37053
rect 50161 36999 50217 37001
rect 50372 36999 50428 37055
rect 50584 36999 50640 37055
rect 50795 36999 50851 37055
rect 51071 36539 51127 36595
rect 51251 36539 51307 36595
rect 51833 36539 51889 36595
rect 52013 36539 52069 36595
rect 52314 36153 52370 36155
rect 52314 36101 52316 36153
rect 52316 36101 52368 36153
rect 52368 36101 52370 36153
rect 52314 36099 52370 36101
rect 52525 36153 52581 36155
rect 52525 36101 52527 36153
rect 52527 36101 52579 36153
rect 52579 36101 52581 36153
rect 52525 36099 52581 36101
rect 52736 36153 52792 36155
rect 52736 36101 52738 36153
rect 52738 36101 52790 36153
rect 52790 36101 52792 36153
rect 52736 36099 52792 36101
rect 52946 36153 53002 36155
rect 52946 36101 52948 36153
rect 52948 36101 53000 36153
rect 53000 36101 53002 36153
rect 52946 36099 53002 36101
rect 53157 36153 53213 36155
rect 53157 36101 53159 36153
rect 53159 36101 53211 36153
rect 53211 36101 53213 36153
rect 53157 36099 53213 36101
rect 53369 36153 53425 36155
rect 53369 36101 53371 36153
rect 53371 36101 53423 36153
rect 53423 36101 53425 36153
rect 53369 36099 53425 36101
rect 53580 36153 53636 36155
rect 53580 36101 53582 36153
rect 53582 36101 53634 36153
rect 53634 36101 53636 36153
rect 53580 36099 53636 36101
rect 53790 36153 53846 36155
rect 53790 36101 53792 36153
rect 53792 36101 53844 36153
rect 53844 36101 53846 36153
rect 53790 36099 53846 36101
rect 54001 36153 54057 36155
rect 54001 36101 54003 36153
rect 54003 36101 54055 36153
rect 54055 36101 54057 36153
rect 54001 36099 54057 36101
rect 54212 36153 54268 36155
rect 54212 36101 54214 36153
rect 54214 36101 54266 36153
rect 54266 36101 54268 36153
rect 54212 36099 54268 36101
rect 56013 44253 56069 44255
rect 56013 44201 56015 44253
rect 56015 44201 56067 44253
rect 56067 44201 56069 44253
rect 56013 44199 56069 44201
rect 56224 44253 56280 44255
rect 56224 44201 56226 44253
rect 56226 44201 56278 44253
rect 56278 44201 56280 44253
rect 56224 44199 56280 44201
rect 56435 44253 56491 44255
rect 56435 44201 56437 44253
rect 56437 44201 56489 44253
rect 56489 44201 56491 44253
rect 56435 44199 56491 44201
rect 56646 44253 56702 44255
rect 56646 44201 56648 44253
rect 56648 44201 56700 44253
rect 56700 44201 56702 44253
rect 56646 44199 56702 44201
rect 56857 44253 56913 44255
rect 56857 44201 56859 44253
rect 56859 44201 56911 44253
rect 56911 44201 56913 44253
rect 56857 44199 56913 44201
rect 57068 44253 57124 44255
rect 57068 44201 57070 44253
rect 57070 44201 57122 44253
rect 57122 44201 57124 44253
rect 57068 44199 57124 44201
rect 57279 44253 57335 44255
rect 57279 44201 57281 44253
rect 57281 44201 57333 44253
rect 57333 44201 57335 44253
rect 57279 44199 57335 44201
rect 54853 43353 54909 43355
rect 54853 43301 54855 43353
rect 54855 43301 54907 43353
rect 54907 43301 54909 43353
rect 54853 43299 54909 43301
rect 55064 43353 55120 43355
rect 55064 43301 55066 43353
rect 55066 43301 55118 43353
rect 55118 43301 55120 43353
rect 55064 43299 55120 43301
rect 55276 43353 55332 43355
rect 55276 43301 55278 43353
rect 55278 43301 55330 43353
rect 55330 43301 55332 43353
rect 55276 43299 55332 43301
rect 55487 43353 55543 43355
rect 55487 43301 55489 43353
rect 55489 43301 55541 43353
rect 55541 43301 55543 43353
rect 55487 43299 55543 43301
rect 56013 42453 56069 42455
rect 56013 42401 56015 42453
rect 56015 42401 56067 42453
rect 56067 42401 56069 42453
rect 56013 42399 56069 42401
rect 56224 42453 56280 42455
rect 56224 42401 56226 42453
rect 56226 42401 56278 42453
rect 56278 42401 56280 42453
rect 56224 42399 56280 42401
rect 56435 42453 56491 42455
rect 56435 42401 56437 42453
rect 56437 42401 56489 42453
rect 56489 42401 56491 42453
rect 56435 42399 56491 42401
rect 56646 42453 56702 42455
rect 56646 42401 56648 42453
rect 56648 42401 56700 42453
rect 56700 42401 56702 42453
rect 56646 42399 56702 42401
rect 56857 42453 56913 42455
rect 56857 42401 56859 42453
rect 56859 42401 56911 42453
rect 56911 42401 56913 42453
rect 56857 42399 56913 42401
rect 57068 42453 57124 42455
rect 57068 42401 57070 42453
rect 57070 42401 57122 42453
rect 57122 42401 57124 42453
rect 57068 42399 57124 42401
rect 57279 42453 57335 42455
rect 57279 42401 57281 42453
rect 57281 42401 57333 42453
rect 57333 42401 57335 42453
rect 57279 42399 57335 42401
rect 54853 41553 54909 41555
rect 54853 41501 54855 41553
rect 54855 41501 54907 41553
rect 54907 41501 54909 41553
rect 54853 41499 54909 41501
rect 55064 41553 55120 41555
rect 55064 41501 55066 41553
rect 55066 41501 55118 41553
rect 55118 41501 55120 41553
rect 55064 41499 55120 41501
rect 55276 41553 55332 41555
rect 55276 41501 55278 41553
rect 55278 41501 55330 41553
rect 55330 41501 55332 41553
rect 55276 41499 55332 41501
rect 55487 41553 55543 41555
rect 55487 41501 55489 41553
rect 55489 41501 55541 41553
rect 55541 41501 55543 41553
rect 55487 41499 55543 41501
rect 56013 40653 56069 40655
rect 56013 40601 56015 40653
rect 56015 40601 56067 40653
rect 56067 40601 56069 40653
rect 56013 40599 56069 40601
rect 56224 40653 56280 40655
rect 56224 40601 56226 40653
rect 56226 40601 56278 40653
rect 56278 40601 56280 40653
rect 56224 40599 56280 40601
rect 56435 40653 56491 40655
rect 56435 40601 56437 40653
rect 56437 40601 56489 40653
rect 56489 40601 56491 40653
rect 56435 40599 56491 40601
rect 56646 40653 56702 40655
rect 56646 40601 56648 40653
rect 56648 40601 56700 40653
rect 56700 40601 56702 40653
rect 56646 40599 56702 40601
rect 56857 40653 56913 40655
rect 56857 40601 56859 40653
rect 56859 40601 56911 40653
rect 56911 40601 56913 40653
rect 56857 40599 56913 40601
rect 57068 40653 57124 40655
rect 57068 40601 57070 40653
rect 57070 40601 57122 40653
rect 57122 40601 57124 40653
rect 57068 40599 57124 40601
rect 57279 40653 57335 40655
rect 57279 40601 57281 40653
rect 57281 40601 57333 40653
rect 57333 40601 57335 40653
rect 57279 40599 57335 40601
rect 54853 39753 54909 39755
rect 54853 39701 54855 39753
rect 54855 39701 54907 39753
rect 54907 39701 54909 39753
rect 54853 39699 54909 39701
rect 55064 39753 55120 39755
rect 55064 39701 55066 39753
rect 55066 39701 55118 39753
rect 55118 39701 55120 39753
rect 55064 39699 55120 39701
rect 55276 39753 55332 39755
rect 55276 39701 55278 39753
rect 55278 39701 55330 39753
rect 55330 39701 55332 39753
rect 55276 39699 55332 39701
rect 55487 39753 55543 39755
rect 55487 39701 55489 39753
rect 55489 39701 55541 39753
rect 55541 39701 55543 39753
rect 55487 39699 55543 39701
rect 56013 38853 56069 38855
rect 56013 38801 56015 38853
rect 56015 38801 56067 38853
rect 56067 38801 56069 38853
rect 56013 38799 56069 38801
rect 56224 38853 56280 38855
rect 56224 38801 56226 38853
rect 56226 38801 56278 38853
rect 56278 38801 56280 38853
rect 56224 38799 56280 38801
rect 56435 38853 56491 38855
rect 56435 38801 56437 38853
rect 56437 38801 56489 38853
rect 56489 38801 56491 38853
rect 56435 38799 56491 38801
rect 56646 38853 56702 38855
rect 56646 38801 56648 38853
rect 56648 38801 56700 38853
rect 56700 38801 56702 38853
rect 56646 38799 56702 38801
rect 56857 38853 56913 38855
rect 56857 38801 56859 38853
rect 56859 38801 56911 38853
rect 56911 38801 56913 38853
rect 56857 38799 56913 38801
rect 57068 38853 57124 38855
rect 57068 38801 57070 38853
rect 57070 38801 57122 38853
rect 57122 38801 57124 38853
rect 57068 38799 57124 38801
rect 57279 38853 57335 38855
rect 57279 38801 57281 38853
rect 57281 38801 57333 38853
rect 57333 38801 57335 38853
rect 57279 38799 57335 38801
rect 54853 37953 54909 37955
rect 54853 37901 54855 37953
rect 54855 37901 54907 37953
rect 54907 37901 54909 37953
rect 54853 37899 54909 37901
rect 55064 37953 55120 37955
rect 55064 37901 55066 37953
rect 55066 37901 55118 37953
rect 55118 37901 55120 37953
rect 55064 37899 55120 37901
rect 55276 37953 55332 37955
rect 55276 37901 55278 37953
rect 55278 37901 55330 37953
rect 55330 37901 55332 37953
rect 55276 37899 55332 37901
rect 55487 37953 55543 37955
rect 55487 37901 55489 37953
rect 55489 37901 55541 37953
rect 55541 37901 55543 37953
rect 55487 37899 55543 37901
rect 56013 37053 56069 37055
rect 56013 37001 56015 37053
rect 56015 37001 56067 37053
rect 56067 37001 56069 37053
rect 56013 36999 56069 37001
rect 56224 37053 56280 37055
rect 56224 37001 56226 37053
rect 56226 37001 56278 37053
rect 56278 37001 56280 37053
rect 56224 36999 56280 37001
rect 56435 37053 56491 37055
rect 56435 37001 56437 37053
rect 56437 37001 56489 37053
rect 56489 37001 56491 37053
rect 56435 36999 56491 37001
rect 56646 37053 56702 37055
rect 56646 37001 56648 37053
rect 56648 37001 56700 37053
rect 56700 37001 56702 37053
rect 56646 36999 56702 37001
rect 56857 37053 56913 37055
rect 56857 37001 56859 37053
rect 56859 37001 56911 37053
rect 56911 37001 56913 37053
rect 56857 36999 56913 37001
rect 57068 37053 57124 37055
rect 57068 37001 57070 37053
rect 57070 37001 57122 37053
rect 57122 37001 57124 37053
rect 57068 36999 57124 37001
rect 57279 37053 57335 37055
rect 57279 37001 57281 37053
rect 57281 37001 57333 37053
rect 57333 37001 57335 37053
rect 57279 36999 57335 37001
rect 54853 36153 54909 36155
rect 54853 36101 54855 36153
rect 54855 36101 54907 36153
rect 54907 36101 54909 36153
rect 54853 36099 54909 36101
rect 55064 36153 55120 36155
rect 55064 36101 55066 36153
rect 55066 36101 55118 36153
rect 55118 36101 55120 36153
rect 55064 36099 55120 36101
rect 55276 36153 55332 36155
rect 55276 36101 55278 36153
rect 55278 36101 55330 36153
rect 55330 36101 55332 36153
rect 55276 36099 55332 36101
rect 55487 36153 55543 36155
rect 55487 36101 55489 36153
rect 55489 36101 55541 36153
rect 55541 36101 55543 36153
rect 55487 36099 55543 36101
rect 27474 33085 27530 33141
rect 27686 33085 27742 33141
rect 27474 32867 27530 32923
rect 27686 32867 27742 32923
rect 27474 32649 27530 32705
rect 27686 32649 27742 32705
rect 27474 32431 27530 32487
rect 27686 32431 27742 32487
rect 27474 31204 27476 31252
rect 27476 31204 27528 31252
rect 27528 31204 27530 31252
rect 27474 31196 27530 31204
rect 27686 31204 27688 31252
rect 27688 31204 27740 31252
rect 27740 31204 27742 31252
rect 27686 31196 27742 31204
rect 27474 30986 27476 31034
rect 27476 30986 27528 31034
rect 27528 30986 27530 31034
rect 27474 30978 27530 30986
rect 27686 30986 27688 31034
rect 27688 30986 27740 31034
rect 27740 30986 27742 31034
rect 27686 30978 27742 30986
rect 27474 30769 27476 30816
rect 27476 30769 27528 30816
rect 27528 30769 27530 30816
rect 27474 30760 27530 30769
rect 27686 30769 27688 30816
rect 27688 30769 27740 30816
rect 27740 30769 27742 30816
rect 27686 30760 27742 30769
rect 27474 30551 27476 30598
rect 27476 30551 27528 30598
rect 27528 30551 27530 30598
rect 27474 30542 27530 30551
rect 27686 30551 27688 30598
rect 27688 30551 27740 30598
rect 27740 30551 27742 30598
rect 27686 30542 27742 30551
rect 27474 26743 27530 26799
rect 27686 26743 27742 26799
rect 27474 26525 27530 26581
rect 27686 26525 27742 26581
rect 27474 24972 27530 25028
rect 27686 24972 27742 25028
rect 27474 24754 27530 24810
rect 27686 24754 27742 24810
rect 27475 22934 27476 22936
rect 27476 22934 27528 22936
rect 27528 22934 27688 22936
rect 27688 22934 27739 22936
rect 27475 22768 27739 22934
rect 27475 22716 27476 22768
rect 27476 22716 27528 22768
rect 27528 22716 27688 22768
rect 27688 22716 27739 22768
rect 27475 22551 27739 22716
rect 27475 22499 27476 22551
rect 27476 22499 27528 22551
rect 27528 22499 27688 22551
rect 27688 22499 27739 22551
rect 27475 22333 27739 22499
rect 27475 22281 27476 22333
rect 27476 22281 27528 22333
rect 27528 22281 27688 22333
rect 27688 22281 27739 22333
rect 27475 22115 27739 22281
rect 27475 22063 27476 22115
rect 27476 22063 27528 22115
rect 27528 22063 27688 22115
rect 27688 22063 27739 22115
rect 27475 22048 27739 22063
rect 27474 16457 27530 16470
rect 27474 16414 27476 16457
rect 27476 16414 27528 16457
rect 27528 16414 27530 16457
rect 27686 16457 27742 16470
rect 27686 16414 27688 16457
rect 27688 16414 27740 16457
rect 27740 16414 27742 16457
rect 27474 16239 27530 16253
rect 27474 16197 27476 16239
rect 27476 16197 27528 16239
rect 27528 16197 27530 16239
rect 27686 16239 27742 16253
rect 27686 16197 27688 16239
rect 27688 16197 27740 16239
rect 27740 16197 27742 16239
rect 27474 16022 27530 16035
rect 27474 15979 27476 16022
rect 27476 15979 27528 16022
rect 27528 15979 27530 16022
rect 27686 16022 27742 16035
rect 27686 15979 27688 16022
rect 27688 15979 27740 16022
rect 27740 15979 27742 16022
rect 27474 15804 27530 15818
rect 27474 15762 27476 15804
rect 27476 15762 27528 15804
rect 27528 15762 27530 15804
rect 27686 15804 27742 15818
rect 27686 15762 27688 15804
rect 27688 15762 27740 15804
rect 27740 15762 27742 15804
rect 27474 15586 27530 15600
rect 27474 15544 27476 15586
rect 27476 15544 27528 15586
rect 27528 15544 27530 15586
rect 27686 15586 27742 15600
rect 27686 15544 27688 15586
rect 27688 15544 27740 15586
rect 27740 15544 27742 15586
rect 27474 15369 27530 15382
rect 27474 15326 27476 15369
rect 27476 15326 27528 15369
rect 27528 15326 27530 15369
rect 27686 15369 27742 15382
rect 27686 15326 27688 15369
rect 27688 15326 27740 15369
rect 27740 15326 27742 15369
rect 27474 15151 27530 15164
rect 27474 15108 27476 15151
rect 27476 15108 27528 15151
rect 27528 15108 27530 15151
rect 27686 15151 27742 15164
rect 27686 15108 27688 15151
rect 27688 15108 27740 15151
rect 27740 15108 27742 15151
rect 27474 14933 27530 14947
rect 27474 14891 27476 14933
rect 27476 14891 27528 14933
rect 27528 14891 27530 14933
rect 27686 14933 27742 14947
rect 27686 14891 27688 14933
rect 27688 14891 27740 14933
rect 27740 14891 27742 14933
rect 27474 14716 27530 14729
rect 27474 14673 27476 14716
rect 27476 14673 27528 14716
rect 27528 14673 27530 14716
rect 27686 14716 27742 14729
rect 27686 14673 27688 14716
rect 27688 14673 27740 14716
rect 27740 14673 27742 14716
rect 27474 14498 27530 14512
rect 27474 14456 27476 14498
rect 27476 14456 27528 14498
rect 27528 14456 27530 14498
rect 27686 14498 27742 14512
rect 27686 14456 27688 14498
rect 27688 14456 27740 14498
rect 27740 14456 27742 14498
rect 27474 14229 27476 14231
rect 27476 14229 27528 14231
rect 27528 14229 27530 14231
rect 27474 14175 27530 14229
rect 27686 14229 27688 14231
rect 27688 14229 27740 14231
rect 27740 14229 27742 14231
rect 27686 14175 27742 14229
rect 27474 14011 27476 14014
rect 27476 14011 27528 14014
rect 27528 14011 27530 14014
rect 27474 13958 27530 14011
rect 27686 14011 27688 14014
rect 27688 14011 27740 14014
rect 27740 14011 27742 14014
rect 27686 13958 27742 14011
rect 27474 13793 27476 13796
rect 27476 13793 27528 13796
rect 27528 13793 27530 13796
rect 27474 13740 27530 13793
rect 27686 13793 27688 13796
rect 27688 13793 27740 13796
rect 27740 13793 27742 13796
rect 27686 13740 27742 13793
rect 27474 13576 27476 13578
rect 27476 13576 27528 13578
rect 27528 13576 27530 13578
rect 27474 13522 27530 13576
rect 27686 13576 27688 13578
rect 27688 13576 27740 13578
rect 27740 13576 27742 13578
rect 27686 13522 27742 13576
rect 27474 13358 27476 13361
rect 27476 13358 27528 13361
rect 27528 13358 27530 13361
rect 27474 13305 27530 13358
rect 27686 13358 27688 13361
rect 27688 13358 27740 13361
rect 27740 13358 27742 13361
rect 27686 13305 27742 13358
rect 27474 11399 27476 11406
rect 27476 11399 27528 11406
rect 27528 11399 27530 11406
rect 27474 11350 27530 11399
rect 27686 11399 27688 11406
rect 27688 11399 27740 11406
rect 27740 11399 27742 11406
rect 27686 11350 27742 11399
rect 27474 11182 27476 11189
rect 27476 11182 27528 11189
rect 27528 11182 27530 11189
rect 27474 11133 27530 11182
rect 27686 11182 27688 11189
rect 27688 11182 27740 11189
rect 27740 11182 27742 11189
rect 27686 11133 27742 11182
rect 27474 10964 27476 10971
rect 27476 10964 27528 10971
rect 27528 10964 27530 10971
rect 27474 10915 27530 10964
rect 27686 10964 27688 10971
rect 27688 10964 27740 10971
rect 27740 10964 27742 10971
rect 27686 10915 27742 10964
rect 27474 10746 27476 10753
rect 27476 10746 27528 10753
rect 27528 10746 27530 10753
rect 27474 10697 27530 10746
rect 27686 10746 27688 10753
rect 27688 10746 27740 10753
rect 27740 10746 27742 10753
rect 27686 10697 27742 10746
rect 27474 10529 27476 10535
rect 27476 10529 27528 10535
rect 27528 10529 27530 10535
rect 27474 10479 27530 10529
rect 27686 10529 27688 10535
rect 27688 10529 27740 10535
rect 27740 10529 27742 10535
rect 27686 10479 27742 10529
rect 27474 10311 27476 10318
rect 27476 10311 27528 10318
rect 27528 10311 27530 10318
rect 27474 10262 27530 10311
rect 27686 10311 27688 10318
rect 27688 10311 27740 10318
rect 27740 10311 27742 10318
rect 27686 10262 27742 10311
rect 57381 33085 57437 33141
rect 57593 33085 57649 33141
rect 57381 32867 57437 32923
rect 57593 32867 57649 32923
rect 57381 32649 57437 32705
rect 57593 32649 57649 32705
rect 57381 32431 57437 32487
rect 57593 32431 57649 32487
rect 57381 31196 57437 31252
rect 57593 31196 57649 31252
rect 57381 30978 57437 31034
rect 57593 30978 57649 31034
rect 57381 30760 57437 30816
rect 57593 30760 57649 30816
rect 57381 30542 57437 30598
rect 57593 30542 57649 30598
rect 57381 26743 57437 26799
rect 57593 26743 57649 26799
rect 57381 26525 57437 26581
rect 57593 26525 57649 26581
rect 57363 22035 57627 22923
rect 57381 16622 57437 16678
rect 57593 16622 57649 16678
rect 57381 16405 57437 16461
rect 57593 16405 57649 16461
rect 57381 16187 57437 16243
rect 57593 16187 57649 16243
rect 57381 15970 57437 16026
rect 57593 15970 57649 16026
rect 57381 15752 57437 15808
rect 57593 15752 57649 15808
rect 57381 15534 57437 15590
rect 57593 15534 57649 15590
rect 57381 15316 57437 15372
rect 57593 15316 57649 15372
rect 57381 15099 57437 15155
rect 57593 15099 57649 15155
rect 57381 14881 57437 14937
rect 57593 14881 57649 14937
rect 57381 14664 57437 14720
rect 57593 14664 57649 14720
rect 57381 11350 57437 11406
rect 57593 11350 57649 11406
rect 57381 11133 57437 11189
rect 57593 11133 57649 11189
rect 57381 10915 57437 10971
rect 57593 10915 57649 10971
rect 57381 10697 57437 10753
rect 57593 10697 57649 10753
rect 57381 10479 57437 10535
rect 57593 10479 57649 10535
rect 57381 10262 57437 10318
rect 57593 10262 57649 10318
rect 51766 9811 51822 9971
rect 49897 8897 50057 8953
rect 27474 7534 27530 7535
rect 27474 7482 27476 7534
rect 27476 7482 27528 7534
rect 27528 7482 27530 7534
rect 27474 7479 27530 7482
rect 27686 7534 27742 7535
rect 27686 7482 27688 7534
rect 27688 7482 27740 7534
rect 27740 7482 27742 7534
rect 27686 7479 27742 7482
rect 27474 7316 27530 7317
rect 27474 7264 27476 7316
rect 27476 7264 27528 7316
rect 27528 7264 27530 7316
rect 27474 7261 27530 7264
rect 27686 7316 27742 7317
rect 27686 7264 27688 7316
rect 27688 7264 27740 7316
rect 27740 7264 27742 7316
rect 27686 7261 27742 7264
rect 27474 7047 27476 7099
rect 27476 7047 27528 7099
rect 27528 7047 27530 7099
rect 27474 7043 27530 7047
rect 27686 7047 27688 7099
rect 27688 7047 27740 7099
rect 27740 7047 27742 7099
rect 27686 7043 27742 7047
rect 28273 6780 28329 6836
rect 28484 6780 28540 6836
rect 28696 6780 28752 6836
rect 28907 6780 28963 6836
rect 28273 6562 28329 6618
rect 28484 6562 28540 6618
rect 28696 6562 28752 6618
rect 28907 6562 28963 6618
rect 28273 6344 28329 6400
rect 28484 6344 28540 6400
rect 28696 6344 28752 6400
rect 28907 6344 28963 6400
rect 27474 6064 27530 6120
rect 27686 6064 27742 6120
rect 27474 5846 27530 5902
rect 27686 5846 27742 5902
rect 26859 4472 26915 4528
rect 27071 4472 27127 4528
rect 26859 4254 26915 4310
rect 27071 4254 27127 4310
rect 27474 3781 27530 3837
rect 27686 3781 27742 3837
rect 27474 3563 27530 3619
rect 27686 3563 27742 3619
rect 28801 3781 28857 3837
rect 28801 3563 28857 3619
rect 57386 8878 57442 8934
rect 57510 8878 57566 8934
rect 57634 8878 57690 8934
rect 57386 8754 57442 8810
rect 57510 8754 57566 8810
rect 57634 8754 57690 8810
rect 57386 8630 57442 8686
rect 57510 8630 57566 8686
rect 57634 8630 57690 8686
rect 57386 8506 57442 8562
rect 57510 8506 57566 8562
rect 57634 8506 57690 8562
rect 57386 8382 57442 8438
rect 57510 8382 57566 8438
rect 57634 8382 57690 8438
rect 57386 8258 57442 8314
rect 57510 8258 57566 8314
rect 57634 8258 57690 8314
rect 57386 8134 57442 8190
rect 57510 8134 57566 8190
rect 57634 8134 57690 8190
rect 57386 8010 57442 8066
rect 57510 8010 57566 8066
rect 57634 8010 57690 8066
rect 57386 7886 57442 7942
rect 57510 7886 57566 7942
rect 57634 7886 57690 7942
rect 57386 7762 57442 7818
rect 57510 7762 57566 7818
rect 57634 7762 57690 7818
rect 57386 7638 57442 7694
rect 57510 7638 57566 7694
rect 57634 7638 57690 7694
rect 57386 7514 57442 7570
rect 57510 7514 57566 7570
rect 57634 7514 57690 7570
rect 57386 7390 57442 7446
rect 57510 7390 57566 7446
rect 57634 7390 57690 7446
rect 57386 7266 57442 7322
rect 57510 7266 57566 7322
rect 57634 7266 57690 7322
rect 57386 7142 57442 7198
rect 57510 7142 57566 7198
rect 57634 7142 57690 7198
rect 56160 6780 56216 6836
rect 56371 6780 56427 6836
rect 56583 6780 56639 6836
rect 56794 6780 56850 6836
rect 56160 6562 56216 6618
rect 56371 6562 56427 6618
rect 56583 6562 56639 6618
rect 56794 6562 56850 6618
rect 56160 6344 56216 6400
rect 56371 6344 56427 6400
rect 56583 6344 56639 6400
rect 56794 6344 56850 6400
rect 57381 6064 57437 6120
rect 57593 6064 57649 6120
rect 57381 5846 57437 5902
rect 57593 5846 57649 5902
rect 43800 2988 43960 3044
rect 48671 2766 48727 2822
rect 48795 2766 48851 2822
rect 48919 2766 48975 2822
rect 48671 2642 48727 2698
rect 48795 2642 48851 2698
rect 48919 2642 48975 2698
rect 48671 2518 48727 2574
rect 48795 2518 48851 2574
rect 48919 2518 48975 2574
rect 49161 2087 49217 2143
rect 49285 2087 49341 2143
rect 49409 2087 49465 2143
rect 49161 1963 49217 2019
rect 49285 1963 49341 2019
rect 49409 1963 49465 2019
rect 49161 1839 49217 1895
rect 49285 1839 49341 1895
rect 49409 1839 49465 1895
rect 57381 3781 57437 3837
rect 57593 3781 57649 3837
rect 57381 3563 57437 3619
rect 57593 3563 57649 3619
rect 57996 33955 58052 34011
rect 58208 33955 58264 34011
rect 57996 33737 58052 33793
rect 58208 33737 58264 33793
rect 57996 33520 58052 33576
rect 58208 33520 58264 33576
rect 57996 33302 58052 33358
rect 58208 33302 58264 33358
rect 57996 33084 58052 33140
rect 58208 33084 58264 33140
rect 57996 32866 58052 32922
rect 58208 32866 58264 32922
rect 57996 32649 58052 32705
rect 58208 32649 58264 32705
rect 57996 32431 58052 32487
rect 58208 32431 58264 32487
rect 57996 32075 57998 32088
rect 57998 32075 58050 32088
rect 58050 32075 58052 32088
rect 57996 32032 58052 32075
rect 58208 32075 58210 32088
rect 58210 32075 58262 32088
rect 58262 32075 58264 32088
rect 58208 32032 58264 32075
rect 57996 31857 57998 31870
rect 57998 31857 58050 31870
rect 58050 31857 58052 31870
rect 57996 31814 58052 31857
rect 58208 31857 58210 31870
rect 58210 31857 58262 31870
rect 58262 31857 58264 31870
rect 58208 31814 58264 31857
rect 57996 31639 57998 31652
rect 57998 31639 58050 31652
rect 58050 31639 58052 31652
rect 57996 31596 58052 31639
rect 58208 31639 58210 31652
rect 58210 31639 58262 31652
rect 58262 31639 58264 31652
rect 58208 31596 58264 31639
rect 57996 29950 58052 29968
rect 57996 29912 57998 29950
rect 57998 29912 58050 29950
rect 58050 29912 58052 29950
rect 58208 29950 58264 29968
rect 58208 29912 58210 29950
rect 58210 29912 58262 29950
rect 58262 29912 58264 29950
rect 57996 29733 58052 29750
rect 57996 29694 57998 29733
rect 57998 29694 58050 29733
rect 58050 29694 58052 29733
rect 58208 29733 58264 29750
rect 58208 29694 58210 29733
rect 58210 29694 58262 29733
rect 58262 29694 58264 29733
rect 57996 29515 58052 29533
rect 57996 29477 57998 29515
rect 57998 29477 58050 29515
rect 58050 29477 58052 29515
rect 58208 29515 58264 29533
rect 58208 29477 58210 29515
rect 58210 29477 58262 29515
rect 58262 29477 58264 29515
rect 57996 29297 58052 29315
rect 57996 29259 57998 29297
rect 57998 29259 58050 29297
rect 58050 29259 58052 29297
rect 58208 29297 58264 29315
rect 58208 29259 58210 29297
rect 58210 29259 58262 29297
rect 58262 29259 58264 29297
rect 57996 29080 58052 29098
rect 57996 29042 57998 29080
rect 57998 29042 58050 29080
rect 58050 29042 58052 29080
rect 58208 29080 58264 29098
rect 58208 29042 58210 29080
rect 58210 29042 58262 29080
rect 58262 29042 58264 29080
rect 57996 28862 58052 28880
rect 57996 28824 57998 28862
rect 57998 28824 58050 28862
rect 58050 28824 58052 28862
rect 58208 28862 58264 28880
rect 58208 28824 58210 28862
rect 58210 28824 58262 28862
rect 58262 28824 58264 28862
rect 57996 28644 58052 28662
rect 57996 28606 57998 28644
rect 57998 28606 58050 28644
rect 58050 28606 58052 28644
rect 58208 28644 58264 28662
rect 58208 28606 58210 28644
rect 58210 28606 58262 28644
rect 58262 28606 58264 28644
rect 57996 28427 58052 28444
rect 57996 28388 57998 28427
rect 57998 28388 58050 28427
rect 58050 28388 58052 28427
rect 58208 28427 58264 28444
rect 58208 28388 58210 28427
rect 58210 28388 58262 28427
rect 58262 28388 58264 28427
rect 57996 28209 58052 28227
rect 57996 28171 57998 28209
rect 57998 28171 58050 28209
rect 58050 28171 58052 28209
rect 58208 28209 58264 28227
rect 58208 28171 58210 28209
rect 58210 28171 58262 28209
rect 58262 28171 58264 28209
rect 57996 27992 58052 28009
rect 57996 27953 57998 27992
rect 57998 27953 58050 27992
rect 58050 27953 58052 27992
rect 58208 27992 58264 28009
rect 58208 27953 58210 27992
rect 58210 27953 58262 27992
rect 58262 27953 58264 27992
rect 57996 27774 58052 27792
rect 57996 27736 57998 27774
rect 57998 27736 58050 27774
rect 58050 27736 58052 27774
rect 58208 27774 58264 27792
rect 58208 27736 58210 27774
rect 58210 27736 58262 27774
rect 58262 27736 58264 27774
rect 57996 27556 58052 27574
rect 57996 27518 57998 27556
rect 57998 27518 58050 27556
rect 58050 27518 58052 27556
rect 58208 27556 58264 27574
rect 58208 27518 58210 27556
rect 58210 27518 58262 27556
rect 58262 27518 58264 27556
rect 58812 44286 58814 44314
rect 58814 44286 58866 44314
rect 58866 44286 58868 44314
rect 58812 44258 58868 44286
rect 58936 44286 58938 44314
rect 58938 44286 58990 44314
rect 58990 44286 58992 44314
rect 58936 44258 58992 44286
rect 59060 44286 59062 44314
rect 59062 44286 59114 44314
rect 59114 44286 59116 44314
rect 59060 44258 59116 44286
rect 59184 44286 59186 44314
rect 59186 44286 59238 44314
rect 59238 44286 59240 44314
rect 59184 44258 59240 44286
rect 59308 44286 59310 44314
rect 59310 44286 59362 44314
rect 59362 44286 59364 44314
rect 59308 44258 59364 44286
rect 59432 44286 59434 44314
rect 59434 44286 59486 44314
rect 59486 44286 59488 44314
rect 59432 44258 59488 44286
rect 58812 44162 58814 44190
rect 58814 44162 58866 44190
rect 58866 44162 58868 44190
rect 58812 44134 58868 44162
rect 58936 44162 58938 44190
rect 58938 44162 58990 44190
rect 58990 44162 58992 44190
rect 58936 44134 58992 44162
rect 59060 44162 59062 44190
rect 59062 44162 59114 44190
rect 59114 44162 59116 44190
rect 59060 44134 59116 44162
rect 59184 44162 59186 44190
rect 59186 44162 59238 44190
rect 59238 44162 59240 44190
rect 59184 44134 59240 44162
rect 59308 44162 59310 44190
rect 59310 44162 59362 44190
rect 59362 44162 59364 44190
rect 59308 44134 59364 44162
rect 59432 44162 59434 44190
rect 59434 44162 59486 44190
rect 59486 44162 59488 44190
rect 59432 44134 59488 44162
rect 58873 31242 58929 31298
rect 58997 31242 59053 31298
rect 59121 31242 59177 31298
rect 59245 31242 59301 31298
rect 59369 31242 59425 31298
rect 58873 31118 58929 31174
rect 58997 31118 59053 31174
rect 59121 31118 59177 31174
rect 59245 31118 59301 31174
rect 59369 31118 59425 31174
rect 58873 30994 58929 31050
rect 58997 30994 59053 31050
rect 59121 30994 59177 31050
rect 59245 30994 59301 31050
rect 59369 30994 59425 31050
rect 58873 30797 58929 30853
rect 58997 30797 59053 30853
rect 59121 30797 59177 30853
rect 59245 30797 59301 30853
rect 59369 30797 59425 30853
rect 58873 30673 58929 30729
rect 58997 30673 59053 30729
rect 59121 30673 59177 30729
rect 59245 30673 59301 30729
rect 59369 30673 59425 30729
rect 58873 30549 58929 30605
rect 58997 30549 59053 30605
rect 59121 30549 59177 30605
rect 59245 30549 59301 30605
rect 59369 30549 59425 30605
rect 58859 28216 58915 28272
rect 58983 28216 59039 28272
rect 59107 28216 59163 28272
rect 59231 28216 59287 28272
rect 59355 28216 59411 28272
rect 58859 28092 58915 28148
rect 58983 28092 59039 28148
rect 59107 28092 59163 28148
rect 59231 28092 59287 28148
rect 59355 28092 59411 28148
rect 58859 27968 58915 28024
rect 58983 27968 59039 28024
rect 59107 27968 59163 28024
rect 59231 27968 59287 28024
rect 59355 27968 59411 28024
rect 58859 27844 58915 27900
rect 58983 27844 59039 27900
rect 59107 27844 59163 27900
rect 59231 27844 59287 27900
rect 59355 27844 59411 27900
rect 58859 27720 58915 27776
rect 58983 27720 59039 27776
rect 59107 27720 59163 27776
rect 59231 27720 59287 27776
rect 59355 27720 59411 27776
rect 58859 27596 58915 27652
rect 58983 27596 59039 27652
rect 59107 27596 59163 27652
rect 59231 27596 59287 27652
rect 59355 27596 59411 27652
rect 58859 27472 58915 27528
rect 58983 27472 59039 27528
rect 59107 27472 59163 27528
rect 59231 27472 59287 27528
rect 59355 27472 59411 27528
rect 58859 27348 58915 27404
rect 58983 27348 59039 27404
rect 59107 27348 59163 27404
rect 59231 27348 59287 27404
rect 59355 27348 59411 27404
rect 58859 27224 58915 27280
rect 58983 27224 59039 27280
rect 59107 27224 59163 27280
rect 59231 27224 59287 27280
rect 59355 27224 59411 27280
rect 58859 27100 58915 27156
rect 58983 27100 59039 27156
rect 59107 27100 59163 27156
rect 59231 27100 59287 27156
rect 59355 27100 59411 27156
rect 58859 26976 58915 27032
rect 58983 26976 59039 27032
rect 59107 26976 59163 27032
rect 59231 26976 59287 27032
rect 59355 26976 59411 27032
rect 58859 26852 58915 26908
rect 58983 26852 59039 26908
rect 59107 26852 59163 26908
rect 59231 26852 59287 26908
rect 59355 26852 59411 26908
rect 58859 26728 58915 26784
rect 58983 26728 59039 26784
rect 59107 26728 59163 26784
rect 59231 26728 59287 26784
rect 59355 26728 59411 26784
rect 58859 26604 58915 26660
rect 58983 26604 59039 26660
rect 59107 26604 59163 26660
rect 59231 26604 59287 26660
rect 59355 26604 59411 26660
rect 58859 26480 58915 26536
rect 58983 26480 59039 26536
rect 59107 26480 59163 26536
rect 59231 26480 59287 26536
rect 59355 26480 59411 26536
rect 57994 24074 58258 24075
rect 57994 24022 57998 24074
rect 57998 24022 58050 24074
rect 58050 24022 58210 24074
rect 58210 24022 58258 24074
rect 57994 23857 58258 24022
rect 57994 23805 57998 23857
rect 57998 23805 58050 23857
rect 58050 23805 58210 23857
rect 58210 23805 58258 23857
rect 57994 23639 58258 23805
rect 57994 23587 57998 23639
rect 57998 23587 58050 23639
rect 58050 23587 58210 23639
rect 58210 23587 58258 23639
rect 57994 23421 58258 23587
rect 57994 23369 57998 23421
rect 57998 23369 58050 23421
rect 58050 23369 58210 23421
rect 58210 23369 58258 23421
rect 57994 23204 58258 23369
rect 57994 23187 57998 23204
rect 57998 23187 58050 23204
rect 58050 23187 58210 23204
rect 58210 23187 58258 23204
rect 58048 20540 58050 20570
rect 58050 20540 58208 20570
rect 58048 20410 58208 20540
rect 58048 20157 58208 20226
rect 58048 20105 58050 20157
rect 58050 20105 58208 20157
rect 58048 20066 58208 20105
rect 57996 13734 58052 13790
rect 58208 13734 58264 13790
rect 57996 13517 58052 13573
rect 58208 13517 58264 13573
rect 57996 13299 58052 13355
rect 58208 13299 58264 13355
rect 57996 13082 58052 13138
rect 58208 13082 58264 13138
rect 57996 12864 58052 12920
rect 58208 12864 58264 12920
rect 57996 12646 58052 12702
rect 58208 12646 58264 12702
rect 57996 12428 58052 12484
rect 58208 12428 58264 12484
rect 57996 12211 58052 12267
rect 58208 12211 58264 12267
rect 57996 11993 58052 12049
rect 58208 11993 58264 12049
rect 57996 11776 58052 11832
rect 58208 11776 58264 11832
rect 57996 9351 58052 9407
rect 58208 9351 58264 9407
rect 57996 9134 58052 9190
rect 58208 9134 58264 9190
rect 57996 8916 58052 8972
rect 58208 8916 58264 8972
rect 57996 8698 58052 8754
rect 58208 8698 58264 8754
rect 57996 8480 58052 8536
rect 58208 8480 58264 8536
rect 57996 8263 58052 8319
rect 58208 8263 58264 8319
rect 57996 5523 57998 5539
rect 57998 5523 58050 5539
rect 58050 5523 58052 5539
rect 57996 5483 58052 5523
rect 58208 5523 58210 5539
rect 58210 5523 58262 5539
rect 58262 5523 58264 5539
rect 58208 5483 58264 5523
rect 57996 5306 57998 5321
rect 57998 5306 58050 5321
rect 58050 5306 58052 5321
rect 57996 5265 58052 5306
rect 58208 5306 58210 5321
rect 58210 5306 58262 5321
rect 58262 5306 58264 5321
rect 58208 5265 58264 5306
rect 57996 4472 58052 4528
rect 58208 4472 58264 4528
rect 57996 4254 58052 4310
rect 58208 4254 58264 4310
<< metal3 >>
rect 1401 45776 2401 46576
rect 2626 45968 3626 46576
rect 4137 45776 5137 46576
rect 5362 45968 6362 46576
rect 6801 45776 7801 46576
rect 8026 45968 9026 46576
rect 9537 45776 10537 46576
rect 10762 45968 11762 46576
rect 12201 45776 13201 46576
rect 13426 45968 14426 46576
rect 14937 45776 15937 46576
rect 16162 45968 17162 46576
rect 17601 45776 18601 46576
rect 18826 45968 19826 46576
rect 20653 45776 21653 46576
rect 22258 45968 23258 46576
rect 23483 45776 24483 46576
rect 25158 45968 26158 46576
rect 26572 45776 27572 46576
rect 27877 45968 28877 46576
rect 29273 45968 30273 46576
rect 30710 45776 31710 46576
rect 32381 45968 33381 46576
rect 34024 45968 35024 46576
rect 35415 45776 36415 46576
rect 36948 45968 37948 46576
rect 38585 45776 39585 46576
rect 39882 45968 40882 46576
rect 41230 45776 42230 46576
rect 42430 45968 43430 46576
rect 43713 45968 44713 46576
rect 45069 45776 46069 46576
rect 46313 45776 47313 46576
rect 47538 45968 48538 46576
rect 48901 45776 49901 46576
rect 50465 45968 51465 46576
rect 52569 45776 53569 46576
rect 54262 45776 55262 46576
rect 55990 45968 56990 46576
rect 57547 45776 58547 46576
rect 58791 45968 59791 46576
rect 60977 45776 61977 46576
rect 62202 45968 63202 46576
rect 63713 45776 64713 46576
rect 64938 45968 65938 46576
rect 66377 45776 67377 46576
rect 67602 45968 68602 46576
rect 69113 45776 70113 46576
rect 70338 45968 71338 46576
rect 71777 45776 72777 46576
rect 73002 45968 74002 46576
rect 74513 45776 75513 46576
rect 75738 45968 76738 46576
rect 77177 45776 78177 46576
rect 78402 45968 79402 46576
rect 80229 45776 81229 46576
rect 81834 45968 82834 46576
rect 83059 45776 84059 46576
rect 84666 45776 85666 46576
rect 0 44776 86372 45776
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44328 27779 44376
rect 57051 44328 86372 44376
rect 0 44314 86372 44328
rect 0 44258 25335 44314
rect 25391 44258 25459 44314
rect 25515 44258 25583 44314
rect 25639 44258 25707 44314
rect 25763 44258 25831 44314
rect 25887 44258 25955 44314
rect 26011 44258 58812 44314
rect 58868 44258 58936 44314
rect 58992 44258 59060 44314
rect 59116 44258 59184 44314
rect 59240 44258 59308 44314
rect 59364 44258 59432 44314
rect 59488 44258 86372 44314
rect 0 44255 86372 44258
rect 0 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 34288 44255
rect 34344 44199 34499 44255
rect 34555 44199 34710 44255
rect 34766 44199 34921 44255
rect 34977 44199 40250 44255
rect 40306 44199 40430 44255
rect 40486 44199 50135 44255
rect 50191 44199 50346 44255
rect 50402 44199 50557 44255
rect 50613 44199 50768 44255
rect 50824 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 86372 44255
rect 0 44190 86372 44199
rect 0 44134 25335 44190
rect 25391 44134 25459 44190
rect 25515 44134 25583 44190
rect 25639 44134 25707 44190
rect 25763 44134 25831 44190
rect 25887 44134 25955 44190
rect 26011 44134 58812 44190
rect 58868 44134 58936 44190
rect 58992 44134 59060 44190
rect 59116 44134 59184 44190
rect 59240 44134 59308 44190
rect 59364 44134 59432 44190
rect 59488 44134 86372 44190
rect 0 44127 86372 44134
rect 0 44076 27779 44127
rect 30402 44126 54622 44127
rect 57051 44076 86372 44127
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 28677 43834 33984 43868
rect 28676 43774 33984 43834
rect 28676 43718 33048 43774
rect 33104 43718 33259 43774
rect 33315 43718 33470 43774
rect 33526 43718 33681 43774
rect 33737 43718 33892 43774
rect 33948 43718 33984 43774
rect 28676 43700 33984 43718
rect 0 42976 1706 43676
rect 28677 43666 33984 43700
rect 36863 43772 42155 43811
rect 36863 43716 36899 43772
rect 36955 43716 37110 43772
rect 37166 43716 37321 43772
rect 37377 43716 37532 43772
rect 37588 43716 41008 43772
rect 41064 43716 41219 43772
rect 41275 43716 41430 43772
rect 41486 43716 41641 43772
rect 41697 43716 41852 43772
rect 41908 43716 42062 43772
rect 42118 43716 42155 43772
rect 36863 43677 42155 43716
rect 42671 43765 43222 43804
rect 42671 43709 42708 43765
rect 42764 43709 42919 43765
rect 42975 43709 43130 43765
rect 43186 43709 43222 43765
rect 42671 43428 43222 43709
rect 51042 43772 61644 43868
rect 51042 43716 51079 43772
rect 51135 43716 51290 43772
rect 51346 43716 51501 43772
rect 51557 43716 51712 43772
rect 51768 43716 51923 43772
rect 51979 43716 61644 43772
rect 51042 43666 61644 43716
rect 25313 43417 59810 43428
rect 25313 43361 26838 43417
rect 26894 43361 26962 43417
rect 27018 43361 27086 43417
rect 27142 43361 59810 43417
rect 25313 43355 59810 43361
rect 25313 43299 29580 43355
rect 29636 43299 29791 43355
rect 29847 43299 30003 43355
rect 30059 43299 30214 43355
rect 30270 43299 30852 43355
rect 30908 43299 31063 43355
rect 31119 43299 31274 43355
rect 31330 43299 31484 43355
rect 31540 43299 31695 43355
rect 31751 43299 31907 43355
rect 31963 43299 32118 43355
rect 32174 43299 32328 43355
rect 32384 43299 32539 43355
rect 32595 43299 32750 43355
rect 32806 43299 35218 43355
rect 35274 43299 35428 43355
rect 35484 43299 35639 43355
rect 35695 43299 35851 43355
rect 35907 43299 36062 43355
rect 36118 43299 36272 43355
rect 36328 43299 39050 43355
rect 39106 43299 39230 43355
rect 39286 43299 40777 43355
rect 40833 43299 40988 43355
rect 41044 43299 41199 43355
rect 41255 43299 44832 43355
rect 44888 43299 45043 43355
rect 45099 43299 45254 43355
rect 45310 43299 48836 43355
rect 48892 43299 49046 43355
rect 49102 43299 49257 43355
rect 49313 43299 49469 43355
rect 49525 43299 49680 43355
rect 49736 43299 49890 43355
rect 49946 43299 52314 43355
rect 52370 43299 52525 43355
rect 52581 43299 52736 43355
rect 52792 43299 52946 43355
rect 53002 43299 53157 43355
rect 53213 43299 53369 43355
rect 53425 43299 53580 43355
rect 53636 43299 53790 43355
rect 53846 43299 54001 43355
rect 54057 43299 54212 43355
rect 54268 43299 54853 43355
rect 54909 43299 55064 43355
rect 55120 43299 55276 43355
rect 55332 43299 55487 43355
rect 55543 43299 59810 43355
rect 25313 43293 59810 43299
rect 25313 43237 26838 43293
rect 26894 43237 26962 43293
rect 27018 43237 27086 43293
rect 27142 43237 59810 43293
rect 25313 43227 59810 43237
rect 30403 43226 54622 43227
rect 36648 43001 40041 43002
rect 25313 42922 34090 42988
rect 25313 42866 33055 42922
rect 33111 42866 33235 42922
rect 33291 42915 34090 42922
rect 33291 42866 33817 42915
rect 25313 42859 33817 42866
rect 33873 42859 33997 42915
rect 34053 42859 34090 42915
rect 36640 42963 40085 43001
rect 36640 42907 36676 42963
rect 36732 42907 39992 42963
rect 40048 42907 40085 42963
rect 36640 42868 40085 42907
rect 48557 42949 48687 42988
rect 48557 42893 48594 42949
rect 48650 42893 48687 42949
rect 25313 42787 34090 42859
rect 30403 42786 34090 42787
rect 0 42576 1014 42776
rect 48557 42770 48687 42893
rect 51034 42915 59810 42988
rect 84666 42976 86372 43676
rect 51034 42859 51071 42915
rect 51127 42859 51251 42915
rect 51307 42859 51833 42915
rect 51889 42859 52013 42915
rect 52069 42859 59810 42915
rect 51034 42787 59810 42859
rect 51034 42786 54622 42787
rect 37852 42732 48687 42770
rect 37852 42676 37889 42732
rect 37945 42676 38069 42732
rect 38125 42676 39773 42732
rect 39829 42731 48687 42732
rect 39829 42676 48594 42731
rect 37852 42675 48594 42676
rect 48650 42675 48687 42731
rect 37852 42637 48687 42675
rect 85358 42576 86372 42776
rect 0 42528 27272 42576
rect 59421 42528 86372 42576
rect 0 42455 86372 42528
rect 0 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 34282 42455
rect 34338 42399 34493 42455
rect 34549 42399 34705 42455
rect 34761 42399 34916 42455
rect 34972 42399 38328 42455
rect 38384 42399 38539 42455
rect 38595 42399 38750 42455
rect 38806 42399 40251 42455
rect 40307 42399 40431 42455
rect 40487 42399 43788 42455
rect 43844 42399 43999 42455
rect 44055 42399 44211 42455
rect 44267 42399 44422 42455
rect 44478 42399 50161 42455
rect 50217 42399 50372 42455
rect 50428 42399 50584 42455
rect 50640 42399 50795 42455
rect 50851 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 86372 42455
rect 0 42327 86372 42399
rect 0 42276 27272 42327
rect 30403 42326 54622 42327
rect 59421 42276 86372 42327
rect 0 42076 1014 42276
rect 37852 42179 48687 42217
rect 37852 42178 48594 42179
rect 37852 42122 37889 42178
rect 37945 42122 38069 42178
rect 38125 42122 39773 42178
rect 39829 42123 48594 42178
rect 48650 42123 48687 42179
rect 39829 42122 48687 42123
rect 37852 42084 48687 42122
rect 25313 41995 34090 42068
rect 25313 41988 33817 41995
rect 25313 41932 33055 41988
rect 33111 41932 33235 41988
rect 33291 41939 33817 41988
rect 33873 41939 33997 41995
rect 34053 41939 34090 41995
rect 33291 41932 34090 41939
rect 0 41176 1706 41876
rect 25313 41866 34090 41932
rect 36640 41947 40085 41986
rect 36640 41891 36676 41947
rect 36732 41891 39992 41947
rect 40048 41891 40085 41947
rect 36640 41853 40085 41891
rect 48557 41961 48687 42084
rect 85358 42076 86372 42276
rect 48557 41905 48594 41961
rect 48650 41905 48687 41961
rect 48557 41866 48687 41905
rect 51034 41995 59810 42068
rect 51034 41939 51071 41995
rect 51127 41939 51251 41995
rect 51307 41939 51833 41995
rect 51889 41939 52013 41995
rect 52069 41939 59810 41995
rect 51034 41866 59810 41939
rect 36648 41852 40041 41853
rect 25313 41555 59810 41628
rect 25313 41499 29580 41555
rect 29636 41499 29791 41555
rect 29847 41499 30003 41555
rect 30059 41499 30214 41555
rect 30270 41499 30852 41555
rect 30908 41499 31063 41555
rect 31119 41499 31274 41555
rect 31330 41499 31484 41555
rect 31540 41499 31695 41555
rect 31751 41499 31907 41555
rect 31963 41499 32118 41555
rect 32174 41499 32328 41555
rect 32384 41499 32539 41555
rect 32595 41499 32750 41555
rect 32806 41499 35218 41555
rect 35274 41499 35428 41555
rect 35484 41499 35639 41555
rect 35695 41499 35851 41555
rect 35907 41499 36062 41555
rect 36118 41499 36272 41555
rect 36328 41499 39050 41555
rect 39106 41499 39230 41555
rect 39286 41499 44832 41555
rect 44888 41499 45043 41555
rect 45099 41499 45254 41555
rect 45310 41499 48836 41555
rect 48892 41499 49046 41555
rect 49102 41499 49257 41555
rect 49313 41499 49469 41555
rect 49525 41499 49680 41555
rect 49736 41499 49890 41555
rect 49946 41499 52314 41555
rect 52370 41499 52525 41555
rect 52581 41499 52736 41555
rect 52792 41499 52946 41555
rect 53002 41499 53157 41555
rect 53213 41499 53369 41555
rect 53425 41499 53580 41555
rect 53636 41499 53790 41555
rect 53846 41499 54001 41555
rect 54057 41499 54212 41555
rect 54268 41499 54853 41555
rect 54909 41499 55064 41555
rect 55120 41499 55276 41555
rect 55332 41499 55487 41555
rect 55543 41499 59810 41555
rect 25313 41427 59810 41499
rect 30403 41426 54622 41427
rect 36648 41201 40041 41202
rect 25313 41122 34090 41188
rect 25313 41066 33055 41122
rect 33111 41066 33235 41122
rect 33291 41115 34090 41122
rect 33291 41066 33817 41115
rect 25313 41059 33817 41066
rect 33873 41059 33997 41115
rect 34053 41059 34090 41115
rect 36640 41163 40085 41201
rect 36640 41107 36676 41163
rect 36732 41107 39992 41163
rect 40048 41107 40085 41163
rect 36640 41068 40085 41107
rect 48557 41149 48687 41188
rect 48557 41093 48594 41149
rect 48650 41093 48687 41149
rect 25313 40987 34090 41059
rect 30403 40986 34090 40987
rect 0 40776 1014 40976
rect 48557 40970 48687 41093
rect 51034 41115 59810 41188
rect 84666 41176 86372 41876
rect 51034 41059 51071 41115
rect 51127 41059 51251 41115
rect 51307 41059 51833 41115
rect 51889 41059 52013 41115
rect 52069 41059 59810 41115
rect 51034 40987 59810 41059
rect 51034 40986 54622 40987
rect 37852 40932 48687 40970
rect 37852 40876 37889 40932
rect 37945 40876 38069 40932
rect 38125 40876 39773 40932
rect 39829 40931 48687 40932
rect 39829 40876 48594 40931
rect 37852 40875 48594 40876
rect 48650 40875 48687 40931
rect 37852 40837 48687 40875
rect 85358 40776 86372 40976
rect 0 40728 27272 40776
rect 59421 40728 86372 40776
rect 0 40655 86372 40728
rect 0 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 34282 40655
rect 34338 40599 34493 40655
rect 34549 40599 34705 40655
rect 34761 40599 34916 40655
rect 34972 40599 38328 40655
rect 38384 40599 38539 40655
rect 38595 40599 38750 40655
rect 38806 40599 40251 40655
rect 40307 40599 40431 40655
rect 40487 40599 43788 40655
rect 43844 40599 43999 40655
rect 44055 40599 44211 40655
rect 44267 40599 44422 40655
rect 44478 40599 50161 40655
rect 50217 40599 50372 40655
rect 50428 40599 50584 40655
rect 50640 40599 50795 40655
rect 50851 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 86372 40655
rect 0 40527 86372 40599
rect 0 40476 27272 40527
rect 30403 40526 54622 40527
rect 59421 40476 86372 40527
rect 0 40276 1014 40476
rect 37852 40379 48687 40417
rect 37852 40378 48594 40379
rect 37852 40322 37889 40378
rect 37945 40322 38069 40378
rect 38125 40322 39773 40378
rect 39829 40323 48594 40378
rect 48650 40323 48687 40379
rect 39829 40322 48687 40323
rect 37852 40284 48687 40322
rect 25313 40195 34090 40268
rect 25313 40188 33817 40195
rect 25313 40132 33055 40188
rect 33111 40132 33235 40188
rect 33291 40139 33817 40188
rect 33873 40139 33997 40195
rect 34053 40139 34090 40195
rect 33291 40132 34090 40139
rect 0 39376 1706 40076
rect 25313 40066 34090 40132
rect 36640 40147 40085 40186
rect 36640 40091 36676 40147
rect 36732 40091 39992 40147
rect 40048 40091 40085 40147
rect 36640 40053 40085 40091
rect 48557 40161 48687 40284
rect 85358 40276 86372 40476
rect 48557 40105 48594 40161
rect 48650 40105 48687 40161
rect 48557 40066 48687 40105
rect 51034 40195 59810 40268
rect 51034 40139 51071 40195
rect 51127 40139 51251 40195
rect 51307 40139 51833 40195
rect 51889 40139 52013 40195
rect 52069 40139 59810 40195
rect 51034 40066 59810 40139
rect 36648 40052 40041 40053
rect 25313 39755 59810 39828
rect 25313 39699 29580 39755
rect 29636 39699 29791 39755
rect 29847 39699 30003 39755
rect 30059 39699 30214 39755
rect 30270 39699 30852 39755
rect 30908 39699 31063 39755
rect 31119 39699 31274 39755
rect 31330 39699 31484 39755
rect 31540 39699 31695 39755
rect 31751 39699 31907 39755
rect 31963 39699 32118 39755
rect 32174 39699 32328 39755
rect 32384 39699 32539 39755
rect 32595 39699 32750 39755
rect 32806 39699 35218 39755
rect 35274 39699 35428 39755
rect 35484 39699 35639 39755
rect 35695 39699 35851 39755
rect 35907 39699 36062 39755
rect 36118 39699 36272 39755
rect 36328 39699 39050 39755
rect 39106 39699 39230 39755
rect 39286 39699 44832 39755
rect 44888 39699 45043 39755
rect 45099 39699 45254 39755
rect 45310 39699 48836 39755
rect 48892 39699 49046 39755
rect 49102 39699 49257 39755
rect 49313 39699 49469 39755
rect 49525 39699 49680 39755
rect 49736 39699 49890 39755
rect 49946 39699 52314 39755
rect 52370 39699 52525 39755
rect 52581 39699 52736 39755
rect 52792 39699 52946 39755
rect 53002 39699 53157 39755
rect 53213 39699 53369 39755
rect 53425 39699 53580 39755
rect 53636 39699 53790 39755
rect 53846 39699 54001 39755
rect 54057 39699 54212 39755
rect 54268 39699 54853 39755
rect 54909 39699 55064 39755
rect 55120 39699 55276 39755
rect 55332 39699 55487 39755
rect 55543 39699 59810 39755
rect 25313 39627 59810 39699
rect 30403 39626 54622 39627
rect 36648 39401 40041 39402
rect 25313 39322 34090 39388
rect 25313 39266 33055 39322
rect 33111 39266 33235 39322
rect 33291 39315 34090 39322
rect 33291 39266 33817 39315
rect 25313 39259 33817 39266
rect 33873 39259 33997 39315
rect 34053 39259 34090 39315
rect 36640 39363 40085 39401
rect 36640 39307 36676 39363
rect 36732 39307 39992 39363
rect 40048 39307 40085 39363
rect 36640 39268 40085 39307
rect 48557 39349 48687 39388
rect 48557 39293 48594 39349
rect 48650 39293 48687 39349
rect 25313 39187 34090 39259
rect 30403 39186 34090 39187
rect 0 38976 1014 39176
rect 48557 39170 48687 39293
rect 51034 39315 59810 39388
rect 84666 39376 86372 40076
rect 51034 39259 51071 39315
rect 51127 39259 51251 39315
rect 51307 39259 51833 39315
rect 51889 39259 52013 39315
rect 52069 39259 59810 39315
rect 51034 39187 59810 39259
rect 51034 39186 54622 39187
rect 37852 39132 48687 39170
rect 37852 39076 37889 39132
rect 37945 39076 38069 39132
rect 38125 39076 39773 39132
rect 39829 39131 48687 39132
rect 39829 39076 48594 39131
rect 37852 39075 48594 39076
rect 48650 39075 48687 39131
rect 37852 39037 48687 39075
rect 85358 38976 86372 39176
rect 0 38928 27272 38976
rect 59421 38928 86372 38976
rect 0 38855 86372 38928
rect 0 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 34282 38855
rect 34338 38799 34493 38855
rect 34549 38799 34705 38855
rect 34761 38799 34916 38855
rect 34972 38799 38328 38855
rect 38384 38799 38539 38855
rect 38595 38799 38750 38855
rect 38806 38799 40251 38855
rect 40307 38799 40431 38855
rect 40487 38799 43788 38855
rect 43844 38799 43999 38855
rect 44055 38799 44211 38855
rect 44267 38799 44422 38855
rect 44478 38799 50161 38855
rect 50217 38799 50372 38855
rect 50428 38799 50584 38855
rect 50640 38799 50795 38855
rect 50851 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 86372 38855
rect 0 38727 86372 38799
rect 0 38676 27272 38727
rect 30403 38726 54622 38727
rect 59421 38676 86372 38727
rect 0 38476 1014 38676
rect 37852 38579 48687 38617
rect 37852 38578 48594 38579
rect 37852 38522 37889 38578
rect 37945 38522 38069 38578
rect 38125 38522 39773 38578
rect 39829 38523 48594 38578
rect 48650 38523 48687 38579
rect 39829 38522 48687 38523
rect 37852 38484 48687 38522
rect 25313 38395 34090 38468
rect 25313 38388 33817 38395
rect 25313 38332 33055 38388
rect 33111 38332 33235 38388
rect 33291 38339 33817 38388
rect 33873 38339 33997 38395
rect 34053 38339 34090 38395
rect 33291 38332 34090 38339
rect 0 37576 1706 38276
rect 25313 38266 34090 38332
rect 36640 38347 40085 38386
rect 36640 38291 36676 38347
rect 36732 38291 39992 38347
rect 40048 38291 40085 38347
rect 36640 38253 40085 38291
rect 48557 38361 48687 38484
rect 85358 38476 86372 38676
rect 48557 38305 48594 38361
rect 48650 38305 48687 38361
rect 48557 38266 48687 38305
rect 51034 38395 59810 38468
rect 51034 38339 51071 38395
rect 51127 38339 51251 38395
rect 51307 38339 51833 38395
rect 51889 38339 52013 38395
rect 52069 38339 59810 38395
rect 51034 38266 59810 38339
rect 36648 38252 40041 38253
rect 25313 37955 59810 38028
rect 25313 37899 29580 37955
rect 29636 37899 29791 37955
rect 29847 37899 30003 37955
rect 30059 37899 30214 37955
rect 30270 37899 30852 37955
rect 30908 37899 31063 37955
rect 31119 37899 31274 37955
rect 31330 37899 31484 37955
rect 31540 37899 31695 37955
rect 31751 37899 31907 37955
rect 31963 37899 32118 37955
rect 32174 37899 32328 37955
rect 32384 37899 32539 37955
rect 32595 37899 32750 37955
rect 32806 37899 35218 37955
rect 35274 37899 35428 37955
rect 35484 37899 35639 37955
rect 35695 37899 35851 37955
rect 35907 37899 36062 37955
rect 36118 37899 36272 37955
rect 36328 37899 39050 37955
rect 39106 37899 39230 37955
rect 39286 37899 44832 37955
rect 44888 37899 45043 37955
rect 45099 37899 45254 37955
rect 45310 37899 48836 37955
rect 48892 37899 49046 37955
rect 49102 37899 49257 37955
rect 49313 37899 49469 37955
rect 49525 37899 49680 37955
rect 49736 37899 49890 37955
rect 49946 37899 52314 37955
rect 52370 37899 52525 37955
rect 52581 37899 52736 37955
rect 52792 37899 52946 37955
rect 53002 37899 53157 37955
rect 53213 37899 53369 37955
rect 53425 37899 53580 37955
rect 53636 37899 53790 37955
rect 53846 37899 54001 37955
rect 54057 37899 54212 37955
rect 54268 37899 54853 37955
rect 54909 37899 55064 37955
rect 55120 37899 55276 37955
rect 55332 37899 55487 37955
rect 55543 37899 59810 37955
rect 25313 37827 59810 37899
rect 30403 37826 54622 37827
rect 36648 37601 40041 37602
rect 25313 37522 34090 37588
rect 25313 37466 33055 37522
rect 33111 37466 33235 37522
rect 33291 37515 34090 37522
rect 33291 37466 33817 37515
rect 25313 37459 33817 37466
rect 33873 37459 33997 37515
rect 34053 37459 34090 37515
rect 36640 37563 40085 37601
rect 36640 37507 36676 37563
rect 36732 37507 39992 37563
rect 40048 37507 40085 37563
rect 36640 37468 40085 37507
rect 48557 37549 48687 37588
rect 48557 37493 48594 37549
rect 48650 37493 48687 37549
rect 25313 37387 34090 37459
rect 30403 37386 34090 37387
rect 0 37176 1014 37376
rect 48557 37370 48687 37493
rect 51034 37515 59810 37588
rect 84666 37576 86372 38276
rect 51034 37459 51071 37515
rect 51127 37459 51251 37515
rect 51307 37459 51833 37515
rect 51889 37459 52013 37515
rect 52069 37459 59810 37515
rect 51034 37387 59810 37459
rect 51034 37386 54622 37387
rect 37852 37332 48687 37370
rect 37852 37276 37889 37332
rect 37945 37276 38069 37332
rect 38125 37276 39773 37332
rect 39829 37331 48687 37332
rect 39829 37276 48594 37331
rect 37852 37275 48594 37276
rect 48650 37275 48687 37331
rect 37852 37237 48687 37275
rect 85358 37176 86372 37376
rect 0 37128 27272 37176
rect 59421 37128 86372 37176
rect 0 37055 86372 37128
rect 0 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 34282 37055
rect 34338 36999 34493 37055
rect 34549 36999 34705 37055
rect 34761 36999 34916 37055
rect 34972 36999 38328 37055
rect 38384 36999 38539 37055
rect 38595 36999 38750 37055
rect 38806 36999 40251 37055
rect 40307 36999 40431 37055
rect 40487 36999 43788 37055
rect 43844 36999 43999 37055
rect 44055 36999 44211 37055
rect 44267 36999 44422 37055
rect 44478 36999 50161 37055
rect 50217 36999 50372 37055
rect 50428 36999 50584 37055
rect 50640 36999 50795 37055
rect 50851 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 86372 37055
rect 0 36927 86372 36999
rect 0 36876 27272 36927
rect 30403 36926 54622 36927
rect 59421 36876 86372 36927
rect 0 36676 1014 36876
rect 37852 36779 48687 36817
rect 37852 36778 48594 36779
rect 37852 36722 37889 36778
rect 37945 36722 38069 36778
rect 38125 36722 39773 36778
rect 39829 36723 48594 36778
rect 48650 36723 48687 36779
rect 39829 36722 48687 36723
rect 37852 36684 48687 36722
rect 25313 36595 34090 36668
rect 25313 36588 33817 36595
rect 25313 36532 33055 36588
rect 33111 36532 33235 36588
rect 33291 36539 33817 36588
rect 33873 36539 33997 36595
rect 34053 36539 34090 36595
rect 33291 36532 34090 36539
rect 0 35776 1706 36476
rect 25313 36466 34090 36532
rect 36640 36547 40085 36586
rect 36640 36491 36676 36547
rect 36732 36491 39992 36547
rect 40048 36491 40085 36547
rect 36640 36453 40085 36491
rect 48557 36561 48687 36684
rect 85358 36676 86372 36876
rect 48557 36505 48594 36561
rect 48650 36505 48687 36561
rect 48557 36466 48687 36505
rect 51034 36595 59810 36668
rect 51034 36539 51071 36595
rect 51127 36539 51251 36595
rect 51307 36539 51833 36595
rect 51889 36539 52013 36595
rect 52069 36539 59810 36595
rect 51034 36466 59810 36539
rect 36648 36452 40041 36453
rect 25313 36218 59810 36228
rect 25313 36162 26838 36218
rect 26894 36162 26962 36218
rect 27018 36162 27086 36218
rect 27142 36162 59810 36218
rect 25313 36155 59810 36162
rect 25313 36099 29580 36155
rect 29636 36099 29791 36155
rect 29847 36099 30003 36155
rect 30059 36099 30214 36155
rect 30270 36099 30852 36155
rect 30908 36099 31063 36155
rect 31119 36099 31274 36155
rect 31330 36099 31484 36155
rect 31540 36099 31695 36155
rect 31751 36099 31907 36155
rect 31963 36099 32118 36155
rect 32174 36099 32328 36155
rect 32384 36099 32539 36155
rect 32595 36099 32750 36155
rect 32806 36099 35218 36155
rect 35274 36099 35428 36155
rect 35484 36099 35639 36155
rect 35695 36099 35851 36155
rect 35907 36099 36062 36155
rect 36118 36099 36272 36155
rect 36328 36099 39050 36155
rect 39106 36099 39230 36155
rect 39286 36099 44832 36155
rect 44888 36099 45043 36155
rect 45099 36099 45254 36155
rect 45310 36099 48836 36155
rect 48892 36099 49046 36155
rect 49102 36099 49257 36155
rect 49313 36099 49469 36155
rect 49525 36099 49680 36155
rect 49736 36099 49890 36155
rect 49946 36099 52314 36155
rect 52370 36099 52525 36155
rect 52581 36099 52736 36155
rect 52792 36099 52946 36155
rect 53002 36099 53157 36155
rect 53213 36099 53369 36155
rect 53425 36099 53580 36155
rect 53636 36099 53790 36155
rect 53846 36099 54001 36155
rect 54057 36099 54212 36155
rect 54268 36099 54853 36155
rect 54909 36099 55064 36155
rect 55120 36099 55276 36155
rect 55332 36099 55487 36155
rect 55543 36099 59810 36155
rect 25313 36094 59810 36099
rect 25313 36038 26838 36094
rect 26894 36038 26962 36094
rect 27018 36038 27086 36094
rect 27142 36038 59810 36094
rect 25313 36027 59810 36038
rect 30403 36026 54622 36027
rect 36863 35881 37743 35920
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 0 35126 24920 35326
rect 0 35016 1014 35126
rect 0 34962 25085 35016
rect 0 34940 27830 34962
rect 0 34884 27447 34940
rect 27503 34884 27571 34940
rect 27627 34884 27695 34940
rect 27751 34884 27830 34940
rect 0 34877 27830 34884
rect 0 34821 25398 34877
rect 25454 34821 25522 34877
rect 25578 34821 25646 34877
rect 25702 34821 25770 34877
rect 25826 34821 25894 34877
rect 25950 34821 27830 34877
rect 0 34816 27830 34821
rect 0 34760 27447 34816
rect 27503 34760 27571 34816
rect 27627 34760 27695 34816
rect 27751 34760 27830 34816
rect 0 34753 27830 34760
rect 0 34697 25398 34753
rect 25454 34697 25522 34753
rect 25578 34697 25646 34753
rect 25702 34697 25770 34753
rect 25826 34697 25894 34753
rect 25950 34697 27830 34753
rect 0 34692 27830 34697
rect 0 34636 27447 34692
rect 27503 34636 27571 34692
rect 27627 34636 27695 34692
rect 27751 34636 27830 34692
rect 0 34629 27830 34636
rect 0 34573 25398 34629
rect 25454 34573 25522 34629
rect 25578 34573 25646 34629
rect 25702 34573 25770 34629
rect 25826 34573 25894 34629
rect 25950 34573 27830 34629
rect 0 34568 27830 34573
rect 0 34536 27447 34568
rect 24942 34512 27447 34536
rect 27503 34512 27571 34568
rect 27627 34512 27695 34568
rect 27751 34512 27830 34568
rect 24942 34490 27830 34512
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 34011 27214 34124
rect 0 33955 26859 34011
rect 26915 33955 27071 34011
rect 27127 33955 27214 34011
rect 0 33793 27214 33955
rect 36863 33927 37743 35825
rect 84666 35776 86372 36476
rect 60549 35298 60639 35370
rect 83360 35298 86372 35326
rect 60549 35158 86372 35298
rect 60549 35086 60639 35158
rect 83360 35126 86372 35158
rect 85358 35016 86372 35126
rect 61311 34962 86372 35016
rect 60510 34536 86372 34962
rect 60510 34490 61754 34536
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 57908 34011 86372 34124
rect 57908 33955 57996 34011
rect 58052 33955 58208 34011
rect 58264 33955 86372 34011
rect 0 33737 26859 33793
rect 26915 33737 27071 33793
rect 27127 33737 27214 33793
rect 0 33576 27214 33737
rect 0 33520 26859 33576
rect 26915 33520 27071 33576
rect 27127 33520 27214 33576
rect 0 33358 27214 33520
rect 0 33302 26859 33358
rect 26915 33302 27071 33358
rect 27127 33302 27214 33358
rect 0 33140 27214 33302
rect 57908 33793 86372 33955
rect 57908 33737 57996 33793
rect 58052 33737 58208 33793
rect 58264 33737 86372 33793
rect 57908 33576 86372 33737
rect 57908 33520 57996 33576
rect 58052 33520 58208 33576
rect 58264 33520 86372 33576
rect 57908 33358 86372 33520
rect 57908 33302 57996 33358
rect 58052 33302 58208 33358
rect 58264 33302 86372 33358
rect 0 33084 26859 33140
rect 26915 33084 27071 33140
rect 27127 33084 27214 33140
rect 0 32922 27214 33084
rect 0 32866 26859 32922
rect 26915 32866 27071 32922
rect 27127 32866 27214 32922
rect 0 32705 27214 32866
rect 0 32649 26859 32705
rect 26915 32649 27071 32705
rect 27127 32649 27214 32705
rect 0 32487 27214 32649
rect 0 32431 26859 32487
rect 26915 32431 27071 32487
rect 27127 32431 27214 32487
rect 0 32318 27214 32431
rect 27387 33141 28929 33263
rect 27387 33085 27474 33141
rect 27530 33085 27686 33141
rect 27742 33085 28929 33141
rect 27387 32923 28929 33085
rect 27387 32867 27474 32923
rect 27530 32867 27686 32923
rect 27742 32867 28929 32923
rect 27387 32705 28929 32867
rect 27387 32649 27474 32705
rect 27530 32649 27686 32705
rect 27742 32649 28929 32705
rect 27387 32487 28929 32649
rect 27387 32431 27474 32487
rect 27530 32431 27686 32487
rect 27742 32431 28929 32487
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 27387 32311 28929 32431
rect 56135 33141 57736 33263
rect 56135 33085 57381 33141
rect 57437 33085 57593 33141
rect 57649 33085 57736 33141
rect 56135 32923 57736 33085
rect 56135 32867 57381 32923
rect 57437 32867 57593 32923
rect 57649 32867 57736 32923
rect 56135 32705 57736 32867
rect 56135 32649 57381 32705
rect 57437 32649 57593 32705
rect 57649 32649 57736 32705
rect 56135 32487 57736 32649
rect 56135 32431 57381 32487
rect 57437 32431 57593 32487
rect 57649 32431 57736 32487
rect 56135 32311 57736 32431
rect 57908 33140 86372 33302
rect 57908 33084 57996 33140
rect 58052 33084 58208 33140
rect 58264 33084 86372 33140
rect 57908 32922 86372 33084
rect 57908 32866 57996 32922
rect 58052 32866 58208 32922
rect 58264 32866 86372 32922
rect 57908 32705 86372 32866
rect 57908 32649 57996 32705
rect 58052 32649 58208 32705
rect 58264 32649 86372 32705
rect 57908 32487 86372 32649
rect 57908 32431 57996 32487
rect 58052 32431 58208 32487
rect 58264 32431 86372 32487
rect 57908 32315 86372 32431
rect 57908 32199 58351 32315
rect 26772 32088 58351 32199
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 26772 31870 58351 32032
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 26772 31652 58351 31814
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 26772 31486 58351 31596
rect 25293 31252 28929 31352
rect 25293 31248 27474 31252
rect 25293 31192 25398 31248
rect 25454 31192 25522 31248
rect 25578 31192 25646 31248
rect 25702 31192 25770 31248
rect 25826 31192 25894 31248
rect 25950 31196 27474 31248
rect 27530 31196 27686 31252
rect 27742 31196 28929 31252
rect 25950 31192 28929 31196
rect 25293 31124 28929 31192
rect 25293 31068 25398 31124
rect 25454 31068 25522 31124
rect 25578 31068 25646 31124
rect 25702 31068 25770 31124
rect 25826 31068 25894 31124
rect 25950 31068 28929 31124
rect 25293 31034 28929 31068
rect 25293 31000 27474 31034
rect 25293 30944 25398 31000
rect 25454 30944 25522 31000
rect 25578 30944 25646 31000
rect 25702 30944 25770 31000
rect 25826 30944 25894 31000
rect 25950 30978 27474 31000
rect 27530 30978 27686 31034
rect 27742 30978 28929 31034
rect 25950 30944 28929 30978
rect 25293 30816 28929 30944
rect 25293 30793 27474 30816
rect 25293 30737 25398 30793
rect 25454 30737 25522 30793
rect 25578 30737 25646 30793
rect 25702 30737 25770 30793
rect 25826 30737 25894 30793
rect 25950 30760 27474 30793
rect 27530 30760 27686 30816
rect 27742 30760 28929 30816
rect 25950 30737 28929 30760
rect 25293 30669 28929 30737
rect 25293 30613 25398 30669
rect 25454 30613 25522 30669
rect 25578 30613 25646 30669
rect 25702 30613 25770 30669
rect 25826 30613 25894 30669
rect 25950 30613 28929 30669
rect 25293 30598 28929 30613
rect 25293 30545 27474 30598
rect 25293 30489 25398 30545
rect 25454 30489 25522 30545
rect 25578 30489 25646 30545
rect 25702 30489 25770 30545
rect 25826 30489 25894 30545
rect 25950 30542 27474 30545
rect 27530 30542 27686 30598
rect 27742 30542 28929 30598
rect 25950 30489 28929 30542
rect 25293 30443 28929 30489
rect 56186 31298 59524 31352
rect 56186 31252 58873 31298
rect 56186 31196 57381 31252
rect 57437 31196 57593 31252
rect 57649 31242 58873 31252
rect 58929 31242 58997 31298
rect 59053 31242 59121 31298
rect 59177 31242 59245 31298
rect 59301 31242 59369 31298
rect 59425 31242 59524 31298
rect 57649 31196 59524 31242
rect 56186 31174 59524 31196
rect 56186 31118 58873 31174
rect 58929 31118 58997 31174
rect 59053 31118 59121 31174
rect 59177 31118 59245 31174
rect 59301 31118 59369 31174
rect 59425 31118 59524 31174
rect 56186 31050 59524 31118
rect 56186 31034 58873 31050
rect 56186 30978 57381 31034
rect 57437 30978 57593 31034
rect 57649 30994 58873 31034
rect 58929 30994 58997 31050
rect 59053 30994 59121 31050
rect 59177 30994 59245 31050
rect 59301 30994 59369 31050
rect 59425 30994 59524 31050
rect 57649 30978 59524 30994
rect 56186 30853 59524 30978
rect 56186 30816 58873 30853
rect 56186 30760 57381 30816
rect 57437 30760 57593 30816
rect 57649 30797 58873 30816
rect 58929 30797 58997 30853
rect 59053 30797 59121 30853
rect 59177 30797 59245 30853
rect 59301 30797 59369 30853
rect 59425 30797 59524 30853
rect 57649 30760 59524 30797
rect 56186 30729 59524 30760
rect 56186 30673 58873 30729
rect 58929 30673 58997 30729
rect 59053 30673 59121 30729
rect 59177 30673 59245 30729
rect 59301 30673 59369 30729
rect 59425 30673 59524 30729
rect 56186 30605 59524 30673
rect 56186 30598 58873 30605
rect 56186 30542 57381 30598
rect 57437 30542 57593 30598
rect 57649 30549 58873 30598
rect 58929 30549 58997 30605
rect 59053 30549 59121 30605
rect 59177 30549 59245 30605
rect 59301 30549 59369 30605
rect 59425 30549 59524 30605
rect 57649 30542 59524 30549
rect 56186 30443 59524 30542
rect 26772 29968 58351 30105
rect 26772 29912 26859 29968
rect 26915 29912 27071 29968
rect 27127 29912 57996 29968
rect 58052 29912 58208 29968
rect 58264 29912 58351 29968
rect 26772 29750 58351 29912
rect 26772 29714 26859 29750
rect 0 29694 26859 29714
rect 26915 29694 27071 29750
rect 27127 29694 57996 29750
rect 58052 29694 58208 29750
rect 58264 29714 58351 29750
rect 84666 29714 86372 32315
rect 58264 29694 86372 29714
rect 0 29533 86372 29694
rect 0 29477 26859 29533
rect 26915 29477 27071 29533
rect 27127 29477 57996 29533
rect 58052 29477 58208 29533
rect 58264 29477 86372 29533
rect 0 29430 86372 29477
rect 26772 29315 58351 29430
rect 26772 29259 26859 29315
rect 26915 29259 27071 29315
rect 27127 29259 57996 29315
rect 58052 29259 58208 29315
rect 58264 29259 58351 29315
rect 26772 29098 58351 29259
rect 26772 29042 26859 29098
rect 26915 29042 27071 29098
rect 27127 29042 57996 29098
rect 58052 29042 58208 29098
rect 58264 29042 58351 29098
rect 26772 28880 58351 29042
rect 26772 28824 26859 28880
rect 26915 28824 27071 28880
rect 27127 28824 57996 28880
rect 58052 28824 58208 28880
rect 58264 28824 58351 28880
rect 26772 28662 58351 28824
rect 26772 28606 26859 28662
rect 26915 28606 27071 28662
rect 27127 28606 57996 28662
rect 58052 28606 58208 28662
rect 58264 28606 58351 28662
rect 26772 28444 58351 28606
rect 0 28282 26070 28416
rect 0 28226 25404 28282
rect 25460 28226 25528 28282
rect 25584 28226 25652 28282
rect 25708 28226 25776 28282
rect 25832 28226 25900 28282
rect 25956 28226 26070 28282
rect 0 28158 26070 28226
rect 0 28102 25404 28158
rect 25460 28102 25528 28158
rect 25584 28102 25652 28158
rect 25708 28102 25776 28158
rect 25832 28102 25900 28158
rect 25956 28102 26070 28158
rect 0 28034 26070 28102
rect 0 27978 25404 28034
rect 25460 27978 25528 28034
rect 25584 27978 25652 28034
rect 25708 27978 25776 28034
rect 25832 27978 25900 28034
rect 25956 27978 26070 28034
rect 0 27910 26070 27978
rect 0 27854 25404 27910
rect 25460 27854 25528 27910
rect 25584 27854 25652 27910
rect 25708 27854 25776 27910
rect 25832 27854 25900 27910
rect 25956 27854 26070 27910
rect 0 27786 26070 27854
rect 0 27730 25404 27786
rect 25460 27730 25528 27786
rect 25584 27730 25652 27786
rect 25708 27730 25776 27786
rect 25832 27730 25900 27786
rect 25956 27730 26070 27786
rect 0 27662 26070 27730
rect 0 27606 25404 27662
rect 25460 27606 25528 27662
rect 25584 27606 25652 27662
rect 25708 27606 25776 27662
rect 25832 27606 25900 27662
rect 25956 27606 26070 27662
rect 0 27538 26070 27606
rect 0 27482 25404 27538
rect 25460 27482 25528 27538
rect 25584 27482 25652 27538
rect 25708 27482 25776 27538
rect 25832 27482 25900 27538
rect 25956 27482 26070 27538
rect 0 27414 26070 27482
rect 0 27358 25404 27414
rect 25460 27358 25528 27414
rect 25584 27358 25652 27414
rect 25708 27358 25776 27414
rect 25832 27358 25900 27414
rect 25956 27358 26070 27414
rect 26772 28388 26859 28444
rect 26915 28388 27071 28444
rect 27127 28388 57996 28444
rect 58052 28388 58208 28444
rect 58264 28388 58351 28444
rect 26772 28227 58351 28388
rect 26772 28171 26859 28227
rect 26915 28171 27071 28227
rect 27127 28171 57996 28227
rect 58052 28171 58208 28227
rect 58264 28171 58351 28227
rect 26772 28009 58351 28171
rect 26772 27953 26859 28009
rect 26915 27953 27071 28009
rect 27127 27953 57996 28009
rect 58052 27953 58208 28009
rect 58264 27953 58351 28009
rect 26772 27792 58351 27953
rect 26772 27736 26859 27792
rect 26915 27736 27071 27792
rect 27127 27736 57996 27792
rect 58052 27736 58208 27792
rect 58264 27736 58351 27792
rect 26772 27574 58351 27736
rect 26772 27518 26859 27574
rect 26915 27518 27071 27574
rect 27127 27518 57996 27574
rect 58052 27518 58208 27574
rect 58264 27518 58351 27574
rect 26772 27382 58351 27518
rect 58785 28272 86372 28416
rect 58785 28216 58859 28272
rect 58915 28216 58983 28272
rect 59039 28216 59107 28272
rect 59163 28216 59231 28272
rect 59287 28216 59355 28272
rect 59411 28216 86372 28272
rect 58785 28148 86372 28216
rect 58785 28092 58859 28148
rect 58915 28092 58983 28148
rect 59039 28092 59107 28148
rect 59163 28092 59231 28148
rect 59287 28092 59355 28148
rect 59411 28092 86372 28148
rect 58785 28024 86372 28092
rect 58785 27968 58859 28024
rect 58915 27968 58983 28024
rect 59039 27968 59107 28024
rect 59163 27968 59231 28024
rect 59287 27968 59355 28024
rect 59411 27968 86372 28024
rect 58785 27900 86372 27968
rect 58785 27844 58859 27900
rect 58915 27844 58983 27900
rect 59039 27844 59107 27900
rect 59163 27844 59231 27900
rect 59287 27844 59355 27900
rect 59411 27844 86372 27900
rect 58785 27776 86372 27844
rect 58785 27720 58859 27776
rect 58915 27720 58983 27776
rect 59039 27720 59107 27776
rect 59163 27720 59231 27776
rect 59287 27720 59355 27776
rect 59411 27720 86372 27776
rect 58785 27652 86372 27720
rect 58785 27596 58859 27652
rect 58915 27596 58983 27652
rect 59039 27596 59107 27652
rect 59163 27596 59231 27652
rect 59287 27596 59355 27652
rect 59411 27596 86372 27652
rect 58785 27528 86372 27596
rect 58785 27472 58859 27528
rect 58915 27472 58983 27528
rect 59039 27472 59107 27528
rect 59163 27472 59231 27528
rect 59287 27472 59355 27528
rect 59411 27472 86372 27528
rect 58785 27404 86372 27472
rect 0 27290 26070 27358
rect 0 27234 25404 27290
rect 25460 27234 25528 27290
rect 25584 27234 25652 27290
rect 25708 27234 25776 27290
rect 25832 27234 25900 27290
rect 25956 27234 26070 27290
rect 0 27166 26070 27234
rect 0 27110 25404 27166
rect 25460 27110 25528 27166
rect 25584 27110 25652 27166
rect 25708 27110 25776 27166
rect 25832 27110 25900 27166
rect 25956 27110 26070 27166
rect 0 27042 26070 27110
rect 0 26986 25404 27042
rect 25460 26986 25528 27042
rect 25584 26986 25652 27042
rect 25708 26986 25776 27042
rect 25832 26986 25900 27042
rect 25956 26986 26070 27042
rect 0 26918 26070 26986
rect 0 26862 25404 26918
rect 25460 26862 25528 26918
rect 25584 26862 25652 26918
rect 25708 26862 25776 26918
rect 25832 26862 25900 26918
rect 25956 26890 26070 26918
rect 58785 27348 58859 27404
rect 58915 27348 58983 27404
rect 59039 27348 59107 27404
rect 59163 27348 59231 27404
rect 59287 27348 59355 27404
rect 59411 27348 86372 27404
rect 58785 27280 86372 27348
rect 58785 27224 58859 27280
rect 58915 27224 58983 27280
rect 59039 27224 59107 27280
rect 59163 27224 59231 27280
rect 59287 27224 59355 27280
rect 59411 27224 86372 27280
rect 58785 27156 86372 27224
rect 58785 27100 58859 27156
rect 58915 27100 58983 27156
rect 59039 27100 59107 27156
rect 59163 27100 59231 27156
rect 59287 27100 59355 27156
rect 59411 27100 86372 27156
rect 58785 27032 86372 27100
rect 58785 26976 58859 27032
rect 58915 26976 58983 27032
rect 59039 26976 59107 27032
rect 59163 26976 59231 27032
rect 59287 26976 59355 27032
rect 59411 26976 86372 27032
rect 58785 26908 86372 26976
rect 58785 26890 58859 26908
rect 25956 26862 27828 26890
rect 0 26799 27828 26862
rect 0 26794 27474 26799
rect 0 26738 25404 26794
rect 25460 26738 25528 26794
rect 25584 26738 25652 26794
rect 25708 26738 25776 26794
rect 25832 26738 25900 26794
rect 25956 26743 27474 26794
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 25956 26738 27828 26743
rect 0 26670 27828 26738
rect 0 26614 25404 26670
rect 25460 26614 25528 26670
rect 25584 26614 25652 26670
rect 25708 26614 25776 26670
rect 25832 26614 25900 26670
rect 25956 26614 27828 26670
rect 0 26581 27828 26614
rect 0 26546 27474 26581
rect 0 26490 25404 26546
rect 25460 26490 25528 26546
rect 25584 26490 25652 26546
rect 25708 26490 25776 26546
rect 25832 26490 25900 26546
rect 25956 26525 27474 26546
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 25956 26490 27828 26525
rect 0 26435 27828 26490
rect 57295 26852 58859 26890
rect 58915 26852 58983 26908
rect 59039 26852 59107 26908
rect 59163 26852 59231 26908
rect 59287 26852 59355 26908
rect 59411 26852 86372 26908
rect 57295 26799 86372 26852
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26784 86372 26799
rect 57649 26743 58859 26784
rect 57295 26728 58859 26743
rect 58915 26728 58983 26784
rect 59039 26728 59107 26784
rect 59163 26728 59231 26784
rect 59287 26728 59355 26784
rect 59411 26728 86372 26784
rect 57295 26660 86372 26728
rect 57295 26604 58859 26660
rect 58915 26604 58983 26660
rect 59039 26604 59107 26660
rect 59163 26604 59231 26660
rect 59287 26604 59355 26660
rect 59411 26604 86372 26660
rect 57295 26581 86372 26604
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26536 86372 26581
rect 57649 26525 58859 26536
rect 57295 26480 58859 26525
rect 58915 26480 58983 26536
rect 59039 26480 59107 26536
rect 59163 26480 59231 26536
rect 59287 26480 59355 26536
rect 59411 26480 86372 26536
rect 57295 26435 86372 26480
rect 1271 26434 27828 26435
rect 61530 26434 84717 26435
rect 1954 26433 2279 26434
rect 12754 26433 13079 26434
rect 61530 26433 61855 26434
rect 72330 26433 72655 26434
rect 23828 26286 26642 26324
rect 23828 26126 26450 26286
rect 26610 26126 26642 26286
rect 23828 26109 26642 26126
rect 23828 25967 26285 26002
rect 23828 25807 26092 25967
rect 26252 25807 26285 25967
rect 23828 25787 26285 25807
rect 23828 25647 25949 25681
rect 23828 25487 25756 25647
rect 25916 25487 25949 25647
rect 23828 25466 25949 25487
rect 23828 25328 25614 25359
rect 23828 25168 25421 25328
rect 25581 25168 25614 25328
rect 23828 25144 25614 25168
rect 27382 25028 29699 25208
rect 27382 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 29699 25028
rect 27382 24810 29699 24972
rect 27382 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 29699 24810
rect 23828 24637 25274 24667
rect 23828 24477 25081 24637
rect 25241 24477 25274 24637
rect 27382 24526 29699 24754
rect 23828 24452 25274 24477
rect 23828 24316 24935 24345
rect 23828 24156 24744 24316
rect 24904 24156 24935 24316
rect 23828 24130 24935 24156
rect 26770 24227 58348 24278
rect 26770 24171 26858 24227
rect 27122 24171 58348 24227
rect 26770 24085 58348 24171
rect 26770 24029 26858 24085
rect 27122 24075 58348 24085
rect 27122 24029 57994 24075
rect 23828 23995 24607 24024
rect 0 23380 1706 23938
rect 23828 23835 24416 23995
rect 24576 23835 24607 23995
rect 23828 23809 24607 23835
rect 26770 23943 57994 24029
rect 26770 23887 26858 23943
rect 27122 23887 57994 23943
rect 26770 23801 57994 23887
rect 26770 23745 26858 23801
rect 27122 23745 57994 23801
rect 24047 23673 24227 23683
rect 24047 23513 24057 23673
rect 24217 23513 24227 23673
rect 24047 23503 24227 23513
rect 26770 23659 57994 23745
rect 26770 23603 26858 23659
rect 27122 23603 57994 23659
rect 26770 23517 57994 23603
rect 26770 23461 26858 23517
rect 27122 23461 57994 23517
rect 26770 23380 57994 23461
rect 0 23375 57994 23380
rect 0 23319 26858 23375
rect 27122 23370 57994 23375
rect 27122 23319 27214 23370
rect 0 23233 27214 23319
rect 0 23177 26858 23233
rect 27122 23177 27214 23233
rect 0 23091 27214 23177
rect 0 23035 26858 23091
rect 27122 23035 27214 23091
rect 0 22938 27214 23035
rect 27387 22936 57677 23199
rect 57908 23187 57994 23370
rect 58258 23380 58348 24075
rect 84666 23380 86372 23938
rect 58258 23187 86372 23380
rect 57908 22938 86372 23187
rect 57908 22937 83763 22938
rect 27387 22282 27475 22936
rect 0 22048 27475 22282
rect 27739 22923 57677 22936
rect 27739 22291 57363 22923
rect 27739 22048 27826 22291
rect 0 21827 27826 22048
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 22035 57363 22291
rect 57627 22282 57677 22923
rect 57627 22035 86372 22282
rect 56078 21827 86372 22035
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 20570 86372 20739
rect 0 20410 26924 20570
rect 27084 20410 58048 20570
rect 58208 20410 86372 20570
rect 0 20226 86372 20410
rect 0 20066 26924 20226
rect 27084 20066 58048 20226
rect 58208 20066 86372 20226
rect 0 19969 86372 20066
rect 0 18016 24250 19969
rect 26435 19692 29403 19731
rect 26435 19532 26465 19692
rect 26625 19532 29403 19692
rect 26435 19502 29403 19532
rect 55720 19502 58817 19731
rect 26077 19347 29403 19391
rect 26077 19187 26107 19347
rect 26267 19187 29403 19347
rect 26077 19162 29403 19187
rect 55720 19162 59177 19391
rect 25742 19027 29403 19051
rect 25742 18867 25771 19027
rect 25931 18867 29403 19027
rect 25742 18822 29403 18867
rect 55720 18822 59515 19051
rect 25406 18684 29403 18711
rect 25406 18524 25434 18684
rect 25594 18524 29403 18684
rect 25406 18482 29403 18524
rect 55720 18482 59846 18711
rect 25066 18350 29403 18371
rect 25066 18190 25094 18350
rect 25254 18190 29403 18350
rect 25066 18142 29403 18190
rect 55720 18142 60184 18371
rect 24730 17977 29403 18031
rect 24730 17817 24757 17977
rect 24917 17817 29403 17977
rect 24730 17802 29403 17817
rect 55720 17802 60525 18031
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 24401 17656 29403 17691
rect 24401 17496 24429 17656
rect 24589 17496 29403 17656
rect 24401 17462 29403 17496
rect 55720 17462 60855 17691
rect 24042 17317 29403 17351
rect 24042 17157 24069 17317
rect 24229 17157 29403 17317
rect 24042 17122 29403 17157
rect 55720 17122 61205 17351
rect 61807 16784 86372 17730
rect 46982 16678 86372 16784
rect 46982 16622 57381 16678
rect 57437 16622 57593 16678
rect 57649 16622 86372 16678
rect 24111 16597 27828 16598
rect 0 16470 27828 16597
rect 0 16414 27474 16470
rect 27530 16414 27686 16470
rect 27742 16414 27828 16470
rect 0 16253 27828 16414
rect 0 16197 27474 16253
rect 27530 16197 27686 16253
rect 27742 16197 27828 16253
rect 0 16035 27828 16197
rect 0 15979 27474 16035
rect 27530 15979 27686 16035
rect 27742 15979 27828 16035
rect 0 15818 27828 15979
rect 0 15762 27474 15818
rect 27530 15762 27686 15818
rect 27742 15762 27828 15818
rect 0 15600 27828 15762
rect 0 15544 27474 15600
rect 27530 15544 27686 15600
rect 27742 15544 27828 15600
rect 0 15382 27828 15544
rect 0 15326 27474 15382
rect 27530 15326 27686 15382
rect 27742 15326 27828 15382
rect 0 15164 27828 15326
rect 0 15108 27474 15164
rect 27530 15108 27686 15164
rect 27742 15108 27828 15164
rect 0 15015 27828 15108
rect 46982 16461 86372 16622
rect 46982 16405 57381 16461
rect 57437 16405 57593 16461
rect 57649 16405 86372 16461
rect 46982 16243 86372 16405
rect 46982 16187 57381 16243
rect 57437 16187 57593 16243
rect 57649 16187 86372 16243
rect 46982 16026 86372 16187
rect 46982 15970 57381 16026
rect 57437 15970 57593 16026
rect 57649 15970 86372 16026
rect 46982 15808 86372 15970
rect 46982 15752 57381 15808
rect 57437 15752 57593 15808
rect 57649 15752 86372 15808
rect 46982 15590 86372 15752
rect 46982 15534 57381 15590
rect 57437 15534 57593 15590
rect 57649 15534 86372 15590
rect 46982 15372 86372 15534
rect 46982 15316 57381 15372
rect 57437 15316 57593 15372
rect 57649 15316 86372 15372
rect 46982 15155 86372 15316
rect 46982 15099 57381 15155
rect 57437 15099 57593 15155
rect 57649 15099 86372 15155
rect 46982 15015 86372 15099
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14947 51760 14966
rect 0 14891 27474 14947
rect 27530 14891 27686 14947
rect 27742 14936 51760 14947
rect 57295 14937 86372 14968
rect 27742 14891 47683 14936
rect 0 14729 47683 14891
rect 0 14673 27474 14729
rect 27530 14673 27686 14729
rect 27742 14673 47683 14729
rect 0 14512 47683 14673
rect 0 14456 27474 14512
rect 27530 14456 27686 14512
rect 27742 14491 47683 14512
rect 57295 14881 57381 14937
rect 57437 14881 57593 14937
rect 57649 14881 86372 14937
rect 57295 14720 86372 14881
rect 57295 14664 57381 14720
rect 57437 14664 57593 14720
rect 57649 14664 86372 14720
rect 27742 14456 45977 14491
rect 0 14329 45977 14456
rect 0 14328 24250 14329
rect 27387 14231 45977 14329
rect 57295 14328 86372 14664
rect 57295 14327 83763 14328
rect 24047 14178 27214 14179
rect 0 14119 27214 14178
rect 0 14063 26859 14119
rect 26915 14063 27071 14119
rect 27127 14063 27214 14119
rect 0 13902 27214 14063
rect 0 13846 26859 13902
rect 26915 13846 27071 13902
rect 27127 13846 27214 13902
rect 0 13684 27214 13846
rect 0 13628 26859 13684
rect 26915 13628 27071 13684
rect 27127 13628 27214 13684
rect 0 13467 27214 13628
rect 0 13461 26859 13467
rect 0 12846 1706 13461
rect 24047 13411 26859 13461
rect 26915 13411 27071 13467
rect 27127 13411 27214 13467
rect 24047 13249 27214 13411
rect 24047 13193 26859 13249
rect 26915 13193 27071 13249
rect 27127 13193 27214 13249
rect 27387 14175 27474 14231
rect 27530 14175 27686 14231
rect 27742 14175 45977 14231
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 27387 14014 45977 14175
rect 27387 13958 27474 14014
rect 27530 13958 27686 14014
rect 27742 13958 45977 14014
rect 27387 13796 45977 13958
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13740 27474 13796
rect 27530 13740 27686 13796
rect 27742 13760 45977 13796
rect 50228 13790 86372 13866
rect 27742 13740 49775 13760
rect 27387 13578 49775 13740
rect 27387 13522 27474 13578
rect 27530 13522 27686 13578
rect 27742 13522 49775 13578
rect 27387 13361 49775 13522
rect 27387 13305 27474 13361
rect 27530 13305 27686 13361
rect 27742 13305 49775 13361
rect 27387 13245 49775 13305
rect 29478 13243 49775 13245
rect 24047 13031 27214 13193
rect 41493 13078 49775 13243
rect 50228 13734 57996 13790
rect 58052 13734 58208 13790
rect 58264 13734 86372 13790
rect 50228 13573 86372 13734
rect 50228 13517 57996 13573
rect 58052 13517 58208 13573
rect 58264 13517 86372 13573
rect 50228 13461 86372 13517
rect 50228 13355 58421 13461
rect 50228 13299 57996 13355
rect 58052 13299 58208 13355
rect 58264 13299 58421 13355
rect 50228 13138 58421 13299
rect 50228 13082 57996 13138
rect 58052 13082 58208 13138
rect 58264 13082 58421 13138
rect 24047 12975 26859 13031
rect 26915 12975 27071 13031
rect 27127 12975 27214 13031
rect 24047 12934 27214 12975
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12813 34761 12846
rect 0 12757 26859 12813
rect 26915 12757 27071 12813
rect 27127 12757 34761 12813
rect 0 12606 34761 12757
rect 50228 12920 58421 13082
rect 50228 12864 57996 12920
rect 58052 12864 58208 12920
rect 58264 12864 58421 12920
rect 50228 12846 58421 12864
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12702 86372 12846
rect 50228 12646 57996 12702
rect 58052 12646 58208 12702
rect 58264 12646 86372 12702
rect 50228 12606 86372 12646
rect 0 12596 86372 12606
rect 0 12540 26859 12596
rect 26915 12540 27071 12596
rect 27127 12540 86372 12596
rect 0 12484 86372 12540
rect 0 12428 57996 12484
rect 58052 12428 58208 12484
rect 58264 12428 86372 12484
rect 0 12378 86372 12428
rect 0 12322 26859 12378
rect 26915 12322 27071 12378
rect 27127 12322 86372 12378
rect 0 12267 86372 12322
rect 0 12211 57996 12267
rect 58052 12211 58208 12267
rect 58264 12211 86372 12267
rect 0 12161 86372 12211
rect 0 12105 26859 12161
rect 26915 12105 27071 12161
rect 27127 12105 86372 12161
rect 0 12049 86372 12105
rect 0 12046 57996 12049
rect 0 12036 24250 12046
rect 26772 11993 57996 12046
rect 58052 11993 58208 12049
rect 58264 12036 86372 12049
rect 58264 12035 84999 12036
rect 58264 11993 58351 12035
rect 26772 11844 58351 11993
rect 29478 11832 58351 11844
rect 29478 11776 57996 11832
rect 58052 11776 58208 11832
rect 58264 11776 58351 11832
rect 29478 11697 58351 11776
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 11406 27828 11491
rect 0 11350 27474 11406
rect 27530 11350 27686 11406
rect 27742 11350 27828 11406
rect 0 11189 27828 11350
rect 0 11133 27474 11189
rect 27530 11133 27686 11189
rect 27742 11133 27828 11189
rect 0 10971 27828 11133
rect 0 10915 27474 10971
rect 27530 10915 27686 10971
rect 27742 10915 27828 10971
rect 0 10753 27828 10915
rect 29478 10756 41353 11697
rect 0 10697 27474 10753
rect 27530 10697 27686 10753
rect 27742 10697 27828 10753
rect 0 10535 27828 10697
rect 0 10479 27474 10535
rect 27530 10479 27686 10535
rect 27742 10479 27828 10535
rect 0 10318 27828 10479
rect 0 10262 27474 10318
rect 27530 10262 27686 10318
rect 27742 10262 27828 10318
rect 0 10176 27828 10262
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 2249 9943 29220 10031
rect 34904 9972 41353 10756
rect 42261 11491 57736 11527
rect 61825 11491 86372 11493
rect 42261 11406 86372 11491
rect 42261 11350 57381 11406
rect 57437 11350 57593 11406
rect 57649 11350 86372 11406
rect 42261 11189 86372 11350
rect 42261 11133 57381 11189
rect 57437 11133 57593 11189
rect 57649 11133 86372 11189
rect 42261 10971 86372 11133
rect 42261 10915 57381 10971
rect 57437 10915 57593 10971
rect 57649 10915 86372 10971
rect 42261 10753 86372 10915
rect 42261 10740 57381 10753
rect 57295 10697 57381 10740
rect 57437 10697 57593 10753
rect 57649 10697 86372 10753
rect 57295 10535 86372 10697
rect 57295 10479 57381 10535
rect 57437 10479 57593 10535
rect 57649 10479 86372 10535
rect 24047 9515 28729 9516
rect 0 9514 1014 9515
rect 2226 9514 28729 9515
rect 0 9407 28729 9514
rect 0 9351 26859 9407
rect 26915 9351 27071 9407
rect 27127 9351 28729 9407
rect 0 9190 28729 9351
rect 29132 9301 29220 9943
rect 41857 9502 51430 10420
rect 57295 10318 86372 10479
rect 57295 10262 57381 10318
rect 57437 10262 57593 10318
rect 57649 10262 86372 10318
rect 51750 10097 54952 10185
rect 57295 10176 86372 10262
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 51750 9971 51838 10097
rect 51750 9811 51766 9971
rect 51822 9811 51838 9971
rect 54864 10028 54952 10097
rect 54864 9940 83193 10028
rect 51750 9791 51838 9811
rect 58688 9681 61743 9777
rect 57909 9515 62278 9516
rect 57909 9514 72434 9515
rect 72602 9514 83234 9515
rect 85358 9514 86372 9515
rect 29132 9213 41655 9301
rect 0 9134 26859 9190
rect 26915 9134 27071 9190
rect 27127 9134 28729 9190
rect 0 8972 28729 9134
rect 0 8916 26859 8972
rect 26915 8916 27071 8972
rect 27127 8916 28729 8972
rect 0 8754 28729 8916
rect 41567 8971 41655 9213
rect 41857 9165 55482 9502
rect 50922 9012 55482 9165
rect 57909 9407 86372 9514
rect 57909 9351 57996 9407
rect 58052 9351 58208 9407
rect 58264 9351 86372 9407
rect 57909 9190 86372 9351
rect 57909 9134 57996 9190
rect 58052 9134 58208 9190
rect 58264 9134 86372 9190
rect 41567 8953 50108 8971
rect 41567 8897 49897 8953
rect 50057 8897 50108 8953
rect 41567 8883 50108 8897
rect 50922 8934 57736 9012
rect 0 8698 26859 8754
rect 26915 8698 27071 8754
rect 27127 8698 28729 8754
rect 0 8536 28729 8698
rect 50922 8878 57386 8934
rect 57442 8878 57510 8934
rect 57566 8878 57634 8934
rect 57690 8878 57736 8934
rect 50922 8810 57736 8878
rect 50922 8754 57386 8810
rect 57442 8754 57510 8810
rect 57566 8754 57634 8810
rect 57690 8754 57736 8810
rect 50922 8686 57736 8754
rect 50922 8630 57386 8686
rect 57442 8630 57510 8686
rect 57566 8630 57634 8686
rect 57690 8630 57736 8686
rect 0 8480 26859 8536
rect 26915 8480 27071 8536
rect 27127 8480 28729 8536
rect 0 8319 28729 8480
rect 0 8263 26859 8319
rect 26915 8263 27071 8319
rect 27127 8263 28729 8319
rect 0 8154 28729 8263
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 28178 7652 28729 8154
rect 29513 7900 41397 8582
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 7535 27828 7595
rect 0 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 0 7317 27828 7479
rect 0 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 0 7099 27828 7261
rect 0 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 28178 7084 34622 7652
rect 0 6982 27828 7043
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 23625 6836 29058 6875
rect 23625 6780 28273 6836
rect 28329 6780 28484 6836
rect 28540 6780 28696 6836
rect 28752 6780 28907 6836
rect 28963 6780 29058 6836
rect 23625 6618 29058 6780
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 8562 57736 8630
rect 50922 8506 57386 8562
rect 57442 8506 57510 8562
rect 57566 8506 57634 8562
rect 57690 8506 57736 8562
rect 50922 8438 57736 8506
rect 50922 8382 57386 8438
rect 57442 8382 57510 8438
rect 57566 8382 57634 8438
rect 57690 8382 57736 8438
rect 50922 8314 57736 8382
rect 50922 8258 57386 8314
rect 57442 8258 57510 8314
rect 57566 8258 57634 8314
rect 57690 8258 57736 8314
rect 50922 8190 57736 8258
rect 50922 8134 57386 8190
rect 57442 8134 57510 8190
rect 57566 8134 57634 8190
rect 57690 8134 57736 8190
rect 57909 8972 86372 9134
rect 57909 8916 57996 8972
rect 58052 8916 58208 8972
rect 58264 8916 86372 8972
rect 57909 8754 86372 8916
rect 57909 8698 57996 8754
rect 58052 8698 58208 8754
rect 58264 8698 86372 8754
rect 57909 8536 86372 8698
rect 57909 8480 57996 8536
rect 58052 8480 58208 8536
rect 58264 8480 86372 8536
rect 57909 8319 86372 8480
rect 57909 8263 57996 8319
rect 58052 8263 58208 8319
rect 58264 8263 86372 8319
rect 57909 8154 86372 8263
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 8066 57736 8134
rect 50922 8010 57386 8066
rect 57442 8010 57510 8066
rect 57566 8010 57634 8066
rect 57690 8010 57736 8066
rect 50922 7942 57736 8010
rect 50922 7886 57386 7942
rect 57442 7886 57510 7942
rect 57566 7886 57634 7942
rect 57690 7886 57736 7942
rect 50922 7818 57736 7886
rect 50922 7762 57386 7818
rect 57442 7762 57510 7818
rect 57566 7762 57634 7818
rect 57690 7762 57736 7818
rect 50922 7694 57736 7762
rect 50922 7638 57386 7694
rect 57442 7638 57510 7694
rect 57566 7638 57634 7694
rect 57690 7638 57736 7694
rect 50922 7596 57736 7638
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7570 86372 7595
rect 50922 7514 57386 7570
rect 57442 7514 57510 7570
rect 57566 7514 57634 7570
rect 57690 7514 86372 7570
rect 50922 7446 86372 7514
rect 50922 7392 57386 7446
rect 34860 7390 57386 7392
rect 57442 7390 57510 7446
rect 57566 7390 57634 7446
rect 57690 7390 86372 7446
rect 34860 7322 86372 7390
rect 34860 7266 57386 7322
rect 57442 7266 57510 7322
rect 57566 7266 57634 7322
rect 57690 7266 86372 7322
rect 34860 7198 86372 7266
rect 34860 7142 57386 7198
rect 57442 7142 57510 7198
rect 57566 7142 57634 7198
rect 57690 7142 86372 7198
rect 34860 7088 86372 7142
rect 23625 6562 28273 6618
rect 28329 6562 28484 6618
rect 28540 6562 28696 6618
rect 28752 6562 28907 6618
rect 28963 6562 29058 6618
rect 34860 6592 55482 7088
rect 59309 6982 86372 7088
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 23625 6400 29058 6562
rect 23625 6344 28273 6400
rect 28329 6344 28484 6400
rect 28540 6344 28696 6400
rect 28752 6344 28907 6400
rect 28963 6344 29058 6400
rect 23625 6306 29058 6344
rect 29458 6199 41397 6573
rect 43655 6291 44077 6379
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 50922 6199 55482 6592
rect 56065 6836 62747 6875
rect 56065 6780 56160 6836
rect 56216 6780 56371 6836
rect 56427 6780 56583 6836
rect 56639 6780 56794 6836
rect 56850 6780 62747 6836
rect 56065 6618 62747 6780
rect 56065 6562 56160 6618
rect 56216 6562 56371 6618
rect 56427 6562 56583 6618
rect 56639 6562 56794 6618
rect 56850 6562 62747 6618
rect 56065 6400 62747 6562
rect 56065 6344 56160 6400
rect 56216 6344 56371 6400
rect 56427 6344 56583 6400
rect 56639 6344 56794 6400
rect 56850 6344 62747 6400
rect 56065 6306 62747 6344
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 0 6120 34622 6177
rect 0 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 34622 6120
rect 0 5902 34622 6064
rect 0 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 34622 5902
rect 0 5766 34622 5846
rect 29458 5665 34622 5766
rect 50922 6120 86372 6198
rect 50922 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 86372 6120
rect 50922 5902 86372 6064
rect 50922 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 86372 5902
rect 50922 5766 86372 5846
rect 23687 5629 27214 5630
rect 0 5539 27214 5629
rect 50922 5605 55482 5766
rect 57909 5629 62429 5630
rect 0 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27214 5539
rect 0 5321 27214 5483
rect 0 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27214 5321
rect 0 5175 27214 5265
rect 57909 5539 86372 5629
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 86372 5539
rect 57909 5321 86372 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 86372 5321
rect 57909 5175 86372 5265
rect 0 5174 24250 5175
rect 61802 5174 86372 5175
rect 0 5173 3011 5174
rect 83361 5173 86372 5174
rect 0 4515 1712 5173
rect 42928 4733 46482 4821
rect 57909 4619 62429 4621
rect 23909 4528 62429 4619
rect 23909 4515 26859 4528
rect 0 4472 26859 4515
rect 26915 4472 27071 4528
rect 27127 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4515 62429 4528
rect 84660 4515 86372 5173
rect 58264 4472 86372 4515
rect 0 4310 86372 4472
rect 0 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 86372 4310
rect 0 4166 86372 4254
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3837 61215 3875
rect 23909 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 28801 3837
rect 28857 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 61215 3837
rect 23909 3772 61215 3781
rect 0 3619 86372 3772
rect 0 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 28801 3619
rect 28857 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 86372 3619
rect 0 3524 86372 3563
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 60886 3420 86372 3524
rect 0 2854 1000 3420
rect 2212 3209 24341 3297
rect 61788 3209 66715 3297
rect 67518 3209 72448 3297
rect 72588 3209 77521 3297
rect 78321 3209 83248 3297
rect 2212 3044 83763 3066
rect 2212 2988 43800 3044
rect 43960 2988 83763 3044
rect 2212 2978 83763 2988
rect 85358 2854 86372 3420
rect 0 2822 86372 2854
rect 0 2766 48671 2822
rect 48727 2766 48795 2822
rect 48851 2766 48919 2822
rect 48975 2766 86372 2822
rect 0 2698 86372 2766
rect 0 2642 48671 2698
rect 48727 2642 48795 2698
rect 48851 2642 48919 2698
rect 48975 2642 86372 2698
rect 0 2574 86372 2642
rect 0 2518 48671 2574
rect 48727 2518 48795 2574
rect 48851 2518 48919 2574
rect 48975 2518 86372 2574
rect 0 2502 86372 2518
rect 0 2143 86372 2232
rect 0 2087 49161 2143
rect 49217 2087 49285 2143
rect 49341 2087 49409 2143
rect 49465 2087 86372 2143
rect 0 2019 86372 2087
rect 0 1963 49161 2019
rect 49217 1963 49285 2019
rect 49341 1963 49409 2019
rect 49465 1963 86372 2019
rect 0 1895 86372 1963
rect 0 1839 49161 1895
rect 49217 1839 49285 1895
rect 49341 1839 49409 1895
rect 49465 1839 86372 1895
rect 0 1232 86372 1839
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
use 64x8M8WM1_PWR_64x8m81  64x8M8WM1_PWR_64x8m81_0
timestamp 1762296095
transform 1 0 0 0 1 0
box 1912 6592 83548 35222
use control_512x8_64x8m81  control_512x8_64x8m81_0
timestamp 1762296095
transform 1 0 27533 0 1 4711
box -3624 -1833 31790 30125
use G_ring_64x8m81  G_ring_64x8m81_0
timestamp 1762296095
transform 1 0 282 0 1 0
box 112 620 85672 45689
use GF018_64x8M8WM1_lef_64x8m81  GF018_64x8M8WM1_lef_64x8m81_0
timestamp 1762296095
transform 1 0 0 0 1 0
box 0 0 86372 46576
use lcol4_64_64x8m81  lcol4_64_64x8m81_0
timestamp 1762296095
transform 1 0 2921 0 1 5019
box -1235 -3394 22810 39307
use M1_PSUB431058998322_64x8m81  M1_PSUB431058998322_64x8m81_0
timestamp 1762296095
transform 1 0 27869 0 1 36019
box 0 0 1 1
use M1_PSUB431058998322_64x8m81  M1_PSUB431058998322_64x8m81_1
timestamp 1762296095
transform 1 0 56655 0 1 36019
box 0 0 1 1
use M1_PSUB431058998323_64x8m81  M1_PSUB431058998323_64x8m81_0
timestamp 1762296095
transform 1 0 57403 0 1 1140
box 0 0 1 1
use M1_PSUB4310589983216_64x8m81  M1_PSUB4310589983216_64x8m81_0
timestamp 1762296095
transform 1 0 34404 0 1 2512
box 0 0 1 1
use M1_PSUB4310589983220_64x8m81  M1_PSUB4310589983220_64x8m81_0
timestamp 1762296095
transform 1 0 53710 0 1 2533
box 0 0 1 1
use M1_PSUB4310589983222_64x8m81  M1_PSUB4310589983222_64x8m81_0
timestamp 1762296095
transform 1 0 27521 0 1 1140
box 0 0 1 1
use M1_PSUB4310589983223_64x8m81  M1_PSUB4310589983223_64x8m81_0
timestamp 1762296095
transform 1 0 27869 0 1 34279
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_0
timestamp 1762296095
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_1
timestamp 1762296095
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_2
timestamp 1762296095
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_3
timestamp 1762296095
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_4
timestamp 1762296095
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_5
timestamp 1762296095
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_6
timestamp 1762296095
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_7
timestamp 1762296095
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_8
timestamp 1762296095
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_64x8m81  M2_M1$$199747628_64x8m81_9
timestamp 1762296095
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M2_M1$$201260076_64x8m81  M2_M1$$201260076_64x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_64x8m81  M2_M1$$201260076_64x8m81_1
timestamp 1762296095
transform 1 0 27608 0 1 19369
box 0 0 1 1
use M2_M1$$201260076_64x8m81  M2_M1$$201260076_64x8m81_2
timestamp 1762296095
transform 1 0 26993 0 1 19369
box 0 0 1 1
use M2_M1$$201261100_64x8m81  M2_M1$$201261100_64x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_64x8m81  M2_M1$$201261100_64x8m81_1
timestamp 1762296095
transform -1 0 57515 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_64x8m81  M2_M1$$201261100_64x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 4126
box 0 0 1 1
use M2_M1$$201261100_64x8m81  M2_M1$$201261100_64x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 4126
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_0
timestamp 1762296095
transform 1 0 72743 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_1
timestamp 1762296095
transform 1 0 72293 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_2
timestamp 1762296095
transform 1 0 62228 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_3
timestamp 1762296095
transform 1 0 49986 0 1 6323
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_4
timestamp 1762296095
transform 1 0 82808 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_5
timestamp 1762296095
transform 1 0 51732 0 1 5173
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_6
timestamp 1762296095
transform 1 0 2652 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_7
timestamp 1762296095
transform 1 0 40701 0 1 3256
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_8
timestamp 1762296095
transform 1 0 23517 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_9
timestamp 1762296095
transform 1 0 13167 0 1 1663
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_10
timestamp 1762296095
transform 1 0 12717 0 1 1663
box 0 0 1 1
use M2_M1431058998324_64x8m81  M2_M1431058998324_64x8m81_0
timestamp 1762296095
transform 1 0 25674 0 1 34822
box 0 0 1 1
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_0
timestamp 1762296095
transform 1 0 60601 0 1 35416
box 0 0 1 1
use M2_M14310589983211_64x8m81  M2_M14310589983211_64x8m81_0
timestamp 1762296095
transform 1 0 25673 0 1 44250
box 0 0 1 1
use M2_M14310589983211_64x8m81  M2_M14310589983211_64x8m81_1
timestamp 1762296095
transform 1 0 59150 0 1 44250
box 0 0 1 1
use M2_M14310589983215_64x8m81  M2_M14310589983215_64x8m81_0
timestamp 1762296095
transform 1 0 48818 0 1 811
box 0 0 1 1
use M2_M14310589983215_64x8m81  M2_M14310589983215_64x8m81_1
timestamp 1762296095
transform 1 0 27599 0 1 34726
box 0 0 1 1
use M2_M14310589983217_64x8m81  M2_M14310589983217_64x8m81_0
timestamp 1762296095
transform 0 -1 29813 1 0 784
box 0 0 1 1
use M2_M14310589983217_64x8m81  M2_M14310589983217_64x8m81_1
timestamp 1762296095
transform 0 -1 29116 1 0 784
box 0 0 1 1
use M2_M14310589983218_64x8m81  M2_M14310589983218_64x8m81_0
timestamp 1762296095
transform 1 0 53933 0 1 824
box 0 0 1 1
use m2m3_64x8m81  m2m3_64x8m81_0
timestamp 1762296095
transform 1 0 58611 0 1 17122
box 0 0 3541 9202
use M3_M2$$201248812_64x8m81  M3_M2$$201248812_64x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 12783
box 0 0 1 1
use M3_M2$$201248812_64x8m81  M3_M2$$201248812_64x8m81_1
timestamp 1762296095
transform -1 0 57515 0 1 15671
box 0 0 1 1
use M3_M2$$201248812_64x8m81  M3_M2$$201248812_64x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 15463
box 0 0 1 1
use M3_M2$$201248812_64x8m81  M3_M2$$201248812_64x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 13112
box 0 0 1 1
use M3_M2$$201249836_64x8m81  M3_M2$$201249836_64x8m81_0
timestamp 1762296095
transform -1 0 57515 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_64x8m81  M3_M2$$201249836_64x8m81_1
timestamp 1762296095
transform -1 0 58130 0 1 8835
box 0 0 1 1
use M3_M2$$201249836_64x8m81  M3_M2$$201249836_64x8m81_2
timestamp 1762296095
transform 1 0 27608 0 1 10834
box 0 0 1 1
use M3_M2$$201249836_64x8m81  M3_M2$$201249836_64x8m81_3
timestamp 1762296095
transform 1 0 26993 0 1 8835
box 0 0 1 1
use M3_M2$$201250860_64x8m81  M3_M2$$201250860_64x8m81_0
timestamp 1762296095
transform -1 0 56505 0 1 6590
box 0 0 1 1
use M3_M2$$201250860_64x8m81  M3_M2$$201250860_64x8m81_1
timestamp 1762296095
transform 1 0 28618 0 1 6590
box 0 0 1 1
use M3_M2$$201251884_64x8m81  M3_M2$$201251884_64x8m81_0
timestamp 1762296095
transform 1 0 37303 0 1 35853
box 0 0 1 1
use M3_M2$$201252908_64x8m81  M3_M2$$201252908_64x8m81_0
timestamp 1762296095
transform 1 0 28829 0 1 3700
box 0 0 1 1
use M3_M2$$201254956_64x8m81  M3_M2$$201254956_64x8m81_0
timestamp 1762296095
transform 1 0 27608 0 1 13768
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_0
timestamp 1762296095
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_1
timestamp 1762296095
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_2
timestamp 1762296095
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_3
timestamp 1762296095
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_4
timestamp 1762296095
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_5
timestamp 1762296095
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_6
timestamp 1762296095
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_7
timestamp 1762296095
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_8
timestamp 1762296095
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_64x8m81  M3_M2$$201258028_64x8m81_9
timestamp 1762296095
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M3_M2$$201412652_64x8m81  M3_M2$$201412652_64x8m81_0
timestamp 1762296095
transform 1 0 27608 0 1 32786
box 0 0 1 1
use M3_M2$$201412652_64x8m81  M3_M2$$201412652_64x8m81_1
timestamp 1762296095
transform 1 0 27608 0 1 30897
box 0 0 1 1
use M3_M2$$201412652_64x8m81  M3_M2$$201412652_64x8m81_2
timestamp 1762296095
transform -1 0 57515 0 1 30897
box 0 0 1 1
use M3_M2$$201412652_64x8m81  M3_M2$$201412652_64x8m81_3
timestamp 1762296095
transform -1 0 57515 0 1 32786
box 0 0 1 1
use M3_M2$$201413676_64x8m81  M3_M2$$201413676_64x8m81_0
timestamp 1762296095
transform 1 0 27608 0 1 7289
box 0 0 1 1
use M3_M2$$201413676_64x8m81  M3_M2$$201413676_64x8m81_1
timestamp 1762296095
transform 1 0 26993 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_64x8m81  M3_M2$$201413676_64x8m81_2
timestamp 1762296095
transform -1 0 58130 0 1 31842
box 0 0 1 1
use M3_M2$$201414700_64x8m81  M3_M2$$201414700_64x8m81_0
timestamp 1762296095
transform 1 0 26993 0 1 33221
box 0 0 1 1
use M3_M2$$201414700_64x8m81  M3_M2$$201414700_64x8m81_1
timestamp 1762296095
transform -1 0 58130 0 1 33221
box 0 0 1 1
use M3_M2$$201415724_64x8m81  M3_M2$$201415724_64x8m81_0
timestamp 1762296095
transform 1 0 26993 0 1 28743
box 0 0 1 1
use M3_M2$$201415724_64x8m81  M3_M2$$201415724_64x8m81_1
timestamp 1762296095
transform -1 0 58130 0 1 28743
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_0
timestamp 1762296095
transform -1 0 58130 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_1
timestamp 1762296095
transform -1 0 57515 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_2
timestamp 1762296095
transform -1 0 58130 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_3
timestamp 1762296095
transform -1 0 57515 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_4
timestamp 1762296095
transform 1 0 27608 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_5
timestamp 1762296095
transform 1 0 26993 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_6
timestamp 1762296095
transform 1 0 27608 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_7
timestamp 1762296095
transform 1 0 26993 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_8
timestamp 1762296095
transform 1 0 27608 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_9
timestamp 1762296095
transform 1 0 27608 0 1 24891
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_10
timestamp 1762296095
transform -1 0 57515 0 1 26662
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_0
timestamp 1762296095
transform 0 -1 49977 1 0 8925
box 0 0 1 1
use M3_M2431058998321_64x8m81  M3_M2431058998321_64x8m81_1
timestamp 1762296095
transform 1 0 51794 0 1 9891
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_0
timestamp 1762296095
transform 1 0 58128 0 1 20490
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_1
timestamp 1762296095
transform 1 0 58128 0 1 20146
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_2
timestamp 1762296095
transform 1 0 25851 0 1 18947
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_3
timestamp 1762296095
transform 1 0 26187 0 1 19267
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_4
timestamp 1762296095
transform 1 0 26545 0 1 19612
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_5
timestamp 1762296095
transform 1 0 24149 0 1 17237
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_6
timestamp 1762296095
transform 1 0 27004 0 1 20490
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_7
timestamp 1762296095
transform 1 0 24509 0 1 17576
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_8
timestamp 1762296095
transform 1 0 27004 0 1 20146
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_9
timestamp 1762296095
transform 1 0 24837 0 1 17897
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_10
timestamp 1762296095
transform 1 0 25174 0 1 18270
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_11
timestamp 1762296095
transform 1 0 25514 0 1 18604
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_12
timestamp 1762296095
transform 1 0 25836 0 1 25567
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_13
timestamp 1762296095
transform 1 0 26172 0 1 25887
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_14
timestamp 1762296095
transform 1 0 26530 0 1 26206
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_15
timestamp 1762296095
transform 1 0 24137 0 1 23593
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_16
timestamp 1762296095
transform 1 0 24496 0 1 23915
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_17
timestamp 1762296095
transform 1 0 24824 0 1 24236
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_18
timestamp 1762296095
transform 1 0 25161 0 1 24557
box 0 0 1 1
use M3_M2431058998325_64x8m81  M3_M2431058998325_64x8m81_19
timestamp 1762296095
transform 1 0 25501 0 1 25248
box 0 0 1 1
use M3_M2431058998326_64x8m81  M3_M2431058998326_64x8m81_0
timestamp 1762296095
transform 1 0 26990 0 1 23631
box 0 0 1 1
use M3_M2431058998327_64x8m81  M3_M2431058998327_64x8m81_0
timestamp 1762296095
transform 1 0 27599 0 1 34726
box 0 0 1 1
use M3_M2431058998328_64x8m81  M3_M2431058998328_64x8m81_0
timestamp 1762296095
transform 1 0 43880 0 1 3016
box 0 0 1 1
use M3_M24310589983210_64x8m81  M3_M24310589983210_64x8m81_0
timestamp 1762296095
transform 1 0 25674 0 1 30641
box 0 0 1 1
use M3_M24310589983210_64x8m81  M3_M24310589983210_64x8m81_1
timestamp 1762296095
transform 1 0 25674 0 1 34725
box 0 0 1 1
use M3_M24310589983210_64x8m81  M3_M24310589983210_64x8m81_2
timestamp 1762296095
transform 1 0 25674 0 1 31096
box 0 0 1 1
use M3_M24310589983210_64x8m81  M3_M24310589983210_64x8m81_3
timestamp 1762296095
transform 1 0 59149 0 1 30701
box 0 0 1 1
use M3_M24310589983210_64x8m81  M3_M24310589983210_64x8m81_4
timestamp 1762296095
transform 1 0 59149 0 1 31146
box 0 0 1 1
use M3_M24310589983212_64x8m81  M3_M24310589983212_64x8m81_0
timestamp 1762296095
transform 1 0 26990 0 1 36128
box 0 0 1 1
use M3_M24310589983212_64x8m81  M3_M24310589983212_64x8m81_1
timestamp 1762296095
transform 1 0 26990 0 1 43327
box 0 0 1 1
use M3_M24310589983213_64x8m81  M3_M24310589983213_64x8m81_0
timestamp 1762296095
transform 1 0 57538 0 1 8038
box 0 0 1 1
use M3_M24310589983214_64x8m81  M3_M24310589983214_64x8m81_0
timestamp 1762296095
transform 1 0 49313 0 1 1991
box 0 0 1 1
use M3_M24310589983214_64x8m81  M3_M24310589983214_64x8m81_1
timestamp 1762296095
transform 1 0 48823 0 1 2670
box 0 0 1 1
use M3_M24310589983219_64x8m81  M3_M24310589983219_64x8m81_0
timestamp 1762296095
transform 1 0 25680 0 1 27386
box 0 0 1 1
use M3_M24310589983219_64x8m81  M3_M24310589983219_64x8m81_1
timestamp 1762296095
transform 1 0 59135 0 1 27376
box 0 0 1 1
use M3_M24310589983221_64x8m81  M3_M24310589983221_64x8m81_0
timestamp 1762296095
transform 1 0 57495 0 1 22479
box 0 0 1 1
use M3_M24310589983221_64x8m81  M3_M24310589983221_64x8m81_1
timestamp 1762296095
transform 1 0 27607 0 1 22492
box 0 0 1 1
use M3_M24310589983221_64x8m81  M3_M24310589983221_64x8m81_2
timestamp 1762296095
transform 1 0 58126 0 1 23631
box 0 0 1 1
use M3_M24310589983224_64x8m81  M3_M24310589983224_64x8m81_0
timestamp 1762296095
transform 1 0 25673 0 1 44224
box 0 0 1 1
use M3_M24310589983224_64x8m81  M3_M24310589983224_64x8m81_1
timestamp 1762296095
transform 1 0 59150 0 1 44224
box 0 0 1 1
use power_a_64x8m81  power_a_64x8m81_0
timestamp 1762296095
transform -1 0 70018 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_1
timestamp 1762296095
transform -1 0 80818 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_2
timestamp 1762296095
transform 1 0 64218 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_3
timestamp 1762296095
transform 1 0 43633 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_4
timestamp 1762296095
transform 1 0 46033 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_5
timestamp 1762296095
transform 1 0 51233 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_6
timestamp 1762296095
transform 1 0 75018 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_7
timestamp 1762296095
transform 1 0 52478 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_8
timestamp 1762296095
transform -1 0 34022 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_9
timestamp 1762296095
transform -1 0 10442 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_10
timestamp 1762296095
transform -1 0 21242 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_11
timestamp 1762296095
transform 1 0 41233 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_12
timestamp 1762296095
transform 1 0 38028 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_13
timestamp 1762296095
transform 1 0 15442 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_14
timestamp 1762296095
transform 1 0 34831 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_15
timestamp 1762296095
transform 1 0 4642 0 1 282
box 0 -282 1000 1000
use power_a_64x8m81  power_a_64x8m81_16
timestamp 1762296095
transform -1 0 32324 0 1 282
box 0 -282 1000 1000
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_0
timestamp 1762296095
transform 1 0 10048 0 1 44146
box -511 630 1714 2430
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_1
timestamp 1762296095
transform 1 0 15448 0 1 44146
box -511 630 1714 2430
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_2
timestamp 1762296095
transform 1 0 4648 0 1 44146
box -511 630 1714 2430
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_3
timestamp 1762296095
transform 1 0 46824 0 1 44146
box -511 630 1714 2430
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_4
timestamp 1762296095
transform 1 0 64224 0 1 44146
box -511 630 1714 2430
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_5
timestamp 1762296095
transform 1 0 69624 0 1 44146
box -511 630 1714 2430
use power_route_01_a_64x8m81  power_route_01_a_64x8m81_6
timestamp 1762296095
transform 1 0 75024 0 1 44146
box -511 630 1714 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_0
timestamp 1762296095
transform -1 0 21142 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_1
timestamp 1762296095
transform -1 0 41719 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_2
timestamp 1762296095
transform -1 0 31199 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_3
timestamp 1762296095
transform -1 0 35904 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_4
timestamp 1762296095
transform -1 0 39074 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_5
timestamp 1762296095
transform -1 0 27061 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_6
timestamp 1762296095
transform -1 0 45558 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_7
timestamp 1762296095
transform -1 0 80718 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_8
timestamp 1762296095
transform -1 0 85155 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_9
timestamp 1762296095
transform -1 0 49390 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_10
timestamp 1762296095
transform -1 0 54751 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_11
timestamp 1762296095
transform -1 0 53058 0 1 44146
box -511 630 489 2430
use power_route_01_b_64x8m81  power_route_01_b_64x8m81_12
timestamp 1762296095
transform -1 0 58036 0 1 44146
box -511 630 489 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_0
timestamp 1762296095
transform -1 0 30987 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_1
timestamp 1762296095
transform -1 0 34095 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_2
timestamp 1762296095
transform -1 0 38662 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_3
timestamp 1762296095
transform -1 0 35738 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_4
timestamp 1762296095
transform -1 0 41596 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_5
timestamp 1762296095
transform -1 0 26872 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_6
timestamp 1762296095
transform -1 0 29591 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_7
timestamp 1762296095
transform -1 0 45427 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_8
timestamp 1762296095
transform -1 0 52179 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_9
timestamp 1762296095
transform -1 0 57704 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_10
timestamp 1762296095
transform -1 0 60505 0 1 44146
box 714 1822 1714 2430
use power_route_01_c_64x8m81  power_route_01_c_64x8m81_11
timestamp 1762296095
transform -1 0 44144 0 1 44146
box 714 1822 1714 2430
use power_route_64_64x8m81  power_route_64_64x8m81_0
timestamp 1762296095
transform 1 0 -1921 0 1 -2063
box 1921 2345 88293 48639
use rcol4_64_64x8m81  rcol4_64_64x8m81_0
timestamp 1762296095
transform 1 0 60511 0 1 5019
box -1090 -3394 25315 39307
use xdec8_64_64x8m81  xdec8_64_64x8m81_0
timestamp 1762296095
transform 1 0 28677 0 1 36127
box 155 -1 27614 8160
<< labels >>
flabel metal3 s 2626 45968 3626 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 42976 1706 43676 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 4642 0 5642 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 5362 45968 6362 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 8026 45968 9026 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 9442 0 10442 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 10762 45968 11762 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 13426 45968 14426 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 15442 0 16442 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 16162 45968 17162 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 18826 45968 19826 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 20242 0 21242 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 41176 1706 41876 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 39376 1706 40076 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 22258 45968 23258 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 25158 45968 26158 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 37576 1706 38276 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 35776 1706 36476 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 8152 1014 9515 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 8152 3011 9514 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 2226 8154 28729 9515 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 8153 24250 9514 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 28178 7084 28729 9516 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 1954 26433 2279 28416 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 24047 8154 28729 9516 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 12754 26433 13079 28416 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 29537 6744 34622 7652 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 28178 7084 34622 7652 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 1401 44776 2401 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 4137 44776 5137 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 6801 44776 7801 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 26435 26070 28416 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 9537 44776 10537 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 12201 44776 13201 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 14937 44776 15937 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 17601 44776 18601 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 20653 44776 21653 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 1271 26434 27828 26890 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 10176 3011 11493 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 2249 10174 24250 11491 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 2229 10175 24250 11491 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 24047 10176 27828 11493 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 34536 1014 35326 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 23483 44776 24483 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 26572 44776 27572 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 30710 44776 31710 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 35126 24920 35326 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 35415 44776 36415 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 34536 25085 35016 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 24942 34490 27830 34962 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 27877 45968 28877 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 29273 45968 30273 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 38585 44776 39585 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 31324 0 32324 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 32381 45968 33381 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 33022 0 34022 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 41230 44776 42230 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 45069 44776 46069 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 46313 44776 47313 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 34024 45968 35024 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 34831 0 35831 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 48901 44776 49901 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 52569 44776 53569 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 36948 45968 37948 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 54262 44776 55262 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 38028 0 39028 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 39882 45968 40882 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 57547 44776 58547 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 41233 0 42233 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 60977 44776 61977 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 42430 45968 43430 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 43633 0 44633 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 43713 45968 44713 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 63713 44776 64713 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 46033 0 47033 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 66377 44776 67377 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 47538 45968 48538 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 69113 44776 70113 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 50465 45968 51465 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 71777 44776 72777 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 74513 44776 75513 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 51233 0 52233 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 77177 44776 78177 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 52478 0 53478 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 80229 44776 81229 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 55990 45968 56990 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 83059 44776 84059 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 58791 45968 59791 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 84666 44776 85666 46576 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 44776 86372 45776 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 84666 42976 86372 43676 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 84666 41176 86372 41876 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 84666 39376 86372 40076 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 62202 45968 63202 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 84666 37576 86372 38276 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 84666 35776 86372 36476 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 64218 0 65218 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 29430 1706 34125 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 64938 45968 65938 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 67602 45968 68602 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 69018 0 70018 932 0 FreeSans 448 180 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 70338 45968 71338 46576 0 FreeSans 448 180 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 73002 45968 74002 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 75018 0 76018 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 75738 45968 76738 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 2095 32315 2188 34126 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 78402 45968 79402 46576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 79818 0 80818 932 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 32315 3011 34125 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 32316 25085 34125 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 81834 45968 82834 46576 0 FreeSans 448 180 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 43876 1014 44576 0 FreeSans 448 180 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 32318 27214 34124 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 26772 31486 58351 32199 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 26772 27382 58351 30105 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 57908 31486 58351 34124 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 61853 32315 72383 34125 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 57908 32315 86372 34124 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 29430 86372 29714 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 84666 29430 86372 34125 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 72653 32315 86372 34125 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 22938 1706 23938 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 22938 27214 23380 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 26770 23370 58348 24278 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 57908 22937 83763 23380 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 57908 22938 86372 23380 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 84666 22938 86372 23938 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 18016 24250 20739 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 29513 19969 55645 21625 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 29521 19969 55645 21707 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 44432 19969 55645 21708 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 44076 27779 44376 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 61825 18015 83763 20739 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 61807 18016 86372 20739 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 19969 86372 20739 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 12036 1706 14178 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 23821 12046 34761 12847 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 13461 27214 14178 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 30402 44126 54622 44328 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 12036 24250 12846 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 24047 12046 27214 14179 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 44127 86372 44328 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 24047 12046 34761 12934 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 34904 9972 41353 12606 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 29478 10756 41353 12606 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 29478 11697 58351 12606 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 26772 11844 58351 12606 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 50228 12035 58421 13866 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 59826 12035 60026 14017 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 50228 13461 86372 13866 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 61807 13461 72429 14178 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 61773 13461 86372 14177 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 57051 44076 86372 44376 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 85358 43876 86372 44576 0 FreeSans 448 180 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 42076 1014 42776 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 42276 27272 42576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 83169 12035 84221 12847 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 83169 13461 84221 14179 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 50228 12036 86372 12846 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 26772 12035 84999 12606 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 30403 42326 54622 42528 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 42327 86372 42528 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 59421 42276 86372 42576 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 84666 12036 86372 14178 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 72607 13461 86372 14178 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 61802 8153 86372 9514 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 85358 42076 86372 42776 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 57909 8154 62278 9516 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 57909 8154 72434 9515 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 0 40276 1014 40976 0 FreeSans 448 180 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 0 40476 27272 40776 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 30403 40526 54622 40728 0 FreeSans 448 0 0 0 VSS
port 27 nsew ground bidirectional
flabel metal3 s 72602 8152 83234 9515 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 61825 8152 86372 9514 0 FreeSans 448 180 0 0 VDD
port 26 nsew power bidirectional
flabel metal3 s 85358 8152 86372 9515 0 FreeSans 448 0 0 0 VDD
port 26 nsew power bidirectional
rlabel metal2 s 27936 0 28160 200 4 CLK
port 8 nsew signal input
rlabel metal2 s 1864 0 2088 200 4 D[0]
port 16 nsew signal input
rlabel metal2 s 30859 0 31083 200 4 A[2]
port 4 nsew signal input
rlabel metal2 s 32552 0 32776 200 4 A[1]
port 5 nsew signal input
rlabel metal2 s 34243 0 34467 200 4 A[0]
port 6 nsew signal input
rlabel metal2 s 14127 0 14351 200 4 Q[2]
port 23 nsew signal output
rlabel metal2 s 22279 0 22503 200 4 Q[3]
port 22 nsew signal output
rlabel metal2 s 50342 0 50566 200 4 CEN
port 7 nsew signal input
rlabel metal2 s 54417 0 54641 200 4 A[5]
port 1 nsew signal input
rlabel metal2 s 55164 0 55388 200 4 A[4]
port 2 nsew signal input
rlabel metal2 s 23404 0 23628 200 4 WEN[3]
port 32 nsew signal input
rlabel metal2 s 83372 0 83596 200 4 D[7]
port 9 nsew signal input
rlabel metal2 s 81855 0 82079 200 4 Q[7]
port 18 nsew signal output
rlabel metal2 s 23795 0 24019 200 4 D[3]
port 13 nsew signal input
rlabel metal2 s 12206 0 12430 200 4 D[1]
port 15 nsew signal input
rlabel metal2 s 13454 0 13678 200 4 D[2]
port 14 nsew signal input
rlabel metal2 s 56265 0 56489 200 4 A[3]
port 3 nsew signal input
rlabel metal2 s 11533 0 11757 200 4 Q[1]
port 24 nsew signal output
rlabel metal2 s 73703 0 73927 200 4 Q[6]
port 19 nsew signal output
rlabel metal2 s 71782 0 72006 200 4 D[5]
port 11 nsew signal input
rlabel metal2 s 62958 0 63182 200 4 Q[4]
port 21 nsew signal output
rlabel metal2 s 72180 0 72404 200 4 WEN[5]
port 30 nsew signal input
rlabel metal2 s 13054 0 13278 200 4 WEN[2]
port 33 nsew signal input
rlabel metal2 s 12604 0 12828 200 4 WEN[1]
port 34 nsew signal input
rlabel metal2 s 62115 0 62339 200 4 WEN[4]
port 31 nsew signal input
rlabel metal2 s 82695 0 82919 200 4 WEN[7]
port 28 nsew signal input
rlabel metal2 s 72630 0 72854 200 4 WEN[6]
port 29 nsew signal input
rlabel metal2 s 61447 0 61671 200 4 D[4]
port 12 nsew signal input
rlabel metal2 s 73030 0 73254 200 4 D[6]
port 10 nsew signal input
rlabel metal2 s 71109 0 71333 200 4 Q[5]
port 20 nsew signal output
rlabel metal2 s 3380 0 3604 200 4 Q[0]
port 25 nsew signal output
rlabel metal2 s 40588 0 40812 200 4 GWEN
port 17 nsew signal input
rlabel metal2 s 2539 0 2763 200 4 WEN[0]
port 35 nsew signal input
rlabel metal3 s 0 4060 1712 5629 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 5173 3011 5629 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 5174 24250 5629 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 4060 24341 4515 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 1 VDD
port 26 nsew power bidirectional
rlabel metal3 s 0 40527 86372 40728 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 38727 86372 38928 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 36927 86372 37128 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60549 35086 60639 35370 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60510 34490 61754 34962 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60549 35158 86372 35298 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61311 34536 86372 35016 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 34536 86372 35326 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 83360 35126 86372 35326 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61530 26433 61855 28416 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 72330 26433 72655 28416 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61530 26434 84717 28416 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28416 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27387 22291 57677 23199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 7088 57736 9012 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 59309 6982 86372 7595 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 7088 62747 7596 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 2502 1000 3772 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 1 VSS
port 27 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 1 VSS
port 27 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 46576
string GDS_END 2322396
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2272184
string LEFclass BLOCK
string LEFsymmetry X Y R90
string path 377.590 4.660 377.590 0.000 
<< end >>
