magic
tech gf180mcuD
magscale 1 10
timestamp 1762296095
<< polysilicon >>
rect 22205 30706 22518 30725
rect 22205 30571 22453 30706
rect 22434 30566 22453 30571
rect 22499 30566 22518 30706
rect 22434 30547 22518 30566
rect 22205 29082 22573 29183
rect 22205 29036 22454 29082
rect 22500 29036 22573 29082
rect 22205 29029 22573 29036
rect 22381 28925 22573 29029
rect 22205 28918 22573 28925
rect 22205 28872 22454 28918
rect 22500 28872 22573 28918
rect 22205 28771 22573 28872
rect 22205 27282 22573 27383
rect 22205 27236 22454 27282
rect 22500 27236 22573 27282
rect 22205 27229 22573 27236
rect 22381 27125 22573 27229
rect 22205 27118 22573 27125
rect 22205 27072 22454 27118
rect 22500 27072 22573 27118
rect 22205 26971 22573 27072
rect 22205 25482 22573 25583
rect 22205 25436 22454 25482
rect 22500 25436 22573 25482
rect 22205 25429 22573 25436
rect 22381 25325 22573 25429
rect 22205 25318 22573 25325
rect 22205 25272 22454 25318
rect 22500 25272 22573 25318
rect 22205 25171 22573 25272
rect 22205 23682 22573 23783
rect 22205 23636 22454 23682
rect 22500 23636 22573 23682
rect 22205 23629 22573 23636
rect 22381 23525 22573 23629
rect 22205 23518 22573 23525
rect 22205 23472 22454 23518
rect 22500 23472 22573 23518
rect 22205 23371 22573 23472
rect 22205 21882 22573 21983
rect 22205 21836 22454 21882
rect 22500 21836 22573 21882
rect 22205 21829 22573 21836
rect 22381 21725 22573 21829
rect 22205 21718 22573 21725
rect 22205 21672 22454 21718
rect 22500 21672 22573 21718
rect 22205 21571 22573 21672
rect 22205 20082 22573 20183
rect 22205 20036 22454 20082
rect 22500 20036 22573 20082
rect 22205 20029 22573 20036
rect 22381 19925 22573 20029
rect 22205 19918 22573 19925
rect 22205 19872 22454 19918
rect 22500 19872 22573 19918
rect 22205 19771 22573 19872
rect 22205 18282 22573 18383
rect 22205 18236 22454 18282
rect 22500 18236 22573 18282
rect 22205 18229 22573 18236
rect 22381 18125 22573 18229
rect 22205 18118 22573 18125
rect 22205 18072 22454 18118
rect 22500 18072 22573 18118
rect 22205 17971 22573 18072
rect 22205 16482 22573 16583
rect 22205 16436 22454 16482
rect 22500 16436 22573 16482
rect 22205 16429 22573 16436
rect 22381 16325 22573 16429
rect 22205 16318 22573 16325
rect 22205 16272 22454 16318
rect 22500 16272 22573 16318
rect 22205 16171 22573 16272
rect 22205 14682 22573 14783
rect 22205 14636 22454 14682
rect 22500 14636 22573 14682
rect 22205 14629 22573 14636
rect 22381 14525 22573 14629
rect 22205 14518 22573 14525
rect 22205 14472 22454 14518
rect 22500 14472 22573 14518
rect 22205 14371 22573 14472
rect 22205 12882 22573 12983
rect 22205 12836 22454 12882
rect 22500 12836 22573 12882
rect 22205 12829 22573 12836
rect 22381 12725 22573 12829
rect 22205 12718 22573 12725
rect 22205 12672 22454 12718
rect 22500 12672 22573 12718
rect 22205 12571 22573 12672
rect 22205 11082 22573 11183
rect 22205 11036 22454 11082
rect 22500 11036 22573 11082
rect 22205 11029 22573 11036
rect 22381 10925 22573 11029
rect 22205 10918 22573 10925
rect 22205 10872 22454 10918
rect 22500 10872 22573 10918
rect 22205 10771 22573 10872
rect 22205 9282 22573 9383
rect 22205 9236 22454 9282
rect 22500 9236 22573 9282
rect 22205 9229 22573 9236
rect 22381 9125 22573 9229
rect 22205 9118 22573 9125
rect 22205 9072 22454 9118
rect 22500 9072 22573 9118
rect 22205 8971 22573 9072
rect 22205 7482 22573 7583
rect 22205 7436 22454 7482
rect 22500 7436 22573 7482
rect 22205 7429 22573 7436
rect 22381 7325 22573 7429
rect 22205 7318 22573 7325
rect 22205 7272 22454 7318
rect 22500 7272 22573 7318
rect 22205 7171 22573 7272
rect 22205 5682 22573 5783
rect 22205 5636 22454 5682
rect 22500 5636 22573 5682
rect 22205 5629 22573 5636
rect 22381 5525 22573 5629
rect 22205 5518 22573 5525
rect 22205 5472 22454 5518
rect 22500 5472 22573 5518
rect 22205 5371 22573 5472
rect 22205 3882 22573 3983
rect 22205 3836 22454 3882
rect 22500 3836 22573 3882
rect 22205 3829 22573 3836
rect 22381 3725 22573 3829
rect 22205 3718 22573 3725
rect 22205 3672 22454 3718
rect 22500 3672 22573 3718
rect 22205 3571 22573 3672
rect 22205 2082 22573 2183
rect 22205 2036 22454 2082
rect 22500 2036 22573 2082
rect 22205 2029 22573 2036
rect 22381 1925 22573 2029
rect 22205 1918 22573 1925
rect 22205 1872 22454 1918
rect 22500 1872 22573 1918
rect 22205 1771 22573 1872
rect 22381 522 22573 568
rect 22381 476 22454 522
rect 22500 476 22573 522
rect 22381 383 22573 476
rect 22205 358 22573 383
rect 22205 312 22454 358
rect 22500 312 22573 358
rect 22205 229 22573 312
<< polycontact >>
rect 22453 30566 22499 30706
rect 22454 29036 22500 29082
rect 22454 28872 22500 28918
rect 22454 27236 22500 27282
rect 22454 27072 22500 27118
rect 22454 25436 22500 25482
rect 22454 25272 22500 25318
rect 22454 23636 22500 23682
rect 22454 23472 22500 23518
rect 22454 21836 22500 21882
rect 22454 21672 22500 21718
rect 22454 20036 22500 20082
rect 22454 19872 22500 19918
rect 22454 18236 22500 18282
rect 22454 18072 22500 18118
rect 22454 16436 22500 16482
rect 22454 16272 22500 16318
rect 22454 14636 22500 14682
rect 22454 14472 22500 14518
rect 22454 12836 22500 12882
rect 22454 12672 22500 12718
rect 22454 11036 22500 11082
rect 22454 10872 22500 10918
rect 22454 9236 22500 9282
rect 22454 9072 22500 9118
rect 22454 7436 22500 7482
rect 22454 7272 22500 7318
rect 22454 5636 22500 5682
rect 22454 5472 22500 5518
rect 22454 3836 22500 3882
rect 22454 3672 22500 3718
rect 22454 2036 22500 2082
rect 22454 1872 22500 1918
rect 22454 476 22500 522
rect 22454 312 22500 358
<< metal1 >>
rect 22438 30706 22514 30717
rect 22438 30705 22453 30706
rect 22499 30705 22514 30706
rect 22438 30445 22450 30705
rect 22502 30445 22514 30705
rect 22438 30433 22514 30445
rect 22413 29110 22537 29150
rect 22413 29058 22449 29110
rect 22501 29058 22537 29110
rect 22413 29036 22454 29058
rect 22500 29036 22537 29058
rect 22413 28918 22537 29036
rect 22413 28892 22454 28918
rect 22500 28892 22537 28918
rect 22413 28840 22449 28892
rect 22501 28840 22537 28892
rect 22413 28800 22537 28840
rect 22413 27310 22537 27350
rect 22413 27258 22449 27310
rect 22501 27258 22537 27310
rect 22413 27236 22454 27258
rect 22500 27236 22537 27258
rect 22413 27118 22537 27236
rect 22413 27092 22454 27118
rect 22500 27092 22537 27118
rect 22413 27040 22449 27092
rect 22501 27040 22537 27092
rect 22413 27000 22537 27040
rect 22413 25514 22537 25554
rect 22413 25462 22449 25514
rect 22501 25462 22537 25514
rect 22413 25436 22454 25462
rect 22500 25436 22537 25462
rect 22413 25318 22537 25436
rect 22413 25296 22454 25318
rect 22500 25296 22537 25318
rect 22413 25244 22449 25296
rect 22501 25244 22537 25296
rect 22413 25204 22537 25244
rect 22413 23710 22537 23750
rect 22413 23658 22449 23710
rect 22501 23658 22537 23710
rect 22413 23636 22454 23658
rect 22500 23636 22537 23658
rect 22413 23518 22537 23636
rect 22413 23492 22454 23518
rect 22500 23492 22537 23518
rect 22413 23440 22449 23492
rect 22501 23440 22537 23492
rect 22413 23400 22537 23440
rect 22413 21914 22537 21954
rect 22413 21862 22449 21914
rect 22501 21862 22537 21914
rect 22413 21836 22454 21862
rect 22500 21836 22537 21862
rect 22413 21718 22537 21836
rect 22413 21696 22454 21718
rect 22500 21696 22537 21718
rect 22413 21644 22449 21696
rect 22501 21644 22537 21696
rect 22413 21604 22537 21644
rect 22413 20110 22537 20150
rect 22413 20058 22449 20110
rect 22501 20058 22537 20110
rect 22413 20036 22454 20058
rect 22500 20036 22537 20058
rect 22413 19918 22537 20036
rect 22413 19892 22454 19918
rect 22500 19892 22537 19918
rect 22413 19840 22449 19892
rect 22501 19840 22537 19892
rect 22413 19800 22537 19840
rect 22413 18314 22537 18354
rect 22413 18262 22449 18314
rect 22501 18262 22537 18314
rect 22413 18236 22454 18262
rect 22500 18236 22537 18262
rect 22413 18118 22537 18236
rect 22413 18096 22454 18118
rect 22500 18096 22537 18118
rect 22413 18044 22449 18096
rect 22501 18044 22537 18096
rect 22413 18004 22537 18044
rect 22413 16510 22537 16550
rect 22413 16458 22449 16510
rect 22501 16458 22537 16510
rect 22413 16436 22454 16458
rect 22500 16436 22537 16458
rect 22413 16318 22537 16436
rect 22413 16292 22454 16318
rect 22500 16292 22537 16318
rect 22413 16240 22449 16292
rect 22501 16240 22537 16292
rect 22413 16200 22537 16240
rect 22413 14714 22537 14754
rect 22413 14662 22449 14714
rect 22501 14662 22537 14714
rect 22413 14636 22454 14662
rect 22500 14636 22537 14662
rect 22413 14518 22537 14636
rect 22413 14496 22454 14518
rect 22500 14496 22537 14518
rect 22413 14444 22449 14496
rect 22501 14444 22537 14496
rect 22413 14404 22537 14444
rect 22413 12910 22537 12950
rect 22413 12858 22449 12910
rect 22501 12858 22537 12910
rect 22413 12836 22454 12858
rect 22500 12836 22537 12858
rect 22413 12718 22537 12836
rect 22413 12692 22454 12718
rect 22500 12692 22537 12718
rect 22413 12640 22449 12692
rect 22501 12640 22537 12692
rect 22413 12600 22537 12640
rect 22413 11114 22537 11154
rect 22413 11062 22449 11114
rect 22501 11062 22537 11114
rect 22413 11036 22454 11062
rect 22500 11036 22537 11062
rect 22413 10918 22537 11036
rect 22413 10896 22454 10918
rect 22500 10896 22537 10918
rect 22413 10844 22449 10896
rect 22501 10844 22537 10896
rect 22413 10804 22537 10844
rect 22413 9310 22537 9350
rect 22413 9258 22449 9310
rect 22501 9258 22537 9310
rect 22413 9236 22454 9258
rect 22500 9236 22537 9258
rect 22413 9118 22537 9236
rect 22413 9092 22454 9118
rect 22500 9092 22537 9118
rect 22413 9040 22449 9092
rect 22501 9040 22537 9092
rect 22413 9000 22537 9040
rect 22413 7514 22537 7554
rect 22413 7462 22449 7514
rect 22501 7462 22537 7514
rect 22413 7436 22454 7462
rect 22500 7436 22537 7462
rect 22413 7318 22537 7436
rect 22413 7296 22454 7318
rect 22500 7296 22537 7318
rect 22413 7244 22449 7296
rect 22501 7244 22537 7296
rect 22413 7204 22537 7244
rect 22413 5710 22537 5750
rect 22413 5658 22449 5710
rect 22501 5658 22537 5710
rect 22413 5636 22454 5658
rect 22500 5636 22537 5658
rect 22413 5518 22537 5636
rect 22413 5492 22454 5518
rect 22500 5492 22537 5518
rect 22413 5440 22449 5492
rect 22501 5440 22537 5492
rect 22413 5400 22537 5440
rect 22413 3914 22537 3954
rect 22413 3862 22449 3914
rect 22501 3862 22537 3914
rect 22413 3836 22454 3862
rect 22500 3836 22537 3862
rect 22413 3718 22537 3836
rect 22413 3696 22454 3718
rect 22500 3696 22537 3718
rect 22413 3644 22449 3696
rect 22501 3644 22537 3696
rect 22413 3604 22537 3644
rect 22413 2110 22537 2150
rect 22413 2058 22449 2110
rect 22501 2058 22537 2110
rect 22413 2036 22454 2058
rect 22500 2036 22537 2058
rect 22413 1918 22537 2036
rect 22413 1892 22454 1918
rect 22500 1892 22537 1918
rect 22413 1840 22449 1892
rect 22501 1840 22537 1892
rect 22413 1800 22537 1840
rect 22421 522 22533 559
rect 22421 476 22454 522
rect 22500 476 22533 522
rect 22421 469 22533 476
rect 22421 313 22447 469
rect 22499 358 22533 469
rect 22421 312 22454 313
rect 22500 312 22533 358
rect 22421 276 22533 312
<< via1 >>
rect 22450 30566 22453 30705
rect 22453 30566 22499 30705
rect 22499 30566 22502 30705
rect 22450 30445 22502 30566
rect 22449 29082 22501 29110
rect 22449 29058 22454 29082
rect 22454 29058 22500 29082
rect 22500 29058 22501 29082
rect 22449 28872 22454 28892
rect 22454 28872 22500 28892
rect 22500 28872 22501 28892
rect 22449 28840 22501 28872
rect 22449 27282 22501 27310
rect 22449 27258 22454 27282
rect 22454 27258 22500 27282
rect 22500 27258 22501 27282
rect 22449 27072 22454 27092
rect 22454 27072 22500 27092
rect 22500 27072 22501 27092
rect 22449 27040 22501 27072
rect 22449 25482 22501 25514
rect 22449 25462 22454 25482
rect 22454 25462 22500 25482
rect 22500 25462 22501 25482
rect 22449 25272 22454 25296
rect 22454 25272 22500 25296
rect 22500 25272 22501 25296
rect 22449 25244 22501 25272
rect 22449 23682 22501 23710
rect 22449 23658 22454 23682
rect 22454 23658 22500 23682
rect 22500 23658 22501 23682
rect 22449 23472 22454 23492
rect 22454 23472 22500 23492
rect 22500 23472 22501 23492
rect 22449 23440 22501 23472
rect 22449 21882 22501 21914
rect 22449 21862 22454 21882
rect 22454 21862 22500 21882
rect 22500 21862 22501 21882
rect 22449 21672 22454 21696
rect 22454 21672 22500 21696
rect 22500 21672 22501 21696
rect 22449 21644 22501 21672
rect 22449 20082 22501 20110
rect 22449 20058 22454 20082
rect 22454 20058 22500 20082
rect 22500 20058 22501 20082
rect 22449 19872 22454 19892
rect 22454 19872 22500 19892
rect 22500 19872 22501 19892
rect 22449 19840 22501 19872
rect 22449 18282 22501 18314
rect 22449 18262 22454 18282
rect 22454 18262 22500 18282
rect 22500 18262 22501 18282
rect 22449 18072 22454 18096
rect 22454 18072 22500 18096
rect 22500 18072 22501 18096
rect 22449 18044 22501 18072
rect 22449 16482 22501 16510
rect 22449 16458 22454 16482
rect 22454 16458 22500 16482
rect 22500 16458 22501 16482
rect 22449 16272 22454 16292
rect 22454 16272 22500 16292
rect 22500 16272 22501 16292
rect 22449 16240 22501 16272
rect 22449 14682 22501 14714
rect 22449 14662 22454 14682
rect 22454 14662 22500 14682
rect 22500 14662 22501 14682
rect 22449 14472 22454 14496
rect 22454 14472 22500 14496
rect 22500 14472 22501 14496
rect 22449 14444 22501 14472
rect 22449 12882 22501 12910
rect 22449 12858 22454 12882
rect 22454 12858 22500 12882
rect 22500 12858 22501 12882
rect 22449 12672 22454 12692
rect 22454 12672 22500 12692
rect 22500 12672 22501 12692
rect 22449 12640 22501 12672
rect 22449 11082 22501 11114
rect 22449 11062 22454 11082
rect 22454 11062 22500 11082
rect 22500 11062 22501 11082
rect 22449 10872 22454 10896
rect 22454 10872 22500 10896
rect 22500 10872 22501 10896
rect 22449 10844 22501 10872
rect 22449 9282 22501 9310
rect 22449 9258 22454 9282
rect 22454 9258 22500 9282
rect 22500 9258 22501 9282
rect 22449 9072 22454 9092
rect 22454 9072 22500 9092
rect 22500 9072 22501 9092
rect 22449 9040 22501 9072
rect 22449 7482 22501 7514
rect 22449 7462 22454 7482
rect 22454 7462 22500 7482
rect 22500 7462 22501 7482
rect 22449 7272 22454 7296
rect 22454 7272 22500 7296
rect 22500 7272 22501 7296
rect 22449 7244 22501 7272
rect 22449 5682 22501 5710
rect 22449 5658 22454 5682
rect 22454 5658 22500 5682
rect 22500 5658 22501 5682
rect 22449 5472 22454 5492
rect 22454 5472 22500 5492
rect 22500 5472 22501 5492
rect 22449 5440 22501 5472
rect 22449 3882 22501 3914
rect 22449 3862 22454 3882
rect 22454 3862 22500 3882
rect 22500 3862 22501 3882
rect 22449 3672 22454 3696
rect 22454 3672 22500 3696
rect 22500 3672 22501 3696
rect 22449 3644 22501 3672
rect 22449 2082 22501 2110
rect 22449 2058 22454 2082
rect 22454 2058 22500 2082
rect 22500 2058 22501 2082
rect 22449 1872 22454 1892
rect 22454 1872 22500 1892
rect 22500 1872 22501 1892
rect 22449 1840 22501 1872
rect 22447 358 22499 469
rect 22447 313 22454 358
rect 22454 313 22499 358
<< metal2 >>
rect 22412 30857 22537 30877
rect 22412 30697 22448 30857
rect 22504 30697 22537 30857
rect 22412 30445 22450 30697
rect 22502 30445 22537 30697
rect 22412 29110 22537 30445
rect 22412 29058 22449 29110
rect 22501 29058 22537 29110
rect 22412 28892 22537 29058
rect 22412 28840 22449 28892
rect 22501 28840 22537 28892
rect 22412 27310 22537 28840
rect 22412 27258 22449 27310
rect 22501 27258 22537 27310
rect 22412 27092 22537 27258
rect 22412 27040 22449 27092
rect 22501 27040 22537 27092
rect 22412 25514 22537 27040
rect 22412 25462 22449 25514
rect 22501 25462 22537 25514
rect 22412 25296 22537 25462
rect 22412 25244 22449 25296
rect 22501 25244 22537 25296
rect 22412 23710 22537 25244
rect 22412 23658 22449 23710
rect 22501 23658 22537 23710
rect 22412 23492 22537 23658
rect 22412 23440 22449 23492
rect 22501 23440 22537 23492
rect 22412 21914 22537 23440
rect 22412 21862 22449 21914
rect 22501 21862 22537 21914
rect 22412 21696 22537 21862
rect 22412 21644 22449 21696
rect 22501 21644 22537 21696
rect 22412 20110 22537 21644
rect 22412 20058 22449 20110
rect 22501 20058 22537 20110
rect 22412 19892 22537 20058
rect 22412 19840 22449 19892
rect 22501 19840 22537 19892
rect 22412 18314 22537 19840
rect 22412 18262 22449 18314
rect 22501 18262 22537 18314
rect 22412 18096 22537 18262
rect 22412 18044 22449 18096
rect 22501 18044 22537 18096
rect 22412 16510 22537 18044
rect 22412 16458 22449 16510
rect 22501 16458 22537 16510
rect 22412 16292 22537 16458
rect 22412 16240 22449 16292
rect 22501 16240 22537 16292
rect 22412 14714 22537 16240
rect 22412 14662 22449 14714
rect 22501 14662 22537 14714
rect 22412 14496 22537 14662
rect 22412 14444 22449 14496
rect 22501 14444 22537 14496
rect 22412 12910 22537 14444
rect 22412 12858 22449 12910
rect 22501 12858 22537 12910
rect 22412 12692 22537 12858
rect 22412 12640 22449 12692
rect 22501 12640 22537 12692
rect 22412 11114 22537 12640
rect 22412 11062 22449 11114
rect 22501 11062 22537 11114
rect 22412 10896 22537 11062
rect 22412 10844 22449 10896
rect 22501 10844 22537 10896
rect 22412 9310 22537 10844
rect 22412 9258 22449 9310
rect 22501 9258 22537 9310
rect 22412 9092 22537 9258
rect 22412 9040 22449 9092
rect 22501 9040 22537 9092
rect 22412 7514 22537 9040
rect 22412 7462 22449 7514
rect 22501 7462 22537 7514
rect 22412 7296 22537 7462
rect 22412 7244 22449 7296
rect 22501 7244 22537 7296
rect 22412 5710 22537 7244
rect 22412 5658 22449 5710
rect 22501 5658 22537 5710
rect 22412 5492 22537 5658
rect 22412 5440 22449 5492
rect 22501 5440 22537 5492
rect 22412 3914 22537 5440
rect 22412 3862 22449 3914
rect 22501 3862 22537 3914
rect 22412 3696 22537 3862
rect 22412 3644 22449 3696
rect 22501 3644 22537 3696
rect 22412 2110 22537 3644
rect 22412 2058 22449 2110
rect 22501 2058 22537 2110
rect 22412 1892 22537 2058
rect 22412 1840 22449 1892
rect 22501 1840 22537 1892
rect 22412 469 22537 1840
rect 22412 313 22447 469
rect 22499 313 22537 469
rect 22412 257 22537 313
rect 22412 97 22445 257
rect 22501 97 22537 257
rect 22412 76 22537 97
<< via2 >>
rect 22448 30705 22504 30857
rect 22448 30697 22450 30705
rect 22450 30697 22502 30705
rect 22502 30697 22504 30705
rect 22445 97 22501 257
<< metal3 >>
rect -636 30857 22538 30877
rect -636 30697 22448 30857
rect 22504 30697 22538 30857
rect -636 30677 22538 30697
rect -636 257 22537 277
rect -636 97 22445 257
rect 22501 97 22537 257
rect -636 77 22537 97
use 018SRAM_cell1_256x8m81  018SRAM_cell1_256x8m81_0
timestamp 1762296095
transform -1 0 22262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_256x8m81  018SRAM_cell1_256x8m81_1
timestamp 1762296095
transform -1 0 22262 0 -1 30777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_0
timestamp 1762296095
transform -1 0 22262 0 1 3777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_1
timestamp 1762296095
transform -1 0 22262 0 -1 5577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_2
timestamp 1762296095
transform -1 0 22262 0 -1 1977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_3
timestamp 1762296095
transform -1 0 22262 0 -1 14577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_4
timestamp 1762296095
transform -1 0 22262 0 -1 12777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_5
timestamp 1762296095
transform -1 0 22262 0 -1 10977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_6
timestamp 1762296095
transform -1 0 22262 0 1 5577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_7
timestamp 1762296095
transform -1 0 22262 0 1 12777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_8
timestamp 1762296095
transform -1 0 22262 0 -1 3777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_9
timestamp 1762296095
transform -1 0 22262 0 -1 7377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_10
timestamp 1762296095
transform -1 0 22262 0 -1 9177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_11
timestamp 1762296095
transform -1 0 22262 0 1 9177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_12
timestamp 1762296095
transform -1 0 22262 0 1 10977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_13
timestamp 1762296095
transform -1 0 22262 0 1 7377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_14
timestamp 1762296095
transform -1 0 22262 0 1 1977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_15
timestamp 1762296095
transform -1 0 22262 0 -1 19977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_16
timestamp 1762296095
transform -1 0 22262 0 1 16377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_17
timestamp 1762296095
transform -1 0 22262 0 1 28977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_18
timestamp 1762296095
transform -1 0 22262 0 1 25377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_19
timestamp 1762296095
transform -1 0 22262 0 1 27177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_20
timestamp 1762296095
transform -1 0 22262 0 1 23577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_21
timestamp 1762296095
transform -1 0 22262 0 1 21777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_22
timestamp 1762296095
transform -1 0 22262 0 1 19977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_23
timestamp 1762296095
transform -1 0 22262 0 1 18177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_24
timestamp 1762296095
transform -1 0 22262 0 -1 21777
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_25
timestamp 1762296095
transform -1 0 22262 0 -1 25377
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_26
timestamp 1762296095
transform -1 0 22262 0 -1 23577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_27
timestamp 1762296095
transform -1 0 22262 0 -1 27177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_28
timestamp 1762296095
transform -1 0 22262 0 -1 28977
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_29
timestamp 1762296095
transform -1 0 22262 0 -1 18177
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_30
timestamp 1762296095
transform -1 0 22262 0 1 14577
box -68 -68 668 968
use 018SRAM_cell1_cutPC_256x8m81  018SRAM_cell1_cutPC_256x8m81_31
timestamp 1762296095
transform -1 0 22262 0 -1 16377
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_0
timestamp 1762296095
transform -1 0 16862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_1
timestamp 1762296095
transform -1 0 17462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_2
timestamp 1762296095
transform -1 0 18662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_3
timestamp 1762296095
transform -1 0 18062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_4
timestamp 1762296095
transform -1 0 19262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_5
timestamp 1762296095
transform -1 0 19862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_6
timestamp 1762296095
transform -1 0 20462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_7
timestamp 1762296095
transform -1 0 21062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_8
timestamp 1762296095
transform -1 0 15662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_9
timestamp 1762296095
transform -1 0 15062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_10
timestamp 1762296095
transform -1 0 14462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_11
timestamp 1762296095
transform -1 0 13862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_12
timestamp 1762296095
transform -1 0 12662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_13
timestamp 1762296095
transform -1 0 13262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_14
timestamp 1762296095
transform -1 0 12062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_15
timestamp 1762296095
transform -1 0 3662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_16
timestamp 1762296095
transform -1 0 3062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_17
timestamp 1762296095
transform -1 0 1862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_18
timestamp 1762296095
transform -1 0 2462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_19
timestamp 1762296095
transform -1 0 1262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_20
timestamp 1762296095
transform -1 0 662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_21
timestamp 1762296095
transform -1 0 6062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_22
timestamp 1762296095
transform -1 0 6662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_23
timestamp 1762296095
transform -1 0 7862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_24
timestamp 1762296095
transform -1 0 7262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_25
timestamp 1762296095
transform -1 0 8462 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_26
timestamp 1762296095
transform -1 0 9062 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_27
timestamp 1762296095
transform -1 0 9662 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_28
timestamp 1762296095
transform -1 0 10262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_29
timestamp 1762296095
transform -1 0 4862 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_30
timestamp 1762296095
transform -1 0 4262 0 1 177
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_31
timestamp 1762296095
transform -1 0 11462 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_0
timestamp 1762296095
transform -1 0 16262 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_1
timestamp 1762296095
transform 1 0 21062 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_2
timestamp 1762296095
transform -1 0 5462 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_3
timestamp 1762296095
transform -1 0 62 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_4
timestamp 1762296095
transform -1 0 10862 0 1 177
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_5
timestamp 1762296095
transform -1 0 62 0 -1 30777
box -68 -68 668 968
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_0
timestamp 1762296095
transform 1 0 22477 0 -1 417
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_1
timestamp 1762296095
transform 1 0 22477 0 -1 12777
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_2
timestamp 1762296095
transform 1 0 22477 0 -1 9177
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_3
timestamp 1762296095
transform 1 0 22477 0 -1 14577
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_4
timestamp 1762296095
transform 1 0 22477 0 -1 10977
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_5
timestamp 1762296095
transform 1 0 22477 0 -1 7377
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_6
timestamp 1762296095
transform 1 0 22477 0 -1 5577
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_7
timestamp 1762296095
transform 1 0 22477 0 -1 1977
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_8
timestamp 1762296095
transform 1 0 22477 0 -1 3777
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_9
timestamp 1762296095
transform 1 0 22477 0 -1 28977
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_10
timestamp 1762296095
transform 1 0 22477 0 -1 25377
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_11
timestamp 1762296095
transform 1 0 22477 0 -1 21777
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_12
timestamp 1762296095
transform 1 0 22477 0 -1 16377
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_13
timestamp 1762296095
transform 1 0 22477 0 -1 18177
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_14
timestamp 1762296095
transform 1 0 22477 0 -1 27177
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_15
timestamp 1762296095
transform 1 0 22477 0 -1 23577
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_16
timestamp 1762296095
transform 1 0 22477 0 -1 19977
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1762296095
transform 1 0 22476 0 1 30636
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1762296095
transform 1 0 22475 0 -1 14579
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1762296095
transform 1 0 22475 0 -1 3779
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1762296095
transform 1 0 22475 0 -1 10979
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1762296095
transform 1 0 22475 0 -1 1975
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_4
timestamp 1762296095
transform 1 0 22475 0 -1 5575
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_5
timestamp 1762296095
transform 1 0 22475 0 -1 9175
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_6
timestamp 1762296095
transform 1 0 22475 0 -1 12775
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_7
timestamp 1762296095
transform 1 0 22475 0 -1 7379
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_8
timestamp 1762296095
transform 1 0 22475 0 -1 21779
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_9
timestamp 1762296095
transform 1 0 22475 0 -1 28975
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_10
timestamp 1762296095
transform 1 0 22475 0 -1 18179
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_11
timestamp 1762296095
transform 1 0 22475 0 -1 25379
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_12
timestamp 1762296095
transform 1 0 22475 0 -1 16375
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_13
timestamp 1762296095
transform 1 0 22475 0 -1 19975
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_14
timestamp 1762296095
transform 1 0 22475 0 -1 23575
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_15
timestamp 1762296095
transform 1 0 22475 0 -1 27175
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_0
timestamp 1762296095
transform 1 0 22476 0 1 30575
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_0
timestamp 1762296095
transform 1 0 22473 0 1 391
box 0 0 1 1
use M3_M2431059087811_256x8m81  M3_M2431059087811_256x8m81_0
timestamp 1762296095
transform 1 0 22473 0 1 177
box 0 0 1 1
use M3_M2431059087811_256x8m81  M3_M2431059087811_256x8m81_1
timestamp 1762296095
transform 1 0 22476 0 1 30777
box 0 0 1 1
use new_dummyrow_unit_01_256x8m81  new_dummyrow_unit_01_256x8m81_0
timestamp 1762296095
transform 1 0 0 0 -1 30954
box -6 109 10930 1145
use new_dummyrow_unit_256x8m81  new_dummyrow_unit_256x8m81_0
timestamp 1762296095
transform 1 0 10800 0 -1 30954
box -6 109 10930 1145
<< labels >>
rlabel metal3 s 22196 1995 22196 1995 4 VSS
rlabel metal3 s 22196 1070 22196 1070 4 VDD
<< properties >>
string GDS_END 1790436
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1780714
<< end >>
